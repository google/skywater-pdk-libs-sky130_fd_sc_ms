* File: sky130_fd_sc_ms__o311a_1.pex.spice
* Created: Wed Sep  2 12:24:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O311A_1%C1 3 7 9 16
r27 15 16 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.525 $Y=1.305
+ $X2=0.58 $Y2=1.305
r28 12 15 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.27 $Y=1.305
+ $X2=0.525 $Y2=1.305
r29 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.305 $X2=0.27 $Y2=1.305
r30 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.14
+ $X2=0.58 $Y2=1.305
r31 5 7 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.58 $Y=1.14 $X2=0.58
+ $Y2=0.69
r32 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.47
+ $X2=0.525 $Y2=1.305
r33 1 3 375.105 $w=1.8e-07 $l=9.65e-07 $layer=POLY_cond $X=0.525 $Y=1.47
+ $X2=0.525 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%B1 3 7 9 12
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.305
+ $X2=1.06 $Y2=1.47
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.305
+ $X2=1.06 $Y2=1.14
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.305 $X2=1.06 $Y2=1.305
r38 9 13 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.305 $X2=1.06
+ $Y2=1.305
r39 7 15 375.105 $w=1.8e-07 $l=9.65e-07 $layer=POLY_cond $X=1.075 $Y=2.435
+ $X2=1.075 $Y2=1.47
r40 3 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.97 $Y=0.69 $X2=0.97
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%A2 3 7 10 11 12 15 16 18 21 31
c70 15 0 1.74145e-20 $X=2.68 $Y=1.61
c71 7 0 4.35611e-20 $X=2.605 $Y=2.435
c72 3 0 1.12678e-19 $X=1.51 $Y=0.69
r73 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.305
+ $X2=1.6 $Y2=1.14
r74 18 31 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.6 $Y=1.305 $X2=1.72
+ $Y2=1.305
r75 18 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.305 $X2=1.6 $Y2=1.305
r76 16 27 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.61
+ $X2=2.68 $Y2=1.775
r77 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.61 $X2=2.68 $Y2=1.61
r78 13 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.68 $Y=2.32 $X2=2.68
+ $Y2=1.61
r79 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.515 $Y=2.405
+ $X2=2.68 $Y2=2.32
r80 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.515 $Y=2.405
+ $X2=1.805 $Y2=2.405
r81 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=2.32
+ $X2=1.805 $Y2=2.405
r82 9 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=1.47 $X2=1.72
+ $Y2=1.305
r83 9 10 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.72 $Y=1.47 $X2=1.72
+ $Y2=2.32
r84 7 27 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.605 $Y=2.435
+ $X2=2.605 $Y2=1.775
r85 3 23 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.51 $Y=0.69 $X2=1.51
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%A3 1 3 4 5 7 10 11 12 13 18 20
c45 18 0 1.74145e-20 $X=2.14 $Y=1.285
c46 11 0 1.12678e-19 $X=2.16 $Y=1.295
r47 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.285
+ $X2=2.14 $Y2=1.45
r48 18 20 52.3316 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.14 $Y=1.285 $X2=2.14
+ $Y2=1.085
r49 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=2.035
r50 11 12 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.14 $Y=1.285
+ $X2=2.14 $Y2=1.665
r51 11 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.285 $X2=2.14 $Y2=1.285
r52 10 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.23 $Y=0.69
+ $X2=2.23 $Y2=1.085
r53 7 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.05 $Y=1.71 $X2=2.05
+ $Y2=1.45
r54 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.975 $Y=1.785
+ $X2=2.05 $Y2=1.71
r55 4 5 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.975 $Y=1.785
+ $X2=1.615 $Y2=1.785
r56 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.525 $Y=1.86
+ $X2=1.615 $Y2=1.785
r57 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.525 $Y=1.86
+ $X2=1.525 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%A1 3 7 8 11 12 13
c38 13 0 1.54042e-19 $X=3.22 $Y=1.12
c39 11 0 1.3462e-19 $X=3.22 $Y=1.285
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.285
+ $X2=3.22 $Y2=1.45
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.285
+ $X2=3.22 $Y2=1.12
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.285 $X2=3.22 $Y2=1.285
r43 8 12 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.12 $Y=1.285 $X2=3.22
+ $Y2=1.285
r44 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.31 $Y=0.69 $X2=3.31
+ $Y2=1.12
r45 3 14 382.879 $w=1.8e-07 $l=9.85e-07 $layer=POLY_cond $X=3.175 $Y=2.435
+ $X2=3.175 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%A_31_387# 1 2 3 12 16 20 26 29 30 31 33 35
+ 36 39 40 41 47 52 53
c122 52 0 1.25197e-19 $X=3.76 $Y=1.515
c123 41 0 4.35611e-20 $X=3.185 $Y=1.705
r124 53 59 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.515
+ $X2=3.76 $Y2=1.68
r125 53 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.515
+ $X2=3.76 $Y2=1.35
r126 52 55 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=3.745 $Y=1.515
+ $X2=3.745 $Y2=1.705
r127 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.515 $X2=3.76 $Y2=1.515
r128 40 55 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.595 $Y=1.705
+ $X2=3.745 $Y2=1.705
r129 40 41 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.595 $Y=1.705
+ $X2=3.185 $Y2=1.705
r130 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=1.79
+ $X2=3.185 $Y2=1.705
r131 38 39 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.1 $Y=1.79
+ $X2=3.1 $Y2=2.785
r132 37 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.87
+ $X2=1.3 $Y2=2.87
r133 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=2.87
+ $X2=3.1 $Y2=2.785
r134 36 37 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=3.015 $Y=2.87
+ $X2=1.465 $Y2=2.87
r135 33 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.785 $X2=1.3
+ $Y2=2.87
r136 33 35 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.3 $Y=2.785
+ $X2=1.3 $Y2=2.08
r137 32 35 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.3 $Y=1.81 $X2=1.3
+ $Y2=2.08
r138 31 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.725
+ $X2=0.665 $Y2=1.725
r139 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.135 $Y=1.725
+ $X2=1.3 $Y2=1.81
r140 30 31 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.135 $Y=1.725
+ $X2=0.75 $Y2=1.725
r141 29 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=1.64
+ $X2=0.665 $Y2=1.725
r142 28 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=0.97
+ $X2=0.665 $Y2=0.885
r143 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.665 $Y=0.97
+ $X2=0.665 $Y2=1.64
r144 24 47 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.365 $Y=0.885
+ $X2=0.665 $Y2=0.885
r145 24 26 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.365 $Y=0.8
+ $X2=0.365 $Y2=0.515
r146 20 22 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.3 $Y=2.08 $X2=0.3
+ $Y2=2.79
r147 18 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.3 $Y=1.725
+ $X2=0.665 $Y2=1.725
r148 18 20 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.3 $Y=1.81 $X2=0.3
+ $Y2=2.08
r149 16 58 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.82 $Y=0.74
+ $X2=3.82 $Y2=1.35
r150 12 59 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.795 $Y=2.4
+ $X2=3.795 $Y2=1.68
r151 3 50 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.935 $X2=1.3 $Y2=2.79
r152 3 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.935 $X2=1.3 $Y2=2.08
r153 2 22 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.935 $X2=0.3 $Y2=2.79
r154 2 20 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.935 $X2=0.3 $Y2=2.08
r155 1 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.37 $X2=0.365 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%VPWR 1 2 9 15 19 21 26 36 37 40 43
r42 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 37 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.52 $Y2=3.33
r47 34 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 27 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r54 27 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.52 $Y2=3.33
r56 26 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r60 21 23 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 19 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 19 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 15 18 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.52 $Y=2.125
+ $X2=3.52 $Y2=2.815
r64 13 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=3.33
r65 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.815
r66 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.8 $Y=2.11 $X2=0.8
+ $Y2=2.79
r67 7 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r68 7 12 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=2.79
r69 2 18 400 $w=1.7e-07 $l=9.994e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.935 $X2=3.52 $Y2=2.815
r70 2 15 400 $w=1.7e-07 $l=3.36861e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.935 $X2=3.52 $Y2=2.125
r71 1 12 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.935 $X2=0.8 $Y2=2.79
r72 1 9 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.935 $X2=0.8 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%X 1 2 9 14 15 16 17 28
c25 17 0 9.42383e-21 $X=3.995 $Y=0.84
c26 16 0 1.54042e-19 $X=4.08 $Y=0.555
r27 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=4.052 $Y=0.948
+ $X2=4.052 $Y2=0.925
r28 17 30 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=4.052 $Y=0.979
+ $X2=4.052 $Y2=1.13
r29 17 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=4.052 $Y=0.979
+ $X2=4.052 $Y2=0.948
r30 17 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=4.052 $Y=0.894
+ $X2=4.052 $Y2=0.925
r31 16 17 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=4.052 $Y=0.515
+ $X2=4.052 $Y2=0.894
r32 15 30 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.15 $Y=1.96
+ $X2=4.15 $Y2=1.13
r33 14 15 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=2.125
+ $X2=4.045 $Y2=1.96
r34 7 14 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.045 $Y=2.15
+ $X2=4.045 $Y2=2.125
r35 7 9 20.1678 $w=3.78e-07 $l=6.65e-07 $layer=LI1_cond $X=4.045 $Y=2.15
+ $X2=4.045 $Y2=2.815
r36 2 14 400 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.02 $Y2=2.125
r37 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.02 $Y2=2.815
r38 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.895
+ $Y=0.37 $X2=4.035 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%A_209_74# 1 2 7 9 13
r19 11 16 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0.445
+ $X2=1.225 $Y2=0.445
r20 11 13 56.7491 $w=3.28e-07 $l=1.625e-06 $layer=LI1_cond $X=1.39 $Y=0.445
+ $X2=3.015 $Y2=0.445
r21 7 16 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0.61
+ $X2=1.225 $Y2=0.445
r22 7 9 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.225 $Y=0.61
+ $X2=1.225 $Y2=0.855
r23 2 13 91 $w=1.7e-07 $l=7.83677e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.37 $X2=3.015 $Y2=0.525
r24 1 16 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.37 $X2=1.225 $Y2=0.515
r25 1 9 182 $w=1.7e-07 $l=5.67913e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.37 $X2=1.225 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_1%VGND 1 2 7 14 15 17 27 28 31
r47 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 28 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r49 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r50 25 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.525
+ $Y2=0
r51 25 27 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=4.08
+ $Y2=0
r52 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r53 23 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r54 19 23 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r55 19 20 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r56 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.525
+ $Y2=0
r57 17 23 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.12
+ $Y2=0
r58 15 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 15 20 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.24
+ $Y2=0
r60 12 14 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.525 $Y=0.78
+ $X2=3.525 $Y2=0.515
r61 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0
r62 11 14 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.515
r63 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.36 $Y=0.865
+ $X2=3.525 $Y2=0.78
r64 7 9 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=3.36 $Y=0.865
+ $X2=1.87 $Y2=0.865
r65 2 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.37 $X2=3.525 $Y2=0.515
r66 1 9 182 $w=1.7e-07 $l=6.21369e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.37 $X2=1.87 $Y2=0.865
.ends


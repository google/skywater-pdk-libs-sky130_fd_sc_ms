* File: sky130_fd_sc_ms__nand4bb_1.spice
* Created: Wed Sep  2 12:14:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4bb_1.pex.spice"
.subckt sky130_fd_sc_ms__nand4bb_1  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_N_M1002_g N_A_27_398#_M1002_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.122187 AS=0.150975 PD=1.025 PS=1.67 NRD=17.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1000 N_A_229_398#_M1000_d N_B_N_M1000_g N_VGND_M1002_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.15055 AS=0.122187 PD=1.69 PS=1.025 NRD=1.08 NRS=15.264 M=1
+ R=3.66667 SA=75000.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1009 A_435_74# N_A_27_398#_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.19585 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1001 A_513_74# N_A_229_398#_M1001_g A_435_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1011 A_627_74# N_C_M1011_g A_513_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75001.1
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g A_627_74# VNB NLOWVT L=0.15 W=0.74 AD=0.266
+ AS=0.1554 PD=2.34 PS=1.16 NRD=23.508 NRS=25.128 M=1 R=4.93333 SA=75001.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_A_N_M1010_g N_A_27_398#_M1010_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1006 N_A_229_398#_M1006_d N_B_N_M1006_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1554 PD=2.24 PS=1.21 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_398#_M1004_g N_Y_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2296 AS=0.3136 PD=1.53 PS=2.8 NRD=15.8191 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_A_229_398#_M1008_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2296 PD=1.44 PS=1.53 NRD=7.8997 NRS=7.0329 M=1 R=6.22222
+ SA=90000.8 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_C_M1007_g N_Y_M1008_d VPB PSHORT L=0.18 W=1.12 AD=0.2072
+ AS=0.1792 PD=1.49 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.3 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_D_M1005_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2072 PD=2.8 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.8 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__nand4bb_1.pxi.spice"
*
.ends
*
*

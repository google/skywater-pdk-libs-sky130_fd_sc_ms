* NGSPICE file created from sky130_fd_sc_ms__mux2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__mux2_1 A0 A1 S VGND VNB VPB VPWR X
M1000 a_304_74# A0 a_226_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=7.85e+11p ps=3.57e+06u
M1001 X a_304_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=8.226e+11p ps=5.83e+06u
M1002 a_443_74# A0 a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=3.1e+06u as=4.033e+11p ps=2.57e+06u
M1003 VPWR S a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 VPWR a_27_112# a_527_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1005 a_527_368# A1 a_304_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND S a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=7.0725e+11p pd=4.91e+06u as=1.5675e+11p ps=1.67e+06u
M1007 a_304_74# A1 a_226_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1008 a_226_74# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_112# a_443_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_304_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1011 a_226_368# S VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__mux2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.180000 2.275000 1.550000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.220000 1.685000 1.550000 ;
        RECT 1.515000 0.810000 2.785000 0.980000 ;
        RECT 1.515000 0.980000 1.685000 1.220000 ;
        RECT 2.455000 0.980000 2.785000 1.550000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.470000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.350000 0.835000 1.780000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795000 1.820000 4.235000 2.980000 ;
        RECT 3.865000 0.350000 4.235000 1.130000 ;
        RECT 4.065000 1.130000 4.235000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.540000 0.445000 1.130000 ;
      RECT 0.115000  1.130000 0.285000 1.950000 ;
      RECT 0.115000  1.950000 0.445000 2.060000 ;
      RECT 0.115000  2.060000 1.320000 2.230000 ;
      RECT 0.115000  2.230000 0.445000 2.700000 ;
      RECT 0.625000  0.085000 1.005000 0.680000 ;
      RECT 0.625000  0.680000 0.835000 1.130000 ;
      RECT 0.650000  2.400000 0.980000 3.245000 ;
      RECT 1.005000  0.850000 1.345000 1.020000 ;
      RECT 1.005000  1.020000 1.175000 1.720000 ;
      RECT 1.005000  1.720000 2.395000 1.890000 ;
      RECT 1.150000  2.230000 1.320000 2.905000 ;
      RECT 1.150000  2.905000 3.125000 3.075000 ;
      RECT 1.175000  0.390000 3.125000 0.640000 ;
      RECT 1.175000  0.640000 1.345000 0.850000 ;
      RECT 2.065000  1.890000 2.395000 2.735000 ;
      RECT 2.955000  0.640000 3.125000 0.980000 ;
      RECT 2.955000  0.980000 3.695000 1.150000 ;
      RECT 2.955000  1.320000 3.355000 1.650000 ;
      RECT 2.955000  1.650000 3.125000 2.905000 ;
      RECT 3.295000  0.085000 3.625000 0.810000 ;
      RECT 3.295000  1.820000 3.625000 3.245000 ;
      RECT 3.525000  1.150000 3.695000 1.300000 ;
      RECT 3.525000  1.300000 3.895000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__mux2_1

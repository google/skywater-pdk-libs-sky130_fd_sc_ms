* File: sky130_fd_sc_ms__a2111oi_2.pex.spice
* Created: Fri Aug 28 16:55:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2111OI_2%D1 3 7 11 13 14 23
c39 23 0 4.04281e-20 $X=1.145 $Y=1.515
c40 11 0 1.08785e-19 $X=1.145 $Y=2.4
r41 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.145 $Y2=1.515
r42 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.515 $X2=1.13 $Y2=1.515
r43 19 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.04 $Y=1.515 $X2=1.13
+ $Y2=1.515
r44 17 19 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.695 $Y=1.515
+ $X2=1.04 $Y2=1.515
r45 14 22 1.87607 $w=4.28e-07 $l=7e-08 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1.13
+ $Y2=1.565
r46 13 22 10.9884 $w=4.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.13 $Y2=1.565
r47 9 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.68
+ $X2=1.145 $Y2=1.515
r48 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.145 $Y=1.68
+ $X2=1.145 $Y2=2.4
r49 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.35
+ $X2=1.04 $Y2=1.515
r50 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.04 $Y=1.35 $X2=1.04
+ $Y2=0.74
r51 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.695 $Y=1.68
+ $X2=0.695 $Y2=1.515
r52 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.695 $Y=1.68
+ $X2=0.695 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%C1 3 5 7 8 10 11 12 13 20
c42 13 0 1.08785e-19 $X=2.64 $Y=1.665
c43 3 0 7.82037e-20 $X=1.58 $Y=0.74
r44 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.515 $X2=1.67 $Y2=1.515
r45 18 20 13.5393 $w=2.67e-07 $l=7.5e-08 $layer=POLY_cond $X=1.595 $Y=1.537
+ $X2=1.67 $Y2=1.537
r46 17 18 2.70787 $w=2.67e-07 $l=1.5e-08 $layer=POLY_cond $X=1.58 $Y=1.537
+ $X2=1.595 $Y2=1.537
r47 12 13 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.64 $Y2=1.565
r48 11 12 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.16 $Y2=1.565
r49 11 21 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.67
+ $Y2=1.565
r50 8 20 67.6966 $w=2.67e-07 $l=4.59483e-07 $layer=POLY_cond $X=2.045 $Y=1.725
+ $X2=1.67 $Y2=1.537
r51 8 10 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.045 $Y=1.725
+ $X2=2.045 $Y2=2.4
r52 5 18 12.032 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=1.595 $Y=1.725
+ $X2=1.595 $Y2=1.537
r53 5 7 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.595 $Y=1.725
+ $X2=1.595 $Y2=2.4
r54 1 17 16.2448 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.58 $Y=1.35
+ $X2=1.58 $Y2=1.537
r55 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.58 $Y=1.35 $X2=1.58
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%B1 1 3 5 8 12 14 15 19 23
r49 21 23 11.857 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.39 $Y=1.367
+ $X2=3.465 $Y2=1.367
r50 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.385 $X2=3.39 $Y2=1.385
r51 18 21 59.2852 $w=3.65e-07 $l=3.75e-07 $layer=POLY_cond $X=3.015 $Y=1.367
+ $X2=3.39 $Y2=1.367
r52 18 19 34.8101 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=3.015 $Y=1.367
+ $X2=2.925 $Y2=1.367
r53 15 22 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=3.39 $Y2=1.365
r54 14 22 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.39 $Y2=1.365
r55 10 23 19.2931 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=3.465 $Y=1.55
+ $X2=3.465 $Y2=1.367
r56 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.465 $Y=1.55
+ $X2=3.465 $Y2=2.4
r57 6 18 19.2931 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=3.015 $Y=1.55
+ $X2=3.015 $Y2=1.367
r58 6 8 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.015 $Y=1.55
+ $X2=3.015 $Y2=2.4
r59 5 19 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.195 $Y=1.26
+ $X2=2.925 $Y2=1.26
r60 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=1.185
+ $X2=2.195 $Y2=1.26
r61 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.12 $Y=1.185
+ $X2=2.12 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%A1 3 7 11 15 17 18 28
r55 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.365 $Y=1.515
+ $X2=4.38 $Y2=1.515
r56 25 27 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=4.13 $Y=1.515
+ $X2=4.365 $Y2=1.515
r57 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.515 $X2=4.13 $Y2=1.515
r58 23 25 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.95 $Y=1.515
+ $X2=4.13 $Y2=1.515
r59 21 23 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.915 $Y=1.515
+ $X2=3.95 $Y2=1.515
r60 18 26 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.13 $Y2=1.565
r61 17 26 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.13
+ $Y2=1.565
r62 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.38 $Y=1.35
+ $X2=4.38 $Y2=1.515
r63 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.38 $Y=1.35
+ $X2=4.38 $Y2=0.74
r64 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.68
+ $X2=4.365 $Y2=1.515
r65 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.365 $Y=1.68
+ $X2=4.365 $Y2=2.4
r66 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.35
+ $X2=3.95 $Y2=1.515
r67 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.95 $Y=1.35 $X2=3.95
+ $Y2=0.74
r68 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.68
+ $X2=3.915 $Y2=1.515
r69 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.915 $Y=1.68
+ $X2=3.915 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%A2 3 7 11 15 17 23 24
c38 7 0 2.06049e-19 $X=4.81 $Y=0.74
r39 24 25 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=5.25 $Y=1.515
+ $X2=5.265 $Y2=1.515
r40 22 24 35.177 $w=3.22e-07 $l=2.35e-07 $layer=POLY_cond $X=5.015 $Y=1.515
+ $X2=5.25 $Y2=1.515
r41 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.015
+ $Y=1.515 $X2=5.015 $Y2=1.515
r42 20 22 29.9379 $w=3.22e-07 $l=2e-07 $layer=POLY_cond $X=4.815 $Y=1.515
+ $X2=5.015 $Y2=1.515
r43 19 20 0.748447 $w=3.22e-07 $l=5e-09 $layer=POLY_cond $X=4.81 $Y=1.515
+ $X2=4.815 $Y2=1.515
r44 17 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.015 $Y=1.665
+ $X2=5.015 $Y2=1.515
r45 13 25 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.68
+ $X2=5.265 $Y2=1.515
r46 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.265 $Y=1.68
+ $X2=5.265 $Y2=2.4
r47 9 24 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.25 $Y=1.35
+ $X2=5.25 $Y2=1.515
r48 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.25 $Y=1.35 $X2=5.25
+ $Y2=0.74
r49 5 19 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.35
+ $X2=4.81 $Y2=1.515
r50 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.81 $Y=1.35 $X2=4.81
+ $Y2=0.74
r51 1 20 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.68
+ $X2=4.815 $Y2=1.515
r52 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.815 $Y=1.68
+ $X2=4.815 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%A_69_368# 1 2 3 12 14 15 18 22 26 28
c32 18 0 4.04281e-20 $X=1.37 $Y=2.115
c33 1 0 1.93692e-19 $X=0.345 $Y=1.84
r34 24 26 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.31 $Y=2.905
+ $X2=2.31 $Y2=2.455
r35 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=2.99
+ $X2=1.37 $Y2=2.99
r36 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.185 $Y=2.99
+ $X2=2.31 $Y2=2.905
r37 22 23 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.185 $Y=2.99
+ $X2=1.455 $Y2=2.99
r38 18 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.37 $Y=2.115 $X2=1.37
+ $Y2=2.815
r39 16 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.905
+ $X2=1.37 $Y2=2.99
r40 16 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.37 $Y=2.905 $X2=1.37
+ $Y2=2.815
r41 14 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=1.37 $Y2=2.99
r42 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=0.555 $Y2=2.99
r43 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.43 $Y=2.905
+ $X2=0.555 $Y2=2.99
r44 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.43 $Y=2.905
+ $X2=0.43 $Y2=2.455
r45 3 26 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=1.84 $X2=2.27 $Y2=2.455
r46 2 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.84 $X2=1.37 $Y2=2.815
r47 2 18 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.84 $X2=1.37 $Y2=2.115
r48 1 12 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.345
+ $Y=1.84 $X2=0.47 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%Y 1 2 3 4 13 14 15 16 21 23 27 29 34 35 36
+ 39 44 45
c71 39 0 4.44094e-20 $X=4.165 $Y=0.872
c72 36 0 7.82037e-20 $X=2.335 $Y=0.872
c73 16 0 1.93692e-19 $X=0.355 $Y=2.035
r74 44 45 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r75 39 42 2.72396 $w=3.28e-07 $l=7.8e-08 $layer=LI1_cond $X=4.165 $Y=0.872
+ $X2=4.165 $Y2=0.95
r76 36 37 7.78772 $w=3.28e-07 $l=2.23e-07 $layer=LI1_cond $X=2.335 $Y=0.872
+ $X2=2.335 $Y2=1.095
r77 32 45 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.95
+ $X2=0.24 $Y2=1.665
r78 31 44 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r79 30 36 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=0.872
+ $X2=2.335 $Y2=0.872
r80 29 39 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=0.872
+ $X2=4.165 $Y2=0.872
r81 29 30 81.153 $w=2.03e-07 $l=1.5e-06 $layer=LI1_cond $X=4 $Y=0.872 $X2=2.5
+ $Y2=0.872
r82 25 36 3.5621 $w=3.28e-07 $l=1.02e-07 $layer=LI1_cond $X=2.335 $Y=0.77
+ $X2=2.335 $Y2=0.872
r83 25 27 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.335 $Y=0.77
+ $X2=2.335 $Y2=0.515
r84 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=1.095
+ $X2=1.325 $Y2=1.095
r85 23 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=1.095
+ $X2=2.335 $Y2=1.095
r86 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.17 $Y=1.095
+ $X2=1.49 $Y2=1.095
r87 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=1.01
+ $X2=1.325 $Y2=1.095
r88 19 21 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.325 $Y=1.01
+ $X2=1.325 $Y2=0.515
r89 16 32 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.035
+ $X2=0.24 $Y2=1.95
r90 15 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=2.035
+ $X2=0.92 $Y2=2.035
r91 15 16 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.755 $Y=2.035
+ $X2=0.355 $Y2=2.035
r92 14 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.095
+ $X2=0.24 $Y2=1.18
r93 13 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=1.095
+ $X2=1.325 $Y2=1.095
r94 13 14 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.16 $Y=1.095
+ $X2=0.355 $Y2=1.095
r95 4 34 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=0.785
+ $Y=1.84 $X2=0.92 $Y2=2.115
r96 3 42 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.37 $X2=4.165 $Y2=0.95
r97 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.195
+ $Y=0.37 $X2=2.335 $Y2=0.515
r98 1 21 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.115
+ $Y=0.37 $X2=1.325 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%A_337_368# 1 2 9 14 16
r23 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=2.035
+ $X2=1.82 $Y2=2.035
r24 9 16 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=3.2 $Y2=1.97
r25 9 10 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=1.985 $Y2=2.035
r26 2 16 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.105
+ $Y=1.84 $X2=3.24 $Y2=1.985
r27 1 14 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.84 $X2=1.82 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%A_533_368# 1 2 3 4 15 17 18 19 22 23 27 29
+ 31 33 38
r55 31 40 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=5.53 $Y=2.12 $X2=5.53
+ $Y2=1.97
r56 31 33 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=5.53 $Y=2.12
+ $X2=5.53 $Y2=2.4
r57 30 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.675 $Y=2.035
+ $X2=4.55 $Y2=2.035
r58 29 40 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=5.53 $Y2=1.97
r59 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=4.675 $Y2=2.035
r60 25 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=2.12
+ $X2=4.55 $Y2=2.035
r61 25 27 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=4.55 $Y=2.12
+ $X2=4.55 $Y2=2.445
r62 24 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.035
+ $X2=3.69 $Y2=2.035
r63 23 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=2.035
+ $X2=4.55 $Y2=2.035
r64 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.425 $Y=2.035
+ $X2=3.855 $Y2=2.035
r65 20 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.69 $Y=2.905 $X2=3.69
+ $Y2=2.815
r66 19 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.12 $X2=3.69
+ $Y2=2.035
r67 19 22 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.69 $Y=2.12
+ $X2=3.69 $Y2=2.815
r68 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=3.69 $Y2=2.905
r69 17 18 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=2.905 $Y2=2.99
r70 13 18 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.765 $Y=2.905
+ $X2=2.905 $Y2=2.99
r71 13 15 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=2.765 $Y=2.905
+ $X2=2.765 $Y2=2.455
r72 4 40 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.84 $X2=5.49 $Y2=1.985
r73 4 33 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.84 $X2=5.49 $Y2=2.4
r74 3 38 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.84 $X2=4.59 $Y2=2.035
r75 3 27 300 $w=1.7e-07 $l=6.69104e-07 $layer=licon1_PDIFF $count=2 $X=4.455
+ $Y=1.84 $X2=4.59 $Y2=2.445
r76 2 36 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=1.84 $X2=3.69 $Y2=2.035
r77 2 22 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=1.84 $X2=3.69 $Y2=2.815
r78 1 15 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.84 $X2=2.79 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%VPWR 1 2 9 13 15 17 22 29 30 33 36
r58 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r59 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r61 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r62 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.04 $Y2=3.33
r63 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.52 $Y2=3.33
r64 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r65 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r67 23 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.14 $Y2=3.33
r68 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.56 $Y2=3.33
r69 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=5.04 $Y2=3.33
r70 22 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 19 20 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 17 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=3.33
+ $X2=4.14 $Y2=3.33
r73 17 19 248.893 $w=1.68e-07 $l=3.815e-06 $layer=LI1_cond $X=4.055 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 15 34 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=4.08 $Y2=3.33
r75 15 20 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=3.33
r77 11 13 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=2.405
r78 7 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=3.245 $X2=4.14
+ $Y2=3.33
r79 7 9 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.14 $Y=3.245 $X2=4.14
+ $Y2=2.455
r80 2 13 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=4.905
+ $Y=1.84 $X2=5.04 $Y2=2.405
r81 1 9 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.005
+ $Y=1.84 $X2=4.14 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%VGND 1 2 3 14 16 20 24 26 28 38 39 42 45
+ 48
r53 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r54 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r56 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r58 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r59 36 48 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.03
+ $Y2=0
r60 36 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.52
+ $Y2=0
r61 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r62 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 32 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r64 31 34 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r65 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r66 29 45 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.83 $Y2=0
r67 29 31 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.16
+ $Y2=0
r68 28 48 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.86 $Y=0 $X2=5.03
+ $Y2=0
r69 28 34 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.86 $Y=0 $X2=4.56
+ $Y2=0
r70 26 35 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r71 26 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r72 22 48 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r73 22 24 19.9983 $w=3.38e-07 $l=5.9e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.675
r74 18 45 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=0.085
+ $X2=1.83 $Y2=0
r75 18 20 19.9983 $w=3.38e-07 $l=5.9e-07 $layer=LI1_cond $X=1.83 $Y=0.085
+ $X2=1.83 $Y2=0.675
r76 17 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.825
+ $Y2=0
r77 16 45 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.83
+ $Y2=0
r78 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=0.99
+ $Y2=0
r79 12 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r80 12 14 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.675
r81 3 24 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.885
+ $Y=0.37 $X2=5.03 $Y2=0.675
r82 2 20 182 $w=1.7e-07 $l=3.82623e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.37 $X2=1.83 $Y2=0.675
r83 1 14 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.37 $X2=0.825 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_2%A_722_74# 1 2 3 10 14 18 19 22
c30 14 0 1.6164e-19 $X=4.595 $Y=0.6
r31 20 22 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.505 $Y=1.01
+ $X2=5.505 $Y2=0.515
r32 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.38 $Y=1.095
+ $X2=5.505 $Y2=1.01
r33 18 19 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.38 $Y=1.095 $X2=4.68
+ $Y2=1.095
r34 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.595 $Y=1.01
+ $X2=4.68 $Y2=1.095
r35 15 17 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.595 $Y=1.01
+ $X2=4.595 $Y2=0.965
r36 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.595 $Y=0.6
+ $X2=4.595 $Y2=0.475
r37 14 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.595 $Y=0.6
+ $X2=4.595 $Y2=0.965
r38 10 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=0.475
+ $X2=4.595 $Y2=0.475
r39 10 12 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=4.51 $Y=0.475
+ $X2=3.735 $Y2=0.475
r40 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.325
+ $Y=0.37 $X2=5.465 $Y2=0.515
r41 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.37 $X2=4.595 $Y2=0.515
r42 2 17 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.37 $X2=4.595 $Y2=0.965
r43 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.61
+ $Y=0.37 $X2=3.735 $Y2=0.515
.ends


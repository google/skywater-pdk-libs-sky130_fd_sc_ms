* File: sky130_fd_sc_ms__a2111oi_2.spice
* Created: Fri Aug 28 16:55:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2111oi_2.pex.spice"
.subckt sky130_fd_sc_ms__a2111oi_2  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_D1_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.2109 PD=1.13 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_C1_M1000_g N_Y_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=5.664 NRS=6.48 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=12.156 M=1 R=4.93333 SA=75001.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_722_74#_M1001_d N_A1_M1001_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1014 N_A_722_74#_M1014_d N_A1_M1014_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_722_74#_M1014_d N_A2_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1073 PD=1.02 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_722_74#_M1013_d N_A2_M1013_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1073 PD=2.01 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_D1_M1003_g N_A_69_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1003_d N_D1_M1004_g N_A_69_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1006 N_A_337_368#_M1006_d N_C1_M1006_g N_A_69_368#_M1004_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1008 N_A_337_368#_M1006_d N_C1_M1008_g N_A_69_368#_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1010 N_A_337_368#_M1010_d N_B1_M1010_g N_A_533_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1011 N_A_337_368#_M1010_d N_B1_M1011_g N_A_533_368#_M1011_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90002 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_533_368#_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1015 N_VPWR_M1012_d N_A1_M1015_g N_A_533_368#_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1002 N_A_533_368#_M1015_s N_A2_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1016 N_A_533_368#_M1016_d N_A2_M1016_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX17_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__a2111oi_2.pxi.spice"
*
.ends
*
*

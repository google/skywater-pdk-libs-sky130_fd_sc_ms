* NGSPICE file created from sky130_fd_sc_ms__nor4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
M1000 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.594e+11p ps=6.85e+06u
M1001 a_347_368# B a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.696e+11p pd=2.9e+06u as=2.688e+11p ps=2.72e+06u
M1002 VGND a_57_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND D_N a_57_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 Y a_57_368# a_449_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.48e+11p pd=3.04e+06u as=4.368e+11p ps=3.02e+06u
M1006 a_263_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.06e+11p ps=3.02e+06u
M1007 a_449_368# C a_347_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR D_N a_57_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


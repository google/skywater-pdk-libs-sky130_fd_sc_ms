* File: sky130_fd_sc_ms__a41oi_4.spice
* Created: Fri Aug 28 17:10:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a41oi_4.pex.spice"
.subckt sky130_fd_sc_ms__a41oi_4  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_B1_M1015_g N_Y_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1032_d N_B1_M1032_g N_Y_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_Y_M1020_d N_A1_M1020_g N_A_325_74#_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1022 N_Y_M1020_d N_A1_M1022_g N_A_325_74#_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2294 PD=1.09 PS=1.36 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1026 N_Y_M1026_d N_A1_M1026_g N_A_325_74#_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2294 PD=1.02 PS=1.36 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1036 N_Y_M1026_d N_A1_M1036_g N_A_325_74#_M1036_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.9
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_852_74#_M1005_d N_A2_M1005_g N_A_325_74#_M1036_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_852_74#_M1005_d N_A2_M1006_g N_A_325_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1023 N_A_852_74#_M1023_d N_A2_M1023_g N_A_325_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1027 N_A_852_74#_M1023_d N_A2_M1027_g N_A_325_74#_M1027_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_1235_74#_M1008_d N_A3_M1008_g N_A_852_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1018 N_A_1235_74#_M1018_d N_A3_M1018_g N_A_852_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1021 N_A_1235_74#_M1018_d N_A3_M1021_g N_A_852_74#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1033 N_A_1235_74#_M1033_d N_A3_M1033_g N_A_852_74#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1004 N_A_1235_74#_M1033_d N_A4_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1016 N_A_1235_74#_M1016_d N_A4_M1016_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1017 N_A_1235_74#_M1016_d N_A4_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1028 N_A_1235_74#_M1028_d N_A4_M1028_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75003.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_27_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.3192 PD=1.435 PS=2.81 NRD=7.0329 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90009.2 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1002_d N_B1_M1007_g N_A_27_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.1792 PD=1.435 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7
+ SB=90008.8 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g N_A_27_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.2
+ SB=90008.3 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1009_d N_B1_M1012_g N_A_27_368#_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90007.8 A=0.2016 P=2.6 MULT=1
MM1000 N_A_27_368#_M1012_s N_A1_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.1
+ SB=90007.4 A=0.2016 P=2.6 MULT=1
MM1010 N_A_27_368#_M1010_d N_A1_M1010_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.6
+ SB=90006.8 A=0.2016 P=2.6 MULT=1
MM1013 N_A_27_368#_M1010_d N_A1_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.182 PD=1.39 PS=1.445 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.1
+ SB=90006.4 A=0.2016 P=2.6 MULT=1
MM1014 N_A_27_368#_M1014_d N_A1_M1014_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.182 PD=1.39 PS=1.445 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90003.6
+ SB=90005.8 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_27_368#_M1014_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1848 AS=0.1512 PD=1.45 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004
+ SB=90005.4 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1003_d N_A2_M1019_g N_A_27_368#_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1848 AS=0.1512 PD=1.45 PS=1.39 NRD=9.6727 NRS=0 M=1 R=6.22222 SA=90004.6
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1024 N_VPWR_M1024_d N_A2_M1024_g N_A_27_368#_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1025 N_VPWR_M1024_d N_A2_M1025_g N_A_27_368#_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90005.5
+ SB=90003.9 A=0.2016 P=2.6 MULT=1
MM1029 N_VPWR_M1029_d N_A3_M1029_g N_A_27_368#_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1030 N_VPWR_M1029_d N_A3_M1030_g N_A_27_368#_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90006.5
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1034 N_VPWR_M1034_d N_A3_M1034_g N_A_27_368#_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.9
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1035 N_VPWR_M1034_d N_A3_M1035_g N_A_27_368#_M1035_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90007.4
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1001_d N_A4_M1001_g N_A_27_368#_M1035_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90007.9
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1011 N_VPWR_M1001_d N_A4_M1011_g N_A_27_368#_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90008.4
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1031 N_VPWR_M1031_d N_A4_M1031_g N_A_27_368#_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90008.8
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1037 N_VPWR_M1031_d N_A4_M1037_g N_A_27_368#_M1037_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90009.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX38_noxref VNB VPB NWDIODE A=19.4556 P=24.64
c_76 VNB 0 1.1015e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a41oi_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_890_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_792_463# a_834_355# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X2 a_303_395# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_2013_409# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_702_463# a_497_395# a_812_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 VPWR a_2013_409# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_124_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 Q a_2013_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR RESET_B a_702_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X9 a_37_78# D a_124_78# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_1353_392# a_303_395# a_1647_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 VPWR a_702_463# a_834_355# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 a_1678_395# a_1353_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X13 VPWR a_303_395# a_497_395# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_37_78# a_497_395# a_702_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 a_37_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X16 a_1827_81# a_1353_392# a_1678_395# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_1353_392# a_497_395# a_1630_493# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X18 a_834_355# a_497_395# a_1353_392# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND RESET_B a_1827_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_1630_493# a_1678_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X21 Q a_2013_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 VGND a_303_395# a_497_395# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR a_1353_392# a_2013_409# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X24 VPWR D a_37_78# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X25 VPWR RESET_B a_1678_395# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X26 a_812_138# a_834_355# a_890_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 Q a_2013_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 VGND a_2013_409# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_303_395# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 a_834_355# a_303_395# a_1353_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X31 a_702_463# a_303_395# a_792_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X32 VGND a_702_463# a_834_355# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 a_2013_409# a_1353_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X34 a_1647_81# a_1678_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 Q a_2013_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_37_78# a_303_395# a_702_463# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VGND a_1353_392# a_2013_409# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 VGND a_2013_409# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

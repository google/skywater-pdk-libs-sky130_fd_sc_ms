* File: sky130_fd_sc_ms__o2bb2a_4.spice
* Created: Fri Aug 28 17:59:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2bb2a_4.pex.spice"
.subckt sky130_fd_sc_ms__o2bb2a_4  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_B1_M1022_g N_A_27_74#_M1022_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1022_d N_B1_M1023_g N_A_27_74#_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.0896 PD=1.06 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.8
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_27_74#_M1023_s N_B2_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1016 N_A_27_74#_M1016_d N_B2_M1016_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0992 AS=0.112 PD=0.95 PS=0.99 NRD=2.808 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_27_74#_M1016_d N_A_476_48#_M1005_g N_A_313_392#_M1005_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0992 AS=0.1008 PD=0.95 PS=0.955 NRD=2.808 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_27_74#_M1019_d N_A_476_48#_M1019_g N_A_313_392#_M1005_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2048 AS=0.1008 PD=1.92 PS=0.955 NRD=6.552 NRS=6.552 M=1
+ R=4.26667 SA=75002.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 A_835_94# N_A2_N_M1020_g N_A_476_48#_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1952 PD=0.88 PS=1.89 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A1_N_M1017_g A_835_94# VNB NLOWVT L=0.15 W=0.64
+ AD=0.157032 AS=0.0768 PD=1.14087 PS=0.88 NRD=19.68 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1004 N_X_M1004_d N_A_313_392#_M1004_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.15725 AS=0.181568 PD=1.165 PS=1.31913 NRD=12.156 NRS=17.016 M=1 R=4.93333
+ SA=75001.1 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1004_d N_A_313_392#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15725 AS=0.1295 PD=1.165 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_313_392#_M1012_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1018 N_X_M1012_d N_A_313_392#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_A_41_392#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1000_d N_B1_M1001_g N_A_41_392#_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 N_A_313_392#_M1006_d N_B2_M1006_g N_A_41_392#_M1001_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_313_392#_M1006_d N_B2_M1009_g N_A_41_392#_M1009_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_476_48#_M1010_g N_A_313_392#_M1010_s VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1428 PD=2.24 PS=1.18 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003.9 A=0.1512 P=2.04 MULT=1
MM1021 N_VPWR_M1021_d N_A_476_48#_M1021_g N_A_313_392#_M1010_s VPB PSHORT L=0.18
+ W=0.84 AD=0.2457 AS=0.1428 PD=1.7 PS=1.18 NRD=55.6919 NRS=14.0658 M=1
+ R=4.66667 SA=90000.7 SB=90003.4 A=0.1512 P=2.04 MULT=1
MM1002 N_A_476_48#_M1002_d N_A2_N_M1002_g N_VPWR_M1021_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2457 PD=1.11 PS=1.7 NRD=0 NRS=55.6919 M=1 R=4.66667
+ SA=90001.3 SB=90002.8 A=0.1512 P=2.04 MULT=1
MM1007 N_VPWR_M1007_d N_A1_N_M1007_g N_A_476_48#_M1002_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2196 AS=0.1134 PD=1.45714 PS=1.11 NRD=48.4029 NRS=0 M=1 R=4.66667
+ SA=90001.8 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1003 N_VPWR_M1007_d N_A_313_392#_M1003_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2928 AS=0.2072 PD=1.94286 PS=1.49 NRD=14.9326 NRS=7.8997 M=1 R=6.22222
+ SA=90001.9 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1011 N_VPWR_M1011_d N_A_313_392#_M1011_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2072 PD=1.44 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.4
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1011_d N_A_313_392#_M1013_g N_X_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.154 PD=1.44 PS=1.395 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1015 N_VPWR_M1015_d N_A_313_392#_M1015_g N_X_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.364 AS=0.154 PD=2.89 PS=1.395 NRD=7.0329 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.0988 P=18.88
c_72 VNB 0 1.74227e-19 $X=0 $Y=0
c_932 A_835_94# 0 2.65681e-20 $X=4.175 $Y=0.47
*
.include "sky130_fd_sc_ms__o2bb2a_4.pxi.spice"
*
.ends
*
*

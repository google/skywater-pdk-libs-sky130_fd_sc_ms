* File: sky130_fd_sc_ms__or2b_4.pxi.spice
* Created: Fri Aug 28 18:07:19 2020
* 
x_PM_SKY130_FD_SC_MS__OR2B_4%A_81_296# N_A_81_296#_M1000_d N_A_81_296#_M1006_d
+ N_A_81_296#_M1001_d N_A_81_296#_M1008_g N_A_81_296#_M1005_g
+ N_A_81_296#_M1010_g N_A_81_296#_M1009_g N_A_81_296#_M1011_g
+ N_A_81_296#_M1012_g N_A_81_296#_M1016_g N_A_81_296#_M1013_g
+ N_A_81_296#_c_123_n N_A_81_296#_c_124_n N_A_81_296#_c_125_n
+ N_A_81_296#_c_126_n N_A_81_296#_c_127_n N_A_81_296#_c_128_n
+ N_A_81_296#_c_129_n N_A_81_296#_c_130_n N_A_81_296#_c_131_n
+ N_A_81_296#_c_132_n N_A_81_296#_c_133_n N_A_81_296#_c_134_n
+ PM_SKY130_FD_SC_MS__OR2B_4%A_81_296#
x_PM_SKY130_FD_SC_MS__OR2B_4%A N_A_M1000_g N_A_M1003_g N_A_c_256_n N_A_M1004_g
+ N_A_M1007_g N_A_c_258_n A A N_A_c_260_n PM_SKY130_FD_SC_MS__OR2B_4%A
x_PM_SKY130_FD_SC_MS__OR2B_4%A_676_48# N_A_676_48#_M1014_d N_A_676_48#_M1015_d
+ N_A_676_48#_M1006_g N_A_676_48#_c_314_n N_A_676_48#_c_315_n
+ N_A_676_48#_M1001_g N_A_676_48#_M1017_g N_A_676_48#_M1002_g
+ N_A_676_48#_c_318_n N_A_676_48#_c_319_n N_A_676_48#_c_320_n
+ N_A_676_48#_c_321_n N_A_676_48#_c_322_n N_A_676_48#_c_323_n
+ N_A_676_48#_c_324_n N_A_676_48#_c_325_n PM_SKY130_FD_SC_MS__OR2B_4%A_676_48#
x_PM_SKY130_FD_SC_MS__OR2B_4%B_N N_B_N_c_400_n N_B_N_M1014_g N_B_N_c_401_n
+ N_B_N_c_402_n N_B_N_c_405_n N_B_N_M1015_g N_B_N_c_403_n B_N B_N N_B_N_c_404_n
+ PM_SKY130_FD_SC_MS__OR2B_4%B_N
x_PM_SKY130_FD_SC_MS__OR2B_4%VPWR N_VPWR_M1008_s N_VPWR_M1009_s N_VPWR_M1016_s
+ N_VPWR_M1004_s N_VPWR_M1015_s N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n
+ N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_446_n VPWR N_VPWR_c_447_n N_VPWR_c_448_n
+ N_VPWR_c_449_n N_VPWR_c_436_n N_VPWR_c_451_n N_VPWR_c_452_n
+ PM_SKY130_FD_SC_MS__OR2B_4%VPWR
x_PM_SKY130_FD_SC_MS__OR2B_4%X N_X_M1005_s N_X_M1012_s N_X_M1008_d N_X_M1011_d
+ N_X_c_514_n N_X_c_515_n N_X_c_516_n N_X_c_521_n N_X_c_517_n N_X_c_522_n
+ N_X_c_523_n N_X_c_518_n N_X_c_519_n N_X_c_524_n X PM_SKY130_FD_SC_MS__OR2B_4%X
x_PM_SKY130_FD_SC_MS__OR2B_4%A_492_392# N_A_492_392#_M1003_d
+ N_A_492_392#_M1001_s N_A_492_392#_M1002_s N_A_492_392#_c_583_n
+ N_A_492_392#_c_584_n N_A_492_392#_c_585_n N_A_492_392#_c_586_n
+ N_A_492_392#_c_587_n N_A_492_392#_c_588_n N_A_492_392#_c_589_n
+ N_A_492_392#_c_590_n PM_SKY130_FD_SC_MS__OR2B_4%A_492_392#
x_PM_SKY130_FD_SC_MS__OR2B_4%VGND N_VGND_M1005_d N_VGND_M1010_d N_VGND_M1013_d
+ N_VGND_M1007_s N_VGND_M1017_s N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n VGND N_VGND_c_643_n
+ N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n N_VGND_c_648_n
+ N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n
+ PM_SKY130_FD_SC_MS__OR2B_4%VGND
cc_1 VNB N_A_81_296#_M1008_g 0.00243092f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A_81_296#_M1005_g 0.0363403f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_A_81_296#_M1010_g 0.021162f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_A_81_296#_M1009_g 0.0015348f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_5 VNB N_A_81_296#_M1011_g 0.00154219f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_6 VNB N_A_81_296#_M1012_g 0.0220733f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_7 VNB N_A_81_296#_M1016_g 0.00167568f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_8 VNB N_A_81_296#_M1013_g 0.0223805f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_9 VNB N_A_81_296#_c_123_n 0.0115322f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.555
cc_10 VNB N_A_81_296#_c_124_n 0.0021705f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.465
cc_11 VNB N_A_81_296#_c_125_n 0.00687872f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.195
cc_12 VNB N_A_81_296#_c_126_n 0.00553968f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.515
cc_13 VNB N_A_81_296#_c_127_n 0.0119082f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.195
cc_14 VNB N_A_81_296#_c_128_n 0.00307801f $X=-0.19 $Y=-0.245 $X2=3.67 $Y2=0.515
cc_15 VNB N_A_81_296#_c_129_n 3.78434e-19 $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.08
cc_16 VNB N_A_81_296#_c_130_n 0.00796175f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.195
cc_17 VNB N_A_81_296#_c_131_n 0.00312763f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.195
cc_18 VNB N_A_81_296#_c_132_n 0.007464f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.28
cc_19 VNB N_A_81_296#_c_133_n 0.00962625f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.465
cc_20 VNB N_A_81_296#_c_134_n 0.0595951f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.465
cc_21 VNB N_A_M1000_g 0.0360123f $X=-0.19 $Y=-0.245 $X2=3.905 $Y2=1.935
cc_22 VNB N_A_M1003_g 0.00382132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_256_n 0.00993221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_M1007_g 0.0365137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_c_258_n 0.006075f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.555
cc_26 VNB A 0.0049455f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_27 VNB N_A_c_260_n 0.0148545f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.63
cc_28 VNB N_A_676_48#_M1006_g 0.0331319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_676_48#_c_314_n 0.0119927f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_30 VNB N_A_676_48#_c_315_n 0.0101155f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_31 VNB N_A_676_48#_M1001_g 0.00403268f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_32 VNB N_A_676_48#_M1017_g 0.035707f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.555
cc_33 VNB N_A_676_48#_c_318_n 0.00374105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_676_48#_c_319_n 0.00141541f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.63
cc_35 VNB N_A_676_48#_c_320_n 0.0385846f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_36 VNB N_A_676_48#_c_321_n 0.0379768f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.63
cc_37 VNB N_A_676_48#_c_322_n 0.00186199f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_38 VNB N_A_676_48#_c_323_n 0.0237469f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_39 VNB N_A_676_48#_c_324_n 0.00618737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_676_48#_c_325_n 0.0121834f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.465
cc_41 VNB N_B_N_c_400_n 0.0204172f $X=-0.19 $Y=-0.245 $X2=2.43 $Y2=0.37
cc_42 VNB N_B_N_c_401_n 0.0538601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_B_N_c_402_n 0.00815644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_B_N_c_403_n 0.00703507f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.63
cc_45 VNB N_B_N_c_404_n 0.0316413f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_46 VNB N_VPWR_c_436_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_514_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_48 VNB N_X_c_515_n 0.0041248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_516_n 0.00156967f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.555
cc_50 VNB N_X_c_517_n 0.0060023f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_51 VNB N_X_c_518_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_52 VNB N_X_c_519_n 0.0182272f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=0.74
cc_53 VNB N_VGND_c_637_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_54 VNB N_VGND_c_638_n 0.0354929f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.555
cc_55 VNB N_VGND_c_639_n 0.00509474f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_56 VNB N_VGND_c_640_n 0.00577125f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_57 VNB N_VGND_c_641_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_58 VNB N_VGND_c_642_n 0.00923674f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_59 VNB N_VGND_c_643_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_60 VNB N_VGND_c_644_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_645_n 0.0193334f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.465
cc_62 VNB N_VGND_c_646_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.195
cc_63 VNB N_VGND_c_647_n 0.0401986f $X=-0.19 $Y=-0.245 $X2=3.67 $Y2=0.515
cc_64 VNB N_VGND_c_648_n 0.324755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_649_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_650_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.195
cc_67 VNB N_VGND_c_651_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_68 VNB N_VGND_c_652_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.465
cc_69 VPB N_A_81_296#_M1008_g 0.0289572f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_70 VPB N_A_81_296#_M1009_g 0.021403f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_71 VPB N_A_81_296#_M1011_g 0.0220397f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_72 VPB N_A_81_296#_M1016_g 0.0236432f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_73 VPB N_A_81_296#_c_129_n 0.00236526f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.08
cc_74 VPB N_A_M1003_g 0.0304936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_M1004_g 0.0276466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB A 0.00637848f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_77 VPB N_A_c_260_n 0.0122605f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.63
cc_78 VPB N_A_676_48#_M1001_g 0.0322072f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_79 VPB N_A_676_48#_M1002_g 0.0259721f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_80 VPB N_A_676_48#_c_321_n 0.0560798f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.63
cc_81 VPB N_A_676_48#_c_322_n 0.00251184f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=0.74
cc_82 VPB N_A_676_48#_c_323_n 0.017365f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=0.74
cc_83 VPB N_B_N_c_405_n 0.0244376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_B_N_c_403_n 0.0288909f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.63
cc_85 VPB B_N 0.00252041f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_86 VPB N_VPWR_c_437_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_87 VPB N_VPWR_c_438_n 0.0576005f $X=-0.19 $Y=1.66 $X2=0.85 $Y2=1.555
cc_88 VPB N_VPWR_c_439_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.63
cc_89 VPB N_VPWR_c_440_n 0.00958622f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.63
cc_90 VPB N_VPWR_c_441_n 0.0153221f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_91 VPB N_VPWR_c_442_n 0.0179486f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_92 VPB N_VPWR_c_443_n 0.0162121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_444_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.555
cc_94 VPB N_VPWR_c_445_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.465
cc_95 VPB N_VPWR_c_446_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.465
cc_96 VPB N_VPWR_c_447_n 0.020445f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=0.515
cc_97 VPB N_VPWR_c_448_n 0.0413605f $X=-0.19 $Y=1.66 $X2=3.63 $Y2=1.11
cc_98 VPB N_VPWR_c_449_n 0.0177091f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=1.465
cc_99 VPB N_VPWR_c_436_n 0.0934715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_451_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.465
cc_101 VPB N_VPWR_c_452_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.465
cc_102 VPB N_X_c_516_n 0.00252674f $X=-0.19 $Y=1.66 $X2=0.85 $Y2=1.555
cc_103 VPB N_X_c_521_n 0.00206342f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_104 VPB N_X_c_522_n 0.00518214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_X_c_523_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_X_c_524_n 8.47995e-19 $X=-0.19 $Y=1.66 $X2=1.88 $Y2=0.74
cc_107 VPB N_A_492_392#_c_583_n 0.00279888f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.63
cc_108 VPB N_A_492_392#_c_584_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_109 VPB N_A_492_392#_c_585_n 0.0146887f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.48
cc_110 VPB N_A_492_392#_c_586_n 0.00345709f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_111 VPB N_A_492_392#_c_587_n 0.00736547f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.555
cc_112 VPB N_A_492_392#_c_588_n 0.00903347f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_113 VPB N_A_492_392#_c_589_n 0.00382309f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_114 VPB N_A_492_392#_c_590_n 0.00954783f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.63
cc_115 N_A_81_296#_M1013_g N_A_M1000_g 0.0123298f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_81_296#_c_125_n N_A_M1000_g 0.0191077f $X=2.475 $Y=1.195 $X2=0 $Y2=0
cc_117 N_A_81_296#_c_126_n N_A_M1000_g 0.00597167f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_118 N_A_81_296#_c_130_n N_A_M1000_g 0.00587547f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_119 N_A_81_296#_M1016_g N_A_M1003_g 0.028323f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_81_296#_c_131_n N_A_c_256_n 0.0068961f $X=2.64 $Y=1.195 $X2=0 $Y2=0
cc_121 N_A_81_296#_c_126_n N_A_M1007_g 0.0105092f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_122 N_A_81_296#_c_127_n N_A_M1007_g 0.0155134f $X=3.505 $Y=1.195 $X2=0 $Y2=0
cc_123 N_A_81_296#_c_128_n N_A_M1007_g 7.89164e-19 $X=3.67 $Y=0.515 $X2=0 $Y2=0
cc_124 N_A_81_296#_c_132_n N_A_M1007_g 8.03754e-19 $X=3.63 $Y=1.28 $X2=0 $Y2=0
cc_125 N_A_81_296#_c_134_n N_A_c_258_n 0.0123298f $X=1.88 $Y=1.465 $X2=0 $Y2=0
cc_126 N_A_81_296#_c_127_n A 0.0325657f $X=3.505 $Y=1.195 $X2=0 $Y2=0
cc_127 N_A_81_296#_c_129_n A 0.00995108f $X=4.04 $Y=2.08 $X2=0 $Y2=0
cc_128 N_A_81_296#_c_130_n A 0.00800544f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_129 N_A_81_296#_c_131_n A 0.0235756f $X=2.64 $Y=1.195 $X2=0 $Y2=0
cc_130 N_A_81_296#_c_127_n N_A_676_48#_M1006_g 0.0126768f $X=3.505 $Y=1.195
+ $X2=0 $Y2=0
cc_131 N_A_81_296#_c_128_n N_A_676_48#_M1006_g 0.0105052f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_132 N_A_81_296#_c_132_n N_A_676_48#_M1006_g 0.00726533f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_133 N_A_81_296#_c_132_n N_A_676_48#_c_314_n 0.00705335f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_134 N_A_81_296#_c_132_n N_A_676_48#_c_315_n 4.99147e-19 $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_135 N_A_81_296#_c_129_n N_A_676_48#_M1001_g 0.0245137f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_136 N_A_81_296#_c_128_n N_A_676_48#_M1017_g 0.00232377f $X=3.67 $Y=0.515
+ $X2=0 $Y2=0
cc_137 N_A_81_296#_c_132_n N_A_676_48#_M1017_g 0.0190269f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_138 N_A_81_296#_c_129_n N_A_676_48#_c_318_n 0.00478313f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_139 N_A_81_296#_c_132_n N_A_676_48#_c_318_n 0.00698284f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_140 N_A_81_296#_c_129_n N_A_676_48#_c_322_n 0.0245536f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_141 N_A_81_296#_c_132_n N_A_676_48#_c_322_n 3.96184e-19 $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_142 N_A_81_296#_c_129_n N_A_676_48#_c_323_n 0.00605141f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_143 N_A_81_296#_c_132_n N_A_676_48#_c_324_n 0.00914716f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_144 N_A_81_296#_c_129_n N_A_676_48#_c_325_n 0.00638285f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_145 N_A_81_296#_c_132_n N_A_676_48#_c_325_n 0.00304884f $X=3.63 $Y=1.28 $X2=0
+ $Y2=0
cc_146 N_A_81_296#_M1008_g N_VPWR_c_438_n 0.020251f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_81_296#_M1009_g N_VPWR_c_438_n 6.46441e-19 $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_148 N_A_81_296#_M1008_g N_VPWR_c_439_n 5.90862e-19 $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_149 N_A_81_296#_M1009_g N_VPWR_c_439_n 0.0152536f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_81_296#_M1011_g N_VPWR_c_439_n 0.00349416f $X=1.395 $Y=2.4 $X2=0
+ $Y2=0
cc_151 N_A_81_296#_M1016_g N_VPWR_c_440_n 0.00311086f $X=1.845 $Y=2.4 $X2=0
+ $Y2=0
cc_152 N_A_81_296#_c_125_n N_VPWR_c_440_n 0.00279228f $X=2.475 $Y=1.195 $X2=0
+ $Y2=0
cc_153 N_A_81_296#_c_130_n N_VPWR_c_440_n 0.00905857f $X=2.06 $Y=1.195 $X2=0
+ $Y2=0
cc_154 N_A_81_296#_M1008_g N_VPWR_c_443_n 0.00460063f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_155 N_A_81_296#_M1009_g N_VPWR_c_443_n 0.00460063f $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_156 N_A_81_296#_M1011_g N_VPWR_c_445_n 0.005209f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_81_296#_M1016_g N_VPWR_c_445_n 0.005209f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_81_296#_M1008_g N_VPWR_c_436_n 0.00908554f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_159 N_A_81_296#_M1009_g N_VPWR_c_436_n 0.00908554f $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_160 N_A_81_296#_M1011_g N_VPWR_c_436_n 0.00982266f $X=1.395 $Y=2.4 $X2=0
+ $Y2=0
cc_161 N_A_81_296#_M1016_g N_VPWR_c_436_n 0.00983045f $X=1.845 $Y=2.4 $X2=0
+ $Y2=0
cc_162 N_A_81_296#_M1005_g N_X_c_514_n 0.00760419f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_81_296#_M1010_g N_X_c_514_n 3.97481e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_81_296#_M1005_g N_X_c_515_n 0.0127847f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_81_296#_M1010_g N_X_c_515_n 0.00591885f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_81_296#_c_124_n N_X_c_515_n 0.00968248f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_167 N_A_81_296#_M1008_g N_X_c_516_n 0.00422544f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A_81_296#_M1005_g N_X_c_516_n 0.00168928f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_81_296#_M1009_g N_X_c_516_n 0.00391396f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A_81_296#_c_124_n N_X_c_516_n 0.0169058f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_171 N_A_81_296#_c_133_n N_X_c_516_n 0.0148528f $X=0.85 $Y=1.465 $X2=0 $Y2=0
cc_172 N_A_81_296#_c_134_n N_X_c_516_n 5.87163e-19 $X=1.88 $Y=1.465 $X2=0 $Y2=0
cc_173 N_A_81_296#_M1008_g N_X_c_521_n 3.79108e-19 $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_81_296#_M1009_g N_X_c_521_n 3.64731e-19 $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_81_296#_M1010_g N_X_c_517_n 0.014308f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_81_296#_M1012_g N_X_c_517_n 0.0125296f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_81_296#_c_124_n N_X_c_517_n 0.066849f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_178 N_A_81_296#_c_126_n N_X_c_517_n 0.00420057f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_179 N_A_81_296#_c_130_n N_X_c_517_n 0.00159809f $X=2.06 $Y=1.195 $X2=0 $Y2=0
cc_180 N_A_81_296#_c_134_n N_X_c_517_n 0.00723585f $X=1.88 $Y=1.465 $X2=0 $Y2=0
cc_181 N_A_81_296#_M1009_g N_X_c_522_n 0.0159541f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_81_296#_M1011_g N_X_c_522_n 0.0142465f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_81_296#_M1016_g N_X_c_522_n 0.00430872f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_81_296#_c_124_n N_X_c_522_n 0.0649634f $X=1.975 $Y=1.465 $X2=0 $Y2=0
cc_185 N_A_81_296#_c_134_n N_X_c_522_n 0.00417362f $X=1.88 $Y=1.465 $X2=0 $Y2=0
cc_186 N_A_81_296#_M1009_g N_X_c_523_n 7.7208e-19 $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_81_296#_M1011_g N_X_c_523_n 0.0145011f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_81_296#_M1016_g N_X_c_523_n 0.0132157f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_81_296#_M1010_g N_X_c_518_n 9.72214e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_81_296#_M1012_g N_X_c_518_n 0.00910117f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_81_296#_M1013_g N_X_c_518_n 4.71232e-19 $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_81_296#_M1005_g N_X_c_519_n 0.0182661f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_81_296#_c_123_n N_X_c_519_n 4.97848e-19 $X=0.495 $Y=1.555 $X2=0 $Y2=0
cc_194 N_A_81_296#_M1008_g N_X_c_524_n 8.3244e-19 $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_81_296#_c_125_n N_A_492_392#_c_583_n 0.00130416f $X=2.475 $Y=1.195
+ $X2=0 $Y2=0
cc_196 N_A_81_296#_c_131_n N_A_492_392#_c_583_n 0.00178483f $X=2.64 $Y=1.195
+ $X2=0 $Y2=0
cc_197 N_A_81_296#_c_127_n N_A_492_392#_c_585_n 0.00530457f $X=3.505 $Y=1.195
+ $X2=0 $Y2=0
cc_198 N_A_81_296#_c_127_n N_A_492_392#_c_586_n 0.00237093f $X=3.505 $Y=1.195
+ $X2=0 $Y2=0
cc_199 N_A_81_296#_c_129_n N_A_492_392#_c_586_n 0.00717766f $X=4.04 $Y=2.08
+ $X2=0 $Y2=0
cc_200 N_A_81_296#_c_132_n N_A_492_392#_c_586_n 0.00708319f $X=3.63 $Y=1.28
+ $X2=0 $Y2=0
cc_201 N_A_81_296#_M1001_d N_A_492_392#_c_588_n 0.00165831f $X=3.905 $Y=1.935
+ $X2=0 $Y2=0
cc_202 N_A_81_296#_c_129_n N_A_492_392#_c_588_n 0.0139027f $X=4.04 $Y=2.08 $X2=0
+ $Y2=0
cc_203 N_A_81_296#_c_130_n N_VGND_M1013_d 0.00184398f $X=2.06 $Y=1.195 $X2=0
+ $Y2=0
cc_204 N_A_81_296#_M1005_g N_VGND_c_638_n 0.00351842f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_81_296#_M1005_g N_VGND_c_639_n 4.94543e-19 $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_81_296#_M1010_g N_VGND_c_639_n 0.00916944f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_81_296#_M1012_g N_VGND_c_639_n 0.00393745f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_81_296#_M1013_g N_VGND_c_640_n 0.00193131f $X=1.88 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_81_296#_c_125_n N_VGND_c_640_n 0.0103909f $X=2.475 $Y=1.195 $X2=0
+ $Y2=0
cc_210 N_A_81_296#_c_126_n N_VGND_c_640_n 0.0229287f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_211 N_A_81_296#_c_130_n N_VGND_c_640_n 0.0132288f $X=2.06 $Y=1.195 $X2=0
+ $Y2=0
cc_212 N_A_81_296#_c_126_n N_VGND_c_641_n 0.0404434f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_213 N_A_81_296#_c_127_n N_VGND_c_641_n 0.0238718f $X=3.505 $Y=1.195 $X2=0
+ $Y2=0
cc_214 N_A_81_296#_c_128_n N_VGND_c_641_n 0.0220066f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_215 N_A_81_296#_c_128_n N_VGND_c_642_n 0.025828f $X=3.67 $Y=0.515 $X2=0 $Y2=0
cc_216 N_A_81_296#_c_132_n N_VGND_c_642_n 0.0132716f $X=3.63 $Y=1.28 $X2=0 $Y2=0
cc_217 N_A_81_296#_M1005_g N_VGND_c_643_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_218 N_A_81_296#_M1010_g N_VGND_c_643_n 0.00383152f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_81_296#_M1012_g N_VGND_c_644_n 0.00434272f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_81_296#_M1013_g N_VGND_c_644_n 0.00461464f $X=1.88 $Y=0.74 $X2=0
+ $Y2=0
cc_221 N_A_81_296#_c_126_n N_VGND_c_645_n 0.0146357f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_222 N_A_81_296#_c_128_n N_VGND_c_646_n 0.0109942f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_223 N_A_81_296#_M1005_g N_VGND_c_648_n 0.00823942f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_224 N_A_81_296#_M1010_g N_VGND_c_648_n 0.0075754f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_81_296#_M1012_g N_VGND_c_648_n 0.00820964f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_81_296#_M1013_g N_VGND_c_648_n 0.00908295f $X=1.88 $Y=0.74 $X2=0
+ $Y2=0
cc_227 N_A_81_296#_c_126_n N_VGND_c_648_n 0.0121141f $X=2.64 $Y=0.515 $X2=0
+ $Y2=0
cc_228 N_A_81_296#_c_128_n N_VGND_c_648_n 0.00904371f $X=3.67 $Y=0.515 $X2=0
+ $Y2=0
cc_229 N_A_M1007_g N_A_676_48#_M1006_g 0.0160624f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_230 A N_A_676_48#_c_315_n 0.00232169f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_231 N_A_c_260_n N_A_676_48#_c_315_n 0.0160624f $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_232 A N_A_676_48#_M1001_g 0.00179782f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_233 N_A_c_260_n N_A_676_48#_M1001_g 0.00197259f $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_234 N_A_M1003_g N_VPWR_c_440_n 0.00885471f $X=2.37 $Y=2.46 $X2=0 $Y2=0
cc_235 N_A_M1004_g N_VPWR_c_441_n 0.00501904f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_236 N_A_M1003_g N_VPWR_c_447_n 0.005209f $X=2.37 $Y=2.46 $X2=0 $Y2=0
cc_237 N_A_M1004_g N_VPWR_c_447_n 0.005209f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_238 N_A_M1003_g N_VPWR_c_436_n 0.00982933f $X=2.37 $Y=2.46 $X2=0 $Y2=0
cc_239 N_A_M1004_g N_VPWR_c_436_n 0.00987399f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_240 N_A_M1000_g N_X_c_517_n 2.21979e-19 $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_241 N_A_M1003_g N_X_c_522_n 6.50767e-19 $X=2.37 $Y=2.46 $X2=0 $Y2=0
cc_242 N_A_M1003_g N_A_492_392#_c_583_n 0.00305947f $X=2.37 $Y=2.46 $X2=0 $Y2=0
cc_243 N_A_c_256_n N_A_492_392#_c_583_n 3.09627e-19 $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A_M1004_g N_A_492_392#_c_583_n 0.0010042f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_245 A N_A_492_392#_c_583_n 0.0204053f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A_c_260_n N_A_492_392#_c_583_n 7.03021e-19 $X=2.865 $Y=1.515 $X2=0
+ $Y2=0
cc_247 N_A_M1003_g N_A_492_392#_c_584_n 0.0107284f $X=2.37 $Y=2.46 $X2=0 $Y2=0
cc_248 N_A_M1004_g N_A_492_392#_c_584_n 0.0130839f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_249 N_A_M1004_g N_A_492_392#_c_585_n 0.0150541f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_250 A N_A_492_392#_c_585_n 0.0359503f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_251 N_A_c_260_n N_A_492_392#_c_585_n 0.00316326f $X=2.865 $Y=1.515 $X2=0
+ $Y2=0
cc_252 N_A_M1004_g N_A_492_392#_c_586_n 8.93544e-19 $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_253 N_A_M1004_g N_A_492_392#_c_587_n 0.00341418f $X=2.82 $Y=2.46 $X2=0 $Y2=0
cc_254 N_A_M1000_g N_VGND_c_640_n 0.0107172f $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_255 N_A_M1007_g N_VGND_c_640_n 6.11496e-19 $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_256 N_A_M1000_g N_VGND_c_641_n 6.29519e-19 $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_257 N_A_M1007_g N_VGND_c_641_n 0.0112125f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_258 N_A_M1000_g N_VGND_c_645_n 0.00383152f $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_259 N_A_M1007_g N_VGND_c_645_n 0.00383152f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_260 N_A_M1000_g N_VGND_c_648_n 0.00758997f $X=2.355 $Y=0.69 $X2=0 $Y2=0
cc_261 N_A_M1007_g N_VGND_c_648_n 0.00758997f $X=2.955 $Y=0.69 $X2=0 $Y2=0
cc_262 N_A_676_48#_M1017_g N_B_N_c_400_n 0.0196085f $X=3.885 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_263 N_A_676_48#_c_319_n N_B_N_c_400_n 0.00686389f $X=4.53 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_264 N_A_676_48#_c_324_n N_B_N_c_400_n 0.00308772f $X=4.46 $Y=1.445 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_676_48#_c_320_n N_B_N_c_401_n 0.0253584f $X=5.405 $Y=0.65 $X2=0 $Y2=0
cc_266 N_A_676_48#_c_321_n N_B_N_c_401_n 0.0196942f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_267 N_A_676_48#_c_324_n N_B_N_c_401_n 0.0113271f $X=4.46 $Y=1.445 $X2=0 $Y2=0
cc_268 N_A_676_48#_c_322_n N_B_N_c_402_n 9.63591e-19 $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_269 N_A_676_48#_c_323_n N_B_N_c_402_n 0.0206255f $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_270 N_A_676_48#_c_324_n N_B_N_c_402_n 0.00296893f $X=4.46 $Y=1.445 $X2=0
+ $Y2=0
cc_271 N_A_676_48#_M1002_g N_B_N_c_403_n 3.61337e-19 $X=4.265 $Y=2.435 $X2=0
+ $Y2=0
cc_272 N_A_676_48#_c_321_n N_B_N_c_403_n 0.00751315f $X=5.49 $Y=2.105 $X2=0
+ $Y2=0
cc_273 N_A_676_48#_c_320_n B_N 0.0282282f $X=5.405 $Y=0.65 $X2=0 $Y2=0
cc_274 N_A_676_48#_c_321_n B_N 0.0517945f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_275 N_A_676_48#_c_323_n B_N 0.00141991f $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_276 N_A_676_48#_c_324_n B_N 0.0330704f $X=4.46 $Y=1.445 $X2=0 $Y2=0
cc_277 N_A_676_48#_c_322_n N_B_N_c_404_n 0.00134012f $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_278 N_A_676_48#_c_323_n N_B_N_c_404_n 0.0149629f $X=4.46 $Y=1.61 $X2=0 $Y2=0
cc_279 N_A_676_48#_c_324_n N_B_N_c_404_n 0.0045702f $X=4.46 $Y=1.445 $X2=0 $Y2=0
cc_280 N_A_676_48#_M1001_g N_VPWR_c_441_n 5.43557e-19 $X=3.815 $Y=2.435 $X2=0
+ $Y2=0
cc_281 N_A_676_48#_M1002_g N_VPWR_c_442_n 0.00217716f $X=4.265 $Y=2.435 $X2=0
+ $Y2=0
cc_282 N_A_676_48#_c_321_n N_VPWR_c_442_n 0.0342803f $X=5.49 $Y=2.105 $X2=0
+ $Y2=0
cc_283 N_A_676_48#_M1001_g N_VPWR_c_448_n 0.00113339f $X=3.815 $Y=2.435 $X2=0
+ $Y2=0
cc_284 N_A_676_48#_M1002_g N_VPWR_c_448_n 0.00115241f $X=4.265 $Y=2.435 $X2=0
+ $Y2=0
cc_285 N_A_676_48#_c_321_n N_VPWR_c_449_n 0.011066f $X=5.49 $Y=2.105 $X2=0 $Y2=0
cc_286 N_A_676_48#_c_321_n N_VPWR_c_436_n 0.00915947f $X=5.49 $Y=2.105 $X2=0
+ $Y2=0
cc_287 N_A_676_48#_c_315_n N_A_492_392#_c_585_n 0.00111948f $X=3.53 $Y=1.52
+ $X2=0 $Y2=0
cc_288 N_A_676_48#_c_315_n N_A_492_392#_c_586_n 0.00633348f $X=3.53 $Y=1.52
+ $X2=0 $Y2=0
cc_289 N_A_676_48#_M1001_g N_A_492_392#_c_586_n 4.69579e-19 $X=3.815 $Y=2.435
+ $X2=0 $Y2=0
cc_290 N_A_676_48#_M1001_g N_A_492_392#_c_588_n 0.016672f $X=3.815 $Y=2.435
+ $X2=0 $Y2=0
cc_291 N_A_676_48#_M1002_g N_A_492_392#_c_588_n 0.0162066f $X=4.265 $Y=2.435
+ $X2=0 $Y2=0
cc_292 N_A_676_48#_M1001_g N_A_492_392#_c_590_n 7.39464e-19 $X=3.815 $Y=2.435
+ $X2=0 $Y2=0
cc_293 N_A_676_48#_M1002_g N_A_492_392#_c_590_n 0.0132212f $X=4.265 $Y=2.435
+ $X2=0 $Y2=0
cc_294 N_A_676_48#_c_322_n N_A_492_392#_c_590_n 0.0228742f $X=4.46 $Y=1.61 $X2=0
+ $Y2=0
cc_295 N_A_676_48#_c_323_n N_A_492_392#_c_590_n 0.00195633f $X=4.46 $Y=1.61
+ $X2=0 $Y2=0
cc_296 N_A_676_48#_M1006_g N_VGND_c_641_n 0.00476029f $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_297 N_A_676_48#_M1006_g N_VGND_c_642_n 5.56357e-19 $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_298 N_A_676_48#_M1017_g N_VGND_c_642_n 0.0117552f $X=3.885 $Y=0.69 $X2=0
+ $Y2=0
cc_299 N_A_676_48#_c_319_n N_VGND_c_642_n 0.0260683f $X=4.53 $Y=0.95 $X2=0 $Y2=0
cc_300 N_A_676_48#_c_324_n N_VGND_c_642_n 0.00351404f $X=4.46 $Y=1.445 $X2=0
+ $Y2=0
cc_301 N_A_676_48#_c_325_n N_VGND_c_642_n 0.00606281f $X=4.175 $Y=1.61 $X2=0
+ $Y2=0
cc_302 N_A_676_48#_M1006_g N_VGND_c_646_n 0.00434272f $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_303 N_A_676_48#_M1017_g N_VGND_c_646_n 0.00383152f $X=3.885 $Y=0.69 $X2=0
+ $Y2=0
cc_304 N_A_676_48#_c_319_n N_VGND_c_647_n 0.00840325f $X=4.53 $Y=0.95 $X2=0
+ $Y2=0
cc_305 N_A_676_48#_c_320_n N_VGND_c_647_n 0.0454555f $X=5.405 $Y=0.65 $X2=0
+ $Y2=0
cc_306 N_A_676_48#_M1006_g N_VGND_c_648_n 0.00820772f $X=3.455 $Y=0.69 $X2=0
+ $Y2=0
cc_307 N_A_676_48#_M1017_g N_VGND_c_648_n 0.0075754f $X=3.885 $Y=0.69 $X2=0
+ $Y2=0
cc_308 N_A_676_48#_c_319_n N_VGND_c_648_n 0.00689675f $X=4.53 $Y=0.95 $X2=0
+ $Y2=0
cc_309 N_A_676_48#_c_320_n N_VGND_c_648_n 0.037886f $X=5.405 $Y=0.65 $X2=0 $Y2=0
cc_310 N_B_N_c_405_n N_VPWR_c_442_n 0.0211243f $X=5.265 $Y=1.88 $X2=0 $Y2=0
cc_311 N_B_N_c_403_n N_VPWR_c_442_n 0.00193159f $X=5.115 $Y=1.58 $X2=0 $Y2=0
cc_312 B_N N_VPWR_c_442_n 0.0233264f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_313 N_B_N_c_405_n N_VPWR_c_449_n 0.00460063f $X=5.265 $Y=1.88 $X2=0 $Y2=0
cc_314 N_B_N_c_405_n N_VPWR_c_436_n 0.00912261f $X=5.265 $Y=1.88 $X2=0 $Y2=0
cc_315 N_B_N_c_405_n N_A_492_392#_c_588_n 6.0406e-19 $X=5.265 $Y=1.88 $X2=0
+ $Y2=0
cc_316 N_B_N_c_405_n N_A_492_392#_c_590_n 3.81037e-19 $X=5.265 $Y=1.88 $X2=0
+ $Y2=0
cc_317 N_B_N_c_400_n N_VGND_c_642_n 0.00676331f $X=4.385 $Y=1.085 $X2=0 $Y2=0
cc_318 N_B_N_c_400_n N_VGND_c_647_n 0.00433139f $X=4.385 $Y=1.085 $X2=0 $Y2=0
cc_319 N_B_N_c_400_n N_VGND_c_648_n 0.00822102f $X=4.385 $Y=1.085 $X2=0 $Y2=0
cc_320 N_VPWR_c_438_n N_X_c_521_n 0.0386303f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_321 N_VPWR_c_439_n N_X_c_521_n 0.0271749f $X=1.17 $Y=2.305 $X2=0 $Y2=0
cc_322 N_VPWR_c_443_n N_X_c_521_n 0.00883494f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_323 N_VPWR_c_436_n N_X_c_521_n 0.0073128f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_324 N_VPWR_M1009_s N_X_c_522_n 0.00165831f $X=1.035 $Y=1.84 $X2=0 $Y2=0
cc_325 N_VPWR_c_439_n N_X_c_522_n 0.0148589f $X=1.17 $Y=2.305 $X2=0 $Y2=0
cc_326 N_VPWR_c_439_n N_X_c_523_n 0.0283501f $X=1.17 $Y=2.305 $X2=0 $Y2=0
cc_327 N_VPWR_c_440_n N_X_c_523_n 0.0339179f $X=2.07 $Y=2.105 $X2=0 $Y2=0
cc_328 N_VPWR_c_445_n N_X_c_523_n 0.0144623f $X=1.985 $Y=3.33 $X2=0 $Y2=0
cc_329 N_VPWR_c_436_n N_X_c_523_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_330 N_VPWR_c_438_n N_X_c_519_n 0.0142765f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_331 N_VPWR_c_438_n N_X_c_524_n 0.00654084f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_332 N_VPWR_c_440_n N_A_492_392#_c_583_n 0.00673913f $X=2.07 $Y=2.105 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_440_n N_A_492_392#_c_584_n 0.0295663f $X=2.07 $Y=2.105 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_441_n N_A_492_392#_c_584_n 0.0234083f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_447_n N_A_492_392#_c_584_n 0.0144623f $X=2.96 $Y=3.33 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_436_n N_A_492_392#_c_584_n 0.0118344f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_M1004_s N_A_492_392#_c_585_n 0.00305629f $X=2.91 $Y=1.96 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_441_n N_A_492_392#_c_585_n 0.0197787f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_441_n N_A_492_392#_c_587_n 0.0416234f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_442_n N_A_492_392#_c_588_n 0.0125436f $X=5.04 $Y=2.125 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_448_n N_A_492_392#_c_588_n 0.0654702f $X=4.875 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_436_n N_A_492_392#_c_588_n 0.0372602f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_441_n N_A_492_392#_c_589_n 0.0124983f $X=3.045 $Y=2.455 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_448_n N_A_492_392#_c_589_n 0.0179217f $X=4.875 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_436_n N_A_492_392#_c_589_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_442_n N_A_492_392#_c_590_n 0.0656669f $X=5.04 $Y=2.125 $X2=0
+ $Y2=0
cc_347 N_X_c_517_n N_VGND_M1010_d 0.00266f $X=1.475 $Y=1.045 $X2=0 $Y2=0
cc_348 N_X_c_514_n N_VGND_c_638_n 0.0216462f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_349 N_X_c_519_n N_VGND_c_638_n 0.0201602f $X=0.545 $Y=1.295 $X2=0 $Y2=0
cc_350 N_X_c_514_n N_VGND_c_639_n 0.0156021f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_351 N_X_c_517_n N_VGND_c_639_n 0.018932f $X=1.475 $Y=1.045 $X2=0 $Y2=0
cc_352 N_X_c_518_n N_VGND_c_639_n 0.0163623f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_353 N_X_c_518_n N_VGND_c_640_n 0.022799f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_354 N_X_c_514_n N_VGND_c_643_n 0.0109942f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_355 N_X_c_518_n N_VGND_c_644_n 0.0145639f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_356 N_X_c_514_n N_VGND_c_648_n 0.00904371f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_357 N_X_c_518_n N_VGND_c_648_n 0.0119984f $X=1.64 $Y=0.515 $X2=0 $Y2=0

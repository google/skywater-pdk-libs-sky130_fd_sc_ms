* File: sky130_fd_sc_ms__dlclkp_4.pex.spice
* Created: Wed Sep  2 12:04:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%A_84_48# 1 2 7 9 12 15 16 18 19 21 23 24 26
+ 28 30 32 36
c92 36 0 6.50014e-20 $X=0.695 $Y=1.385
r93 38 40 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.6 $Y2=1.385
r94 36 40 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.695 $Y=1.385
+ $X2=0.6 $Y2=1.385
r95 35 37 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.707 $Y=1.385
+ $X2=0.707 $Y2=1.55
r96 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.385 $X2=0.695 $Y2=1.385
r97 32 35 3.67446 $w=3.43e-07 $l=1.1e-07 $layer=LI1_cond $X=0.707 $Y=1.275
+ $X2=0.707 $Y2=1.385
r98 28 30 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.605 $Y=2.685
+ $X2=2.15 $Y2=2.685
r99 24 26 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.605 $Y=0.815
+ $X2=2.06 $Y2=0.815
r100 23 28 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.52 $Y=2.52
+ $X2=1.605 $Y2=2.685
r101 22 23 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.52 $Y=2.14
+ $X2=1.52 $Y2=2.52
r102 20 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.52 $Y=0.98
+ $X2=1.605 $Y2=0.815
r103 20 21 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.52 $Y=0.98
+ $X2=1.52 $Y2=1.19
r104 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=2.055
+ $X2=1.52 $Y2=2.14
r105 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.435 $Y=2.055
+ $X2=0.88 $Y2=2.055
r106 17 32 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.88 $Y=1.275
+ $X2=0.707 $Y2=1.275
r107 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.275
+ $X2=1.52 $Y2=1.19
r108 16 17 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.435 $Y=1.275
+ $X2=0.88 $Y2=1.275
r109 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.795 $Y=1.97
+ $X2=0.88 $Y2=2.055
r110 15 37 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.795 $Y=1.97
+ $X2=0.795 $Y2=1.55
r111 10 40 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.55
+ $X2=0.6 $Y2=1.385
r112 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.6 $Y=1.55 $X2=0.6
+ $Y2=2.4
r113 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r114 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=0.74
r115 2 30 600 $w=1.7e-07 $l=8.62047e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.96 $X2=2.15 $Y2=2.685
r116 1 26 182 $w=1.7e-07 $l=5.21368e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.4 $X2=2.06 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%GATE 3 7 9 12
c36 9 0 6.50014e-20 $X=1.2 $Y=1.665
c37 3 0 2.04382e-19 $X=1.34 $Y=2.46
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.635
+ $X2=1.265 $Y2=1.8
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.635
+ $X2=1.265 $Y2=1.47
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.635 $X2=1.265 $Y2=1.635
r41 7 14 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.355 $Y=0.72
+ $X2=1.355 $Y2=1.47
r42 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.34 $Y=2.46 $X2=1.34
+ $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%A_334_54# 1 2 7 9 12 16 21 24 25 27 28 31
+ 32 33 34 35 36 39 43 47 63
c124 43 0 1.38396e-19 $X=4.37 $Y=2.255
c125 39 0 2.3821e-19 $X=3.98 $Y=0.35
c126 34 0 1.60133e-19 $X=4.205 $Y=2.605
c127 28 0 1.41674e-19 $X=2.065 $Y=2.2
c128 24 0 6.27078e-20 $X=1.9 $Y=1.315
c129 21 0 1.80208e-19 $X=3.695 $Y=0.995
r130 62 63 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.585 $Y=1.795
+ $X2=3.695 $Y2=1.795
r131 51 62 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.49 $Y=1.795
+ $X2=3.585 $Y2=1.795
r132 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.795 $X2=3.49 $Y2=1.795
r133 45 47 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.445 $Y=0.515
+ $X2=4.445 $Y2=0.685
r134 41 43 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.37 $Y=2.52
+ $X2=4.37 $Y2=2.255
r135 39 65 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.98 $Y=0.35
+ $X2=3.695 $Y2=0.35
r136 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.98
+ $Y=0.35 $X2=3.98 $Y2=0.35
r137 36 45 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=4.28 $Y=0.385
+ $X2=4.445 $Y2=0.515
r138 36 38 13.2974 $w=2.58e-07 $l=3e-07 $layer=LI1_cond $X=4.28 $Y=0.385
+ $X2=3.98 $Y2=0.385
r139 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.205 $Y=2.605
+ $X2=4.37 $Y2=2.52
r140 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.205 $Y=2.605
+ $X2=3.475 $Y2=2.605
r141 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.39 $Y=2.52
+ $X2=3.475 $Y2=2.605
r142 32 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.39 $Y=2.35
+ $X2=3.39 $Y2=2.52
r143 31 59 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=2.215
+ $X2=2.47 $Y2=2.38
r144 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=2.215 $X2=2.47 $Y2=2.215
r145 28 30 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=2.065 $Y=2.2
+ $X2=2.47 $Y2=2.2
r146 27 32 8.65646 $w=2.42e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.475 $Y=2.2
+ $X2=3.39 $Y2=2.35
r147 27 50 20.4174 $w=2.42e-07 $l=4.05e-07 $layer=LI1_cond $X=3.475 $Y=2.2
+ $X2=3.475 $Y2=1.795
r148 27 30 32.0763 $w=2.98e-07 $l=8.35e-07 $layer=LI1_cond $X=3.305 $Y=2.2
+ $X2=2.47 $Y2=2.2
r149 25 53 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.9 $Y=1.315
+ $X2=1.745 $Y2=1.315
r150 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9
+ $Y=1.315 $X2=1.9 $Y2=1.315
r151 22 28 6.81904 $w=3e-07 $l=2.10357e-07 $layer=LI1_cond $X=1.92 $Y=2.05
+ $X2=2.065 $Y2=2.2
r152 22 24 29.2085 $w=2.88e-07 $l=7.35e-07 $layer=LI1_cond $X=1.92 $Y=2.05
+ $X2=1.92 $Y2=1.315
r153 19 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.63
+ $X2=3.695 $Y2=1.795
r154 19 21 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.695 $Y=1.63
+ $X2=3.695 $Y2=0.995
r155 18 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=0.515
+ $X2=3.695 $Y2=0.35
r156 18 21 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.695 $Y=0.515
+ $X2=3.695 $Y2=0.995
r157 14 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.96
+ $X2=3.585 $Y2=1.795
r158 14 16 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.585 $Y=1.96
+ $X2=3.585 $Y2=2.54
r159 12 59 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.545 $Y=2.75
+ $X2=2.545 $Y2=2.38
r160 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.15
+ $X2=1.745 $Y2=1.315
r161 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.745 $Y=1.15
+ $X2=1.745 $Y2=0.72
r162 2 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=2.11 $X2=4.37 $Y2=2.255
r163 1 47 182 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.37 $X2=4.445 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%A_334_338# 1 2 7 9 10 11 14 19 20 24 29 32
+ 34
c79 29 0 1.02661e-19 $X=3.91 $Y=2.265
c80 20 0 8.09841e-20 $X=2.47 $Y=1.445
r81 31 34 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.91 $Y=1.485 $X2=3.99
+ $Y2=1.485
r82 31 32 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=1.485
+ $X2=3.825 $Y2=1.485
r83 27 29 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.81 $Y=2.265 $X2=3.91
+ $Y2=2.265
r84 24 38 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.47 $Y=1.64
+ $X2=2.47 $Y2=1.765
r85 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.64
+ $X2=2.47 $Y2=1.475
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.64 $X2=2.47 $Y2=1.64
r87 20 23 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.47 $Y=1.445
+ $X2=2.47 $Y2=1.64
r88 19 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=2.18
+ $X2=3.91 $Y2=2.265
r89 18 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.91 $Y=1.61
+ $X2=3.91 $Y2=1.485
r90 18 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.91 $Y=1.61
+ $X2=3.91 $Y2=2.18
r91 17 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=1.445
+ $X2=2.47 $Y2=1.445
r92 17 32 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.635 $Y=1.445
+ $X2=3.825 $Y2=1.445
r93 14 37 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.38 $Y=0.83
+ $X2=2.38 $Y2=1.475
r94 10 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.47 $Y2=1.765
r95 10 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=1.85 $Y2=1.765
r96 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.76 $Y=1.84
+ $X2=1.85 $Y2=1.765
r97 7 9 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=1.76 $Y=1.84 $X2=1.76
+ $Y2=2.46
r98 2 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=2.12 $X2=3.81 $Y2=2.265
r99 1 34 182 $w=1.7e-07 $l=9.23472e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.625 $X2=3.99 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%A_27_74# 1 2 7 9 14 17 21 26 32 34 37 38 39
+ 40 41 42 43 45 47 48 51 55
c142 55 0 1.86552e-19 $X=5.64 $Y=1.465
c143 41 0 9.8676e-20 $X=2.98 $Y=1.02
c144 40 0 1.39534e-19 $X=2.98 $Y=0.425
c145 14 0 8.09841e-20 $X=2.98 $Y=1.155
c146 9 0 1.02661e-19 $X=2.965 $Y=2.75
r147 55 60 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.465
+ $X2=5.64 $Y2=1.63
r148 55 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.465
+ $X2=5.64 $Y2=1.3
r149 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.465 $X2=5.64 $Y2=1.465
r150 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=0.38 $X2=2.98 $Y2=0.38
r151 47 48 6.41202 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.327 $Y=1.985
+ $X2=0.327 $Y2=1.82
r152 42 54 11.8065 $w=3.72e-07 $l=4.76991e-07 $layer=LI1_cond $X=5.26 $Y=1.105
+ $X2=5.532 $Y2=1.465
r153 42 43 137.984 $w=1.68e-07 $l=2.115e-06 $layer=LI1_cond $X=5.26 $Y=1.105
+ $X2=3.145 $Y2=1.105
r154 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.98 $Y=1.02
+ $X2=3.145 $Y2=1.105
r155 40 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.425
+ $X2=2.98 $Y2=0.34
r156 40 41 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.98 $Y=0.425
+ $X2=2.98 $Y2=1.02
r157 38 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0.34
+ $X2=2.98 $Y2=0.34
r158 38 39 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=2.815 $Y=0.34
+ $X2=1.265 $Y2=0.34
r159 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.18 $Y=0.425
+ $X2=1.265 $Y2=0.34
r160 36 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.18 $Y=0.425
+ $X2=1.18 $Y2=0.85
r161 35 45 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.935
+ $X2=0.24 $Y2=0.935
r162 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.095 $Y=0.935
+ $X2=1.18 $Y2=0.85
r163 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=0.935
+ $X2=0.365 $Y2=0.935
r164 30 47 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=0.327 $Y=2.032
+ $X2=0.327 $Y2=1.985
r165 30 32 21.2321 $w=4.23e-07 $l=7.83e-07 $layer=LI1_cond $X=0.327 $Y=2.032
+ $X2=0.327 $Y2=2.815
r166 28 45 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.02
+ $X2=0.24 $Y2=0.935
r167 28 48 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=0.24 $Y=1.02 $X2=0.24
+ $Y2=1.82
r168 24 45 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.85
+ $X2=0.24 $Y2=0.935
r169 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=0.85
+ $X2=0.24 $Y2=0.515
r170 21 60 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.63 $Y=2.4
+ $X2=5.63 $Y2=1.63
r171 17 59 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.55 $Y=0.74
+ $X2=5.55 $Y2=1.3
r172 14 23 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.98 $Y=1.155
+ $X2=2.98 $Y2=1.44
r173 11 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.98 $Y=0.545
+ $X2=2.98 $Y2=0.38
r174 11 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.98 $Y=0.545
+ $X2=2.98 $Y2=1.155
r175 7 23 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.965 $Y=1.53
+ $X2=2.965 $Y2=1.44
r176 7 9 474.226 $w=1.8e-07 $l=1.22e-06 $layer=POLY_cond $X=2.965 $Y=1.53
+ $X2=2.965 $Y2=2.75
r177 2 47 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.84 $X2=0.375 $Y2=1.985
r178 2 32 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=1.84 $X2=0.375 $Y2=2.815
r179 1 45 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.965
r180 1 26 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%CLK 3 7 11 15 17 27 29
c45 27 0 3.6676e-19 $X=4.905 $Y=1.515
c46 11 0 2.98529e-19 $X=5.145 $Y=2.4
r47 28 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.145 $Y=1.515
+ $X2=5.16 $Y2=1.515
r48 26 28 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.905 $Y=1.515
+ $X2=5.145 $Y2=1.515
r49 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.905
+ $Y=1.515 $X2=4.905 $Y2=1.515
r50 24 26 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.73 $Y=1.515
+ $X2=4.905 $Y2=1.515
r51 23 24 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.595 $Y=1.515
+ $X2=4.73 $Y2=1.515
r52 21 27 9.3293 $w=4.18e-07 $l=3.4e-07 $layer=LI1_cond $X=4.565 $Y=1.57
+ $X2=4.905 $Y2=1.57
r53 20 23 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.565 $Y=1.515
+ $X2=4.595 $Y2=1.515
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.565
+ $Y=1.515 $X2=4.565 $Y2=1.515
r55 17 21 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=4.56 $Y=1.57
+ $X2=4.565 $Y2=1.57
r56 13 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.16 $Y=1.35
+ $X2=5.16 $Y2=1.515
r57 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.16 $Y=1.35
+ $X2=5.16 $Y2=0.74
r58 9 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.68
+ $X2=5.145 $Y2=1.515
r59 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.145 $Y=1.68
+ $X2=5.145 $Y2=2.4
r60 5 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.73 $Y=1.35
+ $X2=4.73 $Y2=1.515
r61 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.73 $Y=1.35 $X2=4.73
+ $Y2=0.74
r62 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=1.68
+ $X2=4.595 $Y2=1.515
r63 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.595 $Y=1.68
+ $X2=4.595 $Y2=2.53
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%A_1047_368# 1 2 7 11 15 19 23 25 26 29 33
+ 37 41 49 51 53 55 57 60 68 69
c127 19 0 1.80414e-19 $X=7.2 $Y=2.4
r128 68 69 98.7966 $w=3.3e-07 $l=5.65e-07 $layer=POLY_cond $X=6.185 $Y=0.835
+ $X2=6.185 $Y2=1.4
r129 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.185
+ $Y=0.835 $X2=6.185 $Y2=0.835
r130 65 67 6.55034 $w=5.96e-07 $l=3.2e-07 $layer=LI1_cond $X=5.975 $Y=0.515
+ $X2=5.975 $Y2=0.835
r131 61 69 12.47 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=6.185 $Y=1.54
+ $X2=6.185 $Y2=1.4
r132 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.185
+ $Y=1.515 $X2=6.185 $Y2=1.515
r133 58 60 9.3732 $w=3.73e-07 $l=3.05e-07 $layer=LI1_cond $X=6.162 $Y=1.82
+ $X2=6.162 $Y2=1.515
r134 57 67 7.70783 $w=5.96e-07 $l=3.77081e-07 $layer=LI1_cond $X=6.162 $Y=1.13
+ $X2=5.975 $Y2=0.835
r135 57 60 11.8317 $w=3.73e-07 $l=3.85e-07 $layer=LI1_cond $X=6.162 $Y=1.13
+ $X2=6.162 $Y2=1.515
r136 56 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=1.905
+ $X2=5.405 $Y2=1.905
r137 55 58 8.1532 $w=1.7e-07 $l=2.2553e-07 $layer=LI1_cond $X=5.975 $Y=1.905
+ $X2=6.162 $Y2=1.82
r138 55 56 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.975 $Y=1.905
+ $X2=5.57 $Y2=1.905
r139 51 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=1.99
+ $X2=5.405 $Y2=1.905
r140 51 53 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=5.405 $Y=1.99
+ $X2=5.405 $Y2=2.815
r141 49 50 1.73381 $w=2.78e-07 $l=1e-08 $layer=POLY_cond $X=8.135 $Y=1.54
+ $X2=8.145 $Y2=1.54
r142 48 49 72.8201 $w=2.78e-07 $l=4.2e-07 $layer=POLY_cond $X=7.715 $Y=1.54
+ $X2=8.135 $Y2=1.54
r143 47 48 5.20144 $w=2.78e-07 $l=3e-08 $layer=POLY_cond $X=7.685 $Y=1.54
+ $X2=7.715 $Y2=1.54
r144 45 46 3.21358 $w=2.8e-07 $l=1.5e-08 $layer=POLY_cond $X=7.2 $Y=1.54
+ $X2=7.215 $Y2=1.54
r145 44 45 88.9092 $w=2.8e-07 $l=4.15e-07 $layer=POLY_cond $X=6.785 $Y=1.54
+ $X2=7.2 $Y2=1.54
r146 43 44 10.7119 $w=2.8e-07 $l=5e-08 $layer=POLY_cond $X=6.735 $Y=1.54
+ $X2=6.785 $Y2=1.54
r147 39 50 17.1848 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=8.145 $Y=1.4
+ $X2=8.145 $Y2=1.54
r148 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.145 $Y=1.4
+ $X2=8.145 $Y2=0.74
r149 35 49 12.9618 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=8.135 $Y=1.68
+ $X2=8.135 $Y2=1.54
r150 35 37 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.135 $Y=1.68
+ $X2=8.135 $Y2=2.4
r151 31 48 17.1848 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=7.715 $Y=1.4
+ $X2=7.715 $Y2=1.54
r152 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.715 $Y=1.4
+ $X2=7.715 $Y2=0.74
r153 27 47 12.9618 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=7.685 $Y=1.68
+ $X2=7.685 $Y2=1.54
r154 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.685 $Y=1.68
+ $X2=7.685 $Y2=2.4
r155 26 46 16.0679 $w=2.8e-07 $l=7.5e-08 $layer=POLY_cond $X=7.29 $Y=1.54
+ $X2=7.215 $Y2=1.54
r156 25 47 15.4929 $w=2.8e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=1.54
+ $X2=7.685 $Y2=1.54
r157 25 26 65.3429 $w=2.8e-07 $l=3.05e-07 $layer=POLY_cond $X=7.595 $Y=1.54
+ $X2=7.29 $Y2=1.54
r158 21 46 17.3521 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=7.215 $Y=1.4
+ $X2=7.215 $Y2=1.54
r159 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.215 $Y=1.4
+ $X2=7.215 $Y2=0.74
r160 17 45 13.127 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=7.2 $Y=1.68 $X2=7.2
+ $Y2=1.54
r161 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.2 $Y=1.68 $X2=7.2
+ $Y2=2.4
r162 13 44 17.3521 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=6.785 $Y=1.4
+ $X2=6.785 $Y2=1.54
r163 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.785 $Y=1.4
+ $X2=6.785 $Y2=0.74
r164 9 43 13.127 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=6.735 $Y=1.68
+ $X2=6.735 $Y2=1.54
r165 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.735 $Y=1.68
+ $X2=6.735 $Y2=2.4
r166 8 61 14.6968 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.35 $Y=1.54
+ $X2=6.185 $Y2=1.54
r167 7 43 19.2815 $w=2.8e-07 $l=9e-08 $layer=POLY_cond $X=6.645 $Y=1.54
+ $X2=6.735 $Y2=1.54
r168 7 8 63.2005 $w=2.8e-07 $l=2.95e-07 $layer=POLY_cond $X=6.645 $Y=1.54
+ $X2=6.35 $Y2=1.54
r169 2 63 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.84 $X2=5.405 $Y2=1.985
r170 2 53 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.84 $X2=5.405 $Y2=2.815
r171 1 65 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.625
+ $Y=0.37 $X2=5.765 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 43 48 49
+ 51 52 53 59 70 74 79 85 88 91 95
r102 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r103 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 83 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r107 83 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r108 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 80 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.42 $Y2=3.33
r110 80 82 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 79 94 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.195 $Y=3.33
+ $X2=8.417 $Y2=3.33
r112 79 82 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.195 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 78 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 78 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 75 88 15.3799 $w=1.7e-07 $l=4.43e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.182 $Y2=3.33
r117 75 77 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.625 $Y=3.33
+ $X2=6.96 $Y2=3.33
r118 74 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=7.42 $Y2=3.33
r119 74 77 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 73 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r122 70 88 15.3799 $w=1.7e-07 $l=4.42e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=6.182 $Y2=3.33
r123 70 72 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r125 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 66 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r127 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r128 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 63 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=3.33
+ $X2=3.275 $Y2=3.33
r130 63 65 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.44 $Y=3.33
+ $X2=3.6 $Y2=3.33
r131 62 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=3.275 $Y2=3.33
r134 59 61 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 57 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 53 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 53 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 51 68 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.74 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=3.33
+ $X2=4.905 $Y2=3.33
r141 50 72 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.07 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=3.33
+ $X2=4.905 $Y2=3.33
r143 48 56 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 48 49 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.972 $Y2=3.33
r145 47 61 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.16 $Y=3.33 $X2=1.2
+ $Y2=3.33
r146 47 49 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.972 $Y2=3.33
r147 43 46 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.36 $Y=2.035
+ $X2=8.36 $Y2=2.815
r148 41 94 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.417 $Y2=3.33
r149 41 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.815
r150 37 40 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=7.42 $Y=2.055
+ $X2=7.42 $Y2=2.815
r151 35 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=3.33
r152 35 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=2.815
r153 31 88 3.31993 $w=8.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=3.33
r154 31 33 13.5785 $w=8.83e-07 $l=9.85e-07 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=2.26
r155 27 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=3.245
+ $X2=4.905 $Y2=3.33
r156 27 29 34.5733 $w=3.28e-07 $l=9.9e-07 $layer=LI1_cond $X=4.905 $Y=3.245
+ $X2=4.905 $Y2=2.255
r157 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=3.245
+ $X2=3.275 $Y2=3.33
r158 23 25 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.275 $Y=3.245
+ $X2=3.275 $Y2=3.025
r159 19 49 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.972 $Y=3.245
+ $X2=0.972 $Y2=3.33
r160 19 21 25.6611 $w=3.73e-07 $l=8.35e-07 $layer=LI1_cond $X=0.972 $Y=3.245
+ $X2=0.972 $Y2=2.41
r161 6 46 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.815
r162 6 43 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.035
r163 5 40 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=7.29
+ $Y=1.84 $X2=7.46 $Y2=2.815
r164 5 37 400 $w=1.7e-07 $l=2.87706e-07 $layer=licon1_PDIFF $count=1 $X=7.29
+ $Y=1.84 $X2=7.46 $Y2=2.055
r165 4 33 150 $w=1.7e-07 $l=9.26499e-07 $layer=licon1_PDIFF $count=4 $X=5.72
+ $Y=1.84 $X2=6.46 $Y2=2.26
r166 3 29 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=4.685
+ $Y=2.11 $X2=4.905 $Y2=2.255
r167 2 25 600 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=2.54 $X2=3.275 $Y2=3.025
r168 1 21 300 $w=1.7e-07 $l=6.9401e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=1.84 $X2=0.965 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%GCLK 1 2 3 4 15 21 23 24 25 26 29 35 38 39
+ 40 41
c75 40 0 1.80414e-19 $X=7.92 $Y=1.665
r76 41 44 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=8.4 $Y=1.665
+ $X2=8.015 $Y2=1.665
r77 40 44 3.48671 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=7.88 $Y=1.665
+ $X2=8.015 $Y2=1.665
r78 38 40 2.63492 $w=2.1e-07 $l=1.29132e-07 $layer=LI1_cond $X=7.91 $Y=1.55
+ $X2=7.88 $Y2=1.665
r79 37 39 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=7.91 $Y=1.38
+ $X2=7.89 $Y2=1.295
r80 37 38 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=7.91 $Y=1.38
+ $X2=7.91 $Y2=1.55
r81 33 39 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=1.21 $X2=7.89
+ $Y2=1.295
r82 33 35 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=7.89 $Y=1.21
+ $X2=7.89 $Y2=0.515
r83 29 31 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.87 $Y=1.985
+ $X2=7.87 $Y2=2.815
r84 27 40 2.63492 $w=2.5e-07 $l=1.19896e-07 $layer=LI1_cond $X=7.87 $Y=1.78
+ $X2=7.88 $Y2=1.665
r85 27 29 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=7.87 $Y=1.78
+ $X2=7.87 $Y2=1.985
r86 25 39 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.765 $Y=1.295
+ $X2=7.89 $Y2=1.295
r87 25 26 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.765 $Y=1.295
+ $X2=7.165 $Y2=1.295
r88 23 40 3.48671 $w=1.7e-07 $l=1.49248e-07 $layer=LI1_cond $X=7.745 $Y=1.635
+ $X2=7.88 $Y2=1.665
r89 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.745 $Y=1.635
+ $X2=7.125 $Y2=1.635
r90 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7 $Y=1.21
+ $X2=7.165 $Y2=1.295
r91 19 21 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7 $Y=1.21 $X2=7
+ $Y2=0.515
r92 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.96 $Y=1.985
+ $X2=6.96 $Y2=2.815
r93 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.96 $Y=1.72
+ $X2=7.125 $Y2=1.635
r94 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.96 $Y=1.72
+ $X2=6.96 $Y2=1.985
r95 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.91 $Y2=2.815
r96 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.91 $Y2=1.985
r97 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.84 $X2=6.96 $Y2=2.815
r98 3 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.84 $X2=6.96 $Y2=1.985
r99 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
r100 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.86
+ $Y=0.37 $X2=7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_4%VGND 1 2 3 4 5 6 21 25 29 33 35 37 39 41 46
+ 54 59 64 69 75 78 81 91 95
r98 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r99 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r100 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r102 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 73 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r104 73 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r105 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r106 70 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.46
+ $Y2=0
r107 70 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.585 $Y=0
+ $X2=7.92 $Y2=0
r108 69 94 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.195 $Y=0
+ $X2=8.417 $Y2=0
r109 69 72 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.195 $Y=0
+ $X2=7.92 $Y2=0
r110 68 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r111 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r112 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r113 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.655 $Y=0
+ $X2=6.96 $Y2=0
r114 64 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.46
+ $Y2=0
r115 64 67 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r116 63 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r117 63 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r118 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r119 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=4.945
+ $Y2=0
r120 60 62 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=6
+ $Y2=0
r121 59 88 8.09467 $w=4.93e-07 $l=3.35e-07 $layer=LI1_cond $X=6.407 $Y=0
+ $X2=6.407 $Y2=0.335
r122 59 65 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=6.407 $Y=0
+ $X2=6.655 $Y2=0
r123 59 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r124 59 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.16 $Y=0 $X2=6
+ $Y2=0
r125 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r126 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r127 55 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.48
+ $Y2=0
r128 55 57 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.645 $Y=0
+ $X2=4.56 $Y2=0
r129 54 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=0 $X2=4.945
+ $Y2=0
r130 54 57 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.78 $Y=0 $X2=4.56
+ $Y2=0
r131 53 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r132 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r133 50 53 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r134 50 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r135 49 52 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r136 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r137 47 75 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.925 $Y=0
+ $X2=0.737 $Y2=0
r138 47 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.2
+ $Y2=0
r139 46 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.48
+ $Y2=0
r140 46 52 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.12 $Y2=0
r141 44 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r143 41 75 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.737
+ $Y2=0
r144 41 43 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r145 39 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r146 39 79 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.6
+ $Y2=0
r147 35 94 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.36 $Y=0.085
+ $X2=8.417 $Y2=0
r148 35 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.36 $Y=0.085
+ $X2=8.36 $Y2=0.515
r149 31 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0
r150 31 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0.515
r151 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=0.085
+ $X2=4.945 $Y2=0
r152 27 29 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=4.945 $Y=0.085
+ $X2=4.945 $Y2=0.685
r153 23 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=0.085
+ $X2=3.48 $Y2=0
r154 23 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.48 $Y=0.085
+ $X2=3.48 $Y2=0.765
r155 19 75 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0
r156 19 21 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0.515
r157 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.515
r158 5 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.29
+ $Y=0.37 $X2=7.5 $Y2=0.515
r159 4 88 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.19 $X2=6.405 $Y2=0.335
r160 3 29 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=4.805
+ $Y=0.37 $X2=4.945 $Y2=0.685
r161 2 25 182 $w=1.7e-07 $l=5.07075e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.945 $X2=3.48 $Y2=0.765
r162 1 21 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.735 $Y2=0.515
.ends


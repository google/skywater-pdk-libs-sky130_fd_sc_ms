* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
X0 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 a_357_392# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 a_897_406# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X5 a_796_508# a_897_406# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X6 VPWR a_897_406# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_657_392# a_232_98# a_796_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X8 a_357_392# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_681_74# a_232_98# a_657_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_1139_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_573_392# a_357_392# a_657_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X13 a_897_406# a_657_392# a_1139_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR a_657_392# a_897_406# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 VGND a_27_136# a_681_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_657_392# a_357_392# a_854_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 VPWR a_27_136# a_573_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X18 a_854_74# a_897_406# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 VGND a_897_406# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

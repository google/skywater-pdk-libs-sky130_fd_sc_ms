* File: sky130_fd_sc_ms__o32ai_1.spice
* Created: Fri Aug 28 18:04:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o32ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o32ai_1  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_Y_M1009_d N_B1_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.21645 AS=0.2109 PD=1.325 PS=2.05 NRD=30 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1003_d N_B2_M1003_g N_Y_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.21645 PD=1.09 PS=1.325 NRD=11.34 NRS=19.452 M=1 R=4.93333
+ SA=75000.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A3_M1000_g N_A_27_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1665 AS=0.1295 PD=1.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_74#_M1007_d N_A2_M1007_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1665 PD=1.02 PS=1.19 NRD=0 NRS=16.212 M=1 R=4.93333 SA=75002
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_27_74#_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 A_131_368# N_B1_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3584 PD=1.36 PS=2.88 NRD=11.426 NRS=6.1464 M=1 R=6.22222 SA=90000.2
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_B2_M1008_g A_131_368# VPB PSHORT L=0.18 W=1.12 AD=0.2632
+ AS=0.1344 PD=1.59 PS=1.36 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90000.6 SB=90002
+ A=0.2016 P=2.6 MULT=1
MM1002 A_345_368# N_A3_M1002_g N_Y_M1008_d VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2632 PD=1.51 PS=1.59 NRD=24.6053 NRS=34.2977 M=1 R=6.22222 SA=90001.3
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1005 A_459_368# N_A2_M1005_g A_345_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=24.6053 M=1 R=6.22222 SA=90001.9
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_459_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90002.4 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__o32ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__clkdlyinv5sd2_1.spice
* Created: Fri Aug 28 17:18:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkdlyinv5sd2_1.pex.spice"
.subckt sky130_fd_sc_ms__clkdlyinv5sd2_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_28_74#_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.14805 AS=0.1113 PD=1.125 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_A_288_74#_M1005_d N_A_28_74#_M1005_g N_VGND_M1007_d VNB NLOWVT L=0.18
+ W=0.42 AD=0.1113 AS=0.14805 PD=1.37 PS=1.125 NRD=0 NRS=105.708 M=1 R=2.33333
+ SA=90001 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_A_549_74#_M1000_d N_A_288_74#_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.18
+ W=0.42 AD=0.1113 AS=0.2478 PD=1.37 PS=2.02 NRD=0 NRS=91.428 M=1 R=2.33333
+ SA=90000.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1001 N_VGND_M1001_d N_A_549_74#_M1001_g N_A_682_74#_M1001_s VNB NLOWVT L=0.18
+ W=0.42 AD=0.0966 AS=0.2457 PD=0.88 PS=2.01 NRD=51.42 NRS=91.428 M=1 R=2.33333
+ SA=90000.5 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1002 N_Y_M1002_d N_A_682_74#_M1002_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0966 PD=1.37 PS=0.88 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_28_74#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.338113 AS=0.2968 PD=1.82792 PS=2.77 NRD=2.6201 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1009 N_A_288_74#_M1009_d N_A_28_74#_M1009_g N_VPWR_M1006_d VPB PSHORT L=0.25
+ W=1 AD=0.26 AS=0.301887 PD=2.52 PS=1.63208 NRD=0 NRS=62.0353 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1003 N_A_549_74#_M1003_d N_A_288_74#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.25
+ W=1 AD=0.265 AS=0.52 PD=2.53 PS=3.04 NRD=0 NRS=50.2153 M=1 R=4 SA=125000
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_549_74#_M1004_g N_A_682_74#_M1004_s VPB PSHORT L=0.25
+ W=1 AD=0.231698 AS=0.51 PD=1.49057 PS=3.02 NRD=36.7602 NRS=48.265 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1008 N_Y_M1008_d N_A_682_74#_M1008_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2968 AS=0.259502 PD=2.77 PS=1.66943 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ms__clkdlyinv5sd2_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand3_1.spice
* Created: Fri Aug 28 17:43:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand3_1.pex.spice"
.subckt sky130_fd_sc_ms__nand3_1  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1002 A_155_74# N_C_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1001 A_233_74# N_B_M1001_g A_155_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g A_233_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.2 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_C_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.4032 PD=1.39 PS=2.96 NRD=0 NRS=13.1793 M=1 R=6.22222 SA=90000.3
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_Y_M1003_d VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1512 PD=1.51 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.7 SB=90000.8
+ A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90001.3 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__nand3_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__einvn_8.spice
* Created: Wed Sep  2 12:08:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__einvn_8.pex.spice"
.subckt sky130_fd_sc_ms__einvn_8  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1002 N_A_126_74#_M1002_d N_TE_B_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_293_74#_M1003_d N_A_126_74#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75007 A=0.111 P=1.78 MULT=1
MM1005 N_A_293_74#_M1005_d N_A_126_74#_M1005_g N_VGND_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75006.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_293_74#_M1005_d N_A_126_74#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75006.1 A=0.111 P=1.78 MULT=1
MM1015 N_A_293_74#_M1015_d N_A_126_74#_M1015_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75005.6 A=0.111 P=1.78 MULT=1
MM1016 N_A_293_74#_M1015_d N_A_126_74#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75005.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_293_74#_M1022_d N_A_126_74#_M1022_g N_VGND_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.5 SB=75004.7 A=0.111 P=1.78 MULT=1
MM1029 N_A_293_74#_M1022_d N_A_126_74#_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75004.3 A=0.111 P=1.78 MULT=1
MM1031 N_A_293_74#_M1031_d N_A_126_74#_M1031_g N_VGND_M1029_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.4 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1006 N_Z_M1006_d N_A_M1006_g N_A_293_74#_M1031_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.8
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1011 N_Z_M1006_d N_A_M1011_g N_A_293_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.2
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1013 N_Z_M1013_d N_A_M1013_g N_A_293_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.6
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1014 N_Z_M1013_d N_A_M1014_g N_A_293_74#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75005.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1018 N_Z_M1018_d N_A_M1018_g N_A_293_74#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.6
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1024 N_Z_M1018_d N_A_M1024_g N_A_293_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1027 N_Z_M1027_d N_A_M1027_g N_A_293_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.4
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1030 N_Z_M1027_d N_A_M1030_g N_A_293_74#_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_126_74#_M1009_d N_TE_B_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3696 PD=2.8 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_A_239_368#_M1017_d N_TE_B_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90007.2 A=0.2016 P=2.6 MULT=1
MM1019 N_A_239_368#_M1019_d N_TE_B_M1019_g N_VPWR_M1017_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.7 SB=90006.7 A=0.2016 P=2.6 MULT=1
MM1020 N_A_239_368#_M1019_d N_TE_B_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90006.3 A=0.2016 P=2.6 MULT=1
MM1021 N_A_239_368#_M1021_d N_TE_B_M1021_g N_VPWR_M1020_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.6 SB=90005.8 A=0.2016 P=2.6 MULT=1
MM1023 N_A_239_368#_M1021_d N_TE_B_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.1 SB=90005.3 A=0.2016 P=2.6 MULT=1
MM1025 N_A_239_368#_M1025_d N_TE_B_M1025_g N_VPWR_M1023_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.6 SB=90004.8 A=0.2016 P=2.6 MULT=1
MM1026 N_A_239_368#_M1025_d N_TE_B_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90003 SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1028 N_A_239_368#_M1028_d N_TE_B_M1028_g N_VPWR_M1026_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90003.6 SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1000 N_A_239_368#_M1028_d N_A_M1000_g N_Z_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1001 N_A_239_368#_M1001_d N_A_M1001_g N_Z_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.5
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1004 N_A_239_368#_M1001_d N_A_M1004_g N_Z_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.9
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1007 N_A_239_368#_M1007_d N_A_M1007_g N_Z_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.4
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1010 N_A_239_368#_M1007_d N_A_M1010_g N_Z_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.9
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1012 N_A_239_368#_M1012_d N_A_M1012_g N_Z_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.3
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1032 N_A_239_368#_M1012_d N_A_M1032_g N_Z_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.8
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1033 N_A_239_368#_M1033_d N_A_M1033_g N_Z_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ms__einvn_8.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlrtn_4.pex.spice
* Created: Wed Sep  2 12:05:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRTN_4%D 3 7 9 12
r33 12 15 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.615
+ $X2=0.587 $Y2=1.78
r34 12 14 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.615
+ $X2=0.587 $Y2=1.45
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.615 $X2=0.59 $Y2=1.615
r36 9 13 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.59 $Y2=1.615
r37 7 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.535 $Y=2.39
+ $X2=0.535 $Y2=1.78
r38 3 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=0.955
+ $X2=0.495 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%GATE_N 3 7 9 12
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.615
+ $X2=1.13 $Y2=1.78
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.615
+ $X2=1.13 $Y2=1.45
r39 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.615 $X2=1.13 $Y2=1.615
r40 7 14 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.085 $Y=0.86
+ $X2=1.085 $Y2=1.45
r41 3 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.085 $Y=2.39
+ $X2=1.085 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%A_232_98# 1 2 9 13 17 21 23 24 26 27 32 37
+ 38 41 42 45 46 48 50
c119 24 0 1.26581e-19 $X=2.02 $Y=1.42
r120 48 51 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.662 $Y=1.585
+ $X2=1.662 $Y2=1.75
r121 48 50 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.662 $Y=1.585
+ $X2=1.662 $Y2=1.42
r122 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.585 $X2=1.7 $Y2=1.585
r123 46 51 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.545 $Y=1.95
+ $X2=1.545 $Y2=1.75
r124 45 46 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.387 $Y=2.115
+ $X2=1.387 $Y2=1.95
r125 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=2.195 $X2=4.035 $Y2=2.195
r126 39 41 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.035 $Y=2.6
+ $X2=4.035 $Y2=2.195
r127 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.87 $Y=2.685
+ $X2=4.035 $Y2=2.6
r128 37 38 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=3.87 $Y=2.685
+ $X2=1.63 $Y2=2.685
r129 33 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.545 $Y=1.25
+ $X2=1.545 $Y2=1.42
r130 32 38 9.10402 $w=1.7e-07 $l=2.82319e-07 $layer=LI1_cond $X=1.387 $Y=2.6
+ $X2=1.63 $Y2=2.685
r131 31 45 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=1.387 $Y=2.192
+ $X2=1.387 $Y2=2.115
r132 31 32 10.0619 $w=4.83e-07 $l=4.08e-07 $layer=LI1_cond $X=1.387 $Y=2.192
+ $X2=1.387 $Y2=2.6
r133 27 33 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.46 $Y=1.125
+ $X2=1.545 $Y2=1.25
r134 27 29 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.46 $Y=1.125
+ $X2=1.35 $Y2=1.125
r135 25 42 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.75 $Y=2.195
+ $X2=4.035 $Y2=2.195
r136 25 26 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.75 $Y=2.195
+ $X2=3.66 $Y2=2.195
r137 23 49 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.02 $Y=1.585
+ $X2=1.7 $Y2=1.585
r138 23 24 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.02 $Y=1.585
+ $X2=2.02 $Y2=1.42
r139 19 26 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=2.36
+ $X2=3.66 $Y2=2.195
r140 19 21 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.66 $Y=2.36
+ $X2=3.66 $Y2=2.73
r141 15 26 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.645 $Y=2.03
+ $X2=3.66 $Y2=2.195
r142 15 17 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=3.645 $Y=2.03
+ $X2=3.645 $Y2=0.69
r143 11 24 34.7346 $w=1.65e-07 $l=1.6e-07 $layer=POLY_cond $X=2.18 $Y=1.42
+ $X2=2.02 $Y2=1.42
r144 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.18 $Y=1.42
+ $X2=2.18 $Y2=0.86
r145 7 24 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=2.11 $Y=1.75
+ $X2=2.02 $Y2=1.42
r146 7 9 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.11 $Y=1.75 $X2=2.11
+ $Y2=2.38
r147 2 45 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.175
+ $Y=1.97 $X2=1.31 $Y2=2.115
r148 1 29 182 $w=1.7e-07 $l=6.83429e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.35 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%A_27_136# 1 2 7 9 11 13 15 19 24 25 28 31 33
+ 34
c81 28 0 1.26581e-19 $X=2.655 $Y=1.505
c82 7 0 1.51556e-19 $X=2.73 $Y=1.67
r83 33 34 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=1.95
r84 31 34 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.17 $Y=1.25 $X2=0.17
+ $Y2=1.95
r85 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.505 $X2=2.655 $Y2=1.505
r86 26 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.655 $Y=0.83
+ $X2=2.655 $Y2=1.505
r87 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.49 $Y=0.745
+ $X2=2.655 $Y2=0.83
r88 24 25 133.417 $w=1.68e-07 $l=2.045e-06 $layer=LI1_cond $X=2.49 $Y=0.745
+ $X2=0.445 $Y2=0.745
r89 17 31 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=1.25
r90 17 19 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=0.955
r91 16 25 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.445 $Y2=0.745
r92 16 19 4.00154 $w=3.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.955
r93 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.255 $Y=1.085
+ $X2=3.255 $Y2=0.69
r94 12 29 66.251 $w=2.51e-07 $l=4.19464e-07 $layer=POLY_cond $X=2.82 $Y=1.16
+ $X2=2.655 $Y2=1.505
r95 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.18 $Y=1.16
+ $X2=3.255 $Y2=1.085
r96 11 12 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.18 $Y=1.16
+ $X2=2.82 $Y2=1.16
r97 7 29 35.6167 $w=2.51e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.73 $Y=1.67
+ $X2=2.655 $Y2=1.505
r98 7 9 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.73 $Y=1.67 $X2=2.73
+ $Y2=2.46
r99 2 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.97 $X2=0.31 $Y2=2.115
r100 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%A_348_392# 1 2 9 13 16 17 22 23 24 26 27 32
+ 38
c94 32 0 1.51556e-19 $X=2.12 $Y=1.125
r95 37 38 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=2.175
+ $X2=2.205 $Y2=2.175
r96 35 37 5.51134 $w=5.08e-07 $l=2.35e-07 $layer=LI1_cond $X=1.885 $Y=2.175
+ $X2=2.12 $Y2=2.175
r97 30 32 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=1.965 $Y=1.125
+ $X2=2.12 $Y2=1.125
r98 27 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=1.355
+ $X2=4.095 $Y2=1.19
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=1.355 $X2=4.095 $Y2=1.355
r100 24 26 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=3.36 $Y=1.355
+ $X2=4.095 $Y2=1.355
r101 23 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.61
+ $X2=3.195 $Y2=1.775
r102 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.61 $X2=3.195 $Y2=1.61
r103 20 22 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.195 $Y=1.92
+ $X2=3.195 $Y2=1.61
r104 19 24 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.195 $Y=1.52
+ $X2=3.36 $Y2=1.355
r105 19 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.195 $Y=1.52
+ $X2=3.195 $Y2=1.61
r106 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.03 $Y=2.005
+ $X2=3.195 $Y2=1.92
r107 17 38 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.03 $Y=2.005
+ $X2=2.205 $Y2=2.005
r108 16 37 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.12 $Y=1.92
+ $X2=2.12 $Y2=2.175
r109 15 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=1.25
+ $X2=2.12 $Y2=1.125
r110 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.12 $Y=1.25
+ $X2=2.12 $Y2=1.92
r111 13 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.12 $Y=0.58
+ $X2=4.12 $Y2=1.19
r112 9 41 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=3.12 $Y=2.46
+ $X2=3.12 $Y2=1.775
r113 2 35 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.96 $X2=1.885 $Y2=2.185
r114 1 30 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.49 $X2=1.965 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%A_888_406# 1 2 3 12 16 18 22 24 25 28 32 36
+ 40 44 48 52 55 58 61 66 68 72 81 84 86 87 88 89 91 100
c186 48 0 1.5942e-19 $X=8.985 $Y=2.4
r187 97 98 36.6076 $w=3.16e-07 $l=2.4e-07 $layer=POLY_cond $X=8.435 $Y=1.465
+ $X2=8.675 $Y2=1.465
r188 96 97 28.981 $w=3.16e-07 $l=1.9e-07 $layer=POLY_cond $X=8.245 $Y=1.465
+ $X2=8.435 $Y2=1.465
r189 93 94 18.3038 $w=3.16e-07 $l=1.2e-07 $layer=POLY_cond $X=7.815 $Y=1.465
+ $X2=7.935 $Y2=1.465
r190 88 89 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.725 $Y=1.545
+ $X2=7.895 $Y2=1.545
r191 82 100 11.4399 $w=3.16e-07 $l=7.5e-08 $layer=POLY_cond $X=8.91 $Y=1.465
+ $X2=8.985 $Y2=1.465
r192 82 98 35.8449 $w=3.16e-07 $l=2.35e-07 $layer=POLY_cond $X=8.91 $Y=1.465
+ $X2=8.675 $Y2=1.465
r193 81 82 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.91
+ $Y=1.465 $X2=8.91 $Y2=1.465
r194 79 96 2.28797 $w=3.16e-07 $l=1.5e-08 $layer=POLY_cond $X=8.23 $Y=1.465
+ $X2=8.245 $Y2=1.465
r195 79 94 44.9968 $w=3.16e-07 $l=2.95e-07 $layer=POLY_cond $X=8.23 $Y=1.465
+ $X2=7.935 $Y2=1.465
r196 78 81 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.23 $Y=1.465
+ $X2=8.91 $Y2=1.465
r197 78 89 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.23 $Y=1.465
+ $X2=7.895 $Y2=1.465
r198 78 79 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=1.465 $X2=8.23 $Y2=1.465
r199 75 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.82 $Y=1.705
+ $X2=6.655 $Y2=1.705
r200 75 88 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.82 $Y=1.705
+ $X2=7.725 $Y2=1.705
r201 70 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=1.79
+ $X2=6.655 $Y2=1.705
r202 70 72 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.655 $Y=1.79
+ $X2=6.655 $Y2=2.245
r203 69 84 2.76166 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.835 $Y=1.705
+ $X2=5.662 $Y2=1.705
r204 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=1.705
+ $X2=6.655 $Y2=1.705
r205 68 69 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.49 $Y=1.705
+ $X2=5.835 $Y2=1.705
r206 64 84 3.70735 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=5.75 $Y=1.62
+ $X2=5.662 $Y2=1.705
r207 64 66 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.75 $Y=1.62
+ $X2=5.75 $Y2=0.81
r208 61 86 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=2.03
+ $X2=5.655 $Y2=2.195
r209 60 84 3.70735 $w=2.5e-07 $l=8.84308e-08 $layer=LI1_cond $X=5.655 $Y=1.79
+ $X2=5.662 $Y2=1.705
r210 60 61 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.655 $Y=1.79
+ $X2=5.655 $Y2=2.03
r211 58 92 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=2.195
+ $X2=4.605 $Y2=2.36
r212 58 91 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=2.195
+ $X2=4.605 $Y2=2.03
r213 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.605
+ $Y=2.195 $X2=4.605 $Y2=2.195
r214 55 86 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=2.195
+ $X2=5.655 $Y2=2.195
r215 55 57 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=5.49 $Y=2.195
+ $X2=4.605 $Y2=2.195
r216 50 100 18.3038 $w=3.16e-07 $l=2.16852e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=8.985 $Y2=1.465
r217 50 52 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=9.105 $Y2=0.74
r218 46 100 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.985 $Y=1.63
+ $X2=8.985 $Y2=1.465
r219 46 48 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.985 $Y=1.63
+ $X2=8.985 $Y2=2.4
r220 42 98 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=1.465
r221 42 44 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=0.74
r222 38 97 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.435 $Y=1.63
+ $X2=8.435 $Y2=1.465
r223 38 40 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.435 $Y=1.63
+ $X2=8.435 $Y2=2.4
r224 34 96 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=1.465
r225 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=0.74
r226 30 94 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.935 $Y=1.63
+ $X2=7.935 $Y2=1.465
r227 30 32 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.935 $Y=1.63
+ $X2=7.935 $Y2=2.4
r228 26 93 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=1.3
+ $X2=7.815 $Y2=1.465
r229 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.815 $Y=1.3
+ $X2=7.815 $Y2=0.74
r230 24 93 24.8104 $w=3.16e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.74 $Y=1.555
+ $X2=7.815 $Y2=1.465
r231 24 25 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.74 $Y=1.555
+ $X2=7.575 $Y2=1.555
r232 20 25 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.485 $Y=1.63
+ $X2=7.575 $Y2=1.555
r233 20 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.485 $Y=1.63
+ $X2=7.485 $Y2=2.4
r234 18 54 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.56 $Y=1.825
+ $X2=4.56 $Y2=1.735
r235 18 91 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=4.56 $Y=1.825
+ $X2=4.56 $Y2=2.03
r236 16 54 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=4.545 $Y=0.58
+ $X2=4.545 $Y2=1.735
r237 12 92 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.53 $Y=2.73
+ $X2=4.53 $Y2=2.36
r238 3 72 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=6.47
+ $Y=2.1 $X2=6.655 $Y2=2.245
r239 2 86 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.52
+ $Y=2.1 $X2=5.655 $Y2=2.245
r240 1 66 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.37 $X2=5.75 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%A_642_392# 1 2 9 11 13 16 18 20 21 26 27 28
+ 31 33 34 35 36 44
c116 44 0 1.47145e-19 $X=5.88 $Y=1.455
r117 44 45 6.42163 $w=6.38e-07 $l=8.5e-08 $layer=POLY_cond $X=5.88 $Y=1.455
+ $X2=5.965 $Y2=1.455
r118 43 44 26.0643 $w=6.38e-07 $l=3.45e-07 $layer=POLY_cond $X=5.535 $Y=1.455
+ $X2=5.88 $Y2=1.455
r119 42 43 7.9326 $w=6.38e-07 $l=1.05e-07 $layer=POLY_cond $X=5.43 $Y=1.455
+ $X2=5.535 $Y2=1.455
r120 40 42 28.3307 $w=6.38e-07 $l=3.75e-07 $layer=POLY_cond $X=5.055 $Y=1.455
+ $X2=5.43 $Y2=1.455
r121 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.055
+ $Y=1.285 $X2=5.055 $Y2=1.285
r122 37 39 15.8148 $w=2.7e-07 $l=3.5e-07 $layer=LI1_cond $X=4.985 $Y=0.935
+ $X2=4.985 $Y2=1.285
r123 35 39 2.4733 $w=4.05e-07 $l=5.05272e-08 $layer=LI1_cond $X=5.017 $Y=1.322
+ $X2=4.985 $Y2=1.285
r124 35 36 10.4716 $w=4.03e-07 $l=3.68e-07 $layer=LI1_cond $X=5.017 $Y=1.322
+ $X2=5.017 $Y2=1.69
r125 33 37 3.44395 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.815 $Y=0.935
+ $X2=4.985 $Y2=0.935
r126 33 34 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.815 $Y=0.935
+ $X2=4.07 $Y2=0.935
r127 29 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.905 $Y=0.85
+ $X2=4.07 $Y2=0.935
r128 29 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.905 $Y=0.85
+ $X2=3.905 $Y2=0.565
r129 27 36 8.41448 $w=1.7e-07 $l=2.40778e-07 $layer=LI1_cond $X=4.815 $Y=1.775
+ $X2=5.017 $Y2=1.69
r130 27 28 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=4.815 $Y=1.775
+ $X2=3.7 $Y2=1.775
r131 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=1.86
+ $X2=3.7 $Y2=1.775
r132 25 26 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.615 $Y=1.86
+ $X2=3.615 $Y2=2.26
r133 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=2.345
+ $X2=3.615 $Y2=2.26
r134 21 23 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.53 $Y=2.345
+ $X2=3.345 $Y2=2.345
r135 18 45 37.6732 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.965 $Y=1.12
+ $X2=5.965 $Y2=1.455
r136 18 20 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.965 $Y=1.12
+ $X2=5.965 $Y2=0.69
r137 14 44 32.9664 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=5.88 $Y=1.79
+ $X2=5.88 $Y2=1.455
r138 14 16 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.88 $Y=1.79
+ $X2=5.88 $Y2=2.52
r139 11 43 37.6732 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.535 $Y=1.12
+ $X2=5.535 $Y2=1.455
r140 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.535 $Y=1.12
+ $X2=5.535 $Y2=0.69
r141 7 42 32.9664 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=5.43 $Y=1.79
+ $X2=5.43 $Y2=1.455
r142 7 9 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.43 $Y=1.79 $X2=5.43
+ $Y2=2.52
r143 2 23 600 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.96 $X2=3.345 $Y2=2.345
r144 1 31 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.37 $X2=3.905 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%RESET_B 3 5 7 8 10 13 15 16 17 24
r56 24 26 7.94506 $w=4.55e-07 $l=7.5e-08 $layer=POLY_cond $X=6.825 $Y=1.355
+ $X2=6.9 $Y2=1.355
r57 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.825
+ $Y=1.285 $X2=6.825 $Y2=1.285
r58 22 24 45.5516 $w=4.55e-07 $l=4.3e-07 $layer=POLY_cond $X=6.395 $Y=1.355
+ $X2=6.825 $Y2=1.355
r59 21 22 1.58901 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=6.38 $Y=1.355
+ $X2=6.395 $Y2=1.355
r60 16 17 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.285
+ $X2=7.44 $Y2=1.285
r61 16 25 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.96 $Y=1.285
+ $X2=6.825 $Y2=1.285
r62 15 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.48 $Y=1.285
+ $X2=6.825 $Y2=1.285
r63 11 26 24.5593 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.9 $Y=1.59 $X2=6.9
+ $Y2=1.355
r64 11 13 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=6.9 $Y=1.59 $X2=6.9
+ $Y2=2.52
r65 8 24 29.0417 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.825 $Y=1.12
+ $X2=6.825 $Y2=1.355
r66 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.825 $Y=1.12
+ $X2=6.825 $Y2=0.69
r67 5 22 29.0417 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.395 $Y=1.12
+ $X2=6.395 $Y2=1.355
r68 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.395 $Y=1.12
+ $X2=6.395 $Y2=0.69
r69 1 21 24.5593 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.38 $Y=1.59
+ $X2=6.38 $Y2=1.355
r70 1 3 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=6.38 $Y=1.59 $X2=6.38
+ $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%VPWR 1 2 3 4 5 6 7 26 28 32 36 40 42 44 47
+ 50 54 55 57 58 59 82 87 92 95 97 101
r107 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r108 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r109 94 95 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=3.022
+ $X2=5.32 $Y2=3.022
r110 91 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r111 90 94 1.75222 $w=7.83e-07 $l=1.15e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=5.155 $Y2=3.022
r112 90 92 15.6839 $w=7.83e-07 $l=4.5e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=4.59 $Y2=3.022
r113 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r114 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 85 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 82 100 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=9.045 $Y=3.33
+ $X2=9.322 $Y2=3.33
r118 82 84 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 81 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r120 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 78 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33 $X2=6
+ $Y2=3.33
r123 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 75 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=3.33
+ $X2=6.155 $Y2=3.33
r125 75 77 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.32 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 73 92 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=4.59
+ $Y2=3.33
r127 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 71 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r129 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r130 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r131 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r133 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r134 64 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r135 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r136 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r137 61 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r138 61 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 59 91 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r140 59 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 57 80 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=7.92 $Y2=3.33
r142 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=8.21 $Y2=3.33
r143 56 84 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.88 $Y2=3.33
r144 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.21 $Y2=3.33
r145 54 77 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=6.96 $Y2=3.33
r146 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=7.21 $Y2=3.33
r147 53 80 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.375 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=3.33
+ $X2=7.21 $Y2=3.33
r149 51 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=2.64 $Y2=3.33
r150 50 66 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r151 49 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.585 $Y2=3.33
r152 49 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.255 $Y2=3.33
r153 47 49 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.42 $Y=3.025
+ $X2=2.42 $Y2=3.33
r154 42 100 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=9.21 $Y=3.245
+ $X2=9.322 $Y2=3.33
r155 42 44 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=9.21 $Y=3.245
+ $X2=9.21 $Y2=2.305
r156 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=3.33
r157 38 40 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=2.465
r158 34 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.21 $Y=3.245
+ $X2=7.21 $Y2=3.33
r159 34 36 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=7.21 $Y=3.245
+ $X2=7.21 $Y2=2.245
r160 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=3.33
r161 30 32 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=2.245
r162 28 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=6.155 $Y2=3.33
r163 28 95 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=5.32 $Y2=3.33
r164 24 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r165 24 26 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.115
r166 7 44 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=9.075
+ $Y=1.84 $X2=9.21 $Y2=2.305
r167 6 40 300 $w=1.7e-07 $l=7.11512e-07 $layer=licon1_PDIFF $count=2 $X=8.025
+ $Y=1.84 $X2=8.21 $Y2=2.465
r168 5 36 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=6.99
+ $Y=2.1 $X2=7.21 $Y2=2.245
r169 4 32 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.1 $X2=6.155 $Y2=2.245
r170 3 94 300 $w=1.7e-07 $l=6.58293e-07 $layer=licon1_PDIFF $count=2 $X=4.62
+ $Y=2.52 $X2=5.155 $Y2=2.795
r171 2 47 600 $w=1.7e-07 $l=1.16984e-06 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=1.96 $X2=2.42 $Y2=3.025
r172 1 26 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.625
+ $Y=1.97 $X2=0.81 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%Q 1 2 3 4 13 15 17 21 24 27 31 33 37 43 44
+ 45 55
c74 37 0 1.5942e-19 $X=8.71 $Y=1.885
r75 55 56 6.0176 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.795 $Y=0.965
+ $X2=8.89 $Y2=0.965
r76 44 45 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.36 $Y=1.295
+ $X2=9.36 $Y2=1.665
r77 44 49 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=1.295
+ $X2=9.36 $Y2=1.13
r78 43 49 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.36 $Y=0.965
+ $X2=9.36 $Y2=1.13
r79 43 56 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=9.36 $Y=0.965
+ $X2=8.89 $Y2=0.965
r80 42 45 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=9.36 $Y=1.8
+ $X2=9.36 $Y2=1.665
r81 40 41 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=8.71 $Y=1.985 $X2=8.71
+ $Y2=2.045
r82 37 40 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=8.71 $Y=1.885 $X2=8.71
+ $Y2=1.985
r83 34 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.875 $Y=1.885
+ $X2=8.71 $Y2=1.885
r84 33 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.245 $Y=1.885
+ $X2=9.36 $Y2=1.8
r85 33 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.245 $Y=1.885
+ $X2=8.875 $Y2=1.885
r86 29 56 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=8.89 $Y=0.8 $X2=8.89
+ $Y2=0.965
r87 29 31 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=8.89 $Y=0.8
+ $X2=8.89 $Y2=0.525
r88 25 41 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.71 $Y=2.13
+ $X2=8.71 $Y2=2.045
r89 25 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.71 $Y=2.13
+ $X2=8.71 $Y2=2.4
r90 24 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.125 $Y=1.045
+ $X2=8.795 $Y2=1.045
r91 19 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.03 $Y=0.96
+ $X2=8.125 $Y2=1.045
r92 19 21 25.3923 $w=1.88e-07 $l=4.35e-07 $layer=LI1_cond $X=8.03 $Y=0.96
+ $X2=8.03 $Y2=0.525
r93 18 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=2.045
+ $X2=7.71 $Y2=2.045
r94 17 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.545 $Y=2.045
+ $X2=8.71 $Y2=2.045
r95 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.545 $Y=2.045
+ $X2=7.875 $Y2=2.045
r96 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.71 $Y=2.13 $X2=7.71
+ $Y2=2.045
r97 13 15 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=7.71 $Y=2.13
+ $X2=7.71 $Y2=2.815
r98 4 40 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=1.84 $X2=8.71 $Y2=1.985
r99 4 27 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=8.525
+ $Y=1.84 $X2=8.71 $Y2=2.4
r100 3 36 400 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.84 $X2=7.71 $Y2=2.125
r101 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.84 $X2=7.71 $Y2=2.815
r102 2 56 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.965
r103 2 31 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.525
r104 1 21 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=7.89
+ $Y=0.37 $X2=8.03 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 44 46
+ 49 50 51 53 70 74 79 85 90 96 98 101 104 108
c119 28 0 1.47145e-19 $X=4.76 $Y=0.515
r120 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r121 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r123 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r124 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r125 94 96 6.66521 $w=5.73e-07 $l=5e-09 $layer=LI1_cond $X=3.12 $Y=0.202
+ $X2=3.125 $Y2=0.202
r126 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r127 92 94 3.32822 $w=5.73e-07 $l=1.6e-07 $layer=LI1_cond $X=2.96 $Y=0.202
+ $X2=3.12 $Y2=0.202
r128 89 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r129 88 92 6.65644 $w=5.73e-07 $l=3.2e-07 $layer=LI1_cond $X=2.64 $Y=0.202
+ $X2=2.96 $Y2=0.202
r130 88 90 13.4257 $w=5.73e-07 $l=3.3e-07 $layer=LI1_cond $X=2.64 $Y=0.202
+ $X2=2.31 $Y2=0.202
r131 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r132 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r133 83 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r134 83 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r135 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r136 80 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.46 $Y2=0
r137 80 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.88 $Y2=0
r138 79 107 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=9.377 $Y2=0
r139 79 82 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=8.88 $Y2=0
r140 78 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r141 78 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r142 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r143 75 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0 $X2=7.6
+ $Y2=0
r144 75 77 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.92 $Y2=0
r145 74 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=8.46 $Y2=0
r146 74 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=7.92 $Y2=0
r147 73 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r148 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r149 70 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r150 70 72 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=5.04 $Y2=0
r151 69 95 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=3.12 $Y2=0
r152 68 96 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=4.56 $Y=0
+ $X2=3.125 $Y2=0
r153 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r154 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r155 64 90 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.31
+ $Y2=0
r156 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r157 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r158 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r159 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r160 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r161 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r162 59 61 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r163 56 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r164 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r165 53 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r166 53 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r167 51 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r168 51 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r169 49 68 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.56
+ $Y2=0
r170 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.76
+ $Y2=0
r171 48 72 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.925 $Y=0
+ $X2=5.04 $Y2=0
r172 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0 $X2=4.76
+ $Y2=0
r173 44 107 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.377 $Y2=0
r174 44 46 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.32 $Y2=0.53
r175 40 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=0.085
+ $X2=8.46 $Y2=0
r176 40 42 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.46 $Y=0.085
+ $X2=8.46 $Y2=0.625
r177 36 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0
r178 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0.525
r179 35 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r180 34 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=0 $X2=7.6
+ $Y2=0
r181 34 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.435 $Y=0
+ $X2=6.775 $Y2=0
r182 30 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r183 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.515
r184 26 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0
r185 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0.515
r186 22 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r187 22 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r188 7 46 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.37 $X2=9.32 $Y2=0.53
r189 6 42 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=8.32
+ $Y=0.37 $X2=8.46 $Y2=0.625
r190 5 38 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=7.455
+ $Y=0.37 $X2=7.6 $Y2=0.525
r191 4 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.47
+ $Y=0.37 $X2=6.61 $Y2=0.515
r192 3 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.62
+ $Y=0.37 $X2=4.76 $Y2=0.515
r193 2 92 91 $w=1.7e-07 $l=7.83167e-07 $layer=licon1_NDIFF $count=2 $X=2.255
+ $Y=0.49 $X2=2.96 $Y2=0.325
r194 1 24 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_4%A_1035_74# 1 2 3 12 14 15 17 19 20 22 24
r45 22 29 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=7.075 $Y=0.77 $X2=7.075
+ $Y2=0.86
r46 22 24 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=7.075 $Y=0.77
+ $X2=7.075 $Y2=0.52
r47 21 27 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6.265 $Y=0.86
+ $X2=6.14 $Y2=0.86
r48 20 29 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=6.945 $Y=0.86
+ $X2=7.075 $Y2=0.86
r49 20 21 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.945 $Y=0.86
+ $X2=6.265 $Y2=0.86
r50 17 27 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.14 $Y=0.77 $X2=6.14
+ $Y2=0.86
r51 17 19 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=6.14 $Y=0.77
+ $X2=6.14 $Y2=0.495
r52 16 19 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=6.14 $Y=0.425 $X2=6.14
+ $Y2=0.495
r53 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.015 $Y=0.34
+ $X2=6.14 $Y2=0.425
r54 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.015 $Y=0.34
+ $X2=5.485 $Y2=0.34
r55 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.32 $Y=0.425
+ $X2=5.485 $Y2=0.34
r56 10 12 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=5.32 $Y=0.425 $X2=5.32
+ $Y2=0.495
r57 3 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.37 $X2=7.04 $Y2=0.86
r58 3 24 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.37 $X2=7.04 $Y2=0.52
r59 2 27 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.37 $X2=6.18 $Y2=0.865
r60 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.37 $X2=6.18 $Y2=0.495
r61 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.175
+ $Y=0.37 $X2=5.32 $Y2=0.495
.ends


* NGSPICE file created from sky130_fd_sc_ms__sedfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_2589_508# a_1510_74# a_2403_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.836e+11p ps=2.66e+06u
M1001 a_575_463# DE VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=3.10925e+12p ps=2.772e+07u
M1002 a_135_74# D a_37_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1003 a_661_113# SCE a_1044_125# VNB nlowvt w=420000u l=150000u
+  ad=5.502e+11p pd=5.14e+06u as=8.82e+10p ps=1.26e+06u
M1004 a_129_464# D a_37_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=3.52e+11p ps=3.66e+06u
M1005 a_1074_455# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 VGND DE a_177_290# VNB nlowvt w=420000u l=150000u
+  ad=2.3264e+12p pd=2.159e+07u as=1.197e+11p ps=1.41e+06u
M1007 a_1044_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_545_87# a_2589_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_177_290# a_129_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1313_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1011 a_1510_74# a_1313_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 Q a_2403_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1013 a_2498_74# a_1313_74# a_2403_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.915e+11p ps=1.93e+06u
M1014 VGND a_545_87# a_2498_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1510_74# a_1313_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1016 a_545_87# a_2403_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1017 Q a_2403_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=4.11e+06u as=0p ps=0u
M1018 a_37_464# a_545_87# a_497_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 a_661_113# a_631_87# a_37_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1313_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1021 a_1943_53# a_1756_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.184e+11p pd=2.2e+06u as=0p ps=0u
M1022 a_2403_74# a_1510_74# a_2331_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1023 a_37_464# a_545_87# a_575_463# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR SCE a_631_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1025 VGND a_1943_53# a_1858_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1026 VGND DE a_135_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_661_113# SCE a_37_464# VPB pshort w=640000u l=180000u
+  ad=4.452e+11p pd=4.97e+06u as=0p ps=0u
M1028 a_661_113# a_631_87# a_1074_455# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR DE a_177_290# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1030 a_545_87# a_2403_74# VPWR VPB pshort w=640000u l=180000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1031 a_1858_79# a_1510_74# a_1756_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.6695e+11p ps=1.74e+06u
M1032 VPWR a_2403_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1756_97# a_1510_74# a_661_113# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1034 a_497_113# a_177_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2403_74# a_1313_74# a_2295_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.8e+11p ps=3.56e+06u
M1036 VPWR a_1943_53# a_1902_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1037 VGND a_2403_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1756_97# a_1313_74# a_661_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Q a_2403_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_2403_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Q a_2403_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1902_508# a_1313_74# a_1756_97# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND SCE a_631_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1044 a_2295_392# a_1943_53# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPWR a_2403_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1943_53# a_1756_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1047 a_2331_74# a_1943_53# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__o2bb2a_1.spice
* Created: Wed Sep  2 12:24:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2bb2a_1.pex.spice"
.subckt sky130_fd_sc_ms__o2bb2a_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_83_260#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.202642 AS=0.2109 PD=1.36739 PS=2.05 NRD=19.044 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 A_253_94# N_A1_N_M1003_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.175258 PD=0.88 PS=1.18261 NRD=12.18 NRS=26.244 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1004 N_A_236_384#_M1004_d N_A2_N_M1004_g A_253_94# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.3
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_588_74#_M1006_d N_A_236_384#_M1006_g N_A_83_260#_M1006_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_B2_M1011_g N_A_588_74#_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.0896 PD=1.02 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1009 N_A_588_74#_M1009_d N_B1_M1009_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1216 PD=1.85 PS=1.02 NRD=0 NRS=5.616 M=1 R=4.26667 SA=75001.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A_83_260#_M1002_g N_X_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.243543 AS=0.3136 PD=1.74286 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1000 N_A_236_384#_M1000_d N_A1_N_M1000_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1365 AS=0.182657 PD=1.165 PS=1.30714 NRD=0 NRS=19.1484 M=1
+ R=4.66667 SA=90000.8 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1010 N_VPWR_M1010_d N_A2_N_M1010_g N_A_236_384#_M1000_d VPB PSHORT L=0.18
+ W=0.84 AD=0.4641 AS=0.1365 PD=1.945 PS=1.165 NRD=0 NRS=11.7215 M=1 R=4.66667
+ SA=90001.3 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1007 N_A_83_260#_M1007_d N_A_236_384#_M1007_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.84 AD=0.144809 AS=0.4641 PD=1.21435 PS=1.945 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90002.6 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1005 A_696_384# N_B2_M1005_g N_A_83_260#_M1007_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.172391 PD=1.24 PS=1.44565 NRD=12.7853 NRS=0.9653 M=1 R=5.55556 SA=90002.6
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g A_696_384# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90003 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__o2bb2a_1.pxi.spice"
*
.ends
*
*

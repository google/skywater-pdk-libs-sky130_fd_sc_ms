* File: sky130_fd_sc_ms__clkbuf_4.pxi.spice
* Created: Fri Aug 28 17:17:40 2020
* 
x_PM_SKY130_FD_SC_MS__CLKBUF_4%A_83_270# N_A_83_270#_M1004_d N_A_83_270#_M1005_d
+ N_A_83_270#_M1001_g N_A_83_270#_M1000_g N_A_83_270#_M1007_g
+ N_A_83_270#_M1002_g N_A_83_270#_M1008_g N_A_83_270#_M1003_g
+ N_A_83_270#_M1009_g N_A_83_270#_M1006_g N_A_83_270#_c_67_n N_A_83_270#_c_58_n
+ N_A_83_270#_c_69_n N_A_83_270#_c_59_n N_A_83_270#_c_70_n N_A_83_270#_c_60_n
+ N_A_83_270#_c_61_n N_A_83_270#_c_62_n PM_SKY130_FD_SC_MS__CLKBUF_4%A_83_270#
x_PM_SKY130_FD_SC_MS__CLKBUF_4%A N_A_M1005_g N_A_M1004_g A N_A_c_165_n
+ N_A_c_166_n PM_SKY130_FD_SC_MS__CLKBUF_4%A
x_PM_SKY130_FD_SC_MS__CLKBUF_4%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1006_s
+ N_VPWR_c_200_n N_VPWR_c_201_n N_VPWR_c_202_n N_VPWR_c_203_n N_VPWR_c_204_n
+ N_VPWR_c_205_n VPWR N_VPWR_c_206_n N_VPWR_c_207_n N_VPWR_c_199_n
+ N_VPWR_c_209_n PM_SKY130_FD_SC_MS__CLKBUF_4%VPWR
x_PM_SKY130_FD_SC_MS__CLKBUF_4%X N_X_M1000_s N_X_M1008_s N_X_M1001_d N_X_M1003_d
+ N_X_c_241_n N_X_c_247_n N_X_c_256_n N_X_c_242_n N_X_c_243_n N_X_c_268_n
+ N_X_c_248_n N_X_c_275_n X X X PM_SKY130_FD_SC_MS__CLKBUF_4%X
x_PM_SKY130_FD_SC_MS__CLKBUF_4%VGND N_VGND_M1000_d N_VGND_M1007_d N_VGND_M1009_d
+ N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n
+ N_VGND_c_310_n VGND N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n
+ N_VGND_c_314_n PM_SKY130_FD_SC_MS__CLKBUF_4%VGND
cc_1 VNB N_A_83_270#_M1000_g 0.0542361f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_2 VNB N_A_83_270#_M1007_g 0.0376483f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.58
cc_3 VNB N_A_83_270#_M1008_g 0.0387572f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.58
cc_4 VNB N_A_83_270#_M1009_g 0.0431021f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.58
cc_5 VNB N_A_83_270#_c_58_n 0.00535841f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.665
cc_6 VNB N_A_83_270#_c_59_n 0.0376158f $X=-0.19 $Y=-0.245 $X2=2.71 $Y2=1.58
cc_7 VNB N_A_83_270#_c_60_n 0.00986226f $X=-0.19 $Y=-0.245 $X2=2.605 $Y2=1.665
cc_8 VNB N_A_83_270#_c_61_n 0.0197872f $X=-0.19 $Y=-0.245 $X2=2.71 $Y2=0.645
cc_9 VNB N_A_83_270#_c_62_n 0.0841865f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.515
cc_10 VNB N_A_M1005_g 0.0155743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_M1004_g 0.0337688f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.68
cc_12 VNB N_A_c_165_n 0.0326721f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_13 VNB N_A_c_166_n 0.0049741f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_14 VNB N_VPWR_c_199_n 0.123877f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.515
cc_15 VNB N_X_c_241_n 0.00143018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_X_c_242_n 0.0126859f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_17 VNB N_X_c_243_n 0.00543306f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.58
cc_18 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.68
cc_19 VNB X 0.00447861f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_20 VNB N_VGND_c_305_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_306_n 0.0388367f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_22 VNB N_VGND_c_307_n 0.00964419f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.58
cc_23 VNB N_VGND_c_308_n 0.0170065f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_24 VNB N_VGND_c_309_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.35
cc_25 VNB N_VGND_c_310_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.58
cc_26 VNB N_VGND_c_311_n 0.0189618f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.35
cc_27 VNB N_VGND_c_312_n 0.0199267f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_28 VNB N_VGND_c_313_n 0.185299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_314_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.665
cc_30 VPB N_A_83_270#_M1001_g 0.0257336f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_31 VPB N_A_83_270#_M1002_g 0.020395f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_32 VPB N_A_83_270#_M1003_g 0.020748f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_33 VPB N_A_83_270#_M1006_g 0.0216563f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_34 VPB N_A_83_270#_c_67_n 0.00427588f $X=-0.19 $Y=1.66 $X2=1.685 $Y2=1.55
cc_35 VPB N_A_83_270#_c_58_n 0.00474727f $X=-0.19 $Y=1.66 $X2=2.415 $Y2=1.665
cc_36 VPB N_A_83_270#_c_69_n 0.0531345f $X=-0.19 $Y=1.66 $X2=2.58 $Y2=1.985
cc_37 VPB N_A_83_270#_c_70_n 7.44389e-19 $X=-0.19 $Y=1.66 $X2=1.885 $Y2=1.55
cc_38 VPB N_A_83_270#_c_60_n 0.00423137f $X=-0.19 $Y=1.66 $X2=2.605 $Y2=1.665
cc_39 VPB N_A_83_270#_c_62_n 0.0121059f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.515
cc_40 VPB N_A_M1005_g 0.0287168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_200_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_201_n 0.0637841f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.58
cc_43 VPB N_VPWR_c_202_n 0.0049754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_203_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_204_n 0.0182909f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.68
cc_46 VPB N_VPWR_c_205_n 0.00458862f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_47 VPB N_VPWR_c_206_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.68
cc_48 VPB N_VPWR_c_207_n 0.0193845f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.515
cc_49 VPB N_VPWR_c_199_n 0.0593374f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.515
cc_50 VPB N_VPWR_c_209_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.58 $Y2=1.985
cc_51 VPB N_X_c_241_n 0.00127965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_X_c_247_n 0.00202377f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.58
cc_53 VPB N_X_c_248_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_54 N_A_83_270#_c_58_n N_A_M1005_g 0.0131783f $X=2.415 $Y=1.665 $X2=0 $Y2=0
cc_55 N_A_83_270#_c_69_n N_A_M1005_g 0.0189171f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_56 N_A_83_270#_c_59_n N_A_M1005_g 0.00584384f $X=2.71 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_83_270#_c_70_n N_A_M1005_g 9.26486e-19 $X=1.885 $Y=1.55 $X2=0 $Y2=0
cc_58 N_A_83_270#_c_60_n N_A_M1005_g 0.00446031f $X=2.605 $Y=1.665 $X2=0 $Y2=0
cc_59 N_A_83_270#_c_62_n N_A_M1005_g 0.0231615f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_60 N_A_83_270#_M1009_g N_A_M1004_g 0.0174474f $X=1.84 $Y=0.58 $X2=0 $Y2=0
cc_61 N_A_83_270#_c_59_n N_A_M1004_g 0.00912792f $X=2.71 $Y=1.58 $X2=0 $Y2=0
cc_62 N_A_83_270#_c_61_n N_A_M1004_g 0.00458743f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_63 N_A_83_270#_M1009_g N_A_c_165_n 0.0133899f $X=1.84 $Y=0.58 $X2=0 $Y2=0
cc_64 N_A_83_270#_c_58_n N_A_c_165_n 0.00246626f $X=2.415 $Y=1.665 $X2=0 $Y2=0
cc_65 N_A_83_270#_c_59_n N_A_c_165_n 0.00769124f $X=2.71 $Y=1.58 $X2=0 $Y2=0
cc_66 N_A_83_270#_c_60_n N_A_c_165_n 0.00156619f $X=2.605 $Y=1.665 $X2=0 $Y2=0
cc_67 N_A_83_270#_c_61_n N_A_c_165_n 0.00130341f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_68 N_A_83_270#_c_62_n N_A_c_165_n 0.0039541f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A_83_270#_M1009_g N_A_c_166_n 0.00552999f $X=1.84 $Y=0.58 $X2=0 $Y2=0
cc_70 N_A_83_270#_c_58_n N_A_c_166_n 0.0268738f $X=2.415 $Y=1.665 $X2=0 $Y2=0
cc_71 N_A_83_270#_c_59_n N_A_c_166_n 0.0251396f $X=2.71 $Y=1.58 $X2=0 $Y2=0
cc_72 N_A_83_270#_c_70_n N_A_c_166_n 0.0049623f $X=1.885 $Y=1.55 $X2=0 $Y2=0
cc_73 N_A_83_270#_c_60_n N_A_c_166_n 0.00323807f $X=2.605 $Y=1.665 $X2=0 $Y2=0
cc_74 N_A_83_270#_c_61_n N_A_c_166_n 0.00185729f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_75 N_A_83_270#_c_62_n N_A_c_166_n 4.41551e-19 $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A_83_270#_M1001_g N_VPWR_c_201_n 0.00515532f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_83_270#_M1001_g N_VPWR_c_202_n 5.71655e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_78 N_A_83_270#_M1002_g N_VPWR_c_202_n 0.0129f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_83_270#_M1003_g N_VPWR_c_202_n 0.002979f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_83_270#_M1006_g N_VPWR_c_203_n 0.00306788f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A_83_270#_c_58_n N_VPWR_c_203_n 0.018622f $X=2.415 $Y=1.665 $X2=0 $Y2=0
cc_82 N_A_83_270#_c_69_n N_VPWR_c_203_n 0.0413997f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_83_270#_M1001_g N_VPWR_c_204_n 0.0048691f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_83_270#_M1002_g N_VPWR_c_204_n 0.00460063f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_83_270#_M1003_g N_VPWR_c_206_n 0.005209f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_83_270#_M1006_g N_VPWR_c_206_n 0.005209f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_83_270#_c_69_n N_VPWR_c_207_n 0.01678f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_83_270#_M1001_g N_VPWR_c_199_n 0.00875947f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A_83_270#_M1002_g N_VPWR_c_199_n 0.00908554f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_83_270#_M1003_g N_VPWR_c_199_n 0.00982266f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_83_270#_M1006_g N_VPWR_c_199_n 0.00982832f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_83_270#_c_69_n N_VPWR_c_199_n 0.0138209f $X=2.58 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_83_270#_M1001_g N_X_c_241_n 0.00882232f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A_83_270#_M1000_g N_X_c_241_n 0.010296f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_95 N_A_83_270#_M1007_g N_X_c_241_n 0.00313669f $X=0.94 $Y=0.58 $X2=0 $Y2=0
cc_96 N_A_83_270#_M1002_g N_X_c_241_n 0.00292405f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_83_270#_c_67_n N_X_c_241_n 0.0305337f $X=1.685 $Y=1.55 $X2=0 $Y2=0
cc_98 N_A_83_270#_c_62_n N_X_c_241_n 0.0234504f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A_83_270#_M1001_g N_X_c_247_n 0.0130348f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_83_270#_M1002_g N_X_c_256_n 0.0145311f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_83_270#_M1003_g N_X_c_256_n 0.012931f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_83_270#_c_67_n N_X_c_256_n 0.0404153f $X=1.685 $Y=1.55 $X2=0 $Y2=0
cc_103 N_A_83_270#_c_62_n N_X_c_256_n 5.25301e-19 $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A_83_270#_M1007_g N_X_c_242_n 0.0113002f $X=0.94 $Y=0.58 $X2=0 $Y2=0
cc_105 N_A_83_270#_M1008_g N_X_c_242_n 0.0140197f $X=1.37 $Y=0.58 $X2=0 $Y2=0
cc_106 N_A_83_270#_M1009_g N_X_c_242_n 0.00425798f $X=1.84 $Y=0.58 $X2=0 $Y2=0
cc_107 N_A_83_270#_c_67_n N_X_c_242_n 0.0595809f $X=1.685 $Y=1.55 $X2=0 $Y2=0
cc_108 N_A_83_270#_c_62_n N_X_c_242_n 0.00571564f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A_83_270#_M1007_g N_X_c_243_n 6.3694e-19 $X=0.94 $Y=0.58 $X2=0 $Y2=0
cc_110 N_A_83_270#_M1008_g N_X_c_243_n 0.0106797f $X=1.37 $Y=0.58 $X2=0 $Y2=0
cc_111 N_A_83_270#_M1009_g N_X_c_243_n 0.00541161f $X=1.84 $Y=0.58 $X2=0 $Y2=0
cc_112 N_A_83_270#_M1003_g N_X_c_268_n 8.84614e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_83_270#_M1006_g N_X_c_268_n 0.00246348f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_83_270#_c_67_n N_X_c_268_n 0.0233528f $X=1.685 $Y=1.55 $X2=0 $Y2=0
cc_115 N_A_83_270#_c_62_n N_X_c_268_n 5.94712e-19 $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A_83_270#_M1002_g N_X_c_248_n 6.83718e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_83_270#_M1003_g N_X_c_248_n 0.0124928f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_83_270#_M1006_g N_X_c_248_n 0.0111507f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_83_270#_M1001_g N_X_c_275_n 0.00235661f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_83_270#_c_62_n N_X_c_275_n 0.00288553f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A_83_270#_M1000_g X 0.0154573f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_122 N_A_83_270#_M1007_g X 0.0108162f $X=0.94 $Y=0.58 $X2=0 $Y2=0
cc_123 N_A_83_270#_M1008_g X 6.3694e-19 $X=1.37 $Y=0.58 $X2=0 $Y2=0
cc_124 N_A_83_270#_M1000_g X 0.0116878f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_125 N_A_83_270#_M1007_g X 0.00318666f $X=0.94 $Y=0.58 $X2=0 $Y2=0
cc_126 N_A_83_270#_c_67_n X 0.00106536f $X=1.685 $Y=1.55 $X2=0 $Y2=0
cc_127 N_A_83_270#_c_62_n X 0.0030119f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_83_270#_M1000_g N_VGND_c_306_n 0.00589946f $X=0.51 $Y=0.58 $X2=0
+ $Y2=0
cc_129 N_A_83_270#_M1007_g N_VGND_c_307_n 0.00301336f $X=0.94 $Y=0.58 $X2=0
+ $Y2=0
cc_130 N_A_83_270#_M1008_g N_VGND_c_307_n 0.00301336f $X=1.37 $Y=0.58 $X2=0
+ $Y2=0
cc_131 N_A_83_270#_M1009_g N_VGND_c_308_n 0.00386565f $X=1.84 $Y=0.58 $X2=0
+ $Y2=0
cc_132 N_A_83_270#_c_61_n N_VGND_c_308_n 0.0133724f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_133 N_A_83_270#_c_62_n N_VGND_c_308_n 7.88991e-19 $X=1.855 $Y=1.515 $X2=0
+ $Y2=0
cc_134 N_A_83_270#_M1000_g N_VGND_c_309_n 0.00434272f $X=0.51 $Y=0.58 $X2=0
+ $Y2=0
cc_135 N_A_83_270#_M1007_g N_VGND_c_309_n 0.00434272f $X=0.94 $Y=0.58 $X2=0
+ $Y2=0
cc_136 N_A_83_270#_M1008_g N_VGND_c_311_n 0.00434272f $X=1.37 $Y=0.58 $X2=0
+ $Y2=0
cc_137 N_A_83_270#_M1009_g N_VGND_c_311_n 0.00461464f $X=1.84 $Y=0.58 $X2=0
+ $Y2=0
cc_138 N_A_83_270#_c_61_n N_VGND_c_312_n 0.00934776f $X=2.71 $Y=0.645 $X2=0
+ $Y2=0
cc_139 N_A_83_270#_M1000_g N_VGND_c_313_n 0.00823992f $X=0.51 $Y=0.58 $X2=0
+ $Y2=0
cc_140 N_A_83_270#_M1007_g N_VGND_c_313_n 0.00820284f $X=0.94 $Y=0.58 $X2=0
+ $Y2=0
cc_141 N_A_83_270#_M1008_g N_VGND_c_313_n 0.00820671f $X=1.37 $Y=0.58 $X2=0
+ $Y2=0
cc_142 N_A_83_270#_M1009_g N_VGND_c_313_n 0.00908551f $X=1.84 $Y=0.58 $X2=0
+ $Y2=0
cc_143 N_A_83_270#_c_61_n N_VGND_c_313_n 0.0122187f $X=2.71 $Y=0.645 $X2=0 $Y2=0
cc_144 N_A_M1005_g N_VPWR_c_203_n 0.00318542f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_M1005_g N_VPWR_c_207_n 0.005209f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_M1005_g N_VPWR_c_199_n 0.0098597f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_c_166_n N_X_c_242_n 0.00411964f $X=2.32 $Y=1.245 $X2=0 $Y2=0
cc_148 N_A_M1004_g N_VGND_c_308_n 0.00622707f $X=2.37 $Y=0.58 $X2=0 $Y2=0
cc_149 N_A_c_165_n N_VGND_c_308_n 0.00207081f $X=2.32 $Y=1.245 $X2=0 $Y2=0
cc_150 N_A_c_166_n N_VGND_c_308_n 0.0120196f $X=2.32 $Y=1.245 $X2=0 $Y2=0
cc_151 N_A_M1004_g N_VGND_c_312_n 0.00435951f $X=2.37 $Y=0.58 $X2=0 $Y2=0
cc_152 N_A_M1004_g N_VGND_c_313_n 0.0082442f $X=2.37 $Y=0.58 $X2=0 $Y2=0
cc_153 N_VPWR_c_201_n N_X_c_241_n 0.0045068f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_154 N_VPWR_c_201_n N_X_c_247_n 0.0332863f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_155 N_VPWR_c_202_n N_X_c_247_n 0.0234203f $X=1.18 $Y=2.425 $X2=0 $Y2=0
cc_156 N_VPWR_c_204_n N_X_c_247_n 0.0122283f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_c_199_n N_X_c_247_n 0.00998289f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_158 N_VPWR_M1002_s N_X_c_256_n 0.0031345f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_159 N_VPWR_c_202_n N_X_c_256_n 0.0148589f $X=1.18 $Y=2.425 $X2=0 $Y2=0
cc_160 N_VPWR_c_202_n N_X_c_248_n 0.0243967f $X=1.18 $Y=2.425 $X2=0 $Y2=0
cc_161 N_VPWR_c_203_n N_X_c_248_n 0.0299644f $X=2.08 $Y=2.085 $X2=0 $Y2=0
cc_162 N_VPWR_c_206_n N_X_c_248_n 0.0144623f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_c_199_n N_X_c_248_n 0.0118344f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_164 X N_VGND_c_306_n 0.0179429f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_165 N_X_c_242_n N_VGND_c_307_n 0.0141893f $X=1.42 $Y=1.065 $X2=0 $Y2=0
cc_166 N_X_c_243_n N_VGND_c_307_n 0.0178601f $X=1.585 $Y=0.58 $X2=0 $Y2=0
cc_167 X N_VGND_c_307_n 0.0178601f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_168 N_X_c_243_n N_VGND_c_308_n 0.00316191f $X=1.585 $Y=0.58 $X2=0 $Y2=0
cc_169 X N_VGND_c_309_n 0.0144922f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_170 N_X_c_243_n N_VGND_c_311_n 0.0145639f $X=1.585 $Y=0.58 $X2=0 $Y2=0
cc_171 N_X_c_243_n N_VGND_c_313_n 0.0119984f $X=1.585 $Y=0.58 $X2=0 $Y2=0
cc_172 X N_VGND_c_313_n 0.0118826f $X=0.635 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o2111a_4.spice
* Created: Fri Aug 28 17:51:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2111a_4.pex.spice"
.subckt sky130_fd_sc_ms__o2111a_4  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1010 N_A_27_392#_M1010_d N_D1_M1010_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2146 PD=1.02 PS=2.06 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_392#_M1010_d N_D1_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_287_74#_M1001_d N_C1_M1001_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_287_74#_M1001_d N_C1_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.24285 PD=1.02 PS=2.49 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_287_74#_M1004_d N_B1_M1004_g N_A_477_198#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.21835 PD=1.02 PS=2.21 NRD=0 NRS=6.48 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1026 N_A_287_74#_M1004_d N_B1_M1026_g N_A_477_198#_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_A_477_198#_M1026_s N_A2_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1258 PD=1.02 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1027 N_A_477_198#_M1027_d N_A2_M1027_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2183 AS=0.1258 PD=2.07 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_477_198#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1014 N_A_477_198#_M1005_d N_A1_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1006_d N_A_27_392#_M1006_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1006_d N_A_27_392#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_27_392#_M1012_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1019 N_X_M1012_d N_A_27_392#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D1_M1000_g N_A_27_392#_M1000_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90003.8 A=0.1512 P=2.04 MULT=1
MM1023 N_VPWR_M1000_d N_D1_M1023_g N_A_27_392#_M1023_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.1134 PD=1.21 PS=1.11 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.7
+ SB=90003.3 A=0.1512 P=2.04 MULT=1
MM1024 N_A_27_392#_M1023_s N_C1_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1344 PD=1.11 PS=1.16 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90001.2
+ SB=90002.8 A=0.1512 P=2.04 MULT=1
MM1025 N_A_27_392#_M1025_d N_C1_M1025_g N_VPWR_M1024_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1848 AS=0.1344 PD=1.28 PS=1.16 NRD=18.7544 NRS=0 M=1 R=4.66667 SA=90001.7
+ SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1013 N_VPWR_M1013_d N_B1_M1013_g N_A_27_392#_M1025_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1848 PD=1.11 PS=1.28 NRD=0 NRS=18.7544 M=1 R=4.66667 SA=90002.3
+ SB=90001.7 A=0.1512 P=2.04 MULT=1
MM1020 N_VPWR_M1013_d N_B1_M1020_g N_A_27_392#_M1020_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.179413 PD=1.11 PS=1.28283 NRD=0 NRS=19.1484 M=1 R=4.66667
+ SA=90002.8 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1002 N_A_27_392#_M1020_s N_A2_M1002_g N_A_750_392#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.213587 AS=0.16 PD=1.52717 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90002.8 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_392#_M1003_d N_A2_M1003_g N_A_750_392#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.16 PD=2.56 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90003.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1018 N_A_750_392#_M1018_d N_A1_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.33 PD=1.27 PS=2.66 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.2
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1022 N_A_750_392#_M1018_d N_A1_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.181604 PD=1.27 PS=1.39151 NRD=0 NRS=15.7403 M=1 R=5.55556
+ SA=90000.7 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1022_s N_A_27_392#_M1015_g N_X_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.203396 AS=0.1792 PD=1.55849 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.1 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_A_27_392#_M1016_g N_X_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1016_d N_A_27_392#_M1017_g N_X_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_27_392#_M1021_g N_X_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_78 VNB 0 5.23076e-20 $X=0 $Y=0
c_148 VPB 0 1.58594e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__o2111a_4.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__o21a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.445000 2.275000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.445000 1.505000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.494400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.515000 3.235000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815000 1.720000 5.635000 1.780000 ;
        RECT 3.815000 1.780000 5.145000 1.890000 ;
        RECT 3.815000 1.890000 4.145000 2.980000 ;
        RECT 3.990000 0.330000 4.240000 0.835000 ;
        RECT 3.990000 0.835000 5.135000 1.005000 ;
        RECT 4.815000 1.890000 5.145000 2.980000 ;
        RECT 4.965000 0.350000 5.135000 0.835000 ;
        RECT 4.965000 1.005000 5.135000 1.550000 ;
        RECT 4.965000 1.550000 5.635000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.605000 0.445000 1.105000 ;
      RECT 0.115000  1.105000 2.390000 1.275000 ;
      RECT 0.115000  1.275000 0.445000 1.285000 ;
      RECT 0.115000  1.915000 0.445000 3.245000 ;
      RECT 0.615000  0.085000 0.950000 0.935000 ;
      RECT 0.615000  1.950000 0.865000 2.905000 ;
      RECT 0.615000  2.905000 1.895000 3.075000 ;
      RECT 1.065000  1.950000 3.575000 2.120000 ;
      RECT 1.065000  2.120000 1.395000 2.735000 ;
      RECT 1.130000  0.605000 1.380000 1.105000 ;
      RECT 1.560000  0.085000 1.890000 0.935000 ;
      RECT 1.565000  2.290000 1.895000 2.905000 ;
      RECT 2.060000  0.265000 3.330000 0.435000 ;
      RECT 2.060000  0.435000 2.390000 1.105000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.565000  2.120000 2.895000 2.795000 ;
      RECT 2.570000  0.605000 2.820000 1.175000 ;
      RECT 2.570000  1.175000 4.795000 1.345000 ;
      RECT 3.000000  0.435000 3.330000 1.005000 ;
      RECT 3.135000  2.300000 3.615000 3.245000 ;
      RECT 3.405000  1.345000 4.795000 1.550000 ;
      RECT 3.405000  1.550000 3.575000 1.950000 ;
      RECT 3.560000  0.085000 3.810000 1.005000 ;
      RECT 4.315000  2.060000 4.645000 3.245000 ;
      RECT 4.420000  0.085000 4.785000 0.665000 ;
      RECT 5.315000  0.085000 5.645000 1.130000 ;
      RECT 5.315000  1.950000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__o21a_4
END LIBRARY

* File: sky130_fd_sc_ms__or4_4.spice
* Created: Fri Aug 28 18:09:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4_4.pex.spice"
.subckt sky130_fd_sc_ms__or4_4  VNB VPB B A C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_83_264#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_83_264#_M1007_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75004.6 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1007_d N_A_83_264#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.22385 PD=1.09 PS=1.345 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_83_264#_M1012_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1835 AS=0.22385 PD=1.27 PS=1.345 NRD=16.212 NRS=41.34 M=1 R=4.93333
+ SA=75002 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1004 N_A_83_264#_M1004_d N_B_M1004_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1835 PD=1.02 PS=1.27 NRD=0 NRS=16.212 M=1 R=4.93333 SA=75002.6
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_A_83_264#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.5035 AS=0.1036 PD=2.07 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1015 N_A_83_264#_M1015_d N_C_M1015_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.5035 PD=1.09 PS=2.07 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75004.4
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_D_M1009_g N_A_83_264#_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.3445 AS=0.1295 PD=3.08 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.9
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_A_83_264#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1005_d N_A_83_264#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1008_d N_A_83_264#_M1008_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1008_d N_A_83_264#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1014 N_A_591_392#_M1014_d N_B_M1014_g N_A_499_392#_M1014_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_591_392#_M1014_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1016_d N_A_M1017_g N_A_591_392#_M1017_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1018 N_A_591_392#_M1017_s N_B_M1018_g N_A_499_392#_M1018_s VPB PSHORT L=0.18
+ W=1 AD=0.145 AS=0.16 PD=1.29 PS=1.32 NRD=0.9653 NRS=8.8453 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1003 N_A_499_392#_M1018_s N_C_M1003_g N_A_965_392#_M1003_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_83_264#_M1000_d N_D_M1000_g N_A_965_392#_M1003_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1002 N_A_83_264#_M1000_d N_D_M1002_g N_A_965_392#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90003
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1019 N_A_499_392#_M1019_d N_C_M1019_g N_A_965_392#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.33 AS=0.135 PD=2.66 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90003.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ms__or4_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfxtp_1.spice
* Created: Fri Aug 28 17:25:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfxtp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfxtp_1  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_CLK_M1022_g N_A_27_74#_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1739 AS=0.2109 PD=1.21 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1002 N_A_209_368#_M1002_d N_A_27_74#_M1002_g N_VGND_M1022_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2553 AS=0.1739 PD=2.17 PS=1.21 NRD=9.72 NRS=30.804 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_A_457_503#_M1007_d N_D_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.155625 AS=0.23015 PD=1.215 PS=2.1 NRD=90.144 NRS=140.844 M=1 R=2.8
+ SA=75000.3 SB=75003 A=0.063 P=1.14 MULT=1
MM1017 N_A_564_463#_M1017_d N_A_27_74#_M1017_g N_A_457_503#_M1007_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.07875 AS=0.155625 PD=0.865 PS=1.215 NRD=1.428 NRS=90.144
+ M=1 R=2.8 SA=75000.9 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1016 A_731_101# N_A_209_368#_M1016_g N_A_564_463#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.07875 PD=0.63 PS=0.865 NRD=14.28 NRS=11.424 M=1 R=2.8
+ SA=75001.1 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_713_458#_M1014_g A_731_101# VNB NLOWVT L=0.15 W=0.42
+ AD=0.142713 AS=0.0441 PD=1.07814 PS=0.63 NRD=81.36 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_713_458#_M1004_d N_A_564_463#_M1004_g N_VGND_M1014_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.109062 AS=0.186887 PD=1.025 PS=1.41186 NRD=17.448
+ NRS=38.172 M=1 R=3.66667 SA=75001.7 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1006 N_A_1014_424#_M1006_d N_A_209_368#_M1006_g N_A_713_458#_M1004_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.133928 AS=0.109062 PD=1.17371 PS=1.025 NRD=21.816
+ NRS=0 M=1 R=3.66667 SA=75002.1 SB=75001 A=0.0825 P=1.4 MULT=1
MM1001 A_1168_124# N_A_27_74#_M1001_g N_A_1014_424#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.05565 AS=0.102272 PD=0.685 PS=0.896289 NRD=22.14 NRS=30 M=1 R=2.8
+ SA=75002.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1210_314#_M1021_g A_1168_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.05565 PD=1.41 PS=0.685 NRD=0 NRS=22.14 M=1 R=2.8 SA=75003.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_1014_424#_M1008_g N_A_1210_314#_M1008_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.101153 AS=0.15675 PD=0.925194 PS=1.67 NRD=6.54 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1013 N_Q_M1013_d N_A_1210_314#_M1013_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.136097 PD=2.05 PS=1.24481 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_CLK_M1009_g N_A_27_74#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_A_209_368#_M1010_d N_A_27_74#_M1010_g N_VPWR_M1009_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1020 N_A_457_503#_M1020_d N_D_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=0.42
+ AD=0.09205 AS=0.2909 PD=0.975 PS=2.38 NRD=39.8531 NRS=299.066 M=1 R=2.33333
+ SA=90000.4 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1012 N_A_564_463#_M1012_d N_A_209_368#_M1012_g N_A_457_503#_M1020_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.09205 AS=0.09205 PD=0.975 PS=0.975 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.6 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1015 A_671_503# N_A_27_74#_M1015_g N_A_564_463#_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.09205 PD=0.63 PS=0.975 NRD=23.443 NRS=39.8531 M=1
+ R=2.33333 SA=90000.9 SB=90003 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_713_458#_M1011_g A_671_503# VPB PSHORT L=0.18 W=0.42
+ AD=0.120275 AS=0.0441 PD=1.01 PS=0.63 NRD=108.508 NRS=23.443 M=1 R=2.33333
+ SA=90001.2 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1018 N_A_713_458#_M1018_d N_A_564_463#_M1018_g N_VPWR_M1011_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2205 AS=0.24055 PD=1.365 PS=2.02 NRD=1.1623 NRS=54.2538 M=1
+ R=4.66667 SA=90001 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1003 N_A_1014_424#_M1003_d N_A_27_74#_M1003_g N_A_713_458#_M1018_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1778 AS=0.2205 PD=1.59333 PS=1.365 NRD=0 NRS=56.2829 M=1
+ R=4.66667 SA=90001.7 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1005 A_1121_508# N_A_209_368#_M1005_g N_A_1014_424#_M1003_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09345 AS=0.0889 PD=0.865 PS=0.796667 NRD=78.5636 NRS=39.8531 M=1
+ R=2.33333 SA=90003 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1023 N_VPWR_M1023_d N_A_1210_314#_M1023_g A_1121_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.09345 PD=1.4 PS=0.865 NRD=0 NRS=78.5636 M=1 R=2.33333
+ SA=90003.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_1014_424#_M1000_g N_A_1210_314#_M1000_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.2352 PD=1.23857 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1019 N_Q_M1019_d N_A_1210_314#_M1019_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.196 PD=2.8 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__dfxtp_1.pxi.spice"
*
.ends
*
*

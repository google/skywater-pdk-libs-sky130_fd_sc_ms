* File: sky130_fd_sc_ms__xor2_1.pxi.spice
* Created: Fri Aug 28 18:18:50 2020
* 
x_PM_SKY130_FD_SC_MS__XOR2_1%B N_B_c_70_n N_B_M1001_g N_B_M1002_g N_B_M1005_g
+ N_B_M1006_g N_B_c_66_n B N_B_c_67_n N_B_c_68_n N_B_c_69_n
+ PM_SKY130_FD_SC_MS__XOR2_1%B
x_PM_SKY130_FD_SC_MS__XOR2_1%A N_A_c_133_n N_A_M1000_g N_A_M1008_g N_A_c_135_n
+ N_A_c_136_n N_A_c_137_n N_A_M1003_g N_A_M1004_g N_A_c_140_n A N_A_c_141_n
+ PM_SKY130_FD_SC_MS__XOR2_1%A
x_PM_SKY130_FD_SC_MS__XOR2_1%A_194_125# N_A_194_125#_M1008_d
+ N_A_194_125#_M1001_d N_A_194_125#_M1009_g N_A_194_125#_M1007_g
+ N_A_194_125#_c_191_n N_A_194_125#_c_197_n N_A_194_125#_c_232_n
+ N_A_194_125#_c_208_n N_A_194_125#_c_198_n N_A_194_125#_c_192_n
+ N_A_194_125#_c_200_n N_A_194_125#_c_193_n N_A_194_125#_c_194_n
+ PM_SKY130_FD_SC_MS__XOR2_1%A_194_125#
x_PM_SKY130_FD_SC_MS__XOR2_1%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_277_n
+ N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n VPWR N_VPWR_c_281_n
+ N_VPWR_c_282_n N_VPWR_c_276_n N_VPWR_c_284_n PM_SKY130_FD_SC_MS__XOR2_1%VPWR
x_PM_SKY130_FD_SC_MS__XOR2_1%A_355_368# N_A_355_368#_M1003_s
+ N_A_355_368#_M1006_d N_A_355_368#_c_322_n N_A_355_368#_c_320_n
+ N_A_355_368#_c_321_n PM_SKY130_FD_SC_MS__XOR2_1%A_355_368#
x_PM_SKY130_FD_SC_MS__XOR2_1%X N_X_M1005_d N_X_M1007_d N_X_c_343_n N_X_c_346_n
+ N_X_c_347_n N_X_c_344_n X X N_X_c_350_n X PM_SKY130_FD_SC_MS__XOR2_1%X
x_PM_SKY130_FD_SC_MS__XOR2_1%VGND N_VGND_M1008_s N_VGND_M1002_d N_VGND_M1009_d
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n
+ N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n VGND
+ N_VGND_c_388_n PM_SKY130_FD_SC_MS__XOR2_1%VGND
cc_1 VNB N_B_M1002_g 0.0242428f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=0.9
cc_2 VNB N_B_M1005_g 0.0213738f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_3 VNB N_B_c_66_n 0.0341405f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_4 VNB N_B_c_67_n 0.0228401f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_5 VNB N_B_c_68_n 0.00214447f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_6 VNB N_B_c_69_n 0.0156482f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=1.565
cc_7 VNB N_A_c_133_n 0.0340508f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.845
cc_8 VNB N_A_M1008_g 0.0355836f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=1.35
cc_9 VNB N_A_c_135_n 0.0949481f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_10 VNB N_A_c_136_n 0.0125025f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_11 VNB N_A_c_137_n 0.00596229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1003_g 0.0149528f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_13 VNB N_A_M1004_g 0.0165166f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_14 VNB N_A_c_140_n 0.0616888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_141_n 0.0280619f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_16 VNB N_A_194_125#_M1009_g 0.0223322f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_17 VNB N_A_194_125#_M1007_g 5.19911e-19 $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_18 VNB N_A_194_125#_c_191_n 0.00571579f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=1.53
cc_19 VNB N_A_194_125#_c_192_n 2.29747e-19 $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_20 VNB N_A_194_125#_c_193_n 0.00598789f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.565
cc_21 VNB N_A_194_125#_c_194_n 0.034026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_276_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_343_n 0.0123304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_344_n 0.0241086f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_25 VNB X 0.00313365f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.53
cc_26 VNB N_VGND_c_379_n 0.0193241f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.805
cc_27 VNB N_VGND_c_380_n 0.0506729f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.68
cc_28 VNB N_VGND_c_381_n 0.0138262f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=1.53
cc_29 VNB N_VGND_c_382_n 0.0153054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_383_n 0.0294831f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.605
cc_31 VNB N_VGND_c_384_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_32 VNB N_VGND_c_385_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_33 VNB N_VGND_c_386_n 0.0295747f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.515
cc_34 VNB N_VGND_c_387_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.68 $Y2=1.35
cc_35 VNB N_VGND_c_388_n 0.241744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B_c_70_n 0.0251769f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.845
cc_37 VPB N_B_M1006_g 0.0221579f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_38 VPB N_B_c_66_n 0.0372241f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_39 VPB N_B_c_67_n 0.00551106f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_40 VPB N_B_c_68_n 0.00311346f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_41 VPB N_B_c_69_n 0.00639331f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.565
cc_42 VPB N_A_c_133_n 0.00954348f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.845
cc_43 VPB N_A_M1000_g 0.0303545f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=2.46
cc_44 VPB N_A_M1003_g 0.028563f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_45 VPB N_A_194_125#_M1007_g 0.0271102f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_46 VPB N_A_194_125#_c_191_n 0.00290733f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.53
cc_47 VPB N_A_194_125#_c_197_n 0.0126681f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_48 VPB N_A_194_125#_c_198_n 0.011415f $X=-0.19 $Y=1.66 $X2=1.69 $Y2=1.605
cc_49 VPB N_A_194_125#_c_192_n 0.0013189f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_50 VPB N_A_194_125#_c_200_n 0.00257826f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.68
cc_51 VPB N_VPWR_c_277_n 0.0512407f $X=-0.19 $Y=1.66 $X2=2.59 $Y2=0.805
cc_52 VPB N_VPWR_c_278_n 0.00428891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_279_n 0.0124854f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_54 VPB N_VPWR_c_280_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_55 VPB N_VPWR_c_281_n 0.043458f $X=-0.19 $Y=1.66 $X2=2.68 $Y2=1.515
cc_56 VPB N_VPWR_c_282_n 0.0328281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_276_n 0.0813681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_284_n 0.00805829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_355_368#_c_320_n 0.00941306f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_60 VPB N_A_355_368#_c_321_n 0.00275743f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.53
cc_61 VPB N_X_c_346_n 0.043147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_X_c_347_n 0.0111291f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=1.53
cc_63 VPB N_X_c_344_n 0.0077205f $X=-0.19 $Y=1.66 $X2=1.45 $Y2=1.53
cc_64 N_B_c_66_n N_A_c_133_n 0.0427299f $X=1.45 $Y=1.53 $X2=-0.19 $Y2=-0.245
cc_65 N_B_c_70_n N_A_M1000_g 0.0352137f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_66 N_B_M1002_g N_A_M1008_g 0.00791998f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_67 N_B_M1002_g N_A_c_135_n 0.00897099f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_68 N_B_M1002_g N_A_c_137_n 0.00858201f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_69 N_B_c_67_n N_A_c_137_n 0.0350732f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_70 N_B_M1006_g N_A_M1003_g 0.0389513f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_71 N_B_c_66_n N_A_M1003_g 0.0123464f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_72 N_B_c_68_n N_A_M1003_g 0.00201324f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_73 N_B_c_69_n N_A_M1003_g 0.0231094f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_74 N_B_M1002_g N_A_M1004_g 0.0119366f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_75 N_B_M1005_g N_A_M1004_g 0.0350732f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_76 N_B_M1005_g N_A_194_125#_M1009_g 0.017662f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_77 N_B_c_67_n N_A_194_125#_M1007_g 0.0282217f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B_c_70_n N_A_194_125#_c_191_n 0.00509987f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_79 N_B_M1002_g N_A_194_125#_c_191_n 0.00509445f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_80 N_B_c_66_n N_A_194_125#_c_191_n 0.0107102f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_81 N_B_c_69_n N_A_194_125#_c_191_n 0.0262124f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_82 N_B_c_70_n N_A_194_125#_c_197_n 0.0210178f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_83 N_B_M1002_g N_A_194_125#_c_208_n 0.00436246f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_84 N_B_c_66_n N_A_194_125#_c_208_n 0.0111186f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_85 N_B_c_69_n N_A_194_125#_c_208_n 0.0152632f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_86 N_B_M1006_g N_A_194_125#_c_198_n 0.0125007f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_87 N_B_c_66_n N_A_194_125#_c_198_n 0.00561489f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_88 N_B_c_67_n N_A_194_125#_c_198_n 7.04415e-19 $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B_c_68_n N_A_194_125#_c_198_n 0.023011f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B_c_69_n N_A_194_125#_c_198_n 0.0527539f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_91 N_B_M1006_g N_A_194_125#_c_192_n 0.00357343f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_92 N_B_c_67_n N_A_194_125#_c_192_n 4.25421e-19 $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B_c_68_n N_A_194_125#_c_192_n 0.00947819f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B_c_70_n N_A_194_125#_c_200_n 0.00906611f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_95 N_B_c_66_n N_A_194_125#_c_200_n 0.00895245f $X=1.45 $Y=1.53 $X2=0 $Y2=0
cc_96 N_B_c_69_n N_A_194_125#_c_200_n 0.0149541f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_97 N_B_M1005_g N_A_194_125#_c_193_n 5.92648e-19 $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_98 N_B_c_67_n N_A_194_125#_c_193_n 0.00105206f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_99 N_B_c_68_n N_A_194_125#_c_193_n 0.0243048f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_100 N_B_c_67_n N_A_194_125#_c_194_n 0.0165119f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B_c_68_n N_A_194_125#_c_194_n 3.34415e-19 $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_102 N_B_c_70_n N_VPWR_c_277_n 0.00147226f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_103 N_B_M1006_g N_VPWR_c_278_n 0.00895693f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_104 N_B_c_70_n N_VPWR_c_281_n 0.00349816f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_105 N_B_M1006_g N_VPWR_c_282_n 0.00460063f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_106 N_B_c_70_n N_VPWR_c_276_n 0.00434342f $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_107 N_B_M1006_g N_VPWR_c_276_n 0.00909121f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_108 N_B_M1006_g N_A_355_368#_c_322_n 0.0146331f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_109 N_B_c_70_n N_A_355_368#_c_320_n 9.52434e-19 $X=1.135 $Y=1.845 $X2=0 $Y2=0
cc_110 N_B_M1005_g X 0.0144534f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_111 N_B_M1005_g N_X_c_350_n 0.00594253f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_112 N_B_c_67_n N_X_c_350_n 0.00462664f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_113 N_B_c_68_n N_X_c_350_n 0.0210499f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_VGND_c_381_n 0.00705087f $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_115 N_B_M1005_g N_VGND_c_381_n 0.00272515f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_116 N_B_c_69_n N_VGND_c_381_n 0.0286839f $X=2.515 $Y=1.565 $X2=0 $Y2=0
cc_117 N_B_M1005_g N_VGND_c_382_n 6.01743e-19 $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_118 N_B_M1005_g N_VGND_c_386_n 0.00395427f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_119 N_B_M1002_g N_VGND_c_388_n 9.49986e-19 $X=1.69 $Y=0.9 $X2=0 $Y2=0
cc_120 N_B_M1005_g N_VGND_c_388_n 0.00525227f $X=2.59 $Y=0.805 $X2=0 $Y2=0
cc_121 N_A_c_133_n N_A_194_125#_c_191_n 0.0123983f $X=0.715 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_M1008_g N_A_194_125#_c_191_n 0.00959846f $X=0.895 $Y=0.9 $X2=0 $Y2=0
cc_123 N_A_c_141_n N_A_194_125#_c_191_n 0.034045f $X=0.61 $Y=1.45 $X2=0 $Y2=0
cc_124 N_A_M1000_g N_A_194_125#_c_197_n 0.00706266f $X=0.715 $Y=2.46 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_A_194_125#_c_197_n 0.00418916f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_M1008_g N_A_194_125#_c_232_n 0.00589874f $X=0.895 $Y=0.9 $X2=0 $Y2=0
cc_127 N_A_c_135_n N_A_194_125#_c_232_n 0.00100425f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_128 N_A_c_135_n N_A_194_125#_c_208_n 0.00843612f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_129 N_A_M1003_g N_A_194_125#_c_198_n 0.0149731f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A_M1000_g N_A_194_125#_c_200_n 0.00144094f $X=0.715 $Y=2.46 $X2=0 $Y2=0
cc_131 N_A_M1000_g N_VPWR_c_277_n 0.0206227f $X=0.715 $Y=2.46 $X2=0 $Y2=0
cc_132 N_A_c_140_n N_VPWR_c_277_n 0.00633983f $X=0.625 $Y=1.45 $X2=0 $Y2=0
cc_133 N_A_c_141_n N_VPWR_c_277_n 0.0172437f $X=0.61 $Y=1.45 $X2=0 $Y2=0
cc_134 N_A_M1003_g N_VPWR_c_278_n 0.0158072f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_M1000_g N_VPWR_c_281_n 0.00460063f $X=0.715 $Y=2.46 $X2=0 $Y2=0
cc_136 N_A_M1003_g N_VPWR_c_281_n 0.00490827f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_M1000_g N_VPWR_c_276_n 0.00908371f $X=0.715 $Y=2.46 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_VPWR_c_276_n 0.009739f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_M1003_g N_A_355_368#_c_322_n 0.014915f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_M1003_g N_A_355_368#_c_320_n 4.87455e-19 $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_M1004_g X 0.00192367f $X=2.2 $Y=0.805 $X2=0 $Y2=0
cc_142 N_A_M1004_g N_X_c_350_n 5.78169e-19 $X=2.2 $Y=0.805 $X2=0 $Y2=0
cc_143 N_A_c_136_n N_VGND_c_380_n 0.0232133f $X=0.97 $Y=0.18 $X2=0 $Y2=0
cc_144 N_A_c_140_n N_VGND_c_380_n 0.00360232f $X=0.625 $Y=1.45 $X2=0 $Y2=0
cc_145 N_A_c_141_n N_VGND_c_380_n 0.0484114f $X=0.61 $Y=1.45 $X2=0 $Y2=0
cc_146 N_A_c_135_n N_VGND_c_381_n 0.0226627f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_147 N_A_c_137_n N_VGND_c_381_n 9.38583e-19 $X=2.185 $Y=1.34 $X2=0 $Y2=0
cc_148 N_A_M1004_g N_VGND_c_381_n 0.0204272f $X=2.2 $Y=0.805 $X2=0 $Y2=0
cc_149 N_A_c_136_n N_VGND_c_383_n 0.0292218f $X=0.97 $Y=0.18 $X2=0 $Y2=0
cc_150 N_A_c_135_n N_VGND_c_386_n 0.00486043f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_151 N_A_c_135_n N_VGND_c_388_n 0.0354577f $X=2.125 $Y=0.18 $X2=0 $Y2=0
cc_152 N_A_c_136_n N_VGND_c_388_n 0.0106607f $X=0.97 $Y=0.18 $X2=0 $Y2=0
cc_153 N_A_194_125#_c_198_n N_VPWR_M1003_d 0.00636641f $X=3.025 $Y=2.035 $X2=0
+ $Y2=0
cc_154 N_A_194_125#_c_191_n N_VPWR_c_277_n 4.78303e-19 $X=1.03 $Y=1.95 $X2=0
+ $Y2=0
cc_155 N_A_194_125#_c_197_n N_VPWR_c_277_n 0.0463793f $X=1.36 $Y=2.815 $X2=0
+ $Y2=0
cc_156 N_A_194_125#_c_200_n N_VPWR_c_277_n 0.0093319f $X=1.36 $Y=2.115 $X2=0
+ $Y2=0
cc_157 N_A_194_125#_M1007_g N_VPWR_c_278_n 6.1181e-19 $X=3.255 $Y=2.4 $X2=0
+ $Y2=0
cc_158 N_A_194_125#_c_197_n N_VPWR_c_281_n 0.0252528f $X=1.36 $Y=2.815 $X2=0
+ $Y2=0
cc_159 N_A_194_125#_M1007_g N_VPWR_c_282_n 0.005209f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_194_125#_M1007_g N_VPWR_c_276_n 0.00987919f $X=3.255 $Y=2.4 $X2=0
+ $Y2=0
cc_161 N_A_194_125#_c_197_n N_VPWR_c_276_n 0.0204793f $X=1.36 $Y=2.815 $X2=0
+ $Y2=0
cc_162 N_A_194_125#_c_197_n A_161_392# 0.00897454f $X=1.36 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_194_125#_c_200_n A_161_392# 0.00171724f $X=1.36 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_194_125#_c_198_n N_A_355_368#_M1003_s 0.00745786f $X=3.025 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_165 N_A_194_125#_c_198_n N_A_355_368#_M1006_d 0.00684913f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_166 N_A_194_125#_c_192_n N_A_355_368#_M1006_d 0.0012728f $X=3.11 $Y=1.95
+ $X2=0 $Y2=0
cc_167 N_A_194_125#_c_198_n N_A_355_368#_c_322_n 0.0443799f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_168 N_A_194_125#_c_197_n N_A_355_368#_c_320_n 0.0492555f $X=1.36 $Y=2.815
+ $X2=0 $Y2=0
cc_169 N_A_194_125#_c_198_n N_A_355_368#_c_320_n 0.023114f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_170 N_A_194_125#_M1007_g N_A_355_368#_c_321_n 0.00900562f $X=3.255 $Y=2.4
+ $X2=0 $Y2=0
cc_171 N_A_194_125#_c_198_n N_A_355_368#_c_321_n 0.0195801f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_172 N_A_194_125#_M1009_g N_X_c_343_n 0.0166901f $X=3.16 $Y=0.805 $X2=0 $Y2=0
cc_173 N_A_194_125#_c_193_n N_X_c_343_n 0.0245397f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_174 N_A_194_125#_c_194_n N_X_c_343_n 0.00434404f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_175 N_A_194_125#_M1007_g N_X_c_347_n 0.00200568f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A_194_125#_c_192_n N_X_c_347_n 0.00518253f $X=3.11 $Y=1.95 $X2=0 $Y2=0
cc_177 N_A_194_125#_c_193_n N_X_c_347_n 0.00413233f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_178 N_A_194_125#_c_194_n N_X_c_347_n 0.00114149f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_179 N_A_194_125#_M1009_g N_X_c_344_n 0.00477786f $X=3.16 $Y=0.805 $X2=0 $Y2=0
cc_180 N_A_194_125#_M1007_g N_X_c_344_n 0.00344259f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_194_125#_c_192_n N_X_c_344_n 0.00651142f $X=3.11 $Y=1.95 $X2=0 $Y2=0
cc_182 N_A_194_125#_c_193_n N_X_c_344_n 0.0250916f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_183 N_A_194_125#_c_194_n N_X_c_344_n 0.00231223f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_184 N_A_194_125#_M1009_g X 0.00974015f $X=3.16 $Y=0.805 $X2=0 $Y2=0
cc_185 N_A_194_125#_M1009_g N_VGND_c_382_n 0.00972215f $X=3.16 $Y=0.805 $X2=0
+ $Y2=0
cc_186 N_A_194_125#_c_232_n N_VGND_c_383_n 0.00228482f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_187 N_A_194_125#_c_208_n N_VGND_c_383_n 0.00771542f $X=1.475 $Y=0.875 $X2=0
+ $Y2=0
cc_188 N_A_194_125#_M1009_g N_VGND_c_386_n 0.00441186f $X=3.16 $Y=0.805 $X2=0
+ $Y2=0
cc_189 N_A_194_125#_M1009_g N_VGND_c_388_n 0.0044119f $X=3.16 $Y=0.805 $X2=0
+ $Y2=0
cc_190 N_A_194_125#_c_232_n N_VGND_c_388_n 0.00415706f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_191 N_A_194_125#_c_208_n N_VGND_c_388_n 0.012469f $X=1.475 $Y=0.875 $X2=0
+ $Y2=0
cc_192 N_VPWR_M1003_d N_A_355_368#_c_322_n 0.00621325f $X=2.275 $Y=1.84 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_278_n N_A_355_368#_c_322_n 0.0239701f $X=2.475 $Y=2.815 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_278_n N_A_355_368#_c_320_n 0.01373f $X=2.475 $Y=2.815 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_281_n N_A_355_368#_c_320_n 0.0146513f $X=2.255 $Y=3.33 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_276_n N_A_355_368#_c_320_n 0.0121202f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_278_n N_A_355_368#_c_321_n 0.01373f $X=2.475 $Y=2.815 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_282_n N_A_355_368#_c_321_n 0.0145644f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_276_n N_A_355_368#_c_321_n 0.0119803f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_200 N_VPWR_c_282_n N_X_c_346_n 0.0173129f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_276_n N_X_c_346_n 0.0143301f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_202 N_A_355_368#_c_321_n N_X_c_346_n 0.0202848f $X=3.03 $Y=2.455 $X2=0 $Y2=0
cc_203 N_X_c_343_n N_VGND_M1009_d 0.0136501f $X=3.585 $Y=1.065 $X2=0 $Y2=0
cc_204 N_X_c_344_n N_VGND_M1009_d 3.82603e-19 $X=3.56 $Y=1.82 $X2=0 $Y2=0
cc_205 X N_VGND_c_381_n 0.0229507f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_206 N_X_c_350_n N_VGND_c_381_n 0.00716572f $X=2.747 $Y=0.98 $X2=0 $Y2=0
cc_207 N_X_c_343_n N_VGND_c_382_n 0.0171814f $X=3.585 $Y=1.065 $X2=0 $Y2=0
cc_208 X N_VGND_c_382_n 0.0201618f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_209 X N_VGND_c_386_n 0.0152785f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_210 X N_VGND_c_388_n 0.0155747f $X=2.555 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a211oi_1.pxi.spice
* Created: Fri Aug 28 16:57:05 2020
* 
x_PM_SKY130_FD_SC_MS__A211OI_1%A2 N_A2_M1005_g N_A2_M1003_g A2 N_A2_c_52_n
+ N_A2_c_53_n PM_SKY130_FD_SC_MS__A211OI_1%A2
x_PM_SKY130_FD_SC_MS__A211OI_1%A1 N_A1_M1001_g N_A1_M1000_g A1 N_A1_c_83_n
+ N_A1_c_84_n PM_SKY130_FD_SC_MS__A211OI_1%A1
x_PM_SKY130_FD_SC_MS__A211OI_1%B1 N_B1_M1004_g N_B1_M1002_g B1 N_B1_c_122_n
+ N_B1_c_123_n PM_SKY130_FD_SC_MS__A211OI_1%B1
x_PM_SKY130_FD_SC_MS__A211OI_1%C1 N_C1_c_157_n N_C1_M1007_g N_C1_M1006_g
+ N_C1_c_159_n C1 N_C1_c_161_n PM_SKY130_FD_SC_MS__A211OI_1%C1
x_PM_SKY130_FD_SC_MS__A211OI_1%A_71_368# N_A_71_368#_M1005_s N_A_71_368#_M1000_d
+ N_A_71_368#_c_186_n N_A_71_368#_c_187_n N_A_71_368#_c_193_n
+ N_A_71_368#_c_200_n N_A_71_368#_c_188_n PM_SKY130_FD_SC_MS__A211OI_1%A_71_368#
x_PM_SKY130_FD_SC_MS__A211OI_1%VPWR N_VPWR_M1005_d N_VPWR_c_218_n N_VPWR_c_219_n
+ N_VPWR_c_220_n VPWR N_VPWR_c_221_n N_VPWR_c_217_n
+ PM_SKY130_FD_SC_MS__A211OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A211OI_1%Y N_Y_M1001_d N_Y_M1007_d N_Y_M1006_d N_Y_c_243_n
+ N_Y_c_244_n N_Y_c_249_n N_Y_c_245_n N_Y_c_250_n N_Y_c_246_n Y Y Y N_Y_c_248_n
+ PM_SKY130_FD_SC_MS__A211OI_1%Y
x_PM_SKY130_FD_SC_MS__A211OI_1%VGND N_VGND_M1003_s N_VGND_M1004_d N_VGND_c_294_n
+ N_VGND_c_295_n N_VGND_c_296_n N_VGND_c_297_n VGND N_VGND_c_298_n
+ N_VGND_c_299_n N_VGND_c_300_n N_VGND_c_301_n PM_SKY130_FD_SC_MS__A211OI_1%VGND
cc_1 VNB N_A2_M1003_g 0.03136f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_2 VNB N_A2_c_52_n 0.0349485f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_3 VNB N_A2_c_53_n 0.0052161f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_4 VNB N_A1_M1001_g 0.0248902f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_5 VNB N_A1_c_83_n 0.0262505f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_6 VNB N_A1_c_84_n 0.00166449f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_7 VNB N_B1_M1004_g 0.0261208f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_8 VNB N_B1_c_122_n 0.026255f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_9 VNB N_B1_c_123_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_10 VNB N_C1_c_157_n 0.0234756f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.68
cc_11 VNB N_C1_M1006_g 0.00842224f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_12 VNB N_C1_c_159_n 0.0113697f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB C1 0.0207309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C1_c_161_n 0.0638365f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_15 VNB N_VPWR_c_217_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_243_n 0.00792442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_244_n 0.00317771f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_18 VNB N_Y_c_245_n 0.0204378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_246_n 0.00374926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.0086849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_248_n 0.00924258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_294_n 0.0457851f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_VGND_c_295_n 0.00685406f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_24 VNB N_VGND_c_296_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_25 VNB N_VGND_c_297_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_298_n 0.028216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_299_n 0.0263115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_300_n 0.202322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_301_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A2_M1005_g 0.0288353f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_31 VPB N_A2_c_52_n 0.00618442f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_32 VPB N_A2_c_53_n 0.00630921f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_33 VPB N_A1_M1000_g 0.0226496f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_34 VPB N_A1_c_83_n 0.00561631f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_35 VPB N_A1_c_84_n 0.00200771f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_36 VPB N_B1_M1002_g 0.0215077f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_37 VPB N_B1_c_122_n 0.0055922f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_38 VPB N_B1_c_123_n 0.00525799f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_39 VPB N_C1_M1006_g 0.0308618f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_40 VPB N_A_71_368#_c_186_n 0.00880428f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_41 VPB N_A_71_368#_c_187_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_42 VPB N_A_71_368#_c_188_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.68
cc_43 VPB N_VPWR_c_218_n 0.00958227f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_44 VPB N_VPWR_c_219_n 0.0255159f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_45 VPB N_VPWR_c_220_n 0.00612923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_221_n 0.0510638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_217_n 0.0811476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_Y_c_249_n 0.0398433f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.665
cc_49 VPB N_Y_c_250_n 0.0140179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_Y_c_246_n 0.00115044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 N_A2_M1003_g N_A1_M1001_g 0.0426951f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_52 N_A2_M1005_g N_A1_M1000_g 0.032177f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_53 N_A2_c_53_n N_A1_M1000_g 2.6794e-19 $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_54 N_A2_c_52_n N_A1_c_83_n 0.0426951f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_55 N_A2_c_53_n N_A1_c_83_n 0.00188197f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_56 N_A2_M1005_g N_A1_c_84_n 3.38956e-19 $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A2_c_52_n N_A1_c_84_n 3.80681e-19 $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_58 N_A2_c_53_n N_A1_c_84_n 0.0347534f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_59 N_A2_M1005_g N_A_71_368#_c_186_n 8.8334e-19 $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_60 N_A2_c_52_n N_A_71_368#_c_186_n 7.74224e-19 $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_61 N_A2_c_53_n N_A_71_368#_c_186_n 0.0130747f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_62 N_A2_M1005_g N_A_71_368#_c_187_n 0.0126445f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A2_M1005_g N_A_71_368#_c_193_n 0.0133755f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_64 N_A2_c_53_n N_A_71_368#_c_193_n 0.0126649f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_65 N_A2_M1005_g N_A_71_368#_c_188_n 6.0235e-19 $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A2_M1005_g N_VPWR_c_218_n 0.00340108f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_67 N_A2_M1005_g N_VPWR_c_219_n 0.005209f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_68 N_A2_M1005_g N_VPWR_c_217_n 0.0098676f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A2_M1003_g N_Y_c_243_n 0.0012054f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A2_M1003_g N_Y_c_244_n 0.00134279f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A2_M1003_g N_VGND_c_294_n 0.0188126f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A2_c_52_n N_VGND_c_294_n 0.00136988f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A2_c_53_n N_VGND_c_294_n 0.0143146f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A2_M1003_g N_VGND_c_298_n 0.00383152f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_75 N_A2_M1003_g N_VGND_c_300_n 0.0075694f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A1_M1001_g N_B1_M1004_g 0.0223185f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A1_M1000_g N_B1_M1002_g 0.0153548f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_78 N_A1_c_83_n N_B1_c_122_n 0.0201104f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A1_c_84_n N_B1_c_122_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A1_M1000_g N_B1_c_123_n 5.95548e-19 $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A1_c_83_n N_B1_c_123_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A1_c_84_n N_B1_c_123_n 0.0276387f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A1_M1000_g N_A_71_368#_c_187_n 6.73208e-19 $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A1_M1000_g N_A_71_368#_c_193_n 0.0133755f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A1_c_83_n N_A_71_368#_c_193_n 6.98124e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A1_c_84_n N_A_71_368#_c_193_n 0.0208108f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A1_M1000_g N_A_71_368#_c_200_n 8.8334e-19 $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A1_c_84_n N_A_71_368#_c_200_n 0.00237219f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A1_M1000_g N_A_71_368#_c_188_n 0.0122049f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A1_M1000_g N_VPWR_c_218_n 0.00732726f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A1_M1000_g N_VPWR_c_221_n 0.005209f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A1_M1000_g N_VPWR_c_217_n 0.00982607f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A1_M1001_g N_Y_c_243_n 0.00897846f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A1_c_83_n N_Y_c_243_n 0.00139983f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_95 N_A1_c_84_n N_Y_c_243_n 0.0211742f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A1_M1001_g N_Y_c_244_n 0.0100683f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A1_M1001_g N_VGND_c_294_n 0.00263599f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A1_M1001_g N_VGND_c_295_n 5.90483e-19 $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A1_M1001_g N_VGND_c_298_n 0.00383287f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A1_M1001_g N_VGND_c_300_n 0.00656608f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1004_g N_C1_c_157_n 0.0248511f $X=1.62 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_102 N_B1_M1002_g N_C1_M1006_g 0.0553717f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_103 N_B1_c_123_n N_C1_M1006_g 3.24593e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B1_c_122_n N_C1_c_159_n 0.0206204f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B1_c_123_n N_C1_c_159_n 3.78988e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_106 N_B1_M1002_g N_A_71_368#_c_200_n 0.00323121f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_107 N_B1_c_122_n N_A_71_368#_c_200_n 2.16516e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_c_123_n N_A_71_368#_c_200_n 0.00508185f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_A_71_368#_c_188_n 0.0150131f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_110 N_B1_M1002_g N_VPWR_c_221_n 0.005209f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_111 N_B1_M1002_g N_VPWR_c_217_n 0.00983863f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_112 N_B1_M1004_g N_Y_c_244_n 0.0026934f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B1_M1004_g N_Y_c_245_n 6.39617e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_M1004_g N_Y_c_246_n 0.00296121f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B1_M1002_g N_Y_c_246_n 0.00509978f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B1_c_122_n N_Y_c_246_n 0.00174016f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_117 N_B1_c_123_n N_Y_c_246_n 0.032728f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B1_M1004_g N_Y_c_248_n 0.0217865f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_119 N_B1_c_122_n N_Y_c_248_n 0.00132988f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_120 N_B1_c_123_n N_Y_c_248_n 0.0262137f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_121 N_B1_M1004_g N_VGND_c_295_n 0.00776565f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_122 N_B1_M1004_g N_VGND_c_298_n 0.00383152f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B1_M1004_g N_VGND_c_300_n 0.00378707f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_124 N_C1_M1006_g N_A_71_368#_c_188_n 8.49227e-19 $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_125 N_C1_M1006_g N_VPWR_c_221_n 0.00349816f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_126 N_C1_M1006_g N_VPWR_c_217_n 0.00434046f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_127 N_C1_M1006_g N_Y_c_249_n 0.0225119f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_128 N_C1_c_157_n N_Y_c_245_n 0.00733151f $X=2.16 $Y=1.22 $X2=0 $Y2=0
cc_129 N_C1_M1006_g N_Y_c_250_n 0.00850298f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_130 C1 N_Y_c_250_n 0.00712672f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_131 N_C1_c_161_n N_Y_c_250_n 0.00809123f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_132 N_C1_c_157_n N_Y_c_246_n 9.75292e-19 $X=2.16 $Y=1.22 $X2=0 $Y2=0
cc_133 N_C1_M1006_g N_Y_c_246_n 0.0141712f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_134 N_C1_c_159_n N_Y_c_246_n 0.0106477f $X=2.175 $Y=1.385 $X2=0 $Y2=0
cc_135 C1 N_Y_c_246_n 0.0208673f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_136 N_C1_c_157_n Y 0.0214366f $X=2.16 $Y=1.22 $X2=0 $Y2=0
cc_137 C1 Y 0.00830742f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_138 N_C1_c_161_n Y 0.00747729f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_139 N_C1_c_157_n N_VGND_c_295_n 0.00493436f $X=2.16 $Y=1.22 $X2=0 $Y2=0
cc_140 N_C1_c_157_n N_VGND_c_299_n 0.00434272f $X=2.16 $Y=1.22 $X2=0 $Y2=0
cc_141 N_C1_c_157_n N_VGND_c_300_n 0.00443636f $X=2.16 $Y=1.22 $X2=0 $Y2=0
cc_142 N_A_71_368#_c_193_n N_VPWR_M1005_d 0.00928873f $X=1.305 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_143 N_A_71_368#_c_187_n N_VPWR_c_218_n 0.0266772f $X=0.48 $Y=2.815 $X2=0
+ $Y2=0
cc_144 N_A_71_368#_c_193_n N_VPWR_c_218_n 0.0200142f $X=1.305 $Y=2.035 $X2=0
+ $Y2=0
cc_145 N_A_71_368#_c_188_n N_VPWR_c_218_n 0.0266772f $X=1.47 $Y=2.815 $X2=0
+ $Y2=0
cc_146 N_A_71_368#_c_187_n N_VPWR_c_219_n 0.014549f $X=0.48 $Y=2.815 $X2=0 $Y2=0
cc_147 N_A_71_368#_c_188_n N_VPWR_c_221_n 0.0144436f $X=1.47 $Y=2.815 $X2=0
+ $Y2=0
cc_148 N_A_71_368#_c_187_n N_VPWR_c_217_n 0.0119743f $X=0.48 $Y=2.815 $X2=0
+ $Y2=0
cc_149 N_A_71_368#_c_188_n N_VPWR_c_217_n 0.0118287f $X=1.47 $Y=2.815 $X2=0
+ $Y2=0
cc_150 N_A_71_368#_c_188_n N_Y_c_249_n 0.0163051f $X=1.47 $Y=2.815 $X2=0 $Y2=0
cc_151 N_VPWR_c_221_n N_Y_c_249_n 0.0225756f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_152 N_VPWR_c_217_n N_Y_c_249_n 0.0182633f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_153 N_Y_c_248_n N_VGND_M1004_d 0.00345356f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_154 N_Y_c_243_n N_VGND_c_294_n 0.0123945f $X=1.292 $Y=0.81 $X2=0 $Y2=0
cc_155 N_Y_c_244_n N_VGND_c_294_n 0.0170764f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_156 N_Y_c_244_n N_VGND_c_295_n 0.0118921f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_157 N_Y_c_245_n N_VGND_c_295_n 0.0116858f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_158 N_Y_c_248_n N_VGND_c_295_n 0.0249165f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_159 N_Y_c_244_n N_VGND_c_298_n 0.0182222f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_160 N_Y_c_245_n N_VGND_c_299_n 0.0145369f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_161 N_Y_c_244_n N_VGND_c_300_n 0.0149207f $X=1.315 $Y=0.515 $X2=0 $Y2=0
cc_162 N_Y_c_245_n N_VGND_c_300_n 0.0119879f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_163 Y N_VGND_c_300_n 0.0057112f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_164 N_Y_c_248_n N_VGND_c_300_n 0.00707419f $X=2.045 $Y=0.995 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__sdfrtp_1.pex.spice
* Created: Wed Sep  2 12:30:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%SCE 3 7 11 17 18 19 20 23 24 28 29 30 38 42
+ 44 53 55
c90 38 0 9.7872e-20 $X=0.96 $Y=1.67
c91 24 0 1.56864e-19 $X=2.51 $Y=1.425
c92 23 0 2.15287e-19 $X=2.51 $Y=1.425
r93 44 53 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r94 38 40 6.6128 $w=3.28e-07 $l=4.5e-08 $layer=POLY_cond $X=0.96 $Y=1.67
+ $X2=1.005 $Y2=1.67
r95 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.96
+ $Y=1.67 $X2=0.96 $Y2=1.67
r96 36 38 66.8628 $w=3.28e-07 $l=4.55e-07 $layer=POLY_cond $X=0.505 $Y=1.67
+ $X2=0.96 $Y2=1.67
r97 35 36 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.67
+ $X2=0.505 $Y2=1.67
r98 30 55 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r99 30 53 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r100 30 44 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r101 29 30 13.6623 $w=3.43e-07 $l=4.09e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.609 $Y2=1.662
r102 29 39 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=0.96 $Y2=1.662
r103 28 39 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=1.662
+ $X2=0.96 $Y2=1.662
r104 24 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.425
+ $X2=2.51 $Y2=1.26
r105 23 26 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.535 $Y=1.425
+ $X2=2.535 $Y2=1.575
r106 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.425 $X2=2.51 $Y2=1.425
r107 20 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.345 $Y=1.575
+ $X2=2.535 $Y2=1.575
r108 20 55 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.345 $Y=1.575
+ $X2=1.795 $Y2=1.575
r109 19 42 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.6 $Y=1.05 $X2=2.6
+ $Y2=1.26
r110 18 19 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.625 $Y=0.9
+ $X2=2.625 $Y2=1.05
r111 17 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.65 $Y=0.615
+ $X2=2.65 $Y2=0.9
r112 9 40 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.835
+ $X2=1.005 $Y2=1.67
r113 9 11 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=1.005 $Y=1.835
+ $X2=1.005 $Y2=2.64
r114 5 35 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=1.67
r115 5 7 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.65
r116 1 36 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r117 1 3 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_27_88# 1 2 7 9 12 14 18 21 24 26 30 32 33
+ 35 36 38 39 43
c82 38 0 9.7872e-20 $X=1.21 $Y=1.1
c83 7 0 3.56444e-20 $X=1.485 $Y=0.935
r84 38 41 1.99058 $w=3.28e-07 $l=5.7e-08 $layer=LI1_cond $X=1.21 $Y=1.1 $X2=1.21
+ $Y2=1.157
r85 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.1 $X2=1.21 $Y2=1.1
r86 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.51
+ $Y=1.995 $X2=2.51 $Y2=1.995
r87 30 43 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=2.207 $Y=2.002
+ $X2=2.035 $Y2=2.002
r88 30 32 10.1215 $w=3.43e-07 $l=3.03e-07 $layer=LI1_cond $X=2.207 $Y=2.002
+ $X2=2.51 $Y2=2.002
r89 29 36 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r90 29 43 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=2.035 $Y2=2.09
r91 27 35 1.25797 $w=2.15e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.157
+ $X2=0.24 $Y2=1.157
r92 26 41 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=1.157
+ $X2=1.21 $Y2=1.157
r93 26 27 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=1.157
+ $X2=0.365 $Y2=1.157
r94 22 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r95 22 24 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r96 21 36 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r97 20 35 5.26796 $w=2.1e-07 $l=1.26428e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.157
r98 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265 $X2=0.2
+ $Y2=2.005
r99 16 35 5.26796 $w=2.1e-07 $l=1.07e-07 $layer=LI1_cond $X=0.24 $Y=1.05
+ $X2=0.24 $Y2=1.157
r100 16 18 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=1.05 $X2=0.24
+ $Y2=0.65
r101 12 33 19.4618 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=2.16
+ $X2=2.585 $Y2=1.995
r102 12 14 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2.585 $Y=2.16
+ $X2=2.585 $Y2=2.64
r103 7 39 50.0189 $w=2.65e-07 $l=3.47851e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.21 $Y2=1.1
r104 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r105 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r106 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%D 1 3 5 7 10 13 17 19 22 23 24
c56 17 0 6.10037e-20 $X=1.845 $Y=1.515
c57 5 0 1.54283e-19 $X=1.69 $Y=2.075
r58 22 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=1.935 $Y2=1.265
r59 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=1.935 $Y2=0.935
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r61 19 23 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r62 15 17 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.845 $Y2=1.515
r63 10 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=0.615
+ $X2=1.875 $Y2=0.935
r64 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.44
+ $X2=1.845 $Y2=1.515
r65 7 25 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.845 $Y=1.44
+ $X2=1.845 $Y2=1.265
r66 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=2.075
+ $X2=1.69 $Y2=2.15
r67 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.59 $X2=1.69
+ $Y2=1.515
r68 4 5 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.69 $Y=1.59 $X2=1.69
+ $Y2=2.075
r69 1 13 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.425 $Y=2.15
+ $X2=1.69 $Y2=2.15
r70 1 3 111.128 $w=1.8e-07 $l=4.15e-07 $layer=POLY_cond $X=1.425 $Y=2.225
+ $X2=1.425 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%SCD 3 6 10 11 12 13 17
c41 12 0 1.56864e-19 $X=3.12 $Y=1.665
c42 11 0 9.0609e-20 $X=3.05 $Y=2.245
c43 6 0 1.93733e-19 $X=3.04 $Y=0.615
r44 12 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r45 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.605 $X2=3.05 $Y2=1.605
r46 10 17 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=1.605
r47 10 11 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=2.08
+ $X2=3.05 $Y2=2.245
r48 9 17 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.44
+ $X2=3.05 $Y2=1.605
r49 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.04 $Y=0.615
+ $X2=3.04 $Y2=1.44
r50 3 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.64
+ $X2=3.035 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%CLK 1 3 4 6 7
r56 10 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=1.455 $X2=3.95 $Y2=1.455
r57 7 11 3.23179 $w=6.04e-07 $l=1.6e-07 $layer=LI1_cond $X=4.212 $Y=1.295
+ $X2=4.212 $Y2=1.455
r58 4 13 18.5736 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.645 $Y=1.86
+ $X2=4.645 $Y2=1.575
r59 4 6 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=4.645 $Y=1.86
+ $X2=4.645 $Y2=2.495
r60 1 13 6.80791 $w=3.54e-07 $l=5e-08 $layer=POLY_cond $X=4.595 $Y=1.575
+ $X2=4.645 $Y2=1.575
r61 1 10 87.822 $w=3.54e-07 $l=6.45e-07 $layer=POLY_cond $X=4.595 $Y=1.575
+ $X2=3.95 $Y2=1.575
r62 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.595 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_1037_387# 1 2 9 11 15 17 19 21 24 29 31
+ 32 33 34 36 40 41 42 44 45 46 48 50 51 53 60 65 66 68 73 77
c208 68 0 2.21673e-19 $X=6.065 $Y=1.65
c209 66 0 1.39473e-19 $X=9.33 $Y=1.105
c210 42 0 1.61901e-19 $X=7.22 $Y=0.665
c211 15 0 6.25949e-20 $X=6.525 $Y=0.805
c212 9 0 3.12154e-19 $X=6.135 $Y=2.495
r213 65 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.105
+ $X2=9.085 $Y2=1.105
r214 64 66 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.25 $Y=1.105 $X2=9.33
+ $Y2=1.105
r215 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.25
+ $Y=1.105 $X2=9.25 $Y2=1.105
r216 61 64 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=9.15 $Y=1.105
+ $X2=9.25 $Y2=1.105
r217 59 60 8.01921 $w=4.03e-07 $l=1.55e-07 $layer=LI1_cond $X=5.422 $Y=1.11
+ $X2=5.422 $Y2=1.265
r218 54 77 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=9.81 $Y=2.215
+ $X2=9.89 $Y2=2.215
r219 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.81
+ $Y=2.215 $X2=9.81 $Y2=2.215
r220 51 53 17.8516 $w=2.53e-07 $l=3.95e-07 $layer=LI1_cond $X=9.415 $Y=2.252
+ $X2=9.81 $Y2=2.252
r221 50 51 7.17723 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=9.33 $Y=2.125
+ $X2=9.415 $Y2=2.252
r222 49 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.33 $Y=1.27
+ $X2=9.33 $Y2=1.105
r223 49 50 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=9.33 $Y=1.27
+ $X2=9.33 $Y2=2.125
r224 48 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=0.94
+ $X2=9.15 $Y2=1.105
r225 47 48 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.15 $Y=0.425
+ $X2=9.15 $Y2=0.94
r226 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.065 $Y=0.34
+ $X2=9.15 $Y2=0.425
r227 45 46 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=9.065 $Y=0.34
+ $X2=8.1 $Y2=0.34
r228 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r229 43 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r230 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r231 41 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.22 $Y2=0.665
r232 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.135 $Y=0.58
+ $X2=7.22 $Y2=0.665
r233 39 40 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.135 $Y=0.425
+ $X2=7.135 $Y2=0.58
r234 37 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.71
+ $X2=6.065 $Y2=1.875
r235 37 68 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.065 $Y=1.71
+ $X2=6.065 $Y2=1.65
r236 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.71 $X2=6.065 $Y2=1.71
r237 34 58 16.4 $w=3.05e-07 $l=5.50073e-07 $layer=LI1_cond $X=5.63 $Y=1.71
+ $X2=5.302 $Y2=2.12
r238 34 36 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.63 $Y=1.71
+ $X2=6.065 $Y2=1.71
r239 32 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=7.135 $Y2=0.425
r240 32 33 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.05 $Y=0.34
+ $X2=5.62 $Y2=0.34
r241 31 34 8.63237 $w=3.05e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.63 $Y2=1.71
r242 31 60 17.2525 $w=1.78e-07 $l=2.8e-07 $layer=LI1_cond $X=5.54 $Y=1.545
+ $X2=5.54 $Y2=1.265
r243 29 59 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=5.417 $Y=0.74
+ $X2=5.417 $Y2=1.11
r244 26 33 8.41448 $w=1.7e-07 $l=2.41793e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.62 $Y2=0.34
r245 26 29 8.96345 $w=4.03e-07 $l=3.15e-07 $layer=LI1_cond $X=5.417 $Y=0.425
+ $X2=5.417 $Y2=0.74
r246 22 77 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.89 $Y=2.38
+ $X2=9.89 $Y2=2.215
r247 22 24 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.89 $Y=2.38
+ $X2=9.89 $Y2=2.75
r248 21 73 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.725 $Y=1.16
+ $X2=9.085 $Y2=1.16
r249 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.725 $Y2=1.16
r250 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.65 $Y2=0.69
r251 13 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.525 $Y=1.575
+ $X2=6.525 $Y2=0.805
r252 12 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.65
+ $X2=6.065 $Y2=1.65
r253 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.45 $Y=1.65
+ $X2=6.525 $Y2=1.575
r254 11 12 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=6.45 $Y=1.65
+ $X2=6.23 $Y2=1.65
r255 9 71 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=6.135 $Y=2.495 $X2=6.135
+ $Y2=1.875
r256 2 58 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.935 $X2=5.32 $Y2=2.12
r257 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.595 $X2=5.36 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_1367_93# 1 2 9 13 17 18 20 21 24 26 31 33
c104 17 0 4.99889e-20 $X=7.185 $Y=1.64
c105 9 0 1.55517e-19 $X=6.91 $Y=0.805
r106 34 36 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.91 $Y=1.64
+ $X2=7.06 $Y2=1.64
r107 26 28 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=8.865 $Y=1.88
+ $X2=8.865 $Y2=2.59
r108 24 33 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=8.865 $Y=1.855
+ $X2=8.865 $Y2=1.715
r109 24 26 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=8.865 $Y=1.855
+ $X2=8.865 $Y2=1.88
r110 22 31 12.3649 $w=3.7e-07 $l=4.83348e-07 $layer=LI1_cond $X=8.81 $Y=1.09
+ $X2=8.435 $Y2=0.842
r111 22 33 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.81 $Y=1.09
+ $X2=8.81 $Y2=1.715
r112 20 31 9.03936 $w=3.7e-07 $l=2.32637e-07 $layer=LI1_cond $X=8.27 $Y=1.005
+ $X2=8.435 $Y2=0.842
r113 20 21 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=8.27 $Y=1.005
+ $X2=7.325 $Y2=1.005
r114 18 36 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.185 $Y=1.64
+ $X2=7.06 $Y2=1.64
r115 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.185
+ $Y=1.64 $X2=7.185 $Y2=1.64
r116 15 21 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=7.187 $Y=1.09
+ $X2=7.325 $Y2=1.005
r117 15 17 23.0489 $w=2.73e-07 $l=5.5e-07 $layer=LI1_cond $X=7.187 $Y=1.09
+ $X2=7.187 $Y2=1.64
r118 11 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.06 $Y=1.805
+ $X2=7.06 $Y2=1.64
r119 11 13 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=7.06 $Y=1.805
+ $X2=7.06 $Y2=2.515
r120 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=1.64
r121 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.91 $Y=1.475
+ $X2=6.91 $Y2=0.805
r122 2 28 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=1.735 $X2=8.92 $Y2=2.59
r123 2 26 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=1.735 $X2=8.92 $Y2=1.88
r124 1 31 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.37 $X2=8.435 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%RESET_B 4 7 8 9 10 11 15 16 17 19 22 26 29
+ 32 36 39 41 42 43 44 51 52 56 61 68 69
c225 43 0 1.37312e-19 $X=10.655 $Y=2.035
c226 39 0 6.31244e-20 $X=10.715 $Y=1.375
c227 26 0 5.21422e-20 $X=10.6 $Y=0.58
c228 15 0 1.88097e-19 $X=7.3 $Y=0.805
r229 67 69 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=10.805 $Y=1.985
+ $X2=10.885 $Y2=1.985
r230 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.805
+ $Y=1.985 $X2=10.805 $Y2=1.985
r231 64 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.715 $Y=1.985
+ $X2=10.805 $Y2=1.985
r232 59 61 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=7.685 $Y=1.98
+ $X2=8 $Y2=1.98
r233 57 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.67 $Y=1.98
+ $X2=7.685 $Y2=1.98
r234 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r235 52 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r236 51 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8 $Y=1.98
+ $X2=8 $Y2=1.98
r237 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r238 46 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r239 44 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r240 43 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r241 43 44 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r242 42 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r243 41 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r244 41 42 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r245 37 39 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=10.6 $Y=1.375
+ $X2=10.715 $Y2=1.375
r246 30 69 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.885 $Y=2.15
+ $X2=10.885 $Y2=1.985
r247 30 32 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=10.885 $Y=2.15
+ $X2=10.885 $Y2=2.75
r248 29 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.82
+ $X2=10.715 $Y2=1.985
r249 28 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.45
+ $X2=10.715 $Y2=1.375
r250 28 29 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.715 $Y=1.45
+ $X2=10.715 $Y2=1.82
r251 24 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.6 $Y2=1.375
r252 24 26 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.6 $Y2=0.58
r253 20 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.685 $Y=2.145
+ $X2=7.685 $Y2=1.98
r254 20 22 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.685 $Y=2.145
+ $X2=7.685 $Y2=2.515
r255 19 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.815
+ $X2=7.67 $Y2=1.98
r256 18 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.67 $Y=1.265
+ $X2=7.67 $Y2=1.815
r257 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.595 $Y=1.19
+ $X2=7.67 $Y2=1.265
r258 16 17 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=7.595 $Y=1.19
+ $X2=7.375 $Y2=1.19
r259 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.375 $Y2=1.19
r260 13 15 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.3 $Y=1.115
+ $X2=7.3 $Y2=0.805
r261 12 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.3 $Y=0.255
+ $X2=7.3 $Y2=0.805
r262 11 36 62.2243 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=2.245
r263 11 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.995
+ $X2=3.56 $Y2=1.83
r264 10 55 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.95 $Y2=1.995
r265 10 11 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.695 $Y2=1.995
r266 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=7.3 $Y2=0.255
r267 8 9 1871.6 $w=1.5e-07 $l=3.65e-06 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=3.575 $Y2=0.18
r268 7 36 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.64
+ $X2=3.605 $Y2=2.245
r269 4 35 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.5 $Y=0.615
+ $X2=3.5 $Y2=1.83
r270 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=0.255
+ $X2=3.575 $Y2=0.18
r271 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.5 $Y=0.255 $X2=3.5
+ $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_1234_119# 1 2 3 12 14 18 20 24 27 28 31
+ 32 34 35 38 42
c129 42 0 1.37527e-19 $X=6.795 $Y=2.522
c130 35 0 4.99889e-20 $X=8.15 $Y=1.41
c131 31 0 7.00504e-20 $X=7.58 $Y=2.32
c132 27 0 3.71649e-19 $X=6.795 $Y=2.32
c133 24 0 1.51838e-20 $X=6.71 $Y=0.945
c134 20 0 1.74626e-19 $X=6.71 $Y=2.555
r135 38 40 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=6.307 $Y=0.81
+ $X2=6.307 $Y2=0.945
r136 35 47 16.6207 $w=3.19e-07 $l=1.1e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.52
r137 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.15
+ $Y=1.41 $X2=8.15 $Y2=1.41
r138 32 34 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=7.665 $Y=1.417
+ $X2=8.15 $Y2=1.417
r139 31 45 12.781 $w=3.15e-07 $l=4.22918e-07 $layer=LI1_cond $X=7.58 $Y=2.32
+ $X2=7.91 $Y2=2.532
r140 30 32 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.665 $Y2=1.417
r141 30 31 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.58 $Y2=2.32
r142 29 42 3.64284 $w=2.55e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.88 $Y=2.405
+ $X2=6.795 $Y2=2.522
r143 28 31 5.86024 $w=3.15e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=7.58 $Y2=2.32
r144 28 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=6.88 $Y2=2.405
r145 27 42 2.83584 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=6.795 $Y=2.32
+ $X2=6.795 $Y2=2.522
r146 26 27 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=6.795 $Y=1.03
+ $X2=6.795 $Y2=2.32
r147 25 40 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=6.47 $Y=0.945
+ $X2=6.307 $Y2=0.945
r148 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.71 $Y=0.945
+ $X2=6.795 $Y2=1.03
r149 24 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.71 $Y=0.945
+ $X2=6.47 $Y2=0.945
r150 20 42 3.64284 $w=2.55e-07 $l=1.0015e-07 $layer=LI1_cond $X=6.71 $Y=2.555
+ $X2=6.795 $Y2=2.522
r151 20 22 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=6.71 $Y=2.555
+ $X2=6.415 $Y2=2.555
r152 16 18 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=8.695 $Y=1.595
+ $X2=8.695 $Y2=2.235
r153 15 47 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.52
+ $X2=8.15 $Y2=1.52
r154 14 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.605 $Y=1.52
+ $X2=8.695 $Y2=1.595
r155 14 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.605 $Y=1.52
+ $X2=8.315 $Y2=1.52
r156 10 35 38.5462 $w=3.19e-07 $l=1.96914e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.15 $Y2=1.41
r157 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.22 $Y=1.245
+ $X2=8.22 $Y2=0.69
r158 3 45 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=2.305 $X2=7.91 $Y2=2.53
r159 2 22 600 $w=1.7e-07 $l=3.5242e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=2.285 $X2=6.415 $Y2=2.555
r160 1 38 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.595 $X2=6.31 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_835_93# 1 2 7 9 10 12 14 15 16 17 18 21
+ 25 27 32 33 34 36 39 41 44 47 48 49 50 53 55 59 61 70
c189 70 0 9.23744e-20 $X=5.115 $Y=1.61
c190 55 0 1.88382e-19 $X=4.895 $Y=1.95
c191 39 0 2.96321e-20 $X=9.785 $Y=0.58
c192 33 0 1.09841e-19 $X=9.625 $Y=1.585
c193 21 0 1.51838e-20 $X=6.095 $Y=0.805
c194 16 0 1.72525e-19 $X=5.69 $Y=3.15
r195 71 73 2.03376 $w=4.74e-07 $l=2e-08 $layer=POLY_cond $X=5.115 $Y=1.517
+ $X2=5.095 $Y2=1.517
r196 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.61 $X2=5.115 $Y2=1.61
r197 61 64 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=4.46 $Y=2.06 $X2=4.46
+ $Y2=2.12
r198 57 59 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=4.32 $Y=0.625
+ $X2=4.45 $Y2=0.625
r199 54 66 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=4.895 $Y=1.8
+ $X2=4.895 $Y2=1.622
r200 54 55 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.895 $Y=1.8
+ $X2=4.895 $Y2=1.95
r201 53 70 6.10308 $w=3.53e-07 $l=1.88e-07 $layer=LI1_cond $X=4.927 $Y=1.622
+ $X2=5.115 $Y2=1.622
r202 53 66 1.03882 $w=3.53e-07 $l=3.2e-08 $layer=LI1_cond $X=4.927 $Y=1.622
+ $X2=4.895 $Y2=1.622
r203 52 53 17.4092 $w=2.33e-07 $l=3.55e-07 $layer=LI1_cond $X=4.927 $Y=1.09
+ $X2=4.927 $Y2=1.445
r204 51 61 1.48468 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=2.06
+ $X2=4.46 $Y2=2.06
r205 50 55 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.81 $Y=2.06
+ $X2=4.895 $Y2=1.95
r206 50 51 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=4.81 $Y=2.06
+ $X2=4.585 $Y2=2.06
r207 48 52 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.927 $Y2=1.09
r208 48 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.535 $Y2=1.005
r209 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=0.92
+ $X2=4.535 $Y2=1.005
r210 46 59 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.625
r211 46 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.92
r212 42 44 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=9.7 $Y=1.045
+ $X2=9.785 $Y2=1.045
r213 37 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.785 $Y=0.97
+ $X2=9.785 $Y2=1.045
r214 37 39 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.785 $Y=0.97
+ $X2=9.785 $Y2=0.58
r215 35 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.7 $Y=1.12 $X2=9.7
+ $Y2=1.045
r216 35 36 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.7 $Y=1.12 $X2=9.7
+ $Y2=1.51
r217 33 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.7 $Y2=1.51
r218 33 34 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.235 $Y2=1.585
r219 30 32 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=9.145 $Y=3.075
+ $X2=9.145 $Y2=2.235
r220 29 34 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.145 $Y=1.66
+ $X2=9.235 $Y2=1.585
r221 29 32 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.145 $Y=1.66
+ $X2=9.145 $Y2=2.235
r222 28 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.73 $Y=3.15 $X2=6.64
+ $Y2=3.15
r223 27 30 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.055 $Y=3.15
+ $X2=9.145 $Y2=3.075
r224 27 28 1192.18 $w=1.5e-07 $l=2.325e-06 $layer=POLY_cond $X=9.055 $Y=3.15
+ $X2=6.73 $Y2=3.15
r225 23 41 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.64 $Y=3.075
+ $X2=6.64 $Y2=3.15
r226 23 25 217.677 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=6.64 $Y=3.075
+ $X2=6.64 $Y2=2.515
r227 19 21 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.095 $Y=1.185
+ $X2=6.095 $Y2=0.805
r228 18 76 34.1471 $w=4.74e-07 $l=3.00772e-07 $layer=POLY_cond $X=5.71 $Y=1.26
+ $X2=5.615 $Y2=1.517
r229 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.02 $Y=1.26
+ $X2=6.095 $Y2=1.185
r230 17 18 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.02 $Y=1.26
+ $X2=5.71 $Y2=1.26
r231 15 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=3.15 $X2=6.64
+ $Y2=3.15
r232 15 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.55 $Y=3.15
+ $X2=5.69 $Y2=3.15
r233 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r234 13 76 30.0642 $w=1.5e-07 $l=3.33e-07 $layer=POLY_cond $X=5.615 $Y=1.85
+ $X2=5.615 $Y2=1.517
r235 13 14 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=5.615 $Y=1.85
+ $X2=5.615 $Y2=3.075
r236 10 76 47.7932 $w=4.74e-07 $l=4.7e-07 $layer=POLY_cond $X=5.145 $Y=1.517
+ $X2=5.615 $Y2=1.517
r237 10 71 3.05063 $w=4.74e-07 $l=3e-08 $layer=POLY_cond $X=5.145 $Y=1.517
+ $X2=5.115 $Y2=1.517
r238 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.145 $Y=1.41
+ $X2=5.145 $Y2=0.965
r239 7 73 25.5547 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=5.095 $Y=1.85
+ $X2=5.095 $Y2=1.517
r240 7 9 172.717 $w=1.8e-07 $l=6.45e-07 $layer=POLY_cond $X=5.095 $Y=1.85
+ $X2=5.095 $Y2=2.495
r241 2 64 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.935 $X2=4.42 $Y2=2.12
r242 1 57 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.465 $X2=4.32 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_1997_272# 1 2 9 11 13 15 19 23 25 26 28
+ 33 35 36 38
c110 33 0 6.31244e-20 $X=10.315 $Y=1.525
c111 28 0 1.53844e-19 $X=11.65 $Y=1.445
c112 15 0 6.72618e-20 $X=11.14 $Y=1.53
r113 35 36 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=11.127 $Y=2.75
+ $X2=11.127 $Y2=2.52
r114 30 33 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=1.525
+ $X2=10.315 $Y2=1.525
r115 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.15
+ $Y=1.525 $X2=10.15 $Y2=1.525
r116 27 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.65 $Y=0.925
+ $X2=11.65 $Y2=1.445
r117 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.65 $Y2=0.925
r118 25 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.565 $Y=0.84
+ $X2=11.34 $Y2=0.84
r119 24 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.31 $Y=1.53
+ $X2=11.225 $Y2=1.53
r120 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.565 $Y=1.53
+ $X2=11.65 $Y2=1.445
r121 23 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.565 $Y=1.53
+ $X2=11.31 $Y2=1.53
r122 21 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.225 $Y=1.615
+ $X2=11.225 $Y2=1.53
r123 21 36 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.225 $Y=1.615
+ $X2=11.225 $Y2=2.52
r124 17 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.175 $Y=0.755
+ $X2=11.34 $Y2=0.84
r125 17 19 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=11.175 $Y=0.755
+ $X2=11.175 $Y2=0.58
r126 15 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.14 $Y=1.53
+ $X2=11.225 $Y2=1.53
r127 15 33 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=11.14 $Y=1.53
+ $X2=10.315 $Y2=1.53
r128 11 31 58.2622 $w=3e-07 $l=3.69317e-07 $layer=POLY_cond $X=10.31 $Y=1.84
+ $X2=10.192 $Y2=1.525
r129 11 13 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=10.31 $Y=1.84
+ $X2=10.31 $Y2=2.75
r130 7 31 38.5519 $w=3e-07 $l=1.87029e-07 $layer=POLY_cond $X=10.145 $Y=1.36
+ $X2=10.192 $Y2=1.525
r131 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=10.145 $Y=1.36
+ $X2=10.145 $Y2=0.58
r132 2 35 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=10.975
+ $Y=2.54 $X2=11.11 $Y2=2.75
r133 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.37 $X2=11.175 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_1745_74# 1 2 9 12 15 17 18 19 23 27 29 30
+ 35 37 40 41 43 45 48 50 52
c157 50 0 5.21422e-20 $X=11.23 $Y=1.185
c158 43 0 1.04043e-19 $X=10.23 $Y=2.55
c159 12 0 1.53844e-19 $X=11.32 $Y=1.84
r160 51 56 13.6415 $w=3.18e-07 $l=9e-08 $layer=POLY_cond $X=11.23 $Y=1.145
+ $X2=11.32 $Y2=1.145
r161 50 52 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=11.23 $Y=1.185
+ $X2=11.065 $Y2=1.185
r162 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.23
+ $Y=1.185 $X2=11.23 $Y2=1.185
r163 45 47 9.9702 $w=3.48e-07 $l=2.1e-07 $layer=LI1_cond $X=9.58 $Y=0.56
+ $X2=9.58 $Y2=0.77
r164 42 43 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.23 $Y=1.955
+ $X2=10.23 $Y2=2.55
r165 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=1.87
+ $X2=10.23 $Y2=1.955
r166 40 41 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.145 $Y=1.87
+ $X2=9.755 $Y2=1.87
r167 39 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.755 $Y=1.18
+ $X2=9.67 $Y2=1.18
r168 39 52 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=9.755 $Y=1.18
+ $X2=11.065 $Y2=1.18
r169 37 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.67 $Y=1.785
+ $X2=9.755 $Y2=1.87
r170 36 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.265
+ $X2=9.67 $Y2=1.18
r171 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.67 $Y=1.265
+ $X2=9.67 $Y2=1.785
r172 35 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.67 $Y2=1.18
r173 35 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.67 $Y2=0.77
r174 30 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.145 $Y=2.715
+ $X2=10.23 $Y2=2.55
r175 30 32 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=10.145 $Y=2.715
+ $X2=9.56 $Y2=2.715
r176 25 27 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=11.955 $Y=1.2
+ $X2=11.955 $Y2=0.645
r177 21 23 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=11.92 $Y=1.99
+ $X2=11.92 $Y2=2.54
r178 20 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.425 $Y=1.915
+ $X2=11.335 $Y2=1.915
r179 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.83 $Y=1.915
+ $X2=11.92 $Y2=1.99
r180 19 20 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=11.83 $Y=1.915
+ $X2=11.425 $Y2=1.915
r181 18 56 24.9017 $w=3.18e-07 $l=1.63248e-07 $layer=POLY_cond $X=11.395
+ $Y=1.275 $X2=11.32 $Y2=1.145
r182 17 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.88 $Y=1.275
+ $X2=11.955 $Y2=1.2
r183 17 18 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.88 $Y=1.275
+ $X2=11.395 $Y2=1.275
r184 13 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.335 $Y=1.99
+ $X2=11.335 $Y2=1.915
r185 13 15 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=11.335 $Y=1.99
+ $X2=11.335 $Y2=2.75
r186 12 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.32 $Y=1.84
+ $X2=11.335 $Y2=1.915
r187 11 56 20.3436 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=11.32 $Y=1.35
+ $X2=11.32 $Y2=1.145
r188 11 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=11.32 $Y=1.35
+ $X2=11.32 $Y2=1.84
r189 7 51 40.9245 $w=3.18e-07 $l=3.5812e-07 $layer=POLY_cond $X=10.96 $Y=0.94
+ $X2=11.23 $Y2=1.145
r190 7 9 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.96 $Y=0.94
+ $X2=10.96 $Y2=0.58
r191 2 32 600 $w=1.7e-07 $l=1.13088e-06 $layer=licon1_PDIFF $count=1 $X=9.235
+ $Y=1.735 $X2=9.56 $Y2=2.715
r192 1 45 182 $w=1.7e-07 $l=9.35187e-07 $layer=licon1_NDIFF $count=1 $X=8.725
+ $Y=0.37 $X2=9.57 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_2402_424# 1 2 9 13 15 16 19 23 29 32 33
r45 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.745
+ $Y=1.465 $X2=12.745 $Y2=1.465
r46 27 33 0.189605 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.335 $Y=1.465
+ $X2=12.21 $Y2=1.465
r47 27 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.335 $Y=1.465
+ $X2=12.745 $Y2=1.465
r48 25 33 6.72893 $w=2.37e-07 $l=1.71377e-07 $layer=LI1_cond $X=12.197 $Y=1.63
+ $X2=12.21 $Y2=1.465
r49 25 32 24.0733 $w=2.23e-07 $l=4.7e-07 $layer=LI1_cond $X=12.197 $Y=1.63
+ $X2=12.197 $Y2=2.1
r50 21 33 6.72893 $w=2.37e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=1.3
+ $X2=12.21 $Y2=1.465
r51 21 23 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=12.21 $Y=1.3
+ $X2=12.21 $Y2=0.645
r52 19 32 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.145 $Y=2.265
+ $X2=12.145 $Y2=2.1
r53 15 30 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=12.84 $Y=1.465
+ $X2=12.745 $Y2=1.465
r54 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.84 $Y=1.465
+ $X2=12.93 $Y2=1.465
r55 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.945 $Y=1.3
+ $X2=12.93 $Y2=1.465
r56 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.945 $Y=1.3
+ $X2=12.945 $Y2=0.74
r57 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=12.93 $Y=1.63
+ $X2=12.93 $Y2=1.465
r58 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=12.93 $Y=1.63
+ $X2=12.93 $Y2=2.4
r59 2 19 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.01
+ $Y=2.12 $X2=12.145 $Y2=2.265
r60 1 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=12.03
+ $Y=0.37 $X2=12.17 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 41 45 51
+ 55 61 66 67 69 70 72 73 74 76 81 93 110 116 117 120 123 126 129 132
c161 35 0 1.72525e-19 $X=4.87 $Y=2.885
c162 3 0 1.88382e-19 $X=4.735 $Y=1.935
c163 2 0 1.1782e-19 $X=3.125 $Y=2.32
r164 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r165 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r166 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r167 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r168 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r169 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 117 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r171 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r172 114 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.87 $Y=3.33
+ $X2=12.705 $Y2=3.33
r173 114 116 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=12.87 $Y=3.33
+ $X2=13.2 $Y2=3.33
r174 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r176 110 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.705 $Y2=3.33
r177 110 112 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.24 $Y2=3.33
r178 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r179 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r180 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r181 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r182 103 106 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r183 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r184 102 105 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r185 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r186 100 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.47 $Y2=3.33
r187 100 102 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.88 $Y2=3.33
r188 99 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r189 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r190 95 98 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r191 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r192 93 126 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.372 $Y2=3.33
r193 93 98 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=6.96 $Y2=3.33
r194 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r195 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r196 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r197 89 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r198 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r199 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r200 86 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r201 86 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r202 85 124 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r203 85 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r205 82 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r206 82 84 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r207 81 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r208 81 84 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r209 79 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r210 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r211 76 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r212 76 78 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r213 74 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r214 74 96 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=5.04 $Y2=3.33
r215 72 108 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.28 $Y2=3.33
r216 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.645 $Y2=3.33
r217 71 112 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=11.81 $Y=3.33
+ $X2=12.24 $Y2=3.33
r218 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.81 $Y=3.33
+ $X2=11.645 $Y2=3.33
r219 69 105 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.32 $Y2=3.33
r220 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.485 $Y=3.33
+ $X2=10.61 $Y2=3.33
r221 68 108 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.735 $Y=3.33
+ $X2=11.28 $Y2=3.33
r222 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.735 $Y=3.33
+ $X2=10.61 $Y2=3.33
r223 66 91 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r224 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r225 65 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r226 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r227 61 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.705 $Y=1.985
+ $X2=12.705 $Y2=2.815
r228 59 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.705 $Y=3.245
+ $X2=12.705 $Y2=3.33
r229 59 64 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.705 $Y=3.245
+ $X2=12.705 $Y2=2.815
r230 55 58 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=11.645 $Y=2.265
+ $X2=11.645 $Y2=2.815
r231 53 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.645 $Y=3.245
+ $X2=11.645 $Y2=3.33
r232 53 58 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.645 $Y=3.245
+ $X2=11.645 $Y2=2.815
r233 49 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.61 $Y=3.245
+ $X2=10.61 $Y2=3.33
r234 49 51 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=10.61 $Y=3.245
+ $X2=10.61 $Y2=2.75
r235 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.47 $Y=1.91
+ $X2=8.47 $Y2=2.59
r236 43 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.47 $Y=3.245
+ $X2=8.47 $Y2=3.33
r237 43 48 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.47 $Y=3.245
+ $X2=8.47 $Y2=2.59
r238 42 126 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.372 $Y2=3.33
r239 41 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=3.33
+ $X2=8.47 $Y2=3.33
r240 41 42 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.385 $Y=3.33
+ $X2=7.54 $Y2=3.33
r241 37 126 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.372 $Y=3.245
+ $X2=7.372 $Y2=3.33
r242 37 39 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.372 $Y=3.245
+ $X2=7.372 $Y2=2.825
r243 33 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r244 33 35 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.885
r245 29 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r246 29 31 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.79
r247 25 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r248 25 27 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.465
r249 8 64 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=12.56
+ $Y=1.84 $X2=12.705 $Y2=2.815
r250 8 61 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.56
+ $Y=1.84 $X2=12.705 $Y2=1.985
r251 7 58 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=11.425
+ $Y=2.54 $X2=11.645 $Y2=2.815
r252 7 55 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=11.425
+ $Y=2.54 $X2=11.645 $Y2=2.265
r253 6 51 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=10.4
+ $Y=2.54 $X2=10.57 $Y2=2.75
r254 5 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.735 $X2=8.47 $Y2=2.59
r255 5 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.735 $X2=8.47 $Y2=1.91
r256 4 39 600 $w=1.7e-07 $l=6.20323e-07 $layer=licon1_PDIFF $count=1 $X=7.15
+ $Y=2.305 $X2=7.37 $Y2=2.825
r257 3 35 600 $w=1.7e-07 $l=1.01526e-06 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=1.935 $X2=4.87 $Y2=2.885
r258 2 31 600 $w=1.7e-07 $l=5.33245e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=2.32 $X2=3.26 $Y2=2.79
r259 1 27 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.32 $X2=0.78 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%A_303_464# 1 2 3 4 5 16 20 22 25 28 29 32
+ 35 37 38 39 40 41 43 46 48 54 55
c163 54 0 9.0609e-20 $X=3.83 $Y=2.475
c164 40 0 1.29298e-19 $X=6.37 $Y=2.13
c165 38 0 1.55517e-19 $X=6.37 $Y=1.285
c166 35 0 6.25949e-20 $X=5.887 $Y=1.2
c167 25 0 1.1782e-19 $X=3.53 $Y=2.33
r168 52 54 15.8442 $w=2.31e-07 $l=3e-07 $layer=LI1_cond $X=3.53 $Y=2.48 $X2=3.83
+ $Y2=2.48
r169 48 50 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=0.68
+ $X2=2.435 $Y2=1.005
r170 45 46 11.0435 $w=6.33e-07 $l=2e-07 $layer=LI1_cond $X=2.355 $Y=2.662
+ $X2=2.555 $Y2=2.662
r171 42 43 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.455 $Y=1.37
+ $X2=6.455 $Y2=2.045
r172 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=2.13
+ $X2=6.455 $Y2=2.045
r173 40 41 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=2.13
+ $X2=6.075 $Y2=2.13
r174 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=1.285
+ $X2=6.455 $Y2=1.37
r175 38 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.37 $Y=1.285
+ $X2=5.975 $Y2=1.285
r176 37 57 3.11038 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=5.95 $Y=2.455
+ $X2=5.95 $Y2=2.59
r177 36 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=6.075 $Y2=2.13
r178 36 37 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=5.95 $Y=2.215
+ $X2=5.95 $Y2=2.455
r179 35 39 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.975 $Y2=1.285
r180 35 55 10.4571 $w=1.73e-07 $l=1.65e-07 $layer=LI1_cond $X=5.887 $Y=1.2
+ $X2=5.887 $Y2=1.035
r181 30 55 5.54545 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=5.885 $Y=0.945
+ $X2=5.885 $Y2=1.035
r182 30 32 8.31818 $w=1.78e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=0.945
+ $X2=5.885 $Y2=0.81
r183 29 54 9.46026 $w=2.31e-07 $l=1.93533e-07 $layer=LI1_cond $X=3.995 $Y=2.542
+ $X2=3.83 $Y2=2.48
r184 28 57 3.98589 $w=1.75e-07 $l=1.47054e-07 $layer=LI1_cond $X=5.825 $Y=2.542
+ $X2=5.95 $Y2=2.59
r185 28 29 115.979 $w=1.73e-07 $l=1.83e-06 $layer=LI1_cond $X=5.825 $Y=2.542
+ $X2=3.995 $Y2=2.542
r186 25 52 2.5345 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.53 $Y=2.33 $X2=3.53
+ $Y2=2.48
r187 24 25 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.33
r188 23 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=1.005
+ $X2=2.435 $Y2=1.005
r189 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r190 22 23 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.6 $Y2=1.005
r191 20 52 5.36393 $w=2.31e-07 $l=1.07121e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.53 $Y2=2.48
r192 20 46 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.555 $Y2=2.43
r193 16 45 2.2038 $w=6.33e-07 $l=1.17e-07 $layer=LI1_cond $X=2.238 $Y=2.662
+ $X2=2.355 $Y2=2.662
r194 16 18 11.0755 $w=6.33e-07 $l=5.88e-07 $layer=LI1_cond $X=2.238 $Y=2.662
+ $X2=1.65 $Y2=2.662
r195 5 57 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r196 4 54 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=3.695
+ $Y=2.32 $X2=3.83 $Y2=2.475
r197 3 45 200 $w=1.7e-07 $l=9.09615e-07 $layer=licon1_PDIFF $count=3 $X=1.515
+ $Y=2.32 $X2=2.355 $Y2=2.465
r198 3 18 200 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=3 $X=1.515
+ $Y=2.32 $X2=1.65 $Y2=2.465
r199 2 32 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=5.755
+ $Y=0.595 $X2=5.88 $Y2=0.81
r200 1 48 182 $w=1.7e-07 $l=6.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.405 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%Q 1 2 7 8 9 10 11 12 13 29
r14 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=13.16 $Y=0.965
+ $X2=13.16 $Y2=0.925
r15 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=13.197 $Y=2.405
+ $X2=13.197 $Y2=2.775
r16 11 12 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=13.197 $Y=1.985
+ $X2=13.197 $Y2=2.405
r17 10 11 14.462 $w=2.53e-07 $l=3.2e-07 $layer=LI1_cond $X=13.197 $Y=1.665
+ $X2=13.197 $Y2=1.985
r18 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=13.197 $Y=1.295
+ $X2=13.197 $Y2=1.665
r19 9 45 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=13.197 $Y=1.295
+ $X2=13.197 $Y2=1.13
r20 8 45 5.6192 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=13.16 $Y=0.987
+ $X2=13.16 $Y2=1.13
r21 8 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=13.16 $Y=0.987
+ $X2=13.16 $Y2=0.965
r22 8 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=13.16 $Y=0.902
+ $X2=13.16 $Y2=0.925
r23 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=13.16 $Y=0.515
+ $X2=13.16 $Y2=0.902
r24 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.84 $X2=13.155 $Y2=2.815
r25 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.84 $X2=13.155 $Y2=1.985
r26 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.02
+ $Y=0.37 $X2=13.16 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 47 48
+ 49 51 56 65 69 77 82 89 90 93 96 100 106 109 112
c132 90 0 7.12888e-20 $X=13.2 $Y=0
c133 28 0 1.58089e-19 $X=3.715 $Y=0.565
r134 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r135 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r136 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r137 100 103 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r138 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r139 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r140 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r141 90 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r142 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r143 87 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=12.69 $Y2=0
r144 87 89 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.815 $Y=0
+ $X2=13.2 $Y2=0
r145 86 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r146 86 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r147 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r148 83 109 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=11.737 $Y2=0
r149 83 85 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.905 $Y=0
+ $X2=12.24 $Y2=0
r150 82 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.565 $Y=0
+ $X2=12.69 $Y2=0
r151 82 85 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.565 $Y=0
+ $X2=12.24 $Y2=0
r152 81 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r153 81 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r154 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r155 78 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.525 $Y=0
+ $X2=10.36 $Y2=0
r156 78 80 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=10.525 $Y=0
+ $X2=11.28 $Y2=0
r157 77 109 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.737 $Y2=0
r158 77 80 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.57 $Y=0
+ $X2=11.28 $Y2=0
r159 76 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r160 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r161 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r162 73 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r163 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r164 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r165 70 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r166 70 72 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r167 69 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=10.36 $Y2=0
r168 69 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=9.84 $Y2=0
r169 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r170 65 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r171 65 67 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=7.43 $Y=0 $X2=5.04
+ $Y2=0
r172 64 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r173 64 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r174 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r175 61 96 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.735
+ $Y2=0
r176 61 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.56
+ $Y2=0
r177 60 97 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r178 60 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r179 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r180 57 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r181 57 59 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r182 56 96 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.735
+ $Y2=0
r183 56 59 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=3.59 $Y=0 $X2=1.2
+ $Y2=0
r184 54 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r185 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r186 51 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r187 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r188 49 101 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=7.44 $Y2=0
r189 49 68 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=5.04 $Y2=0
r190 47 63 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r191 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r192 46 67 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r193 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r194 42 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.69 $Y=0.085
+ $X2=12.69 $Y2=0
r195 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.69 $Y=0.085
+ $X2=12.69 $Y2=0.515
r196 38 109 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=11.737 $Y=0.085
+ $X2=11.737 $Y2=0
r197 38 40 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=11.737 $Y=0.085
+ $X2=11.737 $Y2=0.5
r198 34 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0
r199 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0.58
r200 30 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r201 30 32 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.665
r202 26 96 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0
r203 26 28 19.0749 $w=2.88e-07 $l=4.8e-07 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0.565
r204 22 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r205 22 24 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.65
r206 7 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.585
+ $Y=0.37 $X2=12.73 $Y2=0.515
r207 6 40 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=11.59
+ $Y=0.37 $X2=11.735 $Y2=0.5
r208 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.22
+ $Y=0.37 $X2=10.36 $Y2=0.58
r209 4 103 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.595 $X2=7.595 $Y2=0.325
r210 3 32 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.595 $X2=4.87 $Y2=0.665
r211 2 28 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.405 $X2=3.715 $Y2=0.565
r212 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.44 $X2=0.71 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_1%noxref_24 1 2 7 9 14
r32 14 17 7.40856 $w=3.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.235 $Y=0.34
+ $X2=3.235 $Y2=0.565
r33 9 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34 $X2=1.27
+ $Y2=0.55
r34 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34 $X2=1.27
+ $Y2=0.34
r35 7 14 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.06 $Y=0.34 $X2=3.235
+ $Y2=0.34
r36 7 8 106.016 $w=1.68e-07 $l=1.625e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.435 $Y2=0.34
r37 2 17 182 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.405 $X2=3.265 $Y2=0.565
r38 1 12 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends


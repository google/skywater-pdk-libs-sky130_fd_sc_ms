# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a2bb2oi_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__a2bb2oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.262500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.260000 0.435000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.262500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.450000 1.100000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.220000 1.220000 2.755000 1.540000 ;
        RECT 2.525000 1.540000 2.755000 2.150000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.498400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 2.290000 1.780000 2.980000 ;
        RECT 1.610000 1.750000 2.050000 1.920000 ;
        RECT 1.610000 1.920000 2.275000 2.220000 ;
        RECT 1.610000 2.220000 1.780000 2.290000 ;
        RECT 1.880000 0.880000 2.315000 1.050000 ;
        RECT 1.880000 1.050000 2.050000 1.750000 ;
        RECT 2.055000 0.350000 2.315000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.120000  1.950000 0.450000 3.245000 ;
      RECT 0.175000  0.085000 0.425000 1.090000 ;
      RECT 0.605000  0.540000 0.935000 0.960000 ;
      RECT 0.605000  0.960000 1.440000 1.130000 ;
      RECT 0.960000  1.950000 1.440000 2.120000 ;
      RECT 0.960000  2.120000 1.290000 2.980000 ;
      RECT 1.105000  0.085000 1.885000 0.710000 ;
      RECT 1.105000  0.710000 1.710000 0.790000 ;
      RECT 1.270000  1.130000 1.440000 1.220000 ;
      RECT 1.270000  1.220000 1.710000 1.550000 ;
      RECT 1.270000  1.550000 1.440000 1.950000 ;
      RECT 1.980000  2.390000 3.240000 2.560000 ;
      RECT 1.980000  2.560000 2.230000 2.980000 ;
      RECT 2.430000  2.730000 2.790000 2.980000 ;
      RECT 2.430000  2.980000 2.600000 3.245000 ;
      RECT 2.885000  0.085000 3.215000 1.010000 ;
      RECT 2.990000  1.820000 3.240000 2.390000 ;
      RECT 2.990000  2.560000 3.240000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ms__a2bb2oi_1

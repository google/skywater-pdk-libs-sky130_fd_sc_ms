* File: sky130_fd_sc_ms__nand2_2.pxi.spice
* Created: Wed Sep  2 12:12:48 2020
* 
x_PM_SKY130_FD_SC_MS__NAND2_2%B N_B_M1005_g N_B_M1000_g N_B_M1001_g N_B_M1007_g
+ B B N_B_c_48_n PM_SKY130_FD_SC_MS__NAND2_2%B
x_PM_SKY130_FD_SC_MS__NAND2_2%A N_A_M1002_g N_A_M1004_g N_A_M1006_g N_A_M1003_g
+ A N_A_c_86_n N_A_c_87_n PM_SKY130_FD_SC_MS__NAND2_2%A
x_PM_SKY130_FD_SC_MS__NAND2_2%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_M1006_s
+ N_VPWR_c_130_n N_VPWR_c_131_n N_VPWR_c_132_n N_VPWR_c_133_n N_VPWR_c_134_n
+ VPWR N_VPWR_c_135_n N_VPWR_c_136_n N_VPWR_c_137_n N_VPWR_c_129_n
+ PM_SKY130_FD_SC_MS__NAND2_2%VPWR
x_PM_SKY130_FD_SC_MS__NAND2_2%Y N_Y_M1002_d N_Y_M1000_d N_Y_M1004_d N_Y_c_175_n
+ N_Y_c_171_n N_Y_c_179_n N_Y_c_183_n N_Y_c_172_n N_Y_c_173_n N_Y_c_168_n
+ N_Y_c_169_n N_Y_c_191_n Y Y PM_SKY130_FD_SC_MS__NAND2_2%Y
x_PM_SKY130_FD_SC_MS__NAND2_2%A_27_74# N_A_27_74#_M1005_d N_A_27_74#_M1007_d
+ N_A_27_74#_M1003_s N_A_27_74#_c_214_n N_A_27_74#_c_215_n N_A_27_74#_c_216_n
+ N_A_27_74#_c_217_n N_A_27_74#_c_218_n N_A_27_74#_c_219_n
+ PM_SKY130_FD_SC_MS__NAND2_2%A_27_74#
x_PM_SKY130_FD_SC_MS__NAND2_2%VGND N_VGND_M1005_s N_VGND_c_248_n VGND
+ N_VGND_c_249_n N_VGND_c_250_n N_VGND_c_251_n N_VGND_c_252_n
+ PM_SKY130_FD_SC_MS__NAND2_2%VGND
cc_1 VNB N_B_M1005_g 0.0325972f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B_M1007_g 0.0243544f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_3 VNB B 0.00631699f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B_c_48_n 0.0454861f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.515
cc_5 VNB N_A_M1002_g 0.0236545f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_A_M1003_g 0.0267831f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_7 VNB N_A_c_86_n 0.00139482f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_8 VNB N_A_c_87_n 0.0387686f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_9 VNB N_VPWR_c_129_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_Y_c_168_n 0.0105096f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_11 VNB N_Y_c_169_n 0.0025404f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.515
cc_12 VNB Y 0.0241052f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_13 VNB N_A_27_74#_c_214_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_215_n 0.00790826f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_15 VNB N_A_27_74#_c_216_n 0.0116953f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_16 VNB N_A_27_74#_c_217_n 0.0126678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_218_n 0.00217191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_18 VNB N_A_27_74#_c_219_n 0.0161735f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_19 VNB N_VGND_c_248_n 0.00615265f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_20 VNB N_VGND_c_249_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_21 VNB N_VGND_c_250_n 0.0392768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_251_n 0.163114f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_23 VNB N_VGND_c_252_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_24 VPB N_B_M1000_g 0.0263926f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_25 VPB N_B_M1001_g 0.0201415f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_26 VPB B 0.00702098f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_27 VPB N_B_c_48_n 0.0052668f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.515
cc_28 VPB N_A_M1004_g 0.0207341f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_29 VPB N_A_M1006_g 0.0230837f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_30 VPB N_A_c_86_n 0.00251251f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_31 VPB N_A_c_87_n 0.00479899f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_32 VPB N_VPWR_c_130_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_33 VPB N_VPWR_c_131_n 0.0579545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_132_n 0.00273118f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_35 VPB N_VPWR_c_133_n 0.0127942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_134_n 0.0348965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_135_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_38 VPB N_VPWR_c_136_n 0.0167647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_137_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_129_n 0.0572022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_Y_c_171_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_172_n 0.00179776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_Y_c_173_n 0.00793272f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_44 VPB Y 0.0130636f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_45 N_B_M1007_g N_A_M1002_g 0.0220064f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_46 N_B_M1001_g N_A_M1004_g 0.0220064f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_47 B N_A_c_86_n 0.0361808f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_48 N_B_c_48_n N_A_c_86_n 2.85035e-19 $X=0.975 $Y=1.515 $X2=0 $Y2=0
cc_49 B N_A_c_87_n 0.00435599f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_50 N_B_c_48_n N_A_c_87_n 0.0220064f $X=0.975 $Y=1.515 $X2=0 $Y2=0
cc_51 N_B_M1000_g N_VPWR_c_131_n 0.00551672f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_52 N_B_M1000_g N_VPWR_c_132_n 5.60169e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_53 N_B_M1001_g N_VPWR_c_132_n 0.0129287f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_54 N_B_M1000_g N_VPWR_c_135_n 0.005209f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_55 N_B_M1001_g N_VPWR_c_135_n 0.00460063f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_56 N_B_M1000_g N_VPWR_c_129_n 0.00986025f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_57 N_B_M1001_g N_VPWR_c_129_n 0.00908554f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_58 N_B_M1000_g N_Y_c_175_n 0.00364186f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_59 B N_Y_c_175_n 0.0163574f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_60 N_B_c_48_n N_Y_c_175_n 5.54777e-19 $X=0.975 $Y=1.515 $X2=0 $Y2=0
cc_61 N_B_M1000_g N_Y_c_171_n 0.0112102f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_62 N_B_M1001_g N_Y_c_179_n 0.0142777f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_63 B N_Y_c_179_n 0.0327785f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_64 N_B_M1005_g N_A_27_74#_c_214_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_65 N_B_M1005_g N_A_27_74#_c_215_n 0.0184659f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_66 N_B_M1007_g N_A_27_74#_c_215_n 0.013919f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_67 B N_A_27_74#_c_215_n 0.0533206f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_68 N_B_c_48_n N_A_27_74#_c_215_n 0.00359948f $X=0.975 $Y=1.515 $X2=0 $Y2=0
cc_69 N_B_M1007_g N_A_27_74#_c_218_n 0.00106427f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_70 N_B_M1005_g N_VGND_c_248_n 0.0132976f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_71 N_B_M1007_g N_VGND_c_248_n 0.00192886f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_VGND_c_249_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_73 N_B_M1007_g N_VGND_c_250_n 0.00461464f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_74 N_B_M1005_g N_VGND_c_251_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_75 N_B_M1007_g N_VGND_c_251_n 0.00908237f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A_M1004_g N_VPWR_c_132_n 0.0120681f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_VPWR_c_132_n 5.40311e-19 $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_VPWR_c_134_n 5.42556e-19 $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_VPWR_c_134_n 0.0139019f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_M1004_g N_VPWR_c_136_n 0.00490827f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A_M1006_g N_VPWR_c_136_n 0.00460063f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_VPWR_c_129_n 0.00968767f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_VPWR_c_129_n 0.00908554f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_M1004_g N_Y_c_179_n 0.0193471f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_c_86_n N_Y_c_179_n 0.00390336f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A_M1002_g N_Y_c_183_n 0.00543663f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A_M1006_g N_Y_c_173_n 0.0201893f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_c_86_n N_Y_c_173_n 0.00463673f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_Y_c_168_n 0.0178182f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_c_86_n N_Y_c_168_n 0.0021829f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_Y_c_169_n 0.00468846f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_c_86_n N_Y_c_169_n 0.0254953f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_93 N_A_c_87_n N_Y_c_169_n 0.00116051f $X=1.885 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A_c_86_n N_Y_c_191_n 0.0144665f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_95 N_A_c_87_n N_Y_c_191_n 5.53536e-19 $X=1.885 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_M1003_g Y 0.0252898f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_c_86_n Y 0.0263484f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A_M1002_g N_A_27_74#_c_215_n 5.7448e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_M1002_g N_A_27_74#_c_217_n 0.0122924f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_M1003_g N_A_27_74#_c_217_n 0.0121629f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_M1002_g N_A_27_74#_c_219_n 8.69012e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_M1003_g N_A_27_74#_c_219_n 0.00614869f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_VGND_c_250_n 0.00278271f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_M1003_g N_VGND_c_250_n 0.00278266f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_M1002_g N_VGND_c_251_n 0.00354005f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_M1003_g N_VGND_c_251_n 0.00357631f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_107 N_VPWR_c_131_n N_Y_c_171_n 0.0277973f $X=0.285 $Y=1.985 $X2=0 $Y2=0
cc_108 N_VPWR_c_132_n N_Y_c_171_n 0.0234083f $X=1.185 $Y=2.455 $X2=0 $Y2=0
cc_109 N_VPWR_c_135_n N_Y_c_171_n 0.0109793f $X=1.02 $Y=3.33 $X2=0 $Y2=0
cc_110 N_VPWR_c_129_n N_Y_c_171_n 0.00901959f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_111 N_VPWR_M1001_s N_Y_c_179_n 0.00353353f $X=1.05 $Y=1.84 $X2=0 $Y2=0
cc_112 N_VPWR_c_132_n N_Y_c_179_n 0.0170777f $X=1.185 $Y=2.455 $X2=0 $Y2=0
cc_113 N_VPWR_c_132_n N_Y_c_172_n 0.0224803f $X=1.185 $Y=2.455 $X2=0 $Y2=0
cc_114 N_VPWR_c_134_n N_Y_c_172_n 0.0233699f $X=2.095 $Y=2.455 $X2=0 $Y2=0
cc_115 N_VPWR_c_136_n N_Y_c_172_n 0.00749631f $X=1.93 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_c_129_n N_Y_c_172_n 0.0062048f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_117 N_VPWR_M1006_s N_Y_c_173_n 0.00440502f $X=1.96 $Y=1.84 $X2=0 $Y2=0
cc_118 N_VPWR_c_134_n N_Y_c_173_n 0.0237252f $X=2.095 $Y=2.455 $X2=0 $Y2=0
cc_119 N_VPWR_M1006_s Y 0.00185707f $X=1.96 $Y=1.84 $X2=0 $Y2=0
cc_120 N_VPWR_c_131_n N_A_27_74#_c_216_n 0.00901952f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_Y_c_168_n N_A_27_74#_M1003_s 0.00341347f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_122 N_Y_c_169_n N_A_27_74#_c_215_n 0.00997012f $X=1.785 $Y=1.095 $X2=0 $Y2=0
cc_123 N_Y_M1002_d N_A_27_74#_c_217_n 0.00229612f $X=1.48 $Y=0.37 $X2=0 $Y2=0
cc_124 N_Y_c_183_n N_A_27_74#_c_217_n 0.0179413f $X=1.62 $Y=0.86 $X2=0 $Y2=0
cc_125 N_Y_c_168_n N_A_27_74#_c_217_n 0.00352022f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_126 N_Y_c_168_n N_A_27_74#_c_219_n 0.0230579f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_127 N_A_27_74#_c_215_n N_VGND_M1005_s 0.00229612f $X=1.105 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_27_74#_c_214_n N_VGND_c_248_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_215_n N_VGND_c_248_n 0.0194017f $X=1.105 $Y=1.095 $X2=0
+ $Y2=0
cc_130 N_A_27_74#_c_218_n N_VGND_c_248_n 0.00814404f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
cc_131 N_A_27_74#_c_214_n N_VGND_c_249_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_217_n N_VGND_c_250_n 0.066264f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_133 N_A_27_74#_c_218_n N_VGND_c_250_n 0.0121867f $X=1.275 $Y=0.34 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_214_n N_VGND_c_251_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_c_217_n N_VGND_c_251_n 0.0369734f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_136 N_A_27_74#_c_218_n N_VGND_c_251_n 0.00660921f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0

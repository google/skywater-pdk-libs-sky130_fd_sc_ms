* File: sky130_fd_sc_ms__a221oi_1.pxi.spice
* Created: Fri Aug 28 17:01:07 2020
* 
x_PM_SKY130_FD_SC_MS__A221OI_1%C1 N_C1_M1009_g N_C1_M1003_g C1 N_C1_c_58_n
+ N_C1_c_59_n PM_SKY130_FD_SC_MS__A221OI_1%C1
x_PM_SKY130_FD_SC_MS__A221OI_1%B2 N_B2_M1001_g N_B2_M1008_g B2 B2 N_B2_c_86_n
+ PM_SKY130_FD_SC_MS__A221OI_1%B2
x_PM_SKY130_FD_SC_MS__A221OI_1%B1 N_B1_M1000_g N_B1_M1004_g B1 N_B1_c_120_n
+ N_B1_c_121_n PM_SKY130_FD_SC_MS__A221OI_1%B1
x_PM_SKY130_FD_SC_MS__A221OI_1%A1 N_A1_M1002_g N_A1_M1006_g A1 N_A1_c_159_n
+ N_A1_c_160_n PM_SKY130_FD_SC_MS__A221OI_1%A1
x_PM_SKY130_FD_SC_MS__A221OI_1%A2 N_A2_M1007_g N_A2_M1005_g A2 A2 N_A2_c_197_n
+ N_A2_c_198_n PM_SKY130_FD_SC_MS__A221OI_1%A2
x_PM_SKY130_FD_SC_MS__A221OI_1%Y N_Y_M1003_s N_Y_M1000_d N_Y_M1009_s N_Y_c_221_n
+ N_Y_c_222_n Y Y Y Y Y Y N_Y_c_224_n PM_SKY130_FD_SC_MS__A221OI_1%Y
x_PM_SKY130_FD_SC_MS__A221OI_1%A_121_368# N_A_121_368#_M1009_d
+ N_A_121_368#_M1001_d N_A_121_368#_c_258_n N_A_121_368#_c_259_n
+ N_A_121_368#_c_260_n N_A_121_368#_c_267_n
+ PM_SKY130_FD_SC_MS__A221OI_1%A_121_368#
x_PM_SKY130_FD_SC_MS__A221OI_1%A_263_368# N_A_263_368#_M1001_s
+ N_A_263_368#_M1004_d N_A_263_368#_M1005_d N_A_263_368#_c_284_n
+ N_A_263_368#_c_285_n N_A_263_368#_c_291_n N_A_263_368#_c_286_n
+ N_A_263_368#_c_300_n N_A_263_368#_c_287_n N_A_263_368#_c_288_n
+ N_A_263_368#_c_297_n PM_SKY130_FD_SC_MS__A221OI_1%A_263_368#
x_PM_SKY130_FD_SC_MS__A221OI_1%VPWR N_VPWR_M1002_d N_VPWR_c_327_n N_VPWR_c_328_n
+ N_VPWR_c_329_n VPWR N_VPWR_c_330_n N_VPWR_c_326_n
+ PM_SKY130_FD_SC_MS__A221OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A221OI_1%VGND N_VGND_M1003_d N_VGND_M1007_d N_VGND_c_360_n
+ N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n
+ VGND N_VGND_c_366_n N_VGND_c_367_n PM_SKY130_FD_SC_MS__A221OI_1%VGND
cc_1 VNB N_C1_M1003_g 0.031956f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_2 VNB N_C1_c_58_n 0.0539647f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_3 VNB N_C1_c_59_n 0.00305603f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_4 VNB N_B2_M1008_g 0.0236982f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_5 VNB B2 0.00423229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B2_c_86_n 0.0215552f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_7 VNB N_B1_M1000_g 0.0264675f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_8 VNB N_B1_c_120_n 0.0262382f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_9 VNB N_B1_c_121_n 0.00166531f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_10 VNB N_A1_M1006_g 0.0272859f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_11 VNB N_A1_c_159_n 0.0262677f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_12 VNB N_A1_c_160_n 0.00487854f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_13 VNB N_A2_M1005_g 0.00909003f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.74
cc_14 VNB A2 0.0422683f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_15 VNB N_A2_c_197_n 0.033324f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_16 VNB N_A2_c_198_n 0.0204958f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.515
cc_17 VNB N_Y_c_221_n 0.0208183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_222_n 0.00420435f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_19 VNB Y 0.0267465f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.665
cc_20 VNB N_Y_c_224_n 0.0616195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_326_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_360_n 0.00685096f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_VGND_c_361_n 0.0351314f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_24 VNB N_VGND_c_362_n 0.0347153f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_25 VNB N_VGND_c_363_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_364_n 0.0453999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_365_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_366_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_367_n 0.255119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_C1_M1009_g 0.0303189f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_31 VPB N_C1_c_58_n 0.0234117f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_32 VPB N_C1_c_59_n 0.00349083f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_33 VPB N_B2_M1001_g 0.0254389f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_34 VPB B2 0.0121355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_B2_c_86_n 0.0056176f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_36 VPB N_B1_M1004_g 0.0209374f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=0.74
cc_37 VPB N_B1_c_120_n 0.00559219f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_38 VPB N_B1_c_121_n 0.00265226f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_39 VPB N_A1_M1002_g 0.0223107f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_40 VPB N_A1_c_159_n 0.00561942f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_41 VPB N_A1_c_160_n 0.00246017f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_42 VPB N_A2_M1005_g 0.0326315f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=0.74
cc_43 VPB Y 0.0544483f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.665
cc_44 VPB N_A_121_368#_c_258_n 0.0126412f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_45 VPB N_A_121_368#_c_259_n 0.022676f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_46 VPB N_A_121_368#_c_260_n 0.00277569f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_47 VPB N_A_263_368#_c_284_n 0.00241504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_263_368#_c_285_n 0.00755847f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_49 VPB N_A_263_368#_c_286_n 0.0025292f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.665
cc_50 VPB N_A_263_368#_c_287_n 0.0150854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_263_368#_c_288_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_327_n 0.00678734f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=0.74
cc_53 VPB N_VPWR_c_328_n 0.0689094f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_54 VPB N_VPWR_c_329_n 0.00653059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_330_n 0.0255159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_326_n 0.0750005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 N_C1_M1003_g N_B2_M1008_g 0.026363f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_58 N_C1_M1009_g B2 4.41602e-19 $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_59 N_C1_c_58_n B2 0.015868f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_60 N_C1_c_59_n B2 0.0298996f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_61 N_C1_c_58_n N_B2_c_86_n 0.0205274f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_62 N_C1_M1003_g N_Y_c_221_n 0.0116701f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_63 N_C1_M1003_g Y 0.00356034f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_64 N_C1_c_58_n Y 0.0162941f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_65 N_C1_c_59_n Y 0.033251f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_66 N_C1_M1003_g N_Y_c_224_n 0.0140845f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_67 N_C1_c_58_n N_Y_c_224_n 0.0168615f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_68 N_C1_c_59_n N_Y_c_224_n 0.0281815f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_69 N_C1_M1009_g N_A_121_368#_c_258_n 0.0123512f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_70 N_C1_c_58_n N_A_121_368#_c_258_n 0.00263852f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_71 N_C1_c_59_n N_A_121_368#_c_258_n 0.0236659f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_72 N_C1_M1009_g N_A_121_368#_c_260_n 0.00841025f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_73 N_C1_M1009_g N_VPWR_c_328_n 0.00517089f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_74 N_C1_M1009_g N_VPWR_c_326_n 0.00987484f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_75 N_C1_M1003_g N_VGND_c_360_n 0.00601099f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_76 N_C1_M1003_g N_VGND_c_362_n 0.00433162f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_77 N_C1_M1003_g N_VGND_c_367_n 0.00822437f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_78 N_B2_M1008_g N_B1_M1000_g 0.0441025f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_79 N_B2_M1001_g N_B1_M1004_g 0.0340934f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_80 B2 N_B1_M1004_g 3.40762e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_81 B2 N_B1_c_120_n 0.00201442f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_82 N_B2_c_86_n N_B1_c_120_n 0.0441025f $X=1.59 $Y=1.515 $X2=0 $Y2=0
cc_83 N_B2_M1001_g N_B1_c_121_n 3.11382e-19 $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_84 B2 N_B1_c_121_n 0.0366307f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_85 N_B2_c_86_n N_B1_c_121_n 3.7859e-19 $X=1.59 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B2_M1008_g N_Y_c_221_n 0.0143728f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_87 N_B2_c_86_n N_Y_c_221_n 0.0041539f $X=1.59 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B2_M1008_g N_Y_c_224_n 9.00978e-19 $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_89 B2 N_Y_c_224_n 0.0544896f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_90 N_B2_M1001_g N_A_121_368#_c_258_n 0.00483849f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_91 N_B2_M1001_g N_A_121_368#_c_259_n 0.0156736f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_92 N_B2_M1001_g N_A_121_368#_c_267_n 0.0137194f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_93 B2 N_A_263_368#_c_284_n 0.0227263f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_94 N_B2_c_86_n N_A_263_368#_c_284_n 6.7198e-19 $X=1.59 $Y=1.515 $X2=0 $Y2=0
cc_95 N_B2_M1001_g N_A_263_368#_c_291_n 0.0142175f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_96 B2 N_A_263_368#_c_291_n 0.0161329f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_97 N_B2_M1001_g N_VPWR_c_328_n 0.00333896f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_98 N_B2_M1001_g N_VPWR_c_326_n 0.00427929f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_99 N_B2_M1008_g N_VGND_c_360_n 0.0141323f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B2_M1008_g N_VGND_c_364_n 0.00383152f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B2_M1008_g N_VGND_c_367_n 0.0075694f $X=1.68 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B1_M1004_g N_A1_M1002_g 0.0121812f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_103 N_B1_c_121_n N_A1_M1002_g 6.26118e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B1_M1000_g N_A1_M1006_g 0.0173199f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_105 N_B1_c_120_n N_A1_c_159_n 0.0201104f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_106 N_B1_c_121_n N_A1_c_159_n 0.00114936f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B1_c_120_n N_A1_c_160_n 0.00114936f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_c_121_n N_A1_c_160_n 0.0276388f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_109 N_B1_M1000_g N_Y_c_221_n 0.0154892f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_110 N_B1_c_120_n N_Y_c_221_n 0.00136713f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B1_c_121_n N_Y_c_221_n 0.0259226f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B1_M1000_g N_Y_c_222_n 0.00528753f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B1_M1004_g N_A_121_368#_c_259_n 0.00426321f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_114 N_B1_M1004_g N_A_121_368#_c_267_n 0.0082482f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_115 N_B1_M1004_g N_A_263_368#_c_291_n 0.0142101f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B1_c_120_n N_A_263_368#_c_291_n 2.14594e-19 $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_117 N_B1_c_121_n N_A_263_368#_c_291_n 0.0179862f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B1_M1004_g N_A_263_368#_c_286_n 2.32125e-19 $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_119 N_B1_c_120_n N_A_263_368#_c_297_n 2.22404e-19 $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_120 N_B1_c_121_n N_A_263_368#_c_297_n 0.00314801f $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_121 N_B1_M1004_g N_VPWR_c_327_n 5.19999e-19 $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B1_M1004_g N_VPWR_c_328_n 0.00517089f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B1_M1004_g N_VPWR_c_326_n 0.00979075f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B1_M1000_g N_VGND_c_360_n 0.00191029f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_125 N_B1_M1000_g N_VGND_c_364_n 0.00461464f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B1_M1000_g N_VGND_c_367_n 0.00910921f $X=2.04 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_M1002_g N_A2_M1005_g 0.0225279f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A1_c_160_n N_A2_M1005_g 0.00233713f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A1_M1006_g A2 0.00572702f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A1_c_160_n A2 0.0168427f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A1_c_159_n N_A2_c_197_n 0.0432818f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A1_c_160_n N_A2_c_197_n 0.00111347f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A1_M1006_g N_A2_c_198_n 0.0432818f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A1_M1006_g N_Y_c_221_n 0.00555347f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A1_c_159_n N_Y_c_221_n 5.39598e-19 $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A1_c_160_n N_Y_c_221_n 0.00595492f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A1_M1006_g N_Y_c_222_n 0.0103902f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A1_M1002_g N_A_121_368#_c_259_n 3.06664e-19 $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A1_M1002_g N_A_263_368#_c_286_n 2.42757e-19 $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A1_M1002_g N_A_263_368#_c_300_n 0.0153112f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A1_c_159_n N_A_263_368#_c_300_n 6.98124e-19 $X=2.67 $Y=1.515 $X2=0
+ $Y2=0
cc_142 N_A1_c_160_n N_A_263_368#_c_300_n 0.0229716f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A1_M1002_g N_A_263_368#_c_287_n 5.99214e-19 $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A1_M1002_g N_A_263_368#_c_288_n 7.56832e-19 $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A1_M1002_g N_VPWR_c_327_n 0.0113756f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A1_M1002_g N_VPWR_c_328_n 0.00521592f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A1_M1002_g N_VPWR_c_326_n 0.0102937f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A1_M1006_g N_VGND_c_361_n 0.00249753f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A1_M1006_g N_VGND_c_364_n 0.00461464f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A1_M1006_g N_VGND_c_367_n 0.00910921f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_A_263_368#_c_300_n 0.0146034f $X=3.135 $Y=2.4 $X2=0 $Y2=0
cc_152 A2 N_A_263_368#_c_300_n 0.00634715f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A2_M1005_g N_A_263_368#_c_287_n 0.00407495f $X=3.135 $Y=2.4 $X2=0 $Y2=0
cc_154 A2 N_A_263_368#_c_287_n 0.0203808f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_155 N_A2_c_197_n N_A_263_368#_c_287_n 0.00330449f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_156 N_A2_M1005_g N_A_263_368#_c_288_n 0.0129517f $X=3.135 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A2_M1005_g N_VPWR_c_327_n 0.00371878f $X=3.135 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A2_M1005_g N_VPWR_c_330_n 0.005209f $X=3.135 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A2_M1005_g N_VPWR_c_326_n 0.0098676f $X=3.135 $Y=2.4 $X2=0 $Y2=0
cc_160 A2 N_VGND_c_361_n 0.0259761f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A2_c_197_n N_VGND_c_361_n 0.0011179f $X=3.21 $Y=1.385 $X2=0 $Y2=0
cc_162 N_A2_c_198_n N_VGND_c_361_n 0.017286f $X=3.21 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A2_c_198_n N_VGND_c_364_n 0.00383152f $X=3.21 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A2_c_198_n N_VGND_c_367_n 0.0075694f $X=3.21 $Y=1.22 $X2=0 $Y2=0
cc_165 Y N_A_121_368#_c_260_n 0.00345031f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_166 Y N_VPWR_c_328_n 0.011066f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_167 Y N_VPWR_c_326_n 0.00915947f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_168 N_Y_c_221_n N_VGND_M1003_d 0.00320495f $X=2.16 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_169 N_Y_c_221_n N_VGND_c_360_n 0.0227484f $X=2.16 $Y=1.095 $X2=0 $Y2=0
cc_170 N_Y_c_222_n N_VGND_c_360_n 0.00751247f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_171 N_Y_c_224_n N_VGND_c_360_n 0.020732f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_172 N_Y_c_222_n N_VGND_c_361_n 0.0194588f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_173 N_Y_c_224_n N_VGND_c_362_n 0.0428125f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_174 N_Y_c_222_n N_VGND_c_364_n 0.0184284f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_175 N_Y_c_222_n N_VGND_c_367_n 0.0152535f $X=2.375 $Y=0.495 $X2=0 $Y2=0
cc_176 N_Y_c_224_n N_VGND_c_367_n 0.0354986f $X=1.09 $Y=0.765 $X2=0 $Y2=0
cc_177 N_Y_c_221_n A_351_74# 0.00366293f $X=2.16 $Y=1.095 $X2=-0.19 $Y2=-0.245
cc_178 N_A_121_368#_c_259_n N_A_263_368#_M1001_s 0.00239704f $X=1.725 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_179 N_A_121_368#_c_258_n N_A_263_368#_c_284_n 0.00876522f $X=0.74 $Y=2.115
+ $X2=0 $Y2=0
cc_180 N_A_121_368#_c_258_n N_A_263_368#_c_285_n 0.0294464f $X=0.74 $Y=2.115
+ $X2=0 $Y2=0
cc_181 N_A_121_368#_c_259_n N_A_263_368#_c_285_n 0.0185322f $X=1.725 $Y=2.99
+ $X2=0 $Y2=0
cc_182 N_A_121_368#_M1001_d N_A_263_368#_c_291_n 0.00753427f $X=1.755 $Y=1.84
+ $X2=0 $Y2=0
cc_183 N_A_121_368#_c_267_n N_A_263_368#_c_291_n 0.0170259f $X=1.89 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A_121_368#_c_259_n N_A_263_368#_c_286_n 0.00345031f $X=1.725 $Y=2.99
+ $X2=0 $Y2=0
cc_185 N_A_121_368#_c_259_n N_VPWR_c_327_n 0.00259349f $X=1.725 $Y=2.99 $X2=0
+ $Y2=0
cc_186 N_A_121_368#_c_259_n N_VPWR_c_328_n 0.0757767f $X=1.725 $Y=2.99 $X2=0
+ $Y2=0
cc_187 N_A_121_368#_c_260_n N_VPWR_c_328_n 0.0235512f $X=0.905 $Y=2.99 $X2=0
+ $Y2=0
cc_188 N_A_121_368#_c_259_n N_VPWR_c_326_n 0.0426952f $X=1.725 $Y=2.99 $X2=0
+ $Y2=0
cc_189 N_A_121_368#_c_260_n N_VPWR_c_326_n 0.0126924f $X=0.905 $Y=2.99 $X2=0
+ $Y2=0
cc_190 N_A_263_368#_c_300_n N_VPWR_M1002_d 0.00928873f $X=3.195 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_191 N_A_263_368#_c_286_n N_VPWR_c_327_n 0.0536098f $X=2.34 $Y=2.44 $X2=0
+ $Y2=0
cc_192 N_A_263_368#_c_300_n N_VPWR_c_327_n 0.0206577f $X=3.195 $Y=2.035 $X2=0
+ $Y2=0
cc_193 N_A_263_368#_c_288_n N_VPWR_c_327_n 0.026688f $X=3.36 $Y=2.815 $X2=0
+ $Y2=0
cc_194 N_A_263_368#_c_286_n N_VPWR_c_328_n 0.011066f $X=2.34 $Y=2.44 $X2=0 $Y2=0
cc_195 N_A_263_368#_c_288_n N_VPWR_c_330_n 0.014549f $X=3.36 $Y=2.815 $X2=0
+ $Y2=0
cc_196 N_A_263_368#_c_286_n N_VPWR_c_326_n 0.00915947f $X=2.34 $Y=2.44 $X2=0
+ $Y2=0
cc_197 N_A_263_368#_c_288_n N_VPWR_c_326_n 0.0119743f $X=3.36 $Y=2.815 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__dlrbp_2.pex.spice
* Created: Wed Sep  2 12:05:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRBP_2%D 3 7 9 12
c39 12 0 1.09742e-19 $X=0.59 $Y=1.615
r40 12 15 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.615
+ $X2=0.585 $Y2=1.78
r41 12 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.615
+ $X2=0.585 $Y2=1.45
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.615 $X2=0.59 $Y2=1.615
r43 9 13 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.59 $Y2=1.615
r44 7 14 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=1.45
r45 3 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=0.505 $Y=2.38 $X2=0.505
+ $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%GATE 3 6 8 11 13
c38 13 0 2.61276e-20 $X=1.13 $Y=1.22
c39 8 0 1.09742e-19 $X=1.2 $Y=1.295
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.385
+ $X2=1.13 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.385
+ $X2=1.13 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.385 $X2=1.13 $Y2=1.385
r43 8 12 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=1.13 $Y=1.295 $X2=1.13
+ $Y2=1.385
r44 6 14 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=1.125 $Y=2.38
+ $X2=1.125 $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.075 $Y=0.74
+ $X2=1.075 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%A_230_74# 1 2 7 9 11 13 15 16 18 19 20 24 29
+ 30 32 34 35 38 45 48 50 56
c137 34 0 6.32864e-20 $X=3.73 $Y=0.345
c138 30 0 2.61276e-20 $X=2.81 $Y=0.665
c139 19 0 8.05161e-20 $X=3.715 $Y=1.765
c140 16 0 1.64605e-19 $X=3.175 $Y=1.84
r141 49 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.7 $Y=1.505 $X2=1.7
+ $Y2=1.415
r142 48 51 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.505
+ $X2=1.66 $Y2=1.67
r143 48 50 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.505
+ $X2=1.66 $Y2=1.34
r144 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.505 $X2=1.7 $Y2=1.505
r145 43 45 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=2.065
+ $X2=1.54 $Y2=2.065
r146 41 50 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.54 $Y=1.01
+ $X2=1.54 $Y2=1.34
r147 40 41 13.823 $w=4.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.375 $Y=0.665
+ $X2=1.375 $Y2=1.01
r148 38 40 3.58824 $w=4.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.375 $Y=0.515
+ $X2=1.375 $Y2=0.665
r149 35 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=0.345
+ $X2=3.73 $Y2=0.51
r150 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=0.345 $X2=3.73 $Y2=0.345
r151 32 54 18.4631 $w=1.68e-07 $l=2.83e-07 $layer=LI1_cond $X=2.895 $Y=0.382
+ $X2=2.895 $Y2=0.665
r152 32 34 33.8954 $w=2.53e-07 $l=7.5e-07 $layer=LI1_cond $X=2.98 $Y=0.382
+ $X2=3.73 $Y2=0.382
r153 31 40 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.625 $Y=0.665
+ $X2=1.375 $Y2=0.665
r154 30 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.665
+ $X2=2.895 $Y2=0.665
r155 30 31 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=2.81 $Y=0.665
+ $X2=1.625 $Y2=0.665
r156 29 45 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.54 $Y=1.94
+ $X2=1.54 $Y2=2.065
r157 29 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.54 $Y=1.94
+ $X2=1.54 $Y2=1.67
r158 24 62 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.79 $Y=0.83
+ $X2=3.79 $Y2=0.51
r159 22 24 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.79 $Y=1.69
+ $X2=3.79 $Y2=0.83
r160 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=1.765
+ $X2=3.79 $Y2=1.69
r161 19 20 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.715 $Y=1.765
+ $X2=3.265 $Y2=1.765
r162 16 20 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.175 $Y=1.84
+ $X2=3.265 $Y2=1.765
r163 16 18 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.175 $Y=1.84
+ $X2=3.175 $Y2=2.46
r164 13 25 53.0007 $w=1.77e-07 $l=1.94936e-07 $layer=POLY_cond $X=2.175 $Y=1.225
+ $X2=2.185 $Y2=1.415
r165 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.175 $Y=1.225
+ $X2=2.175 $Y2=0.78
r166 9 25 20.0833 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.185 $Y=1.49
+ $X2=2.185 $Y2=1.415
r167 9 11 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.185 $Y=1.49
+ $X2=2.185 $Y2=2.38
r168 8 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.415
+ $X2=1.7 $Y2=1.415
r169 7 25 6.7465 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.095 $Y=1.415
+ $X2=2.185 $Y2=1.415
r170 7 8 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.095 $Y=1.415
+ $X2=1.865 $Y2=1.415
r171 2 43 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.96 $X2=1.375 $Y2=2.105
r172 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.37 $X2=1.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%A_27_112# 1 2 9 13 15 21 22 23 26 27 29 31
+ 32
c85 26 0 9.98003e-21 $X=2.65 $Y=1.635
c86 22 0 1.64605e-19 $X=2.485 $Y=2.445
c87 9 0 1.28743e-19 $X=2.755 $Y=2.46
r88 31 32 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.115
+ $X2=0.265 $Y2=1.95
r89 29 32 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.17 $Y=1.13
+ $X2=0.17 $Y2=1.95
r90 27 35 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.635
+ $X2=2.665 $Y2=1.8
r91 27 34 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.635
+ $X2=2.665 $Y2=1.47
r92 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.635 $X2=2.65 $Y2=1.635
r93 24 26 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=2.645 $Y=2.36
+ $X2=2.645 $Y2=1.635
r94 22 24 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.485 $Y=2.445
+ $X2=2.645 $Y2=2.36
r95 22 23 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.485 $Y=2.445
+ $X2=0.445 $Y2=2.445
r96 21 23 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=2.36
+ $X2=0.445 $Y2=2.445
r97 20 31 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.115
r98 20 21 7.36283 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.36
r99 15 29 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r100 15 17 3.89722 $w=3.6e-07 $l=1.15e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.835
r101 13 34 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.77 $Y=0.72
+ $X2=2.77 $Y2=1.47
r102 9 35 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.755 $Y=2.46
+ $X2=2.755 $Y2=1.8
r103 2 31 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r104 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%A_363_82# 1 2 9 12 14 15 16 19 20 21 24 25
+ 33 35 39 42
c119 39 0 9.98003e-21 $X=3.22 $Y=1.315
c120 35 0 8.05161e-20 $X=3.18 $Y=1.215
c121 15 0 1.28743e-19 $X=2.12 $Y=1.94
r122 39 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.315
+ $X2=3.22 $Y2=1.15
r123 38 40 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.315
+ $X2=3.18 $Y2=1.48
r124 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.315 $X2=3.22 $Y2=1.315
r125 35 38 2.81084 $w=4.08e-07 $l=1e-07 $layer=LI1_cond $X=3.18 $Y=1.215
+ $X2=3.18 $Y2=1.315
r126 31 33 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=1.96 $Y=2.065
+ $X2=2.12 $Y2=2.065
r127 25 44 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.87 $Y=2.215
+ $X2=3.71 $Y2=2.215
r128 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=2.215 $X2=3.87 $Y2=2.215
r129 22 24 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.87 $Y=2.905
+ $X2=3.87 $Y2=2.215
r130 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=3.87 $Y2=2.905
r131 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=3.145 $Y2=2.99
r132 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=2.905
+ $X2=3.145 $Y2=2.99
r133 19 40 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=3.06 $Y=2.905
+ $X2=3.06 $Y2=1.48
r134 17 28 7.83486 $w=3.27e-07 $l=2.95212e-07 $layer=LI1_cond $X=2.205 $Y=1.215
+ $X2=2 $Y2=1.005
r135 16 35 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.975 $Y=1.215
+ $X2=3.18 $Y2=1.215
r136 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.975 $Y=1.215
+ $X2=2.205 $Y2=1.215
r137 15 33 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=1.94
+ $X2=2.12 $Y2=2.065
r138 14 17 5.97199 $w=3.27e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=1.3
+ $X2=2.205 $Y2=1.215
r139 14 15 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.12 $Y=1.3 $X2=2.12
+ $Y2=1.94
r140 10 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=2.38
+ $X2=3.71 $Y2=2.215
r141 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.71 $Y=2.38
+ $X2=3.71 $Y2=2.75
r142 9 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.13 $Y=0.72
+ $X2=3.13 $Y2=1.15
r143 2 31 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=1.96 $X2=1.96 $Y2=2.105
r144 1 28 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.41 $X2=1.96 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%A_821_98# 1 2 7 9 14 18 22 26 30 32 33 36 40
+ 44 46 47 50 54 60 62 64 66 69 70 71 81
c168 71 0 1.03706e-19 $X=5.33 $Y=1.72
c169 62 0 7.12304e-20 $X=5.955 $Y=1.805
c170 47 0 1.21791e-20 $X=5.095 $Y=2.155
c171 26 0 1.93666e-19 $X=6.53 $Y=0.74
c172 7 0 6.32864e-20 $X=4.18 $Y=1.115
r173 83 85 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.1 $Y=1.465
+ $X2=6.155 $Y2=1.465
r174 74 75 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.33 $Y=2.155
+ $X2=5.33 $Y2=2.32
r175 73 74 4.32624 $w=4.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.33 $Y=1.985
+ $X2=5.33 $Y2=2.155
r176 70 73 4.58073 $w=4.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.33 $Y=1.805
+ $X2=5.33 $Y2=1.985
r177 70 71 7.30169 $w=4.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=1.805
+ $X2=5.33 $Y2=1.72
r178 69 71 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.18 $Y=1.13
+ $X2=5.18 $Y2=1.72
r179 67 87 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.53 $Y=1.465
+ $X2=6.605 $Y2=1.465
r180 67 85 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=6.53 $Y=1.465
+ $X2=6.155 $Y2=1.465
r181 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.465 $X2=6.53 $Y2=1.465
r182 64 78 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.04 $Y=1.465
+ $X2=6.04 $Y2=1.805
r183 64 66 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.125 $Y=1.465
+ $X2=6.53 $Y2=1.465
r184 63 70 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=5.565 $Y=1.805
+ $X2=5.33 $Y2=1.805
r185 62 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=1.805
+ $X2=6.04 $Y2=1.805
r186 62 63 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.955 $Y=1.805
+ $X2=5.565 $Y2=1.805
r187 60 75 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.4 $Y=2.4 $X2=5.4
+ $Y2=2.32
r188 52 69 11.1798 $w=4.73e-07 $l=2.37e-07 $layer=LI1_cond $X=5.027 $Y=0.893
+ $X2=5.027 $Y2=1.13
r189 52 54 9.51827 $w=4.73e-07 $l=3.78e-07 $layer=LI1_cond $X=5.027 $Y=0.893
+ $X2=5.027 $Y2=0.515
r190 50 82 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=2.155
+ $X2=4.41 $Y2=2.32
r191 50 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=2.155
+ $X2=4.41 $Y2=1.99
r192 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.41
+ $Y=2.155 $X2=4.41 $Y2=2.155
r193 47 74 2.80859 $w=3.3e-07 $l=2.35e-07 $layer=LI1_cond $X=5.095 $Y=2.155
+ $X2=5.33 $Y2=2.155
r194 47 49 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=5.095 $Y=2.155
+ $X2=4.41 $Y2=2.155
r195 42 44 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.18 $Y=1.19
+ $X2=4.32 $Y2=1.19
r196 38 46 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=7.625 $Y=1.3
+ $X2=7.615 $Y2=1.465
r197 38 40 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.625 $Y=1.3
+ $X2=7.625 $Y2=0.79
r198 34 46 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.63
+ $X2=7.615 $Y2=1.465
r199 34 36 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=7.615 $Y=1.63
+ $X2=7.615 $Y2=2.34
r200 33 87 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.695 $Y=1.465
+ $X2=6.605 $Y2=1.465
r201 32 46 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.525 $Y=1.465
+ $X2=7.615 $Y2=1.465
r202 32 33 145.135 $w=3.3e-07 $l=8.3e-07 $layer=POLY_cond $X=7.525 $Y=1.465
+ $X2=6.695 $Y2=1.465
r203 28 87 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.605 $Y=1.63
+ $X2=6.605 $Y2=1.465
r204 28 30 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.605 $Y=1.63
+ $X2=6.605 $Y2=2.4
r205 24 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.53 $Y=1.3
+ $X2=6.53 $Y2=1.465
r206 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.53 $Y=1.3
+ $X2=6.53 $Y2=0.74
r207 20 85 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.63
+ $X2=6.155 $Y2=1.465
r208 20 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.155 $Y=1.63
+ $X2=6.155 $Y2=2.4
r209 16 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.1 $Y=1.3 $X2=6.1
+ $Y2=1.465
r210 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.1 $Y=1.3 $X2=6.1
+ $Y2=0.74
r211 14 82 167.145 $w=1.8e-07 $l=4.3e-07 $layer=POLY_cond $X=4.365 $Y=2.75
+ $X2=4.365 $Y2=2.32
r212 10 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.32 $Y=1.265
+ $X2=4.32 $Y2=1.19
r213 10 81 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=4.32 $Y=1.265
+ $X2=4.32 $Y2=1.99
r214 7 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.115
+ $X2=4.18 $Y2=1.19
r215 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.18 $Y=1.115 $X2=4.18
+ $Y2=0.83
r216 2 73 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=5.215
+ $Y=1.84 $X2=5.4 $Y2=1.985
r217 2 60 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=5.215
+ $Y=1.84 $X2=5.4 $Y2=2.4
r218 1 54 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.81
+ $Y=0.37 $X2=4.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%A_641_80# 1 2 9 13 15 16 17 23 26 27 28 33
c86 16 0 1.47999e-19 $X=5.035 $Y=1.35
c87 9 0 7.12304e-20 $X=5.125 $Y=2.4
r88 33 36 7.92305 $w=3.18e-07 $l=2.2e-07 $layer=LI1_cond $X=4.765 $Y=1.515
+ $X2=4.765 $Y2=1.735
r89 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.515 $X2=4.77 $Y2=1.515
r90 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.4 $Y=1.735
+ $X2=3.655 $Y2=1.735
r91 28 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=1.735
+ $X2=3.655 $Y2=1.735
r92 27 36 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.605 $Y=1.735
+ $X2=4.765 $Y2=1.735
r93 27 28 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.605 $Y=1.735
+ $X2=3.74 $Y2=1.735
r94 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=1.65
+ $X2=3.655 $Y2=1.735
r95 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.655 $Y=0.96
+ $X2=3.655 $Y2=1.65
r96 21 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=1.82 $X2=3.4
+ $Y2=1.735
r97 21 23 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.4 $Y=1.82 $X2=3.4
+ $Y2=2.11
r98 17 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.57 $Y=0.875
+ $X2=3.655 $Y2=0.96
r99 17 19 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.57 $Y=0.875
+ $X2=3.46 $Y2=0.875
r100 15 34 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=5.035 $Y=1.515
+ $X2=4.77 $Y2=1.515
r101 15 16 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.035 $Y=1.515
+ $X2=5.035 $Y2=1.35
r102 11 16 34.7346 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=5.17 $Y=1.35
+ $X2=5.035 $Y2=1.35
r103 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.17 $Y=1.35
+ $X2=5.17 $Y2=0.74
r104 7 16 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=5.125 $Y=1.68
+ $X2=5.035 $Y2=1.35
r105 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.125 $Y=1.68
+ $X2=5.125 $Y2=2.4
r106 2 23 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=1.96 $X2=3.4 $Y2=2.11
r107 1 19 182 $w=1.7e-07 $l=5.88855e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.4 $X2=3.46 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%RESET_B 3 6 8 11 12 13
c40 13 0 2.71532e-19 $X=5.62 $Y=1.22
c41 12 0 1.47999e-19 $X=5.62 $Y=1.385
c42 6 0 1.21791e-20 $X=5.625 $Y=2.4
r43 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.62 $Y=1.385
+ $X2=5.62 $Y2=1.55
r44 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.62 $Y=1.385
+ $X2=5.62 $Y2=1.22
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.62
+ $Y=1.385 $X2=5.62 $Y2=1.385
r46 8 12 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=5.52 $Y=1.365 $X2=5.62
+ $Y2=1.365
r47 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.625 $Y=2.4
+ $X2=5.625 $Y2=1.55
r48 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.56 $Y=0.74 $X2=5.56
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%A_1449_368# 1 2 9 13 17 21 25 28 31 37 40 41
+ 47
c71 40 0 1.93666e-19 $X=7.41 $Y=1.13
r72 46 47 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.465
+ $X2=8.625 $Y2=1.465
r73 45 46 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.195 $Y=1.465
+ $X2=8.615 $Y2=1.465
r74 44 45 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.165 $Y=1.465
+ $X2=8.195 $Y2=1.465
r75 38 44 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=8.08 $Y=1.465
+ $X2=8.165 $Y2=1.465
r76 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.08
+ $Y=1.465 $X2=8.08 $Y2=1.465
r77 35 41 1.11842 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=7.555 $Y=1.465
+ $X2=7.4 $Y2=1.465
r78 35 37 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=7.555 $Y=1.465
+ $X2=8.08 $Y2=1.465
r79 31 33 26.3947 $w=3.08e-07 $l=7.1e-07 $layer=LI1_cond $X=7.4 $Y=1.985 $X2=7.4
+ $Y2=2.695
r80 29 41 5.44021 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=1.63 $X2=7.4
+ $Y2=1.465
r81 29 31 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=7.4 $Y=1.63 $X2=7.4
+ $Y2=1.985
r82 28 41 5.44021 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=1.3 $X2=7.4
+ $Y2=1.465
r83 28 40 6.31985 $w=3.08e-07 $l=1.7e-07 $layer=LI1_cond $X=7.4 $Y=1.3 $X2=7.4
+ $Y2=1.13
r84 23 40 5.81909 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=0.965
+ $X2=7.41 $Y2=1.13
r85 23 25 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=7.41 $Y=0.965
+ $X2=7.41 $Y2=0.615
r86 19 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=1.465
r87 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=0.74
r88 15 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.63
+ $X2=8.615 $Y2=1.465
r89 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.615 $Y=1.63
+ $X2=8.615 $Y2=2.4
r90 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=1.465
r91 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=0.74
r92 7 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.165 $Y=1.63
+ $X2=8.165 $Y2=1.465
r93 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.165 $Y=1.63
+ $X2=8.165 $Y2=2.4
r94 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.39 $Y2=2.695
r95 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.39 $Y2=1.985
r96 1 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.47 $X2=7.41 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%VPWR 1 2 3 4 5 6 7 26 30 34 40 44 48 50 55
+ 56 58 59 60 62 70 82 86 92 95 98 105 109
r111 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r112 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 98 101 9.62469 $w=6.38e-07 $l=5.15e-07 $layer=LI1_cond $X=4.745 $Y=2.815
+ $X2=4.745 $Y2=3.33
r114 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 90 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 90 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r119 87 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=7.89 $Y2=3.33
r120 87 89 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 86 108 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.937 $Y2=3.33
r122 86 89 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.4 $Y2=3.33
r123 85 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r124 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r125 82 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.89 $Y2=3.33
r126 82 84 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.44 $Y2=3.33
r127 81 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r128 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r129 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r131 75 101 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=4.745 $Y2=3.33
r132 75 77 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=5.52 $Y2=3.33
r133 74 96 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 71 95 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.512 $Y2=3.33
r136 71 73 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 70 101 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.745 $Y2=3.33
r138 70 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 69 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 66 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r144 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r145 63 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r146 63 65 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r147 62 95 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.512 $Y2=3.33
r148 62 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.16 $Y2=3.33
r149 60 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r150 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r151 60 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 58 80 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.665 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=3.33
+ $X2=6.83 $Y2=3.33
r154 57 84 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.995 $Y=3.33
+ $X2=7.44 $Y2=3.33
r155 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.995 $Y=3.33
+ $X2=6.83 $Y2=3.33
r156 55 77 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=5.52 $Y2=3.33
r157 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=5.9 $Y2=3.33
r158 54 80 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.065 $Y=3.33
+ $X2=6.48 $Y2=3.33
r159 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=3.33
+ $X2=5.9 $Y2=3.33
r160 50 53 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.815
r161 48 108 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.937 $Y2=3.33
r162 48 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.88 $Y2=2.815
r163 44 47 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.89 $Y=1.985
+ $X2=7.89 $Y2=2.695
r164 42 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.89 $Y2=3.33
r165 42 47 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.89 $Y2=2.695
r166 38 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=3.33
r167 38 40 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=2.305
r168 34 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.9 $Y=2.145
+ $X2=5.9 $Y2=2.825
r169 32 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=3.245 $X2=5.9
+ $Y2=3.33
r170 32 37 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.9 $Y=3.245
+ $X2=5.9 $Y2=2.825
r171 28 95 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.512 $Y=3.245
+ $X2=2.512 $Y2=3.33
r172 28 30 14.5239 $w=3.63e-07 $l=4.6e-07 $layer=LI1_cond $X=2.512 $Y=3.245
+ $X2=2.512 $Y2=2.785
r173 24 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r174 24 26 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.865
r175 7 53 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.815
r176 7 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=1.985
r177 6 47 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=7.705
+ $Y=1.84 $X2=7.89 $Y2=2.695
r178 6 44 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.705
+ $Y=1.84 $X2=7.89 $Y2=1.985
r179 5 40 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.84 $X2=6.83 $Y2=2.305
r180 4 37 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=5.715
+ $Y=1.84 $X2=5.9 $Y2=2.825
r181 4 34 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=5.715
+ $Y=1.84 $X2=5.9 $Y2=2.145
r182 3 98 600 $w=1.7e-07 $l=4.04784e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=2.54 $X2=4.745 $Y2=2.815
r183 2 30 600 $w=1.7e-07 $l=9.35147e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.96 $X2=2.51 $Y2=2.785
r184 1 26 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.815 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%Q 1 2 9 13 17 18 19 20 23
c53 9 0 1.67826e-19 $X=6.315 $Y=0.515
r54 22 23 25.3036 $w=2.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.96 $Y=1.8
+ $X2=6.96 $Y2=1.295
r55 21 23 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.96 $Y=1.13
+ $X2=6.96 $Y2=1.295
r56 19 21 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.96 $Y2=1.13
r57 19 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.48 $Y2=1.045
r58 17 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.96 $Y2=1.8
r59 17 18 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.465 $Y2=1.885
r60 13 15 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.38 $Y=1.985
+ $X2=6.38 $Y2=2.815
r61 11 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.38 $Y=1.97
+ $X2=6.465 $Y2=1.885
r62 11 13 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.38 $Y=1.97
+ $X2=6.38 $Y2=1.985
r63 7 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.315 $Y=0.96
+ $X2=6.48 $Y2=1.045
r64 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.315 $Y=0.96
+ $X2=6.315 $Y2=0.515
r65 2 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.245
+ $Y=1.84 $X2=6.38 $Y2=2.815
r66 2 13 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.245
+ $Y=1.84 $X2=6.38 $Y2=1.985
r67 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.175
+ $Y=0.37 $X2=6.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%Q_N 1 2 9 13 14 19 25
r31 17 19 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=8.405 $Y=2 $X2=8.405
+ $Y2=2.035
r32 14 17 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=8.405 $Y=1.975
+ $X2=8.405 $Y2=2
r33 14 25 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=8.405 $Y=1.975
+ $X2=8.405 $Y2=1.82
r34 14 22 24.1693 $w=3.58e-07 $l=7.55e-07 $layer=LI1_cond $X=8.405 $Y=2.06
+ $X2=8.405 $Y2=2.815
r35 14 19 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=8.405 $Y=2.06
+ $X2=8.405 $Y2=2.035
r36 13 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.5 $Y=1.13 $X2=8.5
+ $Y2=1.82
r37 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=8.415 $Y=0.96
+ $X2=8.415 $Y2=1.13
r38 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=8.415 $Y=0.96
+ $X2=8.415 $Y2=0.515
r39 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=1.985
r40 2 22 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=2.815
r41 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 47
+ 54 55 57 58 60 61 62 64 91 95 101 104 108
r109 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r110 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r111 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r112 99 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r113 99 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r114 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r115 96 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=7.91 $Y2=0
r116 96 98 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r117 95 107 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.937 $Y2=0
r118 95 98 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=0 $X2=8.4
+ $Y2=0
r119 94 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r120 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 91 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.91 $Y2=0
r122 91 93 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r123 90 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r124 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r125 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r126 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r127 83 86 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r128 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r129 78 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.08 $Y2=0
r130 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r131 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r132 75 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r133 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r134 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r135 72 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r136 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r137 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r138 69 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.79 $Y2=0
r139 69 71 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r140 67 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r141 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r142 64 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.79 $Y2=0
r143 64 66 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r144 62 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r145 62 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r146 62 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r147 60 89 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.65 $Y=0 $X2=6.48
+ $Y2=0
r148 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.65 $Y=0 $X2=6.815
+ $Y2=0
r149 59 93 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.98 $Y=0 $X2=7.44
+ $Y2=0
r150 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.98 $Y=0 $X2=6.815
+ $Y2=0
r151 57 86 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.52
+ $Y2=0
r152 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.775
+ $Y2=0
r153 56 89 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.94 $Y=0 $X2=6.48
+ $Y2=0
r154 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.94 $Y=0 $X2=5.775
+ $Y2=0
r155 55 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.56
+ $Y2=0
r156 54 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.08
+ $Y2=0
r157 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.395
+ $Y2=0
r158 47 74 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.16 $Y2=0
r159 47 51 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=2.472 $Y=0
+ $X2=2.472 $Y2=0.325
r160 47 77 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.472 $Y=0 $X2=2.64
+ $Y2=0
r161 42 107 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.937 $Y2=0
r162 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0.515
r163 38 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r164 38 40 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.615
r165 34 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0.085
+ $X2=6.815 $Y2=0
r166 34 36 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.815 $Y=0.085
+ $X2=6.815 $Y2=0.61
r167 30 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=0.085
+ $X2=5.775 $Y2=0
r168 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.775 $Y=0.085
+ $X2=5.775 $Y2=0.515
r169 26 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=0.085
+ $X2=4.395 $Y2=0
r170 26 28 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.395 $Y=0.085
+ $X2=4.395 $Y2=0.83
r171 22 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r172 22 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.515
r173 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r174 6 40 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.7
+ $Y=0.47 $X2=7.91 $Y2=0.615
r175 5 36 182 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_NDIFF $count=1 $X=6.605
+ $Y=0.37 $X2=6.815 $Y2=0.61
r176 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.635
+ $Y=0.37 $X2=5.775 $Y2=0.515
r177 3 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.255
+ $Y=0.62 $X2=4.395 $Y2=0.83
r178 2 51 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.41 $X2=2.47 $Y2=0.325
r179 1 24 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.56 $X2=0.79 $Y2=0.515
.ends


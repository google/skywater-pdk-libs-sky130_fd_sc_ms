* File: sky130_fd_sc_ms__nand3_2.pex.spice
* Created: Fri Aug 28 17:43:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND3_2%C 1 3 6 8 10 13 15 21 22
c51 22 0 1.28262e-20 $X=0.91 $Y=1.43
c52 21 0 6.03852e-20 $X=0.57 $Y=1.385
c53 13 0 1.85749e-19 $X=0.955 $Y=2.4
r54 22 23 6.39823 $w=3.39e-07 $l=4.5e-08 $layer=POLY_cond $X=0.91 $Y=1.43
+ $X2=0.955 $Y2=1.43
r55 20 22 48.3422 $w=3.39e-07 $l=3.4e-07 $layer=POLY_cond $X=0.57 $Y=1.43
+ $X2=0.91 $Y2=1.43
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.385 $X2=0.57 $Y2=1.385
r57 15 21 10.2785 $w=3.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.57 $Y2=1.365
r58 11 23 17.5597 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.955 $Y=1.64
+ $X2=0.955 $Y2=1.43
r59 11 13 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.955 $Y=1.64
+ $X2=0.955 $Y2=2.4
r60 8 22 21.8644 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.91 $Y=1.22 $X2=0.91
+ $Y2=1.43
r61 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.91 $Y=1.22 $X2=0.91
+ $Y2=0.74
r62 4 20 9.24189 $w=3.39e-07 $l=6.5e-08 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.57 $Y2=1.43
r63 4 17 3.55457 $w=3.39e-07 $l=2.5e-08 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.48 $Y2=1.43
r64 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.4
r65 1 17 21.8644 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.48 $Y=1.22 $X2=0.48
+ $Y2=1.43
r66 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.48 $Y=1.22 $X2=0.48
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%B 3 7 11 15 17 18 20 25 26 28 32 39 44
c92 26 0 1.89089e-19 $X=2.9 $Y=1.485
c93 18 0 1.85749e-19 $X=1.795 $Y=2.035
c94 11 0 2.49691e-20 $X=2.855 $Y=2.4
c95 7 0 6.92032e-20 $X=1.455 $Y=2.4
c96 3 0 6.03852e-20 $X=1.34 $Y=0.74
r97 39 44 0.721711 $w=4.34e-07 $l=8.7178e-08 $layer=LI1_cond $X=1.61 $Y=1.68
+ $X2=1.53 $Y2=1.665
r98 32 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.515
+ $X2=1.43 $Y2=1.68
r99 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.515
+ $X2=1.43 $Y2=1.35
r100 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.515 $X2=1.43 $Y2=1.515
r101 28 44 0.983871 $w=4.34e-07 $l=3.5e-08 $layer=LI1_cond $X=1.53 $Y=1.63
+ $X2=1.53 $Y2=1.665
r102 28 33 3.23272 $w=4.34e-07 $l=1.15e-07 $layer=LI1_cond $X=1.53 $Y=1.63
+ $X2=1.53 $Y2=1.515
r103 28 39 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.61 $Y=1.715
+ $X2=1.61 $Y2=1.68
r104 26 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.9 $Y=1.485
+ $X2=2.9 $Y2=1.65
r105 26 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.9 $Y=1.485
+ $X2=2.9 $Y2=1.32
r106 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.9
+ $Y=1.485 $X2=2.9 $Y2=1.485
r107 22 25 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.74 $Y=1.485
+ $X2=2.9 $Y2=1.485
r108 21 28 7.31957 $w=3.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.61 $Y=1.95
+ $X2=1.61 $Y2=1.715
r109 19 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=1.65
+ $X2=2.74 $Y2=1.485
r110 19 20 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.74 $Y=1.65 $X2=2.74
+ $Y2=1.95
r111 18 21 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.61 $Y2=1.95
r112 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=2.74 $Y2=1.95
r113 17 18 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.655 $Y=2.035
+ $X2=1.795 $Y2=2.035
r114 15 37 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.88 $Y=0.795
+ $X2=2.88 $Y2=1.32
r115 11 38 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.855 $Y=2.4
+ $X2=2.855 $Y2=1.65
r116 7 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=2.4
+ $X2=1.455 $Y2=1.68
r117 3 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.34 $Y=0.74
+ $X2=1.34 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%A 3 7 11 15 17 24 26
c54 24 0 2.83261e-19 $X=2.13 $Y=1.515
c55 11 0 5.74086e-20 $X=2.325 $Y=0.795
r56 25 26 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.325 $Y=1.515
+ $X2=2.405 $Y2=1.515
r57 23 25 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.325 $Y2=1.515
r58 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r59 21 23 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.91 $Y=1.515
+ $X2=2.13 $Y2=1.515
r60 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.895 $Y=1.515
+ $X2=1.91 $Y2=1.515
r61 17 24 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r62 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=1.515
r63 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=2.4
r64 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.35
+ $X2=2.325 $Y2=1.515
r65 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.325 $Y=1.35
+ $X2=2.325 $Y2=0.795
r66 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.68
+ $X2=1.91 $Y2=1.515
r67 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.91 $Y=1.68 $X2=1.91
+ $Y2=2.4
r68 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=1.515
r69 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 45
+ 54 57 61
r54 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r62 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 45 60 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r64 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 41 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.19 $Y2=3.33
r66 41 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r68 40 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 36 51 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r73 36 38 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 35 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.19 $Y2=3.33
r75 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 33 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 33 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 29 32 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=2.815
r80 27 60 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r81 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r82 23 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r83 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.795
r84 19 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r85 19 21 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.795
r86 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r87 13 51 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r88 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r89 4 32 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.815
r90 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=1.985
r91 3 25 600 $w=1.7e-07 $l=1.04112e-06 $layer=licon1_PDIFF $count=1 $X=2 $Y=1.84
+ $X2=2.18 $Y2=2.795
r92 2 21 600 $w=1.7e-07 $l=1.04341e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.795
r93 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r94 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%Y 1 2 3 4 15 19 20 21 23 25 27 30 31 35 41
+ 42
c84 19 0 5.74086e-20 $X=1.945 $Y=1.175
r85 41 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.375
+ $X2=1.68 $Y2=2.46
r86 41 42 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=2.475 $X2=1.68
+ $Y2=2.775
r87 41 46 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.68 $Y=2.475
+ $X2=1.68 $Y2=2.46
r88 35 37 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.11 $Y=1.02
+ $X2=2.11 $Y2=1.175
r89 32 33 3.61166 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=2.375
+ $X2=0.83 $Y2=2.46
r90 30 32 8.80133 $w=5.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.83 $Y=1.985
+ $X2=0.83 $Y2=2.375
r91 30 31 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=1.985
+ $X2=0.83 $Y2=1.82
r92 25 40 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.46 $X2=2.66
+ $Y2=2.375
r93 25 27 15.1525 $w=2.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.66 $Y=2.46
+ $X2=2.66 $Y2=2.815
r94 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.375
+ $X2=1.68 $Y2=2.375
r95 23 40 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=2.66 $Y2=2.375
r96 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=1.845 $Y2=2.375
r97 22 32 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.095 $Y=2.375
+ $X2=0.83 $Y2=2.375
r98 21 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=1.68 $Y2=2.375
r99 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=1.095 $Y2=2.375
r100 19 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=1.175
+ $X2=2.11 $Y2=1.175
r101 19 20 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.945 $Y=1.175
+ $X2=1.095 $Y2=1.175
r102 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.01 $Y=1.26
+ $X2=1.095 $Y2=1.175
r103 17 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.01 $Y=1.26
+ $X2=1.01 $Y2=1.82
r104 15 33 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.73 $Y=2.815
+ $X2=0.73 $Y2=2.46
r105 4 40 600 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.375
r106 4 27 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.815
r107 3 41 300 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.41
r108 2 30 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r109 2 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r110 1 35 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.425 $X2=2.11 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%A_27_74# 1 2 3 12 14 16 20 27 30
c59 27 0 1.28262e-20 $X=1.205 $Y=0.68
r60 27 28 7.32946 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=1.205 $Y=0.68
+ $X2=1.205 $Y2=0.835
r61 26 27 8.74806 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=1.205 $Y=0.495
+ $X2=1.205 $Y2=0.68
r62 20 23 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.265 $Y=0.835
+ $X2=0.265 $Y2=0.895
r63 20 21 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=0.835
+ $X2=0.265 $Y2=0.75
r64 17 27 3.17874 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0.68
+ $X2=1.205 $Y2=0.68
r65 16 30 4.5891 $w=1.7e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.93 $Y=0.68
+ $X2=3.095 $Y2=0.585
r66 16 17 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=2.93 $Y=0.68
+ $X2=1.37 $Y2=0.68
r67 15 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=0.835
+ $X2=0.265 $Y2=0.835
r68 14 28 3.17874 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0.835
+ $X2=1.205 $Y2=0.835
r69 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.04 $Y=0.835
+ $X2=0.43 $Y2=0.835
r70 12 21 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=0.225 $Y=0.515
+ $X2=0.225 $Y2=0.75
r71 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.955
+ $Y=0.425 $X2=3.095 $Y2=0.57
r72 2 26 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.37 $X2=1.125 $Y2=0.495
r73 1 23 182 $w=1.7e-07 $l=5.86409e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.265 $Y2=0.895
r74 1 12 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%VGND 1 6 8 10 20 21 24
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 17 20 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r44 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.695
+ $Y2=0
r46 15 17 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.2
+ $Y2=0
r47 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r48 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.695
+ $Y2=0
r50 10 12 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.24
+ $Y2=0
r51 8 21 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r52 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r53 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r54 4 6 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.495
r55 1 6 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.37 $X2=0.695 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_2%A_283_74# 1 2 11
r16 8 11 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.62 $Y=0.34 $X2=2.6
+ $Y2=0.34
r17 2 11 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.425 $X2=2.6 $Y2=0.34
r18 1 8 182 $w=1.7e-07 $l=2.19488e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.37 $X2=1.62 $Y2=0.34
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_391_368# B2 a_81_48# VPB pshort w=1e+06u l=180000u
+  ad=6.1e+11p pd=5.22e+06u as=3.2e+11p ps=2.64e+06u
M1001 VPWR A2 a_391_368# VPB pshort w=1e+06u l=180000u
+  ad=9.412e+11p pd=8.24e+06u as=0p ps=0u
M1002 VGND a_81_48# X VNB nlowvt w=740000u l=150000u
+  ad=6.808e+11p pd=6.28e+06u as=2.072e+11p ps=2.04e+06u
M1003 a_81_48# B1 a_391_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_304_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1005 X a_81_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 a_491_74# B1 a_81_48# VNB nlowvt w=740000u l=150000u
+  ad=1.85e+11p pd=1.98e+06u as=2.59e+11p ps=2.18e+06u
M1007 VPWR a_81_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_81_48# A1 a_304_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_81_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_391_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_491_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

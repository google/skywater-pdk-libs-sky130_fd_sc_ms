* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 a_1824_97# a_1910_71# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 VGND a_1910_71# a_2313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_639_85# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_27_74# SCE a_669_111# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X4 VGND a_2385_74# a_547_301# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 a_1688_97# a_1295_74# a_1893_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X6 a_1026_125# SCE a_669_111# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_159_404# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X8 VPWR a_1295_74# a_1492_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 a_143_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VPWR DE a_557_463# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X11 VPWR SCD a_1056_455# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X12 VGND a_1295_74# a_1492_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1688_97# a_1492_74# a_1824_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 a_2277_392# a_1295_74# a_2385_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 a_2313_74# a_1492_74# a_2385_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_505_111# a_547_301# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_27_74# a_639_85# a_669_111# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 VGND CLK a_1295_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_1893_508# a_1910_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X20 VGND SCD a_1026_125# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 a_2385_74# a_1492_74# a_2571_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X22 VPWR a_2385_74# a_547_301# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X23 a_117_464# a_159_404# VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X24 a_557_463# a_547_301# a_27_74# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X25 a_1056_455# a_639_85# a_669_111# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X26 a_27_74# D a_143_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 a_159_404# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 a_2571_508# a_547_301# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X29 VPWR a_1910_71# a_2277_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X30 VGND a_1688_97# a_1910_71# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 Q a_2385_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 a_639_85# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X33 Q a_2385_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X34 a_27_74# D a_117_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X35 a_2487_74# a_547_301# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 VGND a_159_404# a_505_111# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 a_669_111# a_1295_74# a_1688_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 a_2385_74# a_1295_74# a_2487_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 VPWR CLK a_1295_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X40 a_669_111# a_1492_74# a_1688_97# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X41 VPWR a_1688_97# a_1910_71# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
.ends

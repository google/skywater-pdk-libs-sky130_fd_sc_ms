* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2_4 A0 A1 S VGND VNB VPB VPWR X
M1000 X a_193_241# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.06535e+12p pd=6.79e+06u as=2.35648e+12p ps=1.609e+07u
M1001 a_709_119# S VGND VNB nlowvt w=640000u l=150000u
+  ad=4.224e+11p pd=3.88e+06u as=1.76805e+12p ps=1.249e+07u
M1002 VGND S a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1003 a_937_119# a_27_368# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.712e+11p pd=3.72e+06u as=0p ps=0u
M1004 X a_193_241# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_939_391# A1 a_193_241# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=9.25e+11p ps=7.85e+06u
M1006 X a_193_241# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=0p ps=0u
M1007 VGND a_27_368# a_937_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_193_241# A1 a_939_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR S a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1010 a_725_391# S VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1011 a_725_391# A0 a_193_241# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_193_241# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR S a_725_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_193_241# A1 a_709_119# VNB nlowvt w=640000u l=150000u
+  ad=9.216e+11p pd=6.72e+06u as=0p ps=0u
M1015 a_939_391# a_27_368# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_193_241# A0 a_725_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_937_119# A0 a_193_241# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_27_368# a_939_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_193_241# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_193_241# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_193_241# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_193_241# A0 a_937_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_193_241# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND S a_709_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_709_119# A1 a_193_241# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

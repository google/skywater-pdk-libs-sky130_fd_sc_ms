# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o31a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o31a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.455000 5.875000 1.785000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.115000 1.455000 6.595000 1.785000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.455000 5.155000 1.785000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.470000 3.235000 2.150000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 0.350000 0.905000 0.960000 ;
        RECT 0.575000 0.960000 1.700000 1.130000 ;
        RECT 0.575000 1.130000 0.835000 1.800000 ;
        RECT 0.575000 1.800000 1.810000 1.970000 ;
        RECT 0.575000 1.970000 0.835000 2.980000 ;
        RECT 1.450000 0.350000 1.700000 0.960000 ;
        RECT 1.480000 1.970000 1.810000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.145000  0.085000 0.395000 1.130000 ;
        RECT 1.085000  0.085000 1.255000 0.790000 ;
        RECT 1.880000  0.085000 2.210000 1.130000 ;
        RECT 3.960000  0.085000 4.210000 0.945000 ;
        RECT 4.820000  0.085000 5.150000 0.945000 ;
        RECT 5.750000  0.085000 6.080000 0.945000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 0.130000 1.820000 0.380000 3.245000 ;
        RECT 1.030000 2.140000 1.280000 3.245000 ;
        RECT 2.010000 1.820000 2.260000 3.245000 ;
        RECT 2.915000 2.715000 3.245000 3.245000 ;
        RECT 5.275000 2.635000 5.605000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.005000 1.300000 2.715000 1.630000 ;
      RECT 2.440000 0.265000 3.780000 0.435000 ;
      RECT 2.440000 0.435000 2.770000 0.960000 ;
      RECT 2.465000 1.630000 2.715000 2.375000 ;
      RECT 2.465000 2.375000 4.255000 2.545000 ;
      RECT 2.465000 2.545000 2.715000 2.980000 ;
      RECT 2.545000 1.130000 3.270000 1.300000 ;
      RECT 2.940000 0.605000 3.270000 1.130000 ;
      RECT 3.450000 0.435000 3.780000 1.115000 ;
      RECT 3.450000 1.115000 6.580000 1.285000 ;
      RECT 3.475000 1.955000 6.605000 2.125000 ;
      RECT 3.475000 2.125000 4.645000 2.205000 ;
      RECT 3.925000 2.545000 4.255000 2.980000 ;
      RECT 4.390000 0.605000 4.640000 1.115000 ;
      RECT 4.435000 2.205000 4.645000 2.980000 ;
      RECT 4.825000 2.295000 6.105000 2.465000 ;
      RECT 4.825000 2.465000 5.075000 2.980000 ;
      RECT 5.320000 0.605000 5.570000 1.115000 ;
      RECT 5.775000 2.465000 6.105000 2.980000 ;
      RECT 6.250000 0.605000 6.580000 1.115000 ;
      RECT 6.275000 2.125000 6.605000 2.980000 ;
  END
END sky130_fd_sc_ms__o31a_4

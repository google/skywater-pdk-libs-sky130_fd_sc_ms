* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_1 A B C VGND VNB VPB VPWR X
X0 a_121_136# B a_233_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_27_398# C VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VGND a_27_398# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_27_398# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_27_398# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 VPWR B a_27_398# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_27_398# A a_121_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_233_136# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

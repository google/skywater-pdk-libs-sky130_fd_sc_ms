* File: sky130_fd_sc_ms__a21oi_4.pex.spice
* Created: Wed Sep  2 11:51:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21OI_4%A2 3 7 11 15 19 23 27 31 33 34 35 53
c86 31 0 7.99896e-20 $X=2.05 $Y=0.74
r87 52 53 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.045 $Y=1.515
+ $X2=2.05 $Y2=1.515
r88 50 52 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.97 $Y=1.515
+ $X2=2.045 $Y2=1.515
r89 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.515 $X2=1.97 $Y2=1.515
r90 48 50 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.62 $Y=1.515
+ $X2=1.97 $Y2=1.515
r91 47 48 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.595 $Y=1.515
+ $X2=1.62 $Y2=1.515
r92 46 47 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.19 $Y=1.515
+ $X2=1.595 $Y2=1.515
r93 45 46 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.145 $Y=1.515
+ $X2=1.19 $Y2=1.515
r94 43 45 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.95 $Y=1.515
+ $X2=1.145 $Y2=1.515
r95 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.515 $X2=0.95 $Y2=1.515
r96 41 43 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.76 $Y=1.515
+ $X2=0.95 $Y2=1.515
r97 39 41 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=0.695 $Y=1.515
+ $X2=0.76 $Y2=1.515
r98 35 51 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.97 $Y2=1.565
r99 34 51 7.77229 $w=4.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.97 $Y2=1.565
r100 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r101 33 44 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.95 $Y2=1.565
r102 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.35
+ $X2=2.05 $Y2=1.515
r103 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.05 $Y=1.35
+ $X2=2.05 $Y2=0.74
r104 25 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.045 $Y=1.68
+ $X2=2.045 $Y2=1.515
r105 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.045 $Y=1.68
+ $X2=2.045 $Y2=2.4
r106 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.62 $Y2=1.515
r107 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.62 $Y2=0.74
r108 17 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.68
+ $X2=1.595 $Y2=1.515
r109 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.595 $Y=1.68
+ $X2=1.595 $Y2=2.4
r110 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=1.515
r111 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=0.74
r112 9 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.68
+ $X2=1.145 $Y2=1.515
r113 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.145 $Y=1.68
+ $X2=1.145 $Y2=2.4
r114 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.76 $Y=1.35
+ $X2=0.76 $Y2=1.515
r115 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.76 $Y=1.35 $X2=0.76
+ $Y2=0.74
r116 1 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.695 $Y=1.68
+ $X2=0.695 $Y2=1.515
r117 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.695 $Y=1.68
+ $X2=0.695 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%A1 3 7 11 15 19 23 27 31 33 34 49 50
c86 31 0 1.19938e-19 $X=3.845 $Y=2.4
c87 19 0 6.95413e-20 $X=3.34 $Y=0.74
c88 11 0 6.95443e-20 $X=2.91 $Y=0.74
c89 7 0 1.53462e-19 $X=2.495 $Y=2.4
c90 3 0 1.9142e-19 $X=2.48 $Y=0.74
r91 48 50 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=1.515
+ $X2=3.845 $Y2=1.515
r92 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.515 $X2=3.77 $Y2=1.515
r93 46 48 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.395 $Y=1.515
+ $X2=3.77 $Y2=1.515
r94 45 46 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.34 $Y=1.515
+ $X2=3.395 $Y2=1.515
r95 43 45 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.09 $Y=1.515
+ $X2=3.34 $Y2=1.515
r96 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.515 $X2=3.09 $Y2=1.515
r97 41 43 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=2.945 $Y=1.515
+ $X2=3.09 $Y2=1.515
r98 40 41 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.91 $Y=1.515
+ $X2=2.945 $Y2=1.515
r99 39 40 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.495 $Y=1.515
+ $X2=2.91 $Y2=1.515
r100 37 39 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.48 $Y=1.515
+ $X2=2.495 $Y2=1.515
r101 34 49 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.77 $Y2=1.565
r102 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r103 33 44 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.09 $Y2=1.565
r104 29 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.68
+ $X2=3.845 $Y2=1.515
r105 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.845 $Y=1.68
+ $X2=3.845 $Y2=2.4
r106 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.77 $Y=1.35
+ $X2=3.77 $Y2=1.515
r107 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.77 $Y=1.35
+ $X2=3.77 $Y2=0.74
r108 21 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.68
+ $X2=3.395 $Y2=1.515
r109 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.395 $Y=1.68
+ $X2=3.395 $Y2=2.4
r110 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.34 $Y=1.35
+ $X2=3.34 $Y2=1.515
r111 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.34 $Y=1.35
+ $X2=3.34 $Y2=0.74
r112 13 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=1.68
+ $X2=2.945 $Y2=1.515
r113 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.945 $Y=1.68
+ $X2=2.945 $Y2=2.4
r114 9 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.35
+ $X2=2.91 $Y2=1.515
r115 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.91 $Y=1.35
+ $X2=2.91 $Y2=0.74
r116 5 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.68
+ $X2=2.495 $Y2=1.515
r117 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.495 $Y=1.68
+ $X2=2.495 $Y2=2.4
r118 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.35
+ $X2=2.48 $Y2=1.515
r119 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.48 $Y=1.35 $X2=2.48
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%B1 1 3 6 10 14 18 20 21 24 26 27 38
c63 38 0 1.19938e-19 $X=5.08 $Y=1.515
r64 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.08
+ $Y=1.515 $X2=5.08 $Y2=1.515
r65 35 37 43.1642 $w=3.35e-07 $l=3e-07 $layer=POLY_cond $X=4.78 $Y=1.56 $X2=5.08
+ $Y2=1.56
r66 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.4
+ $Y=1.515 $X2=4.4 $Y2=1.515
r67 30 32 15.1075 $w=3.35e-07 $l=1.05e-07 $layer=POLY_cond $X=4.295 $Y=1.56
+ $X2=4.4 $Y2=1.56
r68 27 38 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=5.04 $Y=1.565 $X2=5.08
+ $Y2=1.565
r69 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r70 26 33 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.4 $Y2=1.565
r71 22 24 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.645 $Y=1.68
+ $X2=5.645 $Y2=2.4
r72 21 40 25.6873 $w=3.35e-07 $l=9.48683e-08 $layer=POLY_cond $X=5.285 $Y=1.605
+ $X2=5.21 $Y2=1.56
r73 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.555 $Y=1.605
+ $X2=5.645 $Y2=1.68
r74 20 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.555 $Y=1.605
+ $X2=5.285 $Y2=1.605
r75 16 40 21.5811 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.21 $Y=1.35
+ $X2=5.21 $Y2=1.56
r76 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.21 $Y=1.35
+ $X2=5.21 $Y2=0.74
r77 12 40 2.15821 $w=3.35e-07 $l=1.5e-08 $layer=POLY_cond $X=5.195 $Y=1.56
+ $X2=5.21 $Y2=1.56
r78 12 37 16.5463 $w=3.35e-07 $l=1.15e-07 $layer=POLY_cond $X=5.195 $Y=1.56
+ $X2=5.08 $Y2=1.56
r79 12 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.195 $Y=1.68
+ $X2=5.195 $Y2=2.4
r80 8 35 21.5811 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.78 $Y=1.35 $X2=4.78
+ $Y2=1.56
r81 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.78 $Y=1.35 $X2=4.78
+ $Y2=0.74
r82 4 35 5.03582 $w=3.35e-07 $l=3.5e-08 $layer=POLY_cond $X=4.745 $Y=1.56
+ $X2=4.78 $Y2=1.56
r83 4 32 49.6388 $w=3.35e-07 $l=3.45e-07 $layer=POLY_cond $X=4.745 $Y=1.56
+ $X2=4.4 $Y2=1.56
r84 4 6 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.745 $Y=1.68
+ $X2=4.745 $Y2=2.4
r85 1 30 17.2825 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.295 $Y=1.77
+ $X2=4.295 $Y2=1.56
r86 1 3 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=4.295 $Y=1.77 $X2=4.295
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%A_69_368# 1 2 3 4 5 6 7 22 24 26 30 32 34 35
+ 38 40 44 46 47 48 49 52 54 58 65 68 70 73
c98 38 0 1.53462e-19 $X=2.27 $Y=2.465
r99 58 61 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.91 $Y=1.985
+ $X2=5.91 $Y2=2.815
r100 56 61 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.91 $Y=2.905
+ $X2=5.91 $Y2=2.815
r101 55 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=2.99
+ $X2=4.97 $Y2=2.99
r102 54 56 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.785 $Y=2.99
+ $X2=5.91 $Y2=2.905
r103 54 55 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.785 $Y=2.99
+ $X2=5.055 $Y2=2.99
r104 50 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=2.905
+ $X2=4.97 $Y2=2.99
r105 50 52 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.97 $Y=2.905
+ $X2=4.97 $Y2=2.455
r106 48 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=2.99
+ $X2=4.97 $Y2=2.99
r107 48 49 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.885 $Y=2.99
+ $X2=4.155 $Y2=2.99
r108 47 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.03 $Y=2.905
+ $X2=4.155 $Y2=2.99
r109 46 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.46
+ $X2=4.03 $Y2=2.375
r110 46 47 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.03 $Y=2.46
+ $X2=4.03 $Y2=2.905
r111 45 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=2.375
+ $X2=3.17 $Y2=2.375
r112 44 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=2.375
+ $X2=4.03 $Y2=2.375
r113 44 45 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.905 $Y=2.375
+ $X2=3.335 $Y2=2.375
r114 41 68 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.355 $Y=2.375
+ $X2=2.23 $Y2=2.375
r115 40 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=2.375
+ $X2=3.17 $Y2=2.375
r116 40 41 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.005 $Y=2.375
+ $X2=2.355 $Y2=2.375
r117 36 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.46
+ $X2=2.23 $Y2=2.375
r118 36 38 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.23 $Y=2.46
+ $X2=2.23 $Y2=2.465
r119 35 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.29
+ $X2=2.23 $Y2=2.375
r120 34 67 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.035
r121 34 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.29
r122 33 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.37 $Y2=2.035
r123 32 67 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.23 $Y2=2.035
r124 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=1.535 $Y2=2.035
r125 28 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.035
r126 28 30 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.815
r127 27 63 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=0.555 $Y=2.035
+ $X2=0.43 $Y2=1.97
r128 26 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=1.37 $Y2=2.035
r129 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=0.555 $Y2=2.035
r130 22 63 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.43 $Y=2.12 $X2=0.43
+ $Y2=1.97
r131 22 24 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.43 $Y=2.12
+ $X2=0.43 $Y2=2.4
r132 7 61 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.84 $X2=5.87 $Y2=2.815
r133 7 58 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.84 $X2=5.87 $Y2=1.985
r134 6 52 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.835
+ $Y=1.84 $X2=4.97 $Y2=2.455
r135 5 72 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.935
+ $Y=1.84 $X2=4.07 $Y2=2.455
r136 4 70 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.035
+ $Y=1.84 $X2=3.17 $Y2=2.455
r137 3 67 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=1.84 $X2=2.27 $Y2=2.115
r138 3 38 300 $w=1.7e-07 $l=6.89202e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=1.84 $X2=2.27 $Y2=2.465
r139 2 65 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.84 $X2=1.37 $Y2=2.115
r140 2 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.84 $X2=1.37 $Y2=2.815
r141 1 63 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.84 $X2=0.47 $Y2=1.985
r142 1 24 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=0.345
+ $Y=1.84 $X2=0.47 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%VPWR 1 2 3 4 15 19 23 25 29 32 33 35 36 37
+ 46 55 56 59 62
r84 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r85 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r87 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r88 53 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r90 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 50 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.62 $Y2=3.33
r92 50 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 46 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.68 $Y2=3.33
r96 46 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 45 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 37 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 37 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 35 44 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.82 $Y2=3.33
r105 34 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.82 $Y2=3.33
r107 32 40 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.88 $Y2=3.33
r109 31 44 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.88 $Y2=3.33
r111 27 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=3.245
+ $X2=3.62 $Y2=3.33
r112 27 29 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.62 $Y=3.245
+ $X2=3.62 $Y2=2.805
r113 26 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.68 $Y2=3.33
r114 25 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=3.62 $Y2=3.33
r115 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=2.805 $Y2=3.33
r116 21 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r117 21 23 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.805
r118 17 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=3.245
+ $X2=1.82 $Y2=3.33
r119 17 19 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.82 $Y=3.245
+ $X2=1.82 $Y2=2.455
r120 13 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=3.33
r121 13 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=2.455
r122 4 29 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=1.84 $X2=3.62 $Y2=2.805
r123 3 23 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.84 $X2=2.72 $Y2=2.805
r124 2 19 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.84 $X2=1.82 $Y2=2.455
r125 1 15 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.785
+ $Y=1.84 $X2=0.92 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%Y 1 2 3 4 5 6 19 20 21 29 31 33 39 43 44 46
+ 47 48 49 54
c95 47 0 7.99896e-20 $X=2.64 $Y=0.925
r96 48 49 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.665
r97 48 57 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.18
r98 47 54 6.14322 $w=2.42e-07 $l=1.5e-07 $layer=LI1_cond $X=2.652 $Y=1.03
+ $X2=2.652 $Y2=0.88
r99 47 57 6.14322 $w=2.42e-07 $l=1.55885e-07 $layer=LI1_cond $X=2.652 $Y=1.03
+ $X2=2.64 $Y2=1.18
r100 47 54 0.956863 $w=2.55e-07 $l=2e-08 $layer=LI1_cond $X=2.652 $Y=0.86
+ $X2=2.652 $Y2=0.88
r101 41 49 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.64 $Y=1.95
+ $X2=2.64 $Y2=1.665
r102 37 39 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.465 $Y=1.01
+ $X2=5.465 $Y2=0.515
r103 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.685 $Y=2.035
+ $X2=4.52 $Y2=2.035
r104 33 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=5.42 $Y2=2.035
r105 33 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=4.685 $Y2=2.035
r106 32 44 5.43733 $w=2.35e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.65 $Y=1.095
+ $X2=4.525 $Y2=1.03
r107 31 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.34 $Y=1.095
+ $X2=5.465 $Y2=1.01
r108 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.34 $Y=1.095
+ $X2=4.65 $Y2=1.095
r109 27 44 1.12072 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=4.525 $Y=0.88
+ $X2=4.525 $Y2=1.03
r110 27 29 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=4.525 $Y=0.88
+ $X2=4.525 $Y2=0.515
r111 22 47 0.588783 $w=3e-07 $l=1.28e-07 $layer=LI1_cond $X=2.78 $Y=1.03
+ $X2=2.652 $Y2=1.03
r112 22 24 29.7714 $w=2.98e-07 $l=7.75e-07 $layer=LI1_cond $X=2.78 $Y=1.03
+ $X2=3.555 $Y2=1.03
r113 21 44 5.43733 $w=2.35e-07 $l=1.25e-07 $layer=LI1_cond $X=4.4 $Y=1.03
+ $X2=4.525 $Y2=1.03
r114 21 24 32.4605 $w=2.98e-07 $l=8.45e-07 $layer=LI1_cond $X=4.4 $Y=1.03
+ $X2=3.555 $Y2=1.03
r115 20 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.755 $Y=2.035
+ $X2=2.64 $Y2=1.95
r116 19 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=2.035
+ $X2=4.52 $Y2=2.035
r117 19 20 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=4.355 $Y=2.035
+ $X2=2.755 $Y2=2.035
r118 6 46 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.84 $X2=5.42 $Y2=2.115
r119 5 43 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.115
r120 4 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.425 $Y2=0.515
r121 3 29 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.44
+ $Y=0.37 $X2=4.565 $Y2=0.515
r122 2 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.37 $X2=3.555 $Y2=0.965
r123 1 47 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.37 $X2=2.695 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%A_84_74# 1 2 3 4 5 18 20 21 24 26 32 33 34
+ 36 37 42
c72 34 0 6.95443e-20 $X=3.82 $Y=0.34
c73 32 0 6.95413e-20 $X=2.96 $Y=0.34
r74 42 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.985 $Y=0.34
+ $X2=3.985 $Y2=0.53
r75 37 40 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=0.34
+ $X2=3.125 $Y2=0.53
r76 35 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=0.34
+ $X2=3.125 $Y2=0.34
r77 34 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=0.34
+ $X2=3.985 $Y2=0.34
r78 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.82 $Y=0.34
+ $X2=3.29 $Y2=0.34
r79 32 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=0.34
+ $X2=3.125 $Y2=0.34
r80 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.96 $Y=0.34
+ $X2=2.35 $Y2=0.34
r81 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.265 $Y=1.01
+ $X2=2.265 $Y2=0.515
r82 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=0.425
+ $X2=2.35 $Y2=0.34
r83 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.265 $Y=0.425
+ $X2=2.265 $Y2=0.515
r84 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.095
+ $X2=1.405 $Y2=1.095
r85 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.18 $Y=1.095
+ $X2=2.265 $Y2=1.01
r86 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.18 $Y=1.095
+ $X2=1.49 $Y2=1.095
r87 22 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=1.01
+ $X2=1.405 $Y2=1.095
r88 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.405 $Y=1.01
+ $X2=1.405 $Y2=0.515
r89 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=1.095
+ $X2=1.405 $Y2=1.095
r90 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.32 $Y=1.095
+ $X2=0.63 $Y2=1.095
r91 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.505 $Y=1.01
+ $X2=0.63 $Y2=1.095
r92 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.505 $Y=1.01
+ $X2=0.505 $Y2=0.515
r93 5 45 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.37 $X2=3.985 $Y2=0.53
r94 4 40 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=2.985
+ $Y=0.37 $X2=3.125 $Y2=0.53
r95 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.125
+ $Y=0.37 $X2=2.265 $Y2=0.515
r96 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.265
+ $Y=0.37 $X2=1.405 $Y2=0.515
r97 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.42
+ $Y=0.37 $X2=0.545 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_4%VGND 1 2 3 12 14 18 22 24 25 26 32 42 43 46
+ 49
c69 18 0 1.9142e-19 $X=1.835 $Y=0.595
r70 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r71 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r72 43 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r73 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r74 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=4.995
+ $Y2=0
r75 40 42 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=6
+ $Y2=0
r76 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r77 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r79 35 38 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r80 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.835
+ $Y2=0
r82 33 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.16
+ $Y2=0
r83 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.995
+ $Y2=0
r84 32 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.56
+ $Y2=0
r85 30 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r86 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 26 39 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r88 26 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r89 24 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.72
+ $Y2=0
r90 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.975
+ $Y2=0
r91 20 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=0.085
+ $X2=4.995 $Y2=0
r92 20 22 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=4.995 $Y=0.085
+ $X2=4.995 $Y2=0.595
r93 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0
r94 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0.595
r95 15 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.975
+ $Y2=0
r96 14 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.835
+ $Y2=0
r97 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.14
+ $Y2=0
r98 10 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0
r99 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0.595
r100 3 22 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.37 $X2=4.995 $Y2=0.595
r101 2 18 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.37 $X2=1.835 $Y2=0.595
r102 1 12 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.37 $X2=0.975 $Y2=0.595
.ends


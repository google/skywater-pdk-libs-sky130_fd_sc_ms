# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__xnor2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__xnor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.744800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.320000 1.315000 1.650000 ;
        RECT 1.085000 1.650000 1.315000 1.780000 ;
        RECT 4.445000 1.350000 5.835000 1.775000 ;
      LAYER mcon ;
        RECT 1.115000 1.580000 1.285000 1.750000 ;
        RECT 4.475000 1.580000 4.645000 1.750000 ;
      LAYER met1 ;
        RECT 1.055000 1.550000 1.345000 1.595000 ;
        RECT 1.055000 1.595000 4.705000 1.735000 ;
        RECT 1.055000 1.735000 1.345000 1.780000 ;
        RECT 4.415000 1.550000 4.705000 1.595000 ;
        RECT 4.415000 1.735000 4.705000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.744800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 2.155000 1.680000 ;
        RECT 1.985000 1.680000 2.155000 1.945000 ;
        RECT 1.985000 1.945000 6.535000 2.115000 ;
        RECT 6.365000 1.350000 8.155000 1.765000 ;
        RECT 6.365000 1.765000 6.535000 1.945000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.373400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 2.285000 7.655000 2.455000 ;
        RECT 3.035000 0.595000 3.365000 1.010000 ;
        RECT 3.035000 1.010000 8.495000 1.180000 ;
        RECT 4.060000 0.595000 4.390000 1.010000 ;
        RECT 7.325000 1.935000 8.555000 2.105000 ;
        RECT 7.325000 2.105000 7.655000 2.285000 ;
        RECT 7.325000 2.455000 7.655000 2.735000 ;
        RECT 8.225000 2.105000 8.555000 2.735000 ;
        RECT 8.325000 1.180000 8.495000 1.935000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.120000 0.085000 ;
        RECT 0.545000  0.085000 0.875000 0.810000 ;
        RECT 5.070000  0.085000 5.400000 0.500000 ;
        RECT 6.090000  0.085000 6.420000 0.500000 ;
        RECT 7.110000  0.085000 7.475000 0.500000 ;
        RECT 8.165000  0.085000 8.495000 0.500000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.120000 3.415000 ;
        RECT 0.115000 1.820000 0.365000 3.245000 ;
        RECT 1.095000 2.290000 1.265000 3.245000 ;
        RECT 2.000000 2.965000 2.340000 3.245000 ;
        RECT 3.080000 2.965000 3.410000 3.245000 ;
        RECT 5.265000 2.965000 5.600000 3.245000 ;
        RECT 6.340000 2.965000 6.670000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.350000 0.365000 0.980000 ;
      RECT 0.115000 0.980000 1.375000 1.150000 ;
      RECT 0.565000 1.820000 0.895000 1.950000 ;
      RECT 0.565000 1.950000 1.795000 2.120000 ;
      RECT 0.565000 2.120000 0.895000 2.700000 ;
      RECT 1.045000 0.350000 2.305000 0.600000 ;
      RECT 1.045000 0.600000 1.375000 0.980000 ;
      RECT 1.465000 2.120000 1.795000 2.625000 ;
      RECT 1.465000 2.625000 4.590000 2.795000 ;
      RECT 1.545000 0.770000 1.875000 1.010000 ;
      RECT 1.545000 1.010000 2.565000 1.180000 ;
      RECT 2.395000 1.180000 2.565000 1.350000 ;
      RECT 2.395000 1.350000 4.085000 1.680000 ;
      RECT 2.535000 0.255000 4.890000 0.425000 ;
      RECT 2.535000 0.425000 2.865000 0.840000 ;
      RECT 3.535000 0.425000 3.865000 0.840000 ;
      RECT 3.580000 2.795000 4.590000 2.955000 ;
      RECT 4.560000 0.425000 4.890000 0.670000 ;
      RECT 4.560000 0.670000 9.005000 0.840000 ;
      RECT 4.810000 2.625000 7.125000 2.795000 ;
      RECT 4.810000 2.795000 5.060000 2.980000 ;
      RECT 5.580000 0.350000 5.910000 0.670000 ;
      RECT 5.805000 2.795000 6.135000 2.980000 ;
      RECT 6.600000 0.350000 6.930000 0.670000 ;
      RECT 6.875000 2.795000 7.125000 2.905000 ;
      RECT 6.875000 2.905000 9.005000 3.075000 ;
      RECT 7.655000 0.350000 7.985000 0.670000 ;
      RECT 7.855000 2.275000 8.025000 2.905000 ;
      RECT 8.675000 0.350000 9.005000 0.670000 ;
      RECT 8.675000 0.840000 9.005000 1.130000 ;
      RECT 8.755000 1.935000 9.005000 2.905000 ;
  END
END sky130_fd_sc_ms__xnor2_4

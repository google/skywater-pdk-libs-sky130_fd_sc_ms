* File: sky130_fd_sc_ms__fah_1.pex.spice
* Created: Fri Aug 28 17:35:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FAH_1%CI 3 6 8 11 12 13
c42 12 0 1.05236e-19 $X=1.17 $Y=1.575
c43 11 0 4.00034e-20 $X=1.17 $Y=1.575
r44 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.575
+ $X2=1.17 $Y2=1.74
r45 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.575
+ $X2=1.17 $Y2=1.41
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.575 $X2=1.17 $Y2=1.575
r47 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=1.665 $X2=1.17
+ $Y2=1.575
r48 6 14 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.185 $Y=2.4
+ $X2=1.185 $Y2=1.74
r49 3 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.08 $Y=0.98 $X2=1.08
+ $Y2=1.41
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_83_21# 1 2 10 11 13 15 16 18 24 29 30 31 32
+ 33 34 36 37 38 39 42 43 44 45 47 52 56 60 66
c186 52 0 2.42155e-20 $X=4.37 $Y=2.255
c187 45 0 2.4784e-20 $X=5.885 $Y=0.68
c188 33 0 3.05634e-20 $X=3.155 $Y=2.28
c189 30 0 3.87212e-19 $X=2.01 $Y=1.86
c190 24 0 1.37092e-19 $X=1.735 $Y=1.31
r191 60 63 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.05 $Y=0.68
+ $X2=6.05 $Y2=0.775
r192 56 58 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.96 $Y=0.68
+ $X2=4.96 $Y2=0.84
r193 52 54 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.37 $Y=2.255
+ $X2=4.37 $Y2=2.37
r194 47 49 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.24 $Y=2.28 $X2=3.24
+ $Y2=2.37
r195 46 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.68
+ $X2=4.96 $Y2=0.68
r196 45 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.885 $Y=0.68
+ $X2=6.05 $Y2=0.68
r197 45 46 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.885 $Y=0.68
+ $X2=5.045 $Y2=0.68
r198 43 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0.84
+ $X2=4.96 $Y2=0.84
r199 43 44 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.875 $Y=0.84
+ $X2=4.285 $Y2=0.84
r200 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=0.755
+ $X2=4.285 $Y2=0.84
r201 41 42 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.2 $Y=0.425
+ $X2=4.2 $Y2=0.755
r202 40 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.37
+ $X2=3.24 $Y2=2.37
r203 39 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=2.37
+ $X2=4.37 $Y2=2.37
r204 39 40 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.205 $Y=2.37
+ $X2=3.325 $Y2=2.37
r205 37 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=0.34
+ $X2=4.2 $Y2=0.425
r206 37 38 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.115 $Y=0.34
+ $X2=2.765 $Y2=0.34
r207 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.68 $Y=0.425
+ $X2=2.765 $Y2=0.34
r208 35 36 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.68 $Y=0.425
+ $X2=2.68 $Y2=0.9
r209 33 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.28
+ $X2=3.24 $Y2=2.28
r210 33 34 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=3.155 $Y=2.28
+ $X2=2.175 $Y2=2.28
r211 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.595 $Y=0.985
+ $X2=2.68 $Y2=0.9
r212 31 32 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.595 $Y=0.985
+ $X2=2.175 $Y2=0.985
r213 30 66 46.971 $w=5.15e-07 $l=1.65e-07 $layer=POLY_cond $X=1.917 $Y=1.86
+ $X2=1.917 $Y2=1.695
r214 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.01
+ $Y=1.86 $X2=2.01 $Y2=1.86
r215 27 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=2.195
+ $X2=2.175 $Y2=2.28
r216 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.01 $Y=2.195
+ $X2=2.01 $Y2=1.86
r217 26 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=1.07
+ $X2=2.175 $Y2=0.985
r218 26 29 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.01 $Y=1.07
+ $X2=2.01 $Y2=1.86
r219 22 24 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.62 $Y=1.31
+ $X2=1.735 $Y2=1.31
r220 19 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.31
r221 19 66 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.735 $Y=1.385
+ $X2=1.735 $Y2=1.695
r222 18 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.62 $Y=1.235
+ $X2=1.62 $Y2=1.31
r223 17 18 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.62 $Y=0.255
+ $X2=1.62 $Y2=1.235
r224 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.545 $Y=0.18
+ $X2=1.62 $Y2=0.255
r225 15 16 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.545 $Y=0.18
+ $X2=0.565 $Y2=0.18
r226 11 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.375
r227 11 13 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=2.4
r228 10 21 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.49 $Y=0.93
+ $X2=0.49 $Y2=1.375
r229 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.49 $Y=0.255
+ $X2=0.565 $Y2=0.18
r230 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.49 $Y=0.255
+ $X2=0.49 $Y2=0.93
r231 2 52 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.235
+ $Y=2.12 $X2=4.37 $Y2=2.255
r232 1 63 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.625 $X2=6.05 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_410_58# 1 2 9 11 12 13 15 17 18 19 21 23 25
+ 27 29 34 35 38 39
c137 34 0 3.59827e-20 $X=4.88 $Y=1.26
c138 9 0 3.12094e-19 $X=2.125 $Y=0.79
r139 38 39 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=2.465
+ $X2=6.33 $Y2=2.465
r140 33 35 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=1.26
+ $X2=5.13 $Y2=1.26
r141 33 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=1.26
+ $X2=4.88 $Y2=1.26
r142 30 41 12.5376 $w=3.46e-07 $l=9e-08 $layer=POLY_cond $X=2.69 $Y=1.47
+ $X2=2.69 $Y2=1.38
r143 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.47 $X2=2.665 $Y2=1.47
r144 27 39 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.215 $Y=2.405
+ $X2=6.33 $Y2=2.405
r145 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.13 $Y=2.32
+ $X2=5.215 $Y2=2.405
r146 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=1.425
+ $X2=5.13 $Y2=1.26
r147 24 25 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=5.13 $Y=1.425
+ $X2=5.13 $Y2=2.32
r148 23 34 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=3.945 $Y=1.18 $X2=4.88
+ $Y2=1.18
r149 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.86 $Y=1.095
+ $X2=3.945 $Y2=1.18
r150 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.86 $Y=0.765
+ $X2=3.86 $Y2=1.095
r151 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.775 $Y=0.68
+ $X2=3.86 $Y2=0.765
r152 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.775 $Y=0.68
+ $X2=3.105 $Y2=0.68
r153 17 29 14.8322 $w=2.92e-07 $l=4.42674e-07 $layer=LI1_cond $X=3.02 $Y=1.24
+ $X2=2.665 $Y2=1.437
r154 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=0.765
+ $X2=3.105 $Y2=0.68
r155 16 17 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.02 $Y=0.765
+ $X2=3.02 $Y2=1.24
r156 13 30 50.0541 $w=3.46e-07 $l=3.2619e-07 $layer=POLY_cond $X=2.79 $Y=1.75
+ $X2=2.69 $Y2=1.47
r157 13 15 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=2.79 $Y=1.75
+ $X2=2.79 $Y2=2.4
r158 11 41 22.3532 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.5 $Y=1.38
+ $X2=2.69 $Y2=1.38
r159 11 12 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.5 $Y=1.38 $X2=2.2
+ $Y2=1.38
r160 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=1.305
+ $X2=2.2 $Y2=1.38
r161 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.125 $Y=1.305
+ $X2=2.125 $Y2=0.79
r162 2 38 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=6.36
+ $Y=1.865 $X2=6.495 $Y2=2.475
r163 1 33 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=4.905
+ $Y=0.835 $X2=5.045 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_231_132# 1 2 3 4 13 15 18 20 23 28 31 32 33
+ 35 39 42 43 45 48 49 51 52 54 56 57 58 62 67 68 70 71 73 79
c240 68 0 2.42155e-20 $X=4.175 $Y=1.52
c241 67 0 7.86143e-20 $X=4.175 $Y=1.52
c242 57 0 1.55643e-19 $X=1.5 $Y=1.95
c243 56 0 4.00034e-20 $X=1.41 $Y=2.115
c244 33 0 3.05363e-20 $X=3.46 $Y=2.71
c245 23 0 2.93543e-19 $X=1.505 $Y=1.155
r246 78 79 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.96 $Y=2.902
+ $X2=6.125 $Y2=2.902
r247 73 75 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.55 $Y=1.03 $X2=5.55
+ $Y2=1.12
r248 67 70 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=1.6
+ $X2=4.34 $Y2=1.6
r249 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.175
+ $Y=1.52 $X2=4.175 $Y2=1.52
r250 62 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.545 $Y=2.71
+ $X2=3.545 $Y2=2.99
r251 58 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.9 $Y=2.62 $X2=2.9
+ $Y2=2.71
r252 56 57 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.5 $Y=2.115
+ $X2=1.5 $Y2=1.95
r253 53 54 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.915 $Y=2.12
+ $X2=6.915 $Y2=2.905
r254 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.915 $Y2=2.12
r255 51 52 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.225 $Y2=2.035
r256 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=2.99
+ $X2=6.915 $Y2=2.905
r257 49 79 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.83 $Y=2.99
+ $X2=6.125 $Y2=2.99
r258 48 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.14 $Y=1.95
+ $X2=6.225 $Y2=2.035
r259 47 48 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.14 $Y=1.205
+ $X2=6.14 $Y2=1.95
r260 46 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=1.12
+ $X2=5.55 $Y2=1.12
r261 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.055 $Y=1.12
+ $X2=6.14 $Y2=1.205
r262 45 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.055 $Y=1.12
+ $X2=5.715 $Y2=1.12
r263 44 71 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=2.902
+ $X2=4.79 $Y2=2.902
r264 43 78 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=5.953 $Y=2.902
+ $X2=5.96 $Y2=2.902
r265 43 44 36.0097 $w=3.43e-07 $l=1.078e-06 $layer=LI1_cond $X=5.953 $Y=2.902
+ $X2=4.875 $Y2=2.902
r266 42 71 2.87242 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.79 $Y=2.73
+ $X2=4.79 $Y2=2.902
r267 41 42 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=4.79 $Y=1.765
+ $X2=4.79 $Y2=2.73
r268 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.705 $Y=1.68
+ $X2=4.79 $Y2=1.765
r269 39 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.705 $Y=1.68
+ $X2=4.34 $Y2=1.68
r270 36 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=2.99
+ $X2=3.545 $Y2=2.99
r271 35 71 3.6114 $w=2.57e-07 $l=1.23386e-07 $layer=LI1_cond $X=4.705 $Y=2.99
+ $X2=4.79 $Y2=2.902
r272 35 36 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=4.705 $Y=2.99
+ $X2=3.63 $Y2=2.99
r273 34 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=2.71
+ $X2=2.9 $Y2=2.71
r274 33 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.71
+ $X2=3.545 $Y2=2.71
r275 33 34 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.46 $Y=2.71
+ $X2=2.985 $Y2=2.71
r276 31 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=2.62
+ $X2=2.9 $Y2=2.62
r277 31 32 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.815 $Y=2.62
+ $X2=1.675 $Y2=2.62
r278 29 57 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.59 $Y=1.24
+ $X2=1.59 $Y2=1.95
r279 28 32 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.5 $Y=2.535
+ $X2=1.675 $Y2=2.62
r280 27 56 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=1.5 $Y=2.125 $X2=1.5
+ $Y2=2.115
r281 27 28 13.5 $w=3.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.5 $Y=2.125 $X2=1.5
+ $Y2=2.535
r282 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.155
+ $X2=1.59 $Y2=1.24
r283 23 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.505 $Y=1.155
+ $X2=1.31 $Y2=1.155
r284 20 68 81.236 $w=4.45e-07 $l=6.5e-07 $layer=POLY_cond $X=3.525 $Y=1.462
+ $X2=4.175 $Y2=1.462
r285 20 22 17.4857 $w=4.45e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.525 $Y=1.462
+ $X2=3.435 $Y2=1.537
r286 16 22 11.9456 $w=1.8e-07 $l=1.48e-07 $layer=POLY_cond $X=3.435 $Y=1.685
+ $X2=3.435 $Y2=1.537
r287 16 18 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=3.435 $Y=1.685
+ $X2=3.435 $Y2=2.385
r288 13 22 52.5489 $w=2.66e-07 $l=4.17539e-07 $layer=POLY_cond $X=3.145 $Y=1.24
+ $X2=3.435 $Y2=1.537
r289 13 15 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.145 $Y=1.24
+ $X2=3.145 $Y2=0.84
r290 4 78 300 $w=1.7e-07 $l=9.72214e-07 $layer=licon1_PDIFF $count=2 $X=5.295
+ $Y=2.12 $X2=5.96 $Y2=2.815
r291 3 56 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=1.275
+ $Y=1.9 $X2=1.41 $Y2=2.115
r292 2 73 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=5.41
+ $Y=0.625 $X2=5.55 $Y2=1.03
r293 1 25 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.66 $X2=1.31 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_811_379# 1 2 7 9 10 11 13 17 18 19 23 24 26
+ 28 31 33 34 36 41 42 46 49 50 53 56 57
c197 49 0 1.02214e-19 $X=8.78 $Y=2.035
c198 41 0 4.59067e-20 $X=5.785 $Y=1.54
r199 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.925 $Y=2.035
+ $X2=8.925 $Y2=2.035
r200 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r201 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r202 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.78 $Y=2.035
+ $X2=8.925 $Y2=2.035
r203 49 50 3.85519 $w=1.4e-07 $l=3.115e-06 $layer=MET1_cond $X=8.78 $Y=2.035
+ $X2=5.665 $Y2=2.035
r204 46 48 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=10.65 $Y=0.82
+ $X2=10.65 $Y2=1.05
r205 44 57 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.945 $Y=2.565
+ $X2=8.945 $Y2=2.035
r206 42 61 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.785 $Y=1.54
+ $X2=5.785 $Y2=1.715
r207 42 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.785 $Y=1.54
+ $X2=5.785 $Y2=1.375
r208 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.785
+ $Y=1.54 $X2=5.785 $Y2=1.54
r209 38 53 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.52 $Y=1.705
+ $X2=5.52 $Y2=2.035
r210 37 41 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.785 $Y2=1.54
r211 37 38 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.52 $Y2=1.705
r212 36 48 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=10.73 $Y=2.565
+ $X2=10.73 $Y2=1.05
r213 34 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.11 $Y=2.65
+ $X2=8.945 $Y2=2.565
r214 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.645 $Y=2.65
+ $X2=10.73 $Y2=2.565
r215 33 34 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=10.645 $Y=2.65
+ $X2=9.11 $Y2=2.65
r216 29 31 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.655 $Y=1.625
+ $X2=4.83 $Y2=1.625
r217 26 28 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=6.27 $Y=1.79
+ $X2=6.27 $Y2=2.285
r218 25 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.715
+ $X2=5.785 $Y2=1.715
r219 24 26 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.18 $Y=1.715
+ $X2=6.27 $Y2=1.79
r220 24 25 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.18 $Y=1.715
+ $X2=5.95 $Y2=1.715
r221 23 60 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.765 $Y=0.945
+ $X2=5.765 $Y2=1.375
r222 20 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.765 $Y=0.255
+ $X2=5.765 $Y2=0.945
r223 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.69 $Y=0.18
+ $X2=5.765 $Y2=0.255
r224 18 19 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.69 $Y=0.18
+ $X2=4.905 $Y2=0.18
r225 15 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.83 $Y=1.55
+ $X2=4.83 $Y2=1.625
r226 15 17 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.83 $Y=1.55
+ $X2=4.83 $Y2=1.155
r227 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.905 $Y2=0.18
r228 14 17 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.83 $Y2=1.155
r229 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.655 $Y=1.7
+ $X2=4.655 $Y2=1.625
r230 12 13 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.655 $Y=1.7
+ $X2=4.655 $Y2=1.895
r231 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=1.97
+ $X2=4.655 $Y2=1.895
r232 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.58 $Y=1.97
+ $X2=4.235 $Y2=1.97
r233 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.145 $Y=2.045
+ $X2=4.235 $Y2=1.97
r234 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=4.145 $Y=2.045
+ $X2=4.145 $Y2=2.54
r235 2 57 300 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_PDIFF $count=2 $X=8.76
+ $Y=1.87 $X2=8.945 $Y2=2.075
r236 1 46 182 $w=1.7e-07 $l=6.20806e-07 $layer=licon1_NDIFF $count=1 $X=10.18
+ $Y=0.47 $X2=10.65 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_1023_379# 1 2 10 13 15 16 17 19 20 21 25 28
+ 31 34 35 39 43 49 51 52 53 54 57 60 61 66 69
c197 34 0 1.45758e-19 $X=6.9 $Y=0.875
c198 21 0 2.11227e-20 $X=6.34 $Y=1.325
r199 61 70 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.1 $Y=1.665
+ $X2=11.1 $Y2=1.78
r200 61 69 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.1 $Y=1.665
+ $X2=11.1 $Y2=1.55
r201 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.1 $Y=1.665
+ $X2=11.1 $Y2=1.665
r202 57 66 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.55
r203 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.665
+ $X2=6.96 $Y2=1.665
r204 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=1.665
+ $X2=6.96 $Y2=1.665
r205 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.955 $Y=1.665
+ $X2=11.1 $Y2=1.665
r206 53 54 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=10.955 $Y=1.665
+ $X2=7.105 $Y2=1.665
r207 51 66 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=6.955 $Y=1.38
+ $X2=6.955 $Y2=1.55
r208 49 70 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=11.07 $Y=1.98
+ $X2=11.07 $Y2=1.78
r209 45 69 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=11.07 $Y=0.425
+ $X2=11.07 $Y2=1.55
r210 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.985 $Y=0.34
+ $X2=11.07 $Y2=0.425
r211 43 52 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=10.985 $Y=0.34
+ $X2=9.385 $Y2=0.34
r212 39 52 5.72867 $w=1.93e-07 $l=9.7e-08 $layer=LI1_cond $X=9.288 $Y=0.352
+ $X2=9.385 $Y2=0.352
r213 39 41 8.41772 $w=1.93e-07 $l=1.48e-07 $layer=LI1_cond $X=9.288 $Y=0.352
+ $X2=9.14 $Y2=0.352
r214 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.9
+ $Y=0.875 $X2=6.9 $Y2=0.875
r215 32 51 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.9 $Y=1.215
+ $X2=6.9 $Y2=1.38
r216 32 34 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.9 $Y=1.215
+ $X2=6.9 $Y2=0.875
r217 30 35 61.826 $w=3.5e-07 $l=3.75e-07 $layer=POLY_cond $X=6.91 $Y=1.25
+ $X2=6.91 $Y2=0.875
r218 30 31 12.4285 $w=2.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.91 $Y=1.25
+ $X2=6.925 $Y2=1.325
r219 23 25 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=7.025 $Y=3.075
+ $X2=7.025 $Y2=2.285
r220 22 31 12.4285 $w=2.65e-07 $l=1.32288e-07 $layer=POLY_cond $X=7.025 $Y=1.4
+ $X2=6.925 $Y2=1.325
r221 22 25 344.008 $w=1.8e-07 $l=8.85e-07 $layer=POLY_cond $X=7.025 $Y=1.4
+ $X2=7.025 $Y2=2.285
r222 20 31 13.6393 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.735 $Y=1.325
+ $X2=6.925 $Y2=1.325
r223 20 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.735 $Y=1.325
+ $X2=6.34 $Y2=1.325
r224 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.265 $Y=1.25
+ $X2=6.34 $Y2=1.325
r225 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.265 $Y=1.25
+ $X2=6.265 $Y2=0.855
r226 15 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.935 $Y=3.15
+ $X2=7.025 $Y2=3.075
r227 15 16 840.936 $w=1.5e-07 $l=1.64e-06 $layer=POLY_cond $X=6.935 $Y=3.15
+ $X2=5.295 $Y2=3.15
r228 11 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.335 $Y=1.895
+ $X2=5.335 $Y2=1.97
r229 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.335 $Y=1.895
+ $X2=5.335 $Y2=0.945
r230 8 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.205 $Y=3.075
+ $X2=5.295 $Y2=3.15
r231 8 10 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=5.205 $Y=3.075
+ $X2=5.205 $Y2=2.54
r232 7 28 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=5.205 $Y=1.97
+ $X2=5.335 $Y2=1.97
r233 7 10 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.205 $Y=2.045
+ $X2=5.205 $Y2=2.54
r234 2 49 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=10.935
+ $Y=1.84 $X2=11.07 $Y2=1.98
r235 1 41 182 $w=1.7e-07 $l=3.48569e-07 $layer=licon1_NDIFF $count=1 $X=8.84
+ $Y=0.47 $X2=9.14 $Y2=0.365
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_879_55# 1 2 3 12 16 18 20 21 25 27 31 36 38
+ 41 44 45 49 55 56 57 58 61 63 65 67 69 77
c187 61 0 2.52778e-19 $X=8.675 $Y=1.545
c188 27 0 3.59827e-20 $X=7.235 $Y=0.34
r189 68 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.31 $Y=1.385
+ $X2=10.475 $Y2=1.385
r190 68 74 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=10.31 $Y=1.385
+ $X2=10.105 $Y2=1.385
r191 67 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.31 $Y=1.385
+ $X2=10.31 $Y2=1.22
r192 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.31
+ $Y=1.385 $X2=10.31 $Y2=1.385
r193 61 73 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.545
+ $X2=8.675 $Y2=1.71
r194 61 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.545
+ $X2=8.675 $Y2=1.38
r195 60 63 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=8.675 $Y=1.545
+ $X2=8.89 $Y2=1.545
r196 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.675
+ $Y=1.545 $X2=8.675 $Y2=1.545
r197 56 58 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=7.415 $Y=1.95
+ $X2=7.415 $Y2=1.13
r198 55 56 6.19221 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=7.335 $Y=2.05
+ $X2=7.335 $Y2=1.95
r199 49 52 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.58 $Y=0.34 $X2=4.58
+ $Y2=0.42
r200 47 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.23 $Y=0.79
+ $X2=10.23 $Y2=1.22
r201 46 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.975 $Y=0.705
+ $X2=8.89 $Y2=0.705
r202 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=0.705
+ $X2=10.23 $Y2=0.79
r203 45 46 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=10.145 $Y=0.705
+ $X2=8.975 $Y2=0.705
r204 44 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.89 $Y=1.38
+ $X2=8.89 $Y2=1.545
r205 43 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=0.79
+ $X2=8.89 $Y2=0.705
r206 43 44 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.89 $Y=0.79
+ $X2=8.89 $Y2=1.38
r207 42 57 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.565 $Y=0.705
+ $X2=7.4 $Y2=0.705
r208 41 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.805 $Y=0.705
+ $X2=8.89 $Y2=0.705
r209 41 42 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=8.805 $Y=0.705
+ $X2=7.565 $Y2=0.705
r210 38 58 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=0.965
+ $X2=7.4 $Y2=1.13
r211 37 57 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.79 $X2=7.4
+ $Y2=0.705
r212 37 38 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.4 $Y=0.79
+ $X2=7.4 $Y2=0.965
r213 34 57 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.62 $X2=7.4
+ $Y2=0.705
r214 34 36 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.4 $Y=0.62
+ $X2=7.4 $Y2=0.515
r215 33 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.4 $Y=0.425 $X2=7.4
+ $Y2=0.515
r216 29 55 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=7.335 $Y=2.115
+ $X2=7.335 $Y2=2.05
r217 29 31 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=7.335 $Y=2.115
+ $X2=7.335 $Y2=2.76
r218 28 49 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.705 $Y=0.34
+ $X2=4.58 $Y2=0.34
r219 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.235 $Y=0.34
+ $X2=7.4 $Y2=0.425
r220 27 28 165.059 $w=1.68e-07 $l=2.53e-06 $layer=LI1_cond $X=7.235 $Y=0.34
+ $X2=4.705 $Y2=0.34
r221 23 25 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=10.845 $Y=1.55
+ $X2=10.845 $Y2=2.26
r222 21 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=10.755 $Y=1.475
+ $X2=10.845 $Y2=1.55
r223 21 77 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.755 $Y=1.475
+ $X2=10.475 $Y2=1.475
r224 18 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.105 $Y=1.22
+ $X2=10.105 $Y2=1.385
r225 18 20 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.105 $Y=1.22
+ $X2=10.105 $Y2=0.79
r226 16 72 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.765 $Y=0.79
+ $X2=8.765 $Y2=1.38
r227 12 73 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=8.67 $Y=2.29
+ $X2=8.67 $Y2=1.71
r228 3 55 300 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_PDIFF $count=2 $X=7.115
+ $Y=1.865 $X2=7.335 $Y2=2.05
r229 3 31 600 $w=1.7e-07 $l=9.98962e-07 $layer=licon1_PDIFF $count=1 $X=7.115
+ $Y=1.865 $X2=7.335 $Y2=2.76
r230 2 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.255
+ $Y=0.37 $X2=7.4 $Y2=0.515
r231 1 52 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.275 $X2=4.54 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%B 1 3 6 8 11 12 13 17 18 20 22 25 30 31 32 34
+ 35 42
c130 35 0 1.50564e-19 $X=9.36 $Y=1.295
c131 8 0 1.01602e-19 $X=8.055 $Y=1.635
c132 6 0 1.45758e-19 $X=7.615 $Y=0.74
r133 40 42 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.31 $Y=1.385
+ $X2=9.515 $Y2=1.385
r134 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.31
+ $Y=1.385 $X2=9.31 $Y2=1.385
r135 37 40 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=9.17 $Y=1.385
+ $X2=9.31 $Y2=1.385
r136 35 41 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.31 $Y=1.295
+ $X2=9.31 $Y2=1.385
r137 33 34 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=11.292 $Y=1.35
+ $X2=11.292 $Y2=1.5
r138 30 34 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=11.295 $Y=2.26
+ $X2=11.295 $Y2=1.5
r139 28 30 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=11.295 $Y=3.075
+ $X2=11.295 $Y2=2.26
r140 25 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.275 $Y=0.79
+ $X2=11.275 $Y2=1.35
r141 20 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.515 $Y=1.22
+ $X2=9.515 $Y2=1.385
r142 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.515 $Y=1.22
+ $X2=9.515 $Y2=0.79
r143 19 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.26 $Y=3.15 $X2=9.17
+ $Y2=3.15
r144 18 28 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.205 $Y=3.15
+ $X2=11.295 $Y2=3.075
r145 18 19 997.33 $w=1.5e-07 $l=1.945e-06 $layer=POLY_cond $X=11.205 $Y=3.15
+ $X2=9.26 $Y2=3.15
r146 15 32 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.17 $Y=3.075
+ $X2=9.17 $Y2=3.15
r147 15 17 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=9.17 $Y=3.075
+ $X2=9.17 $Y2=2.29
r148 14 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.17 $Y=1.55
+ $X2=9.17 $Y2=1.385
r149 14 17 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=9.17 $Y=1.55
+ $X2=9.17 $Y2=2.29
r150 12 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.08 $Y=3.15 $X2=9.17
+ $Y2=3.15
r151 12 13 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=9.08 $Y=3.15
+ $X2=8.205 $Y2=3.15
r152 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.13 $Y=3.075
+ $X2=8.205 $Y2=3.15
r153 10 11 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=8.13 $Y=1.71
+ $X2=8.13 $Y2=3.075
r154 9 31 6.66866 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=7.69 $Y=1.635
+ $X2=7.58 $Y2=1.635
r155 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.055 $Y=1.635
+ $X2=8.13 $Y2=1.71
r156 8 9 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=8.055 $Y=1.635
+ $X2=7.69 $Y2=1.635
r157 4 31 18.8402 $w=1.65e-07 $l=9.08295e-08 $layer=POLY_cond $X=7.615 $Y=1.56
+ $X2=7.58 $Y2=1.635
r158 4 6 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.615 $Y=1.56
+ $X2=7.615 $Y2=0.74
r159 1 31 18.8402 $w=1.65e-07 $l=8.44097e-08 $layer=POLY_cond $X=7.56 $Y=1.71
+ $X2=7.58 $Y2=1.635
r160 1 3 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=7.56 $Y=1.71
+ $X2=7.56 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_2342_48# 1 2 7 9 12 15 16 20 24 28 32 35 36
+ 37
c78 28 0 1.0013e-19 $X=12.415 $Y=1.215
r79 35 36 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=13.65 $Y=2.135
+ $X2=13.65 $Y2=1.97
r80 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.415
+ $Y=1.385 $X2=12.415 $Y2=1.385
r81 28 31 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.415 $Y=1.215
+ $X2=12.415 $Y2=1.385
r82 26 37 3.55013 $w=2.62e-07 $l=1.28662e-07 $layer=LI1_cond $X=13.745 $Y=1.3
+ $X2=13.652 $Y2=1.215
r83 26 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.745 $Y=1.3
+ $X2=13.745 $Y2=1.97
r84 22 37 3.55013 $w=2.62e-07 $l=8.5e-08 $layer=LI1_cond $X=13.652 $Y=1.13
+ $X2=13.652 $Y2=1.215
r85 22 24 19.9649 $w=3.53e-07 $l=6.15e-07 $layer=LI1_cond $X=13.652 $Y=1.13
+ $X2=13.652 $Y2=0.515
r86 18 35 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=13.65 $Y=2.15
+ $X2=13.65 $Y2=2.135
r87 18 20 21.2882 $w=3.58e-07 $l=6.65e-07 $layer=LI1_cond $X=13.65 $Y=2.15
+ $X2=13.65 $Y2=2.815
r88 17 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.58 $Y=1.215
+ $X2=12.415 $Y2=1.215
r89 16 37 2.9446 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=13.475 $Y=1.215
+ $X2=13.652 $Y2=1.215
r90 16 17 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=13.475 $Y=1.215
+ $X2=12.58 $Y2=1.215
r91 14 32 91.8022 $w=3.3e-07 $l=5.25e-07 $layer=POLY_cond $X=11.89 $Y=1.385
+ $X2=12.415 $Y2=1.385
r92 14 15 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.89 $Y=1.385
+ $X2=11.8 $Y2=1.385
r93 10 15 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=11.8 $Y=1.55
+ $X2=11.8 $Y2=1.385
r94 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=11.8 $Y=1.55
+ $X2=11.8 $Y2=2.4
r95 7 15 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=11.785 $Y=1.22
+ $X2=11.8 $Y2=1.385
r96 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.785 $Y=1.22
+ $X2=11.785 $Y2=0.74
r97 2 35 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.96 $X2=13.635 $Y2=2.135
r98 2 20 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.96 $X2=13.635 $Y2=2.815
r99 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.37 $X2=13.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A 3 7 11 15 17 24 26
c47 26 0 1.0013e-19 $X=13.425 $Y=1.635
r48 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=13.41 $Y=1.635
+ $X2=13.425 $Y2=1.635
r49 23 25 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=13.325 $Y=1.635
+ $X2=13.41 $Y2=1.635
r50 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.325
+ $Y=1.635 $X2=13.325 $Y2=1.635
r51 21 23 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=12.91 $Y=1.635
+ $X2=13.325 $Y2=1.635
r52 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.895 $Y=1.635
+ $X2=12.91 $Y2=1.635
r53 17 24 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=13.2 $Y=1.635
+ $X2=13.325 $Y2=1.635
r54 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.425 $Y=1.47
+ $X2=13.425 $Y2=1.635
r55 13 15 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=13.425 $Y=1.47
+ $X2=13.425 $Y2=0.69
r56 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.41 $Y=1.8
+ $X2=13.41 $Y2=1.635
r57 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=13.41 $Y=1.8
+ $X2=13.41 $Y2=2.46
r58 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.91 $Y=1.8
+ $X2=12.91 $Y2=1.635
r59 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=12.91 $Y=1.8 $X2=12.91
+ $Y2=2.46
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.895 $Y=1.47
+ $X2=12.895 $Y2=1.635
r61 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.895 $Y=1.47
+ $X2=12.895 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%SUM 1 2 7 8 9 10 11 18
r17 10 11 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=2.405
+ $X2=0.277 $Y2=2.775
r18 9 10 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=0.277 $Y=1.985
+ $X2=0.277 $Y2=2.405
r19 8 9 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.985
r20 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.665
r21 7 18 20.2968 $w=3.33e-07 $l=5.9e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=0.705
r22 2 11 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r23 2 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r24 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.56 $X2=0.275 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%VPWR 1 2 3 4 5 20 24 28 31 36 43 44 45 47 55
+ 67 73 74 77 80 87 90
c131 80 0 3.05634e-20 $X=3.11 $Y=3.05
r132 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r133 87 88 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r135 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r136 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r137 71 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.3 $Y=3.33
+ $X2=13.175 $Y2=3.33
r138 71 73 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=13.3 $Y=3.33
+ $X2=13.68 $Y2=3.33
r139 70 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r140 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r141 67 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.05 $Y=3.33
+ $X2=13.175 $Y2=3.33
r142 67 69 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=13.05 $Y=3.33
+ $X2=12.72 $Y2=3.33
r143 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r144 66 88 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=7.92 $Y2=3.33
r145 65 66 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r146 63 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8 $Y=3.33 $X2=7.835
+ $Y2=3.33
r147 63 65 245.305 $w=1.68e-07 $l=3.76e-06 $layer=LI1_cond $X=8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r148 62 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r149 61 62 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r150 59 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r151 58 61 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r152 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r153 56 58 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 55 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.67 $Y=3.33
+ $X2=7.835 $Y2=3.33
r155 55 61 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.67 $Y=3.33
+ $X2=7.44 $Y2=3.33
r156 54 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r157 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r158 51 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r159 51 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r160 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r161 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r162 48 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r163 48 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r164 47 56 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=3.112 $Y=3.33
+ $X2=3.29 $Y2=3.33
r165 47 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r166 47 80 9.08969 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=3.112 $Y=3.33
+ $X2=3.112 $Y2=3.05
r167 47 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=2.64 $Y2=3.33
r168 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r169 45 59 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=3.6 $Y2=3.33
r170 43 65 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=11.76 $Y2=3.33
r171 43 44 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=12.12 $Y2=3.33
r172 42 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.29 $Y=3.33
+ $X2=12.72 $Y2=3.33
r173 42 44 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.29 $Y=3.33
+ $X2=12.12 $Y2=3.33
r174 36 39 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=13.175 $Y=2.135
+ $X2=13.175 $Y2=2.815
r175 34 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.175 $Y=3.245
+ $X2=13.175 $Y2=3.33
r176 34 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.175 $Y=3.245
+ $X2=13.175 $Y2=2.815
r177 31 33 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=12.12 $Y=2.615
+ $X2=12.12 $Y2=2.955
r178 29 44 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.12 $Y=3.245
+ $X2=12.12 $Y2=3.33
r179 29 33 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=12.12 $Y=3.245
+ $X2=12.12 $Y2=2.955
r180 28 41 8.27282 $w=3.4e-07 $l=2.25e-07 $layer=LI1_cond $X=12.12 $Y=2.5
+ $X2=12.12 $Y2=2.275
r181 28 31 3.89797 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=12.12 $Y=2.5
+ $X2=12.12 $Y2=2.615
r182 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.835 $Y=1.93
+ $X2=7.835 $Y2=2.76
r183 22 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=3.33
r184 22 27 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=2.76
r185 18 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r186 18 20 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r187 5 39 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=13
+ $Y=1.96 $X2=13.135 $Y2=2.815
r188 5 36 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=13
+ $Y=1.96 $X2=13.135 $Y2=2.135
r189 4 41 600 $w=1.7e-07 $l=5.35817e-07 $layer=licon1_PDIFF $count=1 $X=11.89
+ $Y=1.84 $X2=12.115 $Y2=2.275
r190 4 33 600 $w=1.7e-07 $l=1.22233e-06 $layer=licon1_PDIFF $count=1 $X=11.89
+ $Y=1.84 $X2=12.115 $Y2=2.955
r191 4 31 600 $w=1.7e-07 $l=8.80341e-07 $layer=licon1_PDIFF $count=1 $X=11.89
+ $Y=1.84 $X2=12.115 $Y2=2.615
r192 3 27 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=7.65
+ $Y=1.785 $X2=7.835 $Y2=2.76
r193 3 24 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.65
+ $Y=1.785 $X2=7.835 $Y2=1.93
r194 2 80 600 $w=1.7e-07 $l=1.32e-06 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.11 $Y2=3.05
r195 1 20 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%COUT 1 2 8 9 10 12 14 17 20 21 23
c72 17 0 1.13036e-19 $X=1.07 $Y=2.035
c73 12 0 1.68941e-19 $X=1.07 $Y=2.905
r74 23 28 7.38421 $w=3.8e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=0.65 $X2=1.91
+ $Y2=0.65
r75 20 21 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.975
+ $X2=2.315 $Y2=2.975
r76 15 17 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.75 $Y=2.035
+ $X2=1.07 $Y2=2.035
r77 14 21 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.155 $Y=2.99
+ $X2=2.315 $Y2=2.99
r78 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=2.905
+ $X2=1.155 $Y2=2.99
r79 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=2.12
+ $X2=1.07 $Y2=2.035
r80 11 12 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.07 $Y=2.12
+ $X2=1.07 $Y2=2.905
r81 9 23 9.3947 $w=3.8e-07 $l=2.43926e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=1.68 $Y2=0.65
r82 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=0.835 $Y2=0.815
r83 8 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.95 $X2=0.75
+ $Y2=2.035
r84 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=0.9
+ $X2=0.835 $Y2=0.815
r85 7 8 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=0.75 $Y=0.9 $X2=0.75
+ $Y2=1.95
r86 2 20 600 $w=1.7e-07 $l=1.19029e-06 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.84 $X2=2.48 $Y2=2.96
r87 1 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.42 $X2=1.91 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_644_104# 1 2 3 11 14 17 20 21 27 28 31
c99 31 0 3.05363e-20 $X=3.36 $Y=1.855
c100 21 0 7.86143e-20 $X=3.265 $Y=1.665
r101 31 33 13.9377 $w=3.37e-07 $l=3.85e-07 $layer=LI1_cond $X=3.36 $Y=1.855
+ $X2=3.745 $Y2=1.855
r102 28 35 6.65862 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=6.495 $Y=1.665
+ $X2=6.495 $Y2=1.55
r103 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r104 24 31 8.68843 $w=3.37e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.855
+ $X2=3.36 $Y2=1.855
r105 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r106 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r107 20 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r108 20 21 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=3.265 $Y2=1.665
r109 17 19 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=1.02
+ $X2=3.44 $Y2=1.185
r110 14 35 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.48 $Y=0.875
+ $X2=6.48 $Y2=1.55
r111 11 31 4.74843 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.36 $Y=1.58
+ $X2=3.36 $Y2=1.855
r112 11 19 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.36 $Y=1.58
+ $X2=3.36 $Y2=1.185
r113 3 33 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.885 $X2=3.745 $Y2=2.03
r114 2 14 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.535 $X2=6.48 $Y2=0.875
r115 1 17 182 $w=1.7e-07 $l=6e-07 $layer=licon1_NDIFF $count=1 $X=3.22 $Y=0.52
+ $X2=3.44 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_1660_374# 1 2 3 4 16 17 18 19 22 25 32 35 36
c89 32 0 1.01602e-19 $X=8.47 $Y=1.045
r90 35 36 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.39 $Y=2.045
+ $X2=8.39 $Y2=1.88
r91 29 32 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=8.255 $Y=1.085
+ $X2=8.47 $Y2=1.085
r92 28 37 5.67621 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=11.572 $Y=0.965
+ $X2=11.572 $Y2=1.13
r93 25 28 15.4806 $w=3.33e-07 $l=4.5e-07 $layer=LI1_cond $X=11.572 $Y=0.515
+ $X2=11.572 $Y2=0.965
r94 20 22 29.7038 $w=3.53e-07 $l=9.15e-07 $layer=LI1_cond $X=11.562 $Y=2.905
+ $X2=11.562 $Y2=1.99
r95 19 37 5.79584 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=11.562 $Y=1.307
+ $X2=11.562 $Y2=1.13
r96 19 22 22.1724 $w=3.53e-07 $l=6.83e-07 $layer=LI1_cond $X=11.562 $Y=1.307
+ $X2=11.562 $Y2=1.99
r97 17 20 7.97992 $w=1.7e-07 $l=2.15346e-07 $layer=LI1_cond $X=11.385 $Y=2.99
+ $X2=11.562 $Y2=2.905
r98 17 18 181.043 $w=1.68e-07 $l=2.775e-06 $layer=LI1_cond $X=11.385 $Y=2.99
+ $X2=8.61 $Y2=2.99
r99 16 18 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=8.39 $Y=2.905
+ $X2=8.61 $Y2=2.99
r100 15 35 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=8.39 $Y=2.1
+ $X2=8.39 $Y2=2.045
r101 15 16 21.0845 $w=4.38e-07 $l=8.05e-07 $layer=LI1_cond $X=8.39 $Y=2.1
+ $X2=8.39 $Y2=2.905
r102 13 29 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.255 $Y=1.21
+ $X2=8.255 $Y2=1.085
r103 13 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.255 $Y=1.21
+ $X2=8.255 $Y2=1.88
r104 4 22 300 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=2 $X=11.385
+ $Y=1.84 $X2=11.545 $Y2=1.99
r105 3 35 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=8.3
+ $Y=1.87 $X2=8.445 $Y2=2.045
r106 2 28 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=11.35
+ $Y=0.47 $X2=11.57 $Y2=0.965
r107 2 25 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=11.35
+ $Y=0.47 $X2=11.57 $Y2=0.515
r108 1 32 182 $w=1.7e-07 $l=6.43428e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.47 $X2=8.47 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%A_1852_374# 1 2 3 4 15 18 19 20 21 22 25 27 29
+ 31 36 37 39 47
r102 45 47 10.1363 $w=5.88e-07 $l=5e-07 $layer=LI1_cond $X=9.81 $Y=2.1 $X2=10.31
+ $Y2=2.1
r103 43 45 6.68993 $w=5.88e-07 $l=3.3e-07 $layer=LI1_cond $X=9.48 $Y=2.1
+ $X2=9.81 $Y2=2.1
r104 40 49 7.22832 $w=3.46e-07 $l=2.05e-07 $layer=LI1_cond $X=12.62 $Y=2.035
+ $X2=12.62 $Y2=1.83
r105 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.52 $Y=2.035
+ $X2=12.52 $Y2=2.035
r106 36 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.375 $Y=2.035
+ $X2=12.52 $Y2=2.035
r107 36 37 2.35148 $w=1.4e-07 $l=1.9e-06 $layer=MET1_cond $X=12.375 $Y=2.035
+ $X2=10.475 $Y2=2.035
r108 33 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.33 $Y=2.035
+ $X2=10.33 $Y2=2.035
r109 31 37 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=10.36 $Y=2.035
+ $X2=10.475 $Y2=2.035
r110 31 33 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=10.36 $Y=2.035
+ $X2=10.33 $Y2=2.035
r111 27 40 4.40751 $w=3.46e-07 $l=1.5411e-07 $layer=LI1_cond $X=12.685 $Y=2.16
+ $X2=12.62 $Y2=2.035
r112 27 29 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=12.685 $Y=2.16
+ $X2=12.685 $Y2=2.815
r113 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.64 $Y=0.79
+ $X2=12.64 $Y2=0.515
r114 21 49 3.38667 $w=2.2e-07 $l=2.3e-07 $layer=LI1_cond $X=12.39 $Y=1.83
+ $X2=12.62 $Y2=1.83
r115 21 22 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=12.39 $Y=1.83
+ $X2=12.08 $Y2=1.83
r116 19 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.475 $Y=0.875
+ $X2=12.64 $Y2=0.79
r117 19 20 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.475 $Y=0.875
+ $X2=12.08 $Y2=0.875
r118 18 22 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.995 $Y=1.72
+ $X2=12.08 $Y2=1.83
r119 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.995 $Y=0.96
+ $X2=12.08 $Y2=0.875
r120 17 18 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=11.995 $Y=0.96
+ $X2=11.995 $Y2=1.72
r121 13 45 4.13774 $w=3.3e-07 $l=2.95e-07 $layer=LI1_cond $X=9.81 $Y=1.805
+ $X2=9.81 $Y2=2.1
r122 13 15 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=9.81 $Y=1.805
+ $X2=9.81 $Y2=1.045
r123 4 40 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.96 $X2=12.685 $Y2=2.135
r124 4 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.96 $X2=12.685 $Y2=2.815
r125 3 47 150 $w=1.7e-07 $l=1.09886e-06 $layer=licon1_PDIFF $count=4 $X=9.26
+ $Y=1.87 $X2=10.31 $Y2=1.97
r126 3 43 300 $w=1.7e-07 $l=2.6533e-07 $layer=licon1_PDIFF $count=2 $X=9.26
+ $Y=1.87 $X2=9.48 $Y2=1.97
r127 2 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.495
+ $Y=0.37 $X2=12.64 $Y2=0.515
r128 1 15 182 $w=1.7e-07 $l=6.7611e-07 $layer=licon1_NDIFF $count=1 $X=9.59
+ $Y=0.47 $X2=9.81 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 56 70 76 77 80 83 86
r120 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r121 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r122 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 77 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r124 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r125 74 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.14 $Y2=0
r126 74 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.68 $Y2=0
r127 73 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r128 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r129 70 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=13.14 $Y2=0
r130 70 72 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=12.72 $Y2=0
r131 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r132 68 69 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r133 66 69 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=11.76 $Y2=0
r134 66 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r135 65 68 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=11.76
+ $Y2=0
r136 65 66 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r137 63 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r138 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r139 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r140 61 62 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r141 58 61 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=7.44
+ $Y2=0
r142 58 59 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r143 56 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r144 56 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r145 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r146 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r147 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r148 52 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r149 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r150 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r151 49 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r152 49 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r153 47 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r154 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r155 44 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r156 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r157 42 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r158 42 59 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=2.64
+ $Y2=0
r159 40 68 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=11.76 $Y2=0
r160 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=12.08 $Y2=0
r161 39 72 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=12.245 $Y=0
+ $X2=12.72 $Y2=0
r162 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=0
+ $X2=12.08 $Y2=0
r163 37 54 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.16
+ $Y2=0
r164 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.34
+ $Y2=0
r165 36 58 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.425 $Y=0
+ $X2=2.64 $Y2=0
r166 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.34
+ $Y2=0
r167 32 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0
r168 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0.515
r169 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.08 $Y=0.085
+ $X2=12.08 $Y2=0
r170 28 30 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.08 $Y=0.085
+ $X2=12.08 $Y2=0.455
r171 24 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r172 24 26 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.365
r173 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0
r174 20 22 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0.565
r175 16 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r176 16 18 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.475
r177 5 34 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=12.97
+ $Y=0.37 $X2=13.14 $Y2=0.515
r178 4 30 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=11.86
+ $Y=0.37 $X2=12.08 $Y2=0.455
r179 3 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.69
+ $Y=0.37 $X2=7.91 $Y2=0.365
r180 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.42 $X2=2.34 $Y2=0.565
r181 1 18 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.56 $X2=0.785 $Y2=0.475
.ends


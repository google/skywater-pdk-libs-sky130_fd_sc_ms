* File: sky130_fd_sc_ms__nor4b_1.spice
* Created: Fri Aug 28 17:49:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4b_1.pex.spice"
.subckt sky130_fd_sc_ms__nor4b_1  VNB VPB D_N A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_D_N_M1004_g N_A_57_368#_M1004_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.11874 AS=0.15675 PD=0.989147 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.15976 PD=1.02 PS=1.33085 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_Y_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.1591
+ AS=0.1036 PD=1.17 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1591 PD=1.02 PS=1.17 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.6 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_57_368#_M1002_g N_Y_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_D_N_M1008_g N_A_57_368#_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.174 AS=0.2352 PD=1.29429 PS=2.24 NRD=26.9693 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1006 A_263_368# N_A_M1006_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.232 PD=1.36 PS=1.72571 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1001 A_347_368# N_B_M1001_g A_263_368# VPB PSHORT L=0.18 W=1.12 AD=0.1848
+ AS=0.1344 PD=1.45 PS=1.36 NRD=19.3454 NRS=11.426 M=1 R=6.22222 SA=90001
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1007 A_449_368# N_C_M1007_g A_347_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1848 PD=1.51 PS=1.45 NRD=24.6053 NRS=19.3454 M=1 R=6.22222 SA=90001.5
+ SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_A_57_368#_M1005_g A_449_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.448 AS=0.2184 PD=3.04 PS=1.51 NRD=20.2122 NRS=24.6053 M=1 R=6.22222
+ SA=90002.1 SB=90000.3 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__nor4b_1.pxi.spice"
*
.ends
*
*

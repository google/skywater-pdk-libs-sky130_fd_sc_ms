* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_755_74# a_797_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_565_392# a_243_394# a_640_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 a_640_74# a_364_120# a_750_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X3 Q a_797_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR GATE a_243_394# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 a_938_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VGND GATE a_243_394# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND a_797_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_364_120# a_243_394# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X9 Q a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_797_48# a_640_74# a_938_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VPWR a_640_74# a_797_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X12 VGND a_797_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_27_126# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X14 a_797_48# a_640_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X15 VGND RESET_B a_938_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 VPWR a_797_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 Q a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 Q a_797_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR RESET_B a_797_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X20 a_750_508# a_797_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X21 a_559_74# a_364_120# a_640_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 VPWR a_797_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 a_27_126# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X24 VPWR a_27_126# a_565_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X25 a_364_120# a_243_394# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_938_74# a_640_74# a_797_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 VGND a_27_126# a_559_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 a_797_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X29 a_640_74# a_243_394# a_755_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

* File: sky130_fd_sc_ms__a221oi_1.pex.spice
* Created: Wed Sep  2 11:52:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A221OI_1%C1 3 7 9 13 14
c27 14 0 1.63146e-19 $X=0.71 $Y=1.515
r28 13 15 64.567 $w=3.21e-07 $l=4.3e-07 $layer=POLY_cond $X=0.71 $Y=1.515
+ $X2=1.14 $Y2=1.515
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.515 $X2=0.71 $Y2=1.515
r30 11 13 29.2804 $w=3.21e-07 $l=1.95e-07 $layer=POLY_cond $X=0.515 $Y=1.515
+ $X2=0.71 $Y2=1.515
r31 9 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=1.515
r32 5 15 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.35
+ $X2=1.14 $Y2=1.515
r33 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.14 $Y=1.35 $X2=1.14
+ $Y2=0.74
r34 1 11 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.68
+ $X2=0.515 $Y2=1.515
r35 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.515 $Y=1.68
+ $X2=0.515 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%B2 3 7 9 10 14
c35 14 0 1.63146e-19 $X=1.59 $Y=1.515
r36 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.515
+ $X2=1.59 $Y2=1.68
r37 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.515
+ $X2=1.59 $Y2=1.35
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.59
+ $Y=1.515 $X2=1.59 $Y2=1.515
r39 10 15 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.59
+ $Y2=1.565
r40 9 15 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1.59
+ $Y2=1.565
r41 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.68 $Y=0.74 $X2=1.68
+ $Y2=1.35
r42 3 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.665 $Y=2.4
+ $X2=1.665 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%B1 3 7 9 12 13
c39 7 0 1.10616e-19 $X=2.115 $Y=2.4
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r44 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.115 $Y=2.4
+ $X2=2.115 $Y2=1.68
r45 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.04 $Y=0.74 $X2=2.04
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%A1 3 7 9 12 13
c37 13 0 1.10616e-19 $X=2.67 $Y=1.515
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.515
+ $X2=2.67 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.515
+ $X2=2.67 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.515 $X2=2.67 $Y2=1.515
r41 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.515
r42 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.76 $Y=0.74 $X2=2.76
+ $Y2=1.35
r43 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.595 $Y=2.4
+ $X2=2.595 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%A2 3 6 8 9 13 15
r26 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.385
+ $X2=3.21 $Y2=1.55
r27 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.385
+ $X2=3.21 $Y2=1.22
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.385 $X2=3.21 $Y2=1.385
r29 9 14 12.1474 $w=3.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.21
+ $Y2=1.365
r30 8 14 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=1.365 $X2=3.21
+ $Y2=1.365
r31 6 16 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.135 $Y=2.4
+ $X2=3.135 $Y2=1.55
r32 3 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.12 $Y=0.74 $X2=3.12
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%Y 1 2 3 10 14 16 18 19 20 21 22 51
r37 50 51 11.617 $w=8.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0.765
+ $X2=1.09 $Y2=0.765
r38 48 50 9.72714 $w=8.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.25 $Y=0.765
+ $X2=0.925 $Y2=0.765
r39 30 48 7.92413 $w=2.5e-07 $l=4.15e-07 $layer=LI1_cond $X=0.25 $Y=1.18
+ $X2=0.25 $Y2=0.765
r40 21 22 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.775
r41 20 21 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.25 $Y=1.985
+ $X2=0.25 $Y2=2.405
r42 19 20 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=1.985
r43 18 19 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r44 18 30 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.18
r45 16 48 0.144106 $w=8.28e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0.765
+ $X2=0.25 $Y2=0.765
r46 12 14 14.3014 $w=4.13e-07 $l=5.15e-07 $layer=LI1_cond $X=2.367 $Y=1.01
+ $X2=2.367 $Y2=0.495
r47 10 12 8.50155 $w=1.7e-07 $l=2.45854e-07 $layer=LI1_cond $X=2.16 $Y=1.095
+ $X2=2.367 $Y2=1.01
r48 10 51 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=2.16 $Y=1.095
+ $X2=1.09 $Y2=1.095
r49 3 22 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.29 $Y2=2.815
r50 3 20 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.29 $Y2=1.985
r51 2 14 91 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=2 $X=2.115
+ $Y=0.37 $X2=2.375 $Y2=0.495
r52 1 50 45.5 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_NDIFF $count=4 $X=0.46
+ $Y=0.37 $X2=0.925 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%A_121_368# 1 2 9 13 14 17
r26 15 17 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.89 $Y=2.905
+ $X2=1.89 $Y2=2.4
r27 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=2.99
+ $X2=1.89 $Y2=2.905
r28 13 14 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.725 $Y=2.99
+ $X2=0.905 $Y2=2.99
r29 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.74 $Y=2.115 $X2=0.74
+ $Y2=2.815
r30 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.74 $Y=2.905
+ $X2=0.905 $Y2=2.99
r31 7 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.74 $Y=2.905 $X2=0.74
+ $Y2=2.815
r32 2 17 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=1.755
+ $Y=1.84 $X2=1.89 $Y2=2.4
r33 1 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.74 $Y2=2.815
r34 1 9 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.74 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%A_263_368# 1 2 3 10 12 14 18 20 22 24 29
r42 22 31 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=3.36 $Y=2.12 $X2=3.36
+ $Y2=1.97
r43 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.36 $Y=2.12
+ $X2=3.36 $Y2=2.815
r44 21 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=2.38 $Y2=2.035
r45 20 31 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=3.36 $Y2=1.97
r46 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=2.505 $Y2=2.035
r47 16 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=2.38 $Y2=2.035
r48 16 18 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=2.38 $Y2=2.44
r49 15 27 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.545 $Y=2.035
+ $X2=1.41 $Y2=2.035
r50 14 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=2.38 $Y2=2.035
r51 14 15 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=1.545 $Y2=2.035
r52 10 27 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=2.12 $X2=1.41
+ $Y2=2.035
r53 10 12 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.41 $Y=2.12
+ $X2=1.41 $Y2=2.57
r54 3 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.84 $X2=3.36 $Y2=1.985
r55 3 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.84 $X2=3.36 $Y2=2.815
r56 2 29 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.84 $X2=2.34 $Y2=2.035
r57 2 18 300 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_PDIFF $count=2 $X=2.205
+ $Y=1.84 $X2=2.34 $Y2=2.44
r58 1 27 600 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=2.035
r59 1 12 600 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%VPWR 1 6 9 10 11 21 22
r34 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r35 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r36 18 19 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 14 18 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 14 15 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 11 15 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 9 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 9 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.675 $Y=3.33 $X2=2.85
+ $Y2=3.33
r43 8 21 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 8 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.025 $Y=3.33 $X2=2.85
+ $Y2=3.33
r45 4 10 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245 $X2=2.85
+ $Y2=3.33
r46 4 6 27.8233 $w=3.48e-07 $l=8.45e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.4
r47 1 6 300 $w=1.7e-07 $l=6.37181e-07 $layer=licon1_PDIFF $count=2 $X=2.685
+ $Y=1.84 $X2=2.85 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A221OI_1%VGND 1 2 9 13 16 17 19 20 21 37 38
r34 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r35 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r36 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r38 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r39 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r40 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r42 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r43 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 21 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r45 21 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r46 19 34 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.12
+ $Y2=0
r47 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.335
+ $Y2=0
r48 18 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.6 $Y2=0
r49 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.335
+ $Y2=0
r50 16 28 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.2
+ $Y2=0
r51 16 17 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.445
+ $Y2=0
r52 15 31 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.68
+ $Y2=0
r53 15 17 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.445
+ $Y2=0
r54 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0
r55 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0.515
r56 7 17 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=0.085
+ $X2=1.445 $Y2=0
r57 7 9 18.3768 $w=3.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.445 $Y=0.085
+ $X2=1.445 $Y2=0.675
r58 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.195
+ $Y=0.37 $X2=3.335 $Y2=0.515
r59 1 9 182 $w=1.7e-07 $l=4.03949e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.37 $X2=1.445 $Y2=0.675
.ends


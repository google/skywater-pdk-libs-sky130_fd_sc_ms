* File: sky130_fd_sc_ms__o31a_4.pxi.spice
* Created: Wed Sep  2 12:25:42 2020
* 
x_PM_SKY130_FD_SC_MS__O31A_4%A_86_260# N_A_86_260#_M1009_s N_A_86_260#_M1002_d
+ N_A_86_260#_M1012_d N_A_86_260#_M1007_g N_A_86_260#_M1003_g
+ N_A_86_260#_M1006_g N_A_86_260#_M1008_g N_A_86_260#_M1018_g
+ N_A_86_260#_M1011_g N_A_86_260#_M1020_g N_A_86_260#_M1014_g
+ N_A_86_260#_c_138_n N_A_86_260#_c_139_n N_A_86_260#_c_149_n
+ N_A_86_260#_c_150_n N_A_86_260#_c_140_n N_A_86_260#_c_151_n
+ N_A_86_260#_c_141_n N_A_86_260#_c_142_n N_A_86_260#_c_157_p
+ N_A_86_260#_c_152_n N_A_86_260#_c_143_n N_A_86_260#_c_144_n
+ PM_SKY130_FD_SC_MS__O31A_4%A_86_260#
x_PM_SKY130_FD_SC_MS__O31A_4%B1 N_B1_M1002_g N_B1_c_264_n N_B1_M1009_g
+ N_B1_M1004_g N_B1_M1023_g B1 B1 N_B1_c_268_n N_B1_c_269_n
+ PM_SKY130_FD_SC_MS__O31A_4%B1
x_PM_SKY130_FD_SC_MS__O31A_4%A3 N_A3_M1012_g N_A3_M1021_g N_A3_M1013_g
+ N_A3_M1022_g A3 A3 A3 A3 N_A3_c_324_n PM_SKY130_FD_SC_MS__O31A_4%A3
x_PM_SKY130_FD_SC_MS__O31A_4%A1 N_A1_M1016_g N_A1_M1000_g N_A1_M1019_g
+ N_A1_M1001_g A1 N_A1_c_377_n N_A1_c_378_n PM_SKY130_FD_SC_MS__O31A_4%A1
x_PM_SKY130_FD_SC_MS__O31A_4%A2 N_A2_c_426_n N_A2_M1005_g N_A2_M1010_g
+ N_A2_c_429_n N_A2_c_430_n N_A2_M1015_g N_A2_M1017_g A2 N_A2_c_433_n
+ PM_SKY130_FD_SC_MS__O31A_4%A2
x_PM_SKY130_FD_SC_MS__O31A_4%VPWR N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_M1014_d
+ N_VPWR_M1004_s N_VPWR_M1000_d N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n
+ VPWR N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n
+ N_VPWR_c_486_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ PM_SKY130_FD_SC_MS__O31A_4%VPWR
x_PM_SKY130_FD_SC_MS__O31A_4%X N_X_M1003_s N_X_M1018_s N_X_M1007_s N_X_M1011_s
+ N_X_c_581_n N_X_c_576_n N_X_c_577_n N_X_c_582_n X X X X X X X X X
+ PM_SKY130_FD_SC_MS__O31A_4%X
x_PM_SKY130_FD_SC_MS__O31A_4%A_699_392# N_A_699_392#_M1012_s
+ N_A_699_392#_M1013_s N_A_699_392#_M1015_d N_A_699_392#_c_640_n
+ N_A_699_392#_c_641_n N_A_699_392#_c_642_n N_A_699_392#_c_643_n
+ N_A_699_392#_c_644_n N_A_699_392#_c_645_n
+ PM_SKY130_FD_SC_MS__O31A_4%A_699_392#
x_PM_SKY130_FD_SC_MS__O31A_4%A_971_392# N_A_971_392#_M1005_s
+ N_A_971_392#_M1001_s N_A_971_392#_c_694_n N_A_971_392#_c_687_n
+ N_A_971_392#_c_690_n N_A_971_392#_c_688_n
+ PM_SKY130_FD_SC_MS__O31A_4%A_971_392#
x_PM_SKY130_FD_SC_MS__O31A_4%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_M1020_d
+ N_VGND_M1021_d N_VGND_M1010_d N_VGND_M1019_d N_VGND_c_712_n N_VGND_c_713_n
+ N_VGND_c_714_n N_VGND_c_715_n N_VGND_c_716_n N_VGND_c_717_n N_VGND_c_718_n
+ N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n N_VGND_c_722_n VGND
+ N_VGND_c_723_n N_VGND_c_724_n N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n
+ N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n PM_SKY130_FD_SC_MS__O31A_4%VGND
x_PM_SKY130_FD_SC_MS__O31A_4%A_492_125# N_A_492_125#_M1009_d
+ N_A_492_125#_M1023_d N_A_492_125#_M1022_s N_A_492_125#_M1016_s
+ N_A_492_125#_M1017_s N_A_492_125#_c_808_n N_A_492_125#_c_809_n
+ N_A_492_125#_c_810_n N_A_492_125#_c_811_n N_A_492_125#_c_812_n
+ N_A_492_125#_c_813_n N_A_492_125#_c_814_n N_A_492_125#_c_815_n
+ N_A_492_125#_c_816_n N_A_492_125#_c_817_n N_A_492_125#_c_818_n
+ N_A_492_125#_c_819_n N_A_492_125#_c_820_n
+ PM_SKY130_FD_SC_MS__O31A_4%A_492_125#
cc_1 VNB N_A_86_260#_M1007_g 0.00949968f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_2 VNB N_A_86_260#_M1003_g 0.0260209f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_3 VNB N_A_86_260#_M1006_g 0.0210733f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.74
cc_4 VNB N_A_86_260#_M1008_g 0.0015344f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_5 VNB N_A_86_260#_M1018_g 0.0210988f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_6 VNB N_A_86_260#_M1011_g 0.00154196f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_7 VNB N_A_86_260#_M1020_g 0.0250096f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=0.74
cc_8 VNB N_A_86_260#_M1014_g 0.00168479f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_9 VNB N_A_86_260#_c_138_n 0.0189554f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.42
cc_10 VNB N_A_86_260#_c_139_n 0.0151647f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=1.465
cc_11 VNB N_A_86_260#_c_140_n 0.0033999f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=1.215
cc_12 VNB N_A_86_260#_c_141_n 0.00272643f $X=-0.19 $Y=-0.245 $X2=3.105 $Y2=0.77
cc_13 VNB N_A_86_260#_c_142_n 0.00351491f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=1.3
cc_14 VNB N_A_86_260#_c_143_n 0.0122613f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.465
cc_15 VNB N_A_86_260#_c_144_n 0.0636314f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.465
cc_16 VNB N_B1_M1002_g 0.00200761f $X=-0.19 $Y=-0.245 $X2=3.955 $Y2=1.96
cc_17 VNB N_B1_c_264_n 0.010089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_M1009_g 0.0234854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_M1023_g 0.023331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.00140579f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.42
cc_21 VNB N_B1_c_268_n 0.0143854f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.63
cc_22 VNB N_B1_c_269_n 0.0218147f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_23 VNB N_A3_M1021_g 0.0221804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A3_M1022_g 0.0209132f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_25 VNB A3 0.00920475f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.3
cc_26 VNB N_A3_c_324_n 0.0257987f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_27 VNB N_A1_M1016_g 0.0191469f $X=-0.19 $Y=-0.245 $X2=3.955 $Y2=1.96
cc_28 VNB N_A1_M1019_g 0.0200124f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_29 VNB N_A1_c_377_n 0.00143943f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_30 VNB N_A1_c_378_n 0.0279499f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_31 VNB N_A2_c_426_n 0.00583194f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=0.625
cc_32 VNB N_A2_M1005_g 0.0105049f $X=-0.19 $Y=-0.245 $X2=3.955 $Y2=1.96
cc_33 VNB N_A2_M1010_g 0.0273481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_429_n 0.101926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_430_n 0.0124157f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.54
cc_36 VNB N_A2_M1017_g 0.0461536f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.42
cc_37 VNB A2 0.0112145f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.3
cc_38 VNB N_A2_c_433_n 0.0197857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_486_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_576_n 0.00426489f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_41 VNB N_X_c_577_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.42
cc_42 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB X 6.83523e-19 $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.3
cc_44 VNB X 0.00241697f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_45 VNB N_VGND_c_712_n 0.011635f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.42
cc_46 VNB N_VGND_c_713_n 0.0505972f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.74
cc_47 VNB N_VGND_c_714_n 0.00728606f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_48 VNB N_VGND_c_715_n 0.0172342f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_49 VNB N_VGND_c_716_n 0.0125309f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_50 VNB N_VGND_c_717_n 0.00373475f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=0.74
cc_51 VNB N_VGND_c_718_n 0.0081779f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_52 VNB N_VGND_c_719_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.42
cc_53 VNB N_VGND_c_720_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=1.465
cc_54 VNB N_VGND_c_721_n 0.0157641f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.465
cc_55 VNB N_VGND_c_722_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.465
cc_56 VNB N_VGND_c_723_n 0.0177297f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.105
cc_57 VNB N_VGND_c_724_n 0.0432711f $X=-0.19 $Y=-0.245 $X2=2.63 $Y2=2.815
cc_58 VNB N_VGND_c_725_n 0.0171291f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=2.46
cc_59 VNB N_VGND_c_726_n 0.0199127f $X=-0.19 $Y=-0.245 $X2=4.09 $Y2=2.46
cc_60 VNB N_VGND_c_727_n 0.382101f $X=-0.19 $Y=-0.245 $X2=4.09 $Y2=2.46
cc_61 VNB N_VGND_c_728_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.465
cc_62 VNB N_VGND_c_729_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.465
cc_63 VNB N_VGND_c_730_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_492_125#_c_808_n 0.007888f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.42
cc_65 VNB N_A_492_125#_c_809_n 0.0224913f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.3
cc_66 VNB N_A_492_125#_c_810_n 0.00508483f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.74
cc_67 VNB N_A_492_125#_c_811_n 0.00701587f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_68 VNB N_A_492_125#_c_812_n 0.00257879f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_69 VNB N_A_492_125#_c_813_n 0.00404805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_492_125#_c_814_n 0.00299721f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_71 VNB N_A_492_125#_c_815_n 0.00366864f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.63
cc_72 VNB N_A_492_125#_c_816_n 0.00252922f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.3
cc_73 VNB N_A_492_125#_c_817_n 0.0145756f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=0.74
cc_74 VNB N_A_492_125#_c_818_n 0.0232757f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_75 VNB N_A_492_125#_c_819_n 0.00210347f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.42
cc_76 VNB N_A_492_125#_c_820_n 0.00228969f $X=-0.19 $Y=-0.245 $X2=2.465
+ $Y2=1.465
cc_77 VPB N_A_86_260#_M1007_g 0.0274048f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.4
cc_78 VPB N_A_86_260#_M1008_g 0.0214037f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_79 VPB N_A_86_260#_M1011_g 0.0220386f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=2.4
cc_80 VPB N_A_86_260#_M1014_g 0.0237294f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_81 VPB N_A_86_260#_c_149_n 0.00203102f $X=-0.19 $Y=1.66 $X2=2.63 $Y2=2.105
cc_82 VPB N_A_86_260#_c_150_n 0.00202354f $X=-0.19 $Y=1.66 $X2=2.63 $Y2=2.815
cc_83 VPB N_A_86_260#_c_151_n 0.011168f $X=-0.19 $Y=1.66 $X2=3.925 $Y2=2.46
cc_84 VPB N_A_86_260#_c_152_n 0.00231117f $X=-0.19 $Y=1.66 $X2=4.09 $Y2=2.46
cc_85 VPB N_B1_M1002_g 0.0295631f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=1.96
cc_86 VPB N_B1_M1004_g 0.0244252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB B1 0.00400555f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.42
cc_88 VPB N_B1_c_269_n 0.0286336f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_89 VPB N_A3_M1012_g 0.0256795f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=1.96
cc_90 VPB N_A3_M1013_g 0.0225377f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.4
cc_91 VPB A3 0.00849667f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.3
cc_92 VPB N_A3_c_324_n 0.0156204f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_93 VPB N_A1_M1000_g 0.0225089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A1_M1001_g 0.0235204f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.74
cc_95 VPB N_A1_c_377_n 8.74948e-19 $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_96 VPB N_A1_c_378_n 0.0180575f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_97 VPB N_A2_M1005_g 0.0287094f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=1.96
cc_98 VPB N_A2_M1015_g 0.0318458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB A2 0.00710695f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.3
cc_100 VPB N_A2_c_433_n 0.012984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_487_n 0.0111306f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.74
cc_102 VPB N_VPWR_c_488_n 0.0638588f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.42
cc_103 VPB N_VPWR_c_489_n 0.0049754f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.63
cc_104 VPB N_VPWR_c_490_n 0.0118948f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.3
cc_105 VPB N_VPWR_c_491_n 0.0103514f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=2.4
cc_106 VPB N_VPWR_c_492_n 0.00635773f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_107 VPB N_VPWR_c_493_n 0.0184472f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_108 VPB N_VPWR_c_494_n 0.00458862f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_109 VPB N_VPWR_c_495_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_496_n 0.0186844f $X=-0.19 $Y=1.66 $X2=2.59 $Y2=1.63
cc_111 VPB N_VPWR_c_497_n 0.0582525f $X=-0.19 $Y=1.66 $X2=2.59 $Y2=2.815
cc_112 VPB N_VPWR_c_498_n 0.0325002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_486_n 0.0847647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_500_n 0.0047828f $X=-0.19 $Y=1.66 $X2=4.09 $Y2=2.46
cc_115 VPB N_VPWR_c_501_n 0.00612837f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.465
cc_116 VPB N_VPWR_c_502_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.465
cc_117 VPB N_X_c_581_n 0.00510549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_X_c_582_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB X 0.00132696f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_120 VPB X 0.00206901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_699_392#_c_640_n 0.00801296f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.54
cc_122 VPB N_A_699_392#_c_641_n 0.00216001f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.74
cc_123 VPB N_A_699_392#_c_642_n 0.0104158f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.42
cc_124 VPB N_A_699_392#_c_643_n 0.00977958f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.3
cc_125 VPB N_A_699_392#_c_644_n 0.0351596f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=0.74
cc_126 VPB N_A_699_392#_c_645_n 0.001972f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_127 VPB N_A_971_392#_c_687_n 0.00202379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_971_392#_c_688_n 0.00275667f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.42
cc_129 N_A_86_260#_M1014_g N_B1_M1002_g 0.0255846f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A_86_260#_c_139_n N_B1_M1002_g 0.00732671f $X=2.465 $Y=1.465 $X2=0
+ $Y2=0
cc_131 N_A_86_260#_c_149_n N_B1_M1002_g 0.0133856f $X=2.63 $Y=2.105 $X2=0 $Y2=0
cc_132 N_A_86_260#_c_150_n N_B1_M1002_g 0.00572734f $X=2.63 $Y=2.815 $X2=0 $Y2=0
cc_133 N_A_86_260#_c_157_p N_B1_M1002_g 0.00207369f $X=2.63 $Y=2.46 $X2=0 $Y2=0
cc_134 N_A_86_260#_c_139_n N_B1_c_264_n 0.00665072f $X=2.465 $Y=1.465 $X2=0
+ $Y2=0
cc_135 N_A_86_260#_c_142_n N_B1_c_264_n 9.5723e-19 $X=2.465 $Y=1.3 $X2=0 $Y2=0
cc_136 N_A_86_260#_c_144_n N_B1_c_264_n 0.00669127f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_137 N_A_86_260#_c_140_n N_B1_M1009_g 0.0183346f $X=2.94 $Y=1.215 $X2=0 $Y2=0
cc_138 N_A_86_260#_c_142_n N_B1_M1009_g 0.00794685f $X=2.465 $Y=1.3 $X2=0 $Y2=0
cc_139 N_A_86_260#_c_151_n N_B1_M1004_g 0.0173779f $X=3.925 $Y=2.46 $X2=0 $Y2=0
cc_140 N_A_86_260#_c_140_n N_B1_M1023_g 0.00360052f $X=2.94 $Y=1.215 $X2=0 $Y2=0
cc_141 N_A_86_260#_c_141_n N_B1_M1023_g 0.00594662f $X=3.105 $Y=0.77 $X2=0 $Y2=0
cc_142 N_A_86_260#_c_149_n B1 0.0299118f $X=2.63 $Y=2.105 $X2=0 $Y2=0
cc_143 N_A_86_260#_c_140_n B1 0.0289054f $X=2.94 $Y=1.215 $X2=0 $Y2=0
cc_144 N_A_86_260#_c_151_n B1 0.017729f $X=3.925 $Y=2.46 $X2=0 $Y2=0
cc_145 N_A_86_260#_c_142_n B1 0.0117228f $X=2.465 $Y=1.3 $X2=0 $Y2=0
cc_146 N_A_86_260#_c_140_n N_B1_c_268_n 0.0020338f $X=2.94 $Y=1.215 $X2=0 $Y2=0
cc_147 N_A_86_260#_c_142_n N_B1_c_268_n 0.0119589f $X=2.465 $Y=1.3 $X2=0 $Y2=0
cc_148 N_A_86_260#_c_149_n N_B1_c_269_n 0.00276789f $X=2.63 $Y=2.105 $X2=0 $Y2=0
cc_149 N_A_86_260#_c_140_n N_B1_c_269_n 0.00118356f $X=2.94 $Y=1.215 $X2=0 $Y2=0
cc_150 N_A_86_260#_c_151_n N_B1_c_269_n 0.00527458f $X=3.925 $Y=2.46 $X2=0 $Y2=0
cc_151 N_A_86_260#_c_151_n N_A3_M1012_g 0.0117172f $X=3.925 $Y=2.46 $X2=0 $Y2=0
cc_152 N_A_86_260#_c_152_n N_A3_M1012_g 0.0205284f $X=4.09 $Y=2.46 $X2=0 $Y2=0
cc_153 N_A_86_260#_c_152_n N_A3_M1013_g 0.00781286f $X=4.09 $Y=2.46 $X2=0 $Y2=0
cc_154 N_A_86_260#_c_151_n N_VPWR_M1004_s 0.00567487f $X=3.925 $Y=2.46 $X2=0
+ $Y2=0
cc_155 N_A_86_260#_M1007_g N_VPWR_c_488_n 0.00517052f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_86_260#_M1007_g N_VPWR_c_489_n 6.24656e-19 $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_86_260#_M1008_g N_VPWR_c_489_n 0.0152854f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_86_260#_M1011_g N_VPWR_c_489_n 0.00349416f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_86_260#_M1014_g N_VPWR_c_490_n 0.00357619f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_86_260#_c_139_n N_VPWR_c_490_n 0.0202614f $X=2.465 $Y=1.465 $X2=0
+ $Y2=0
cc_161 N_A_86_260#_c_149_n N_VPWR_c_490_n 0.0220111f $X=2.63 $Y=2.105 $X2=0
+ $Y2=0
cc_162 N_A_86_260#_c_150_n N_VPWR_c_490_n 0.0140997f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_163 N_A_86_260#_c_150_n N_VPWR_c_491_n 0.00940654f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_164 N_A_86_260#_c_151_n N_VPWR_c_491_n 0.021375f $X=3.925 $Y=2.46 $X2=0 $Y2=0
cc_165 N_A_86_260#_M1007_g N_VPWR_c_493_n 0.00515235f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_86_260#_M1008_g N_VPWR_c_493_n 0.00460063f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A_86_260#_M1011_g N_VPWR_c_495_n 0.005209f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A_86_260#_M1014_g N_VPWR_c_495_n 0.005209f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_86_260#_c_150_n N_VPWR_c_496_n 0.0109793f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_170 N_A_86_260#_c_152_n N_VPWR_c_497_n 0.0143411f $X=4.09 $Y=2.46 $X2=0 $Y2=0
cc_171 N_A_86_260#_M1007_g N_VPWR_c_486_n 0.00967715f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_86_260#_M1008_g N_VPWR_c_486_n 0.00908554f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A_86_260#_M1011_g N_VPWR_c_486_n 0.00982266f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_86_260#_M1014_g N_VPWR_c_486_n 0.00983127f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_86_260#_c_150_n N_VPWR_c_486_n 0.00901959f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_176 N_A_86_260#_c_151_n N_VPWR_c_486_n 0.030885f $X=3.925 $Y=2.46 $X2=0 $Y2=0
cc_177 N_A_86_260#_c_152_n N_VPWR_c_486_n 0.0117867f $X=4.09 $Y=2.46 $X2=0 $Y2=0
cc_178 N_A_86_260#_M1008_g N_X_c_581_n 0.0165554f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_86_260#_M1011_g N_X_c_581_n 0.0142852f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_86_260#_M1014_g N_X_c_581_n 0.00312116f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_86_260#_c_139_n N_X_c_581_n 0.0624639f $X=2.465 $Y=1.465 $X2=0 $Y2=0
cc_182 N_A_86_260#_c_149_n N_X_c_581_n 5.06195e-19 $X=2.63 $Y=2.105 $X2=0 $Y2=0
cc_183 N_A_86_260#_c_144_n N_X_c_581_n 0.00423276f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_184 N_A_86_260#_M1006_g N_X_c_576_n 0.01265f $X=0.955 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_86_260#_M1018_g N_X_c_576_n 0.0121615f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_86_260#_c_139_n N_X_c_576_n 0.0538252f $X=2.465 $Y=1.465 $X2=0 $Y2=0
cc_187 N_A_86_260#_c_144_n N_X_c_576_n 0.00516417f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_188 N_A_86_260#_M1006_g N_X_c_577_n 6.43273e-19 $X=0.955 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_86_260#_M1018_g N_X_c_577_n 0.00867431f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_86_260#_M1020_g N_X_c_577_n 3.97481e-19 $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_86_260#_M1008_g N_X_c_582_n 7.71145e-19 $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_86_260#_M1011_g N_X_c_582_n 0.0144894f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_86_260#_M1014_g N_X_c_582_n 0.013233f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_86_260#_M1003_g X 0.00783249f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_86_260#_M1006_g X 0.00874985f $X=0.955 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_86_260#_M1018_g X 6.3164e-19 $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_86_260#_M1003_g X 0.00209097f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_86_260#_M1006_g X 0.00132316f $X=0.955 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_86_260#_M1007_g X 0.0134878f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_86_260#_M1003_g X 0.00866064f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_86_260#_M1006_g X 0.00443027f $X=0.955 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_86_260#_c_138_n X 0.0104392f $X=0.52 $Y=1.42 $X2=0 $Y2=0
cc_203 N_A_86_260#_c_139_n X 0.0260905f $X=2.465 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_86_260#_c_143_n X 0.0130055f $X=0.88 $Y=1.465 $X2=0 $Y2=0
cc_205 N_A_86_260#_c_144_n X 0.00527186f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_206 N_A_86_260#_M1007_g X 0.00333871f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_86_260#_M1007_g X 0.0138065f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_86_260#_M1008_g X 3.7104e-19 $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_86_260#_c_151_n N_A_699_392#_M1012_s 0.00757695f $X=3.925 $Y=2.46
+ $X2=-0.19 $Y2=-0.245
cc_210 N_A_86_260#_M1012_d N_A_699_392#_c_640_n 0.00167813f $X=3.955 $Y=1.96
+ $X2=0 $Y2=0
cc_211 N_A_86_260#_c_151_n N_A_699_392#_c_640_n 0.0286378f $X=3.925 $Y=2.46
+ $X2=0 $Y2=0
cc_212 N_A_86_260#_c_152_n N_A_699_392#_c_640_n 0.0174794f $X=4.09 $Y=2.46 $X2=0
+ $Y2=0
cc_213 N_A_86_260#_c_152_n N_A_699_392#_c_641_n 0.0162641f $X=4.09 $Y=2.46 $X2=0
+ $Y2=0
cc_214 N_A_86_260#_M1003_g N_VGND_c_713_n 0.00647381f $X=0.525 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_86_260#_M1006_g N_VGND_c_714_n 0.002905f $X=0.955 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_86_260#_M1018_g N_VGND_c_714_n 0.00291178f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_86_260#_M1018_g N_VGND_c_715_n 6.16597e-19 $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_86_260#_M1020_g N_VGND_c_715_n 0.0151659f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_86_260#_c_139_n N_VGND_c_715_n 0.028354f $X=2.465 $Y=1.465 $X2=0
+ $Y2=0
cc_220 N_A_86_260#_c_144_n N_VGND_c_715_n 0.00277945f $X=1.87 $Y=1.465 $X2=0
+ $Y2=0
cc_221 N_A_86_260#_M1003_g N_VGND_c_719_n 0.00434272f $X=0.525 $Y=0.74 $X2=0
+ $Y2=0
cc_222 N_A_86_260#_M1006_g N_VGND_c_719_n 0.00434272f $X=0.955 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_86_260#_M1018_g N_VGND_c_723_n 0.00434272f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_86_260#_M1020_g N_VGND_c_723_n 0.00383152f $X=1.83 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_86_260#_M1003_g N_VGND_c_727_n 0.0082404f $X=0.525 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_86_260#_M1006_g N_VGND_c_727_n 0.00820433f $X=0.955 $Y=0.74 $X2=0
+ $Y2=0
cc_227 N_A_86_260#_M1018_g N_VGND_c_727_n 0.00820769f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_86_260#_M1020_g N_VGND_c_727_n 0.0075754f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_86_260#_c_142_n N_A_492_125#_M1009_d 0.00486326f $X=2.465 $Y=1.3
+ $X2=-0.19 $Y2=-0.245
cc_230 N_A_86_260#_M1020_g N_A_492_125#_c_808_n 0.00104088f $X=1.83 $Y=0.74
+ $X2=0 $Y2=0
cc_231 N_A_86_260#_c_139_n N_A_492_125#_c_808_n 0.00127831f $X=2.465 $Y=1.465
+ $X2=0 $Y2=0
cc_232 N_A_86_260#_c_140_n N_A_492_125#_c_808_n 2.62997e-19 $X=2.94 $Y=1.215
+ $X2=0 $Y2=0
cc_233 N_A_86_260#_c_141_n N_A_492_125#_c_808_n 0.0141109f $X=3.105 $Y=0.77
+ $X2=0 $Y2=0
cc_234 N_A_86_260#_c_142_n N_A_492_125#_c_808_n 0.0191947f $X=2.465 $Y=1.3 $X2=0
+ $Y2=0
cc_235 N_A_86_260#_c_141_n N_A_492_125#_c_809_n 0.0259178f $X=3.105 $Y=0.77
+ $X2=0 $Y2=0
cc_236 N_A_86_260#_M1020_g N_A_492_125#_c_810_n 5.82409e-19 $X=1.83 $Y=0.74
+ $X2=0 $Y2=0
cc_237 N_A_86_260#_c_141_n N_A_492_125#_c_811_n 0.0190383f $X=3.105 $Y=0.77
+ $X2=0 $Y2=0
cc_238 N_A_86_260#_c_140_n N_A_492_125#_c_813_n 0.00711695f $X=2.94 $Y=1.215
+ $X2=0 $Y2=0
cc_239 B1 N_A3_M1012_g 0.00442778f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B1_c_269_n N_A3_M1012_g 5.6578e-19 $X=3.32 $Y=1.635 $X2=0 $Y2=0
cc_241 N_B1_M1023_g N_A3_M1021_g 0.0201055f $X=3.32 $Y=0.945 $X2=0 $Y2=0
cc_242 N_B1_M1023_g A3 0.00408488f $X=3.32 $Y=0.945 $X2=0 $Y2=0
cc_243 B1 A3 0.0198498f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_244 N_B1_M1023_g N_A3_c_324_n 0.0113055f $X=3.32 $Y=0.945 $X2=0 $Y2=0
cc_245 B1 N_A3_c_324_n 2.27913e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_246 B1 N_VPWR_M1004_s 0.00374091f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_247 N_B1_M1002_g N_VPWR_c_490_n 0.00844293f $X=2.405 $Y=2.46 $X2=0 $Y2=0
cc_248 N_B1_M1002_g N_VPWR_c_491_n 4.26426e-19 $X=2.405 $Y=2.46 $X2=0 $Y2=0
cc_249 N_B1_M1004_g N_VPWR_c_491_n 0.00897501f $X=2.855 $Y=2.46 $X2=0 $Y2=0
cc_250 N_B1_M1002_g N_VPWR_c_496_n 0.005209f $X=2.405 $Y=2.46 $X2=0 $Y2=0
cc_251 N_B1_M1004_g N_VPWR_c_496_n 0.00460063f $X=2.855 $Y=2.46 $X2=0 $Y2=0
cc_252 N_B1_M1002_g N_VPWR_c_486_n 0.00983239f $X=2.405 $Y=2.46 $X2=0 $Y2=0
cc_253 N_B1_M1004_g N_VPWR_c_486_n 0.00447027f $X=2.855 $Y=2.46 $X2=0 $Y2=0
cc_254 N_B1_M1004_g N_A_699_392#_c_640_n 0.00239877f $X=2.855 $Y=2.46 $X2=0
+ $Y2=0
cc_255 B1 N_A_699_392#_c_640_n 0.0134747f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_256 N_B1_M1009_g N_VGND_c_715_n 0.00510703f $X=2.84 $Y=0.945 $X2=0 $Y2=0
cc_257 N_B1_c_264_n N_A_492_125#_c_808_n 0.00120332f $X=2.495 $Y=1.545 $X2=0
+ $Y2=0
cc_258 N_B1_M1009_g N_A_492_125#_c_808_n 0.00770967f $X=2.84 $Y=0.945 $X2=0
+ $Y2=0
cc_259 N_B1_M1023_g N_A_492_125#_c_808_n 5.99032e-19 $X=3.32 $Y=0.945 $X2=0
+ $Y2=0
cc_260 N_B1_M1009_g N_A_492_125#_c_809_n 0.00676567f $X=2.84 $Y=0.945 $X2=0
+ $Y2=0
cc_261 N_B1_M1023_g N_A_492_125#_c_809_n 0.00661564f $X=3.32 $Y=0.945 $X2=0
+ $Y2=0
cc_262 N_B1_M1023_g N_A_492_125#_c_811_n 0.00641777f $X=3.32 $Y=0.945 $X2=0
+ $Y2=0
cc_263 N_B1_M1023_g N_A_492_125#_c_813_n 0.00113032f $X=3.32 $Y=0.945 $X2=0
+ $Y2=0
cc_264 A3 N_A1_c_377_n 0.0197842f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_265 A3 N_A1_c_378_n 0.0114116f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_266 N_A3_M1022_g N_A2_c_426_n 0.00688379f $X=4.34 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_267 A3 N_A2_M1005_g 0.0178412f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_268 N_A3_c_324_n N_A2_M1005_g 0.0315281f $X=4.315 $Y=1.62 $X2=0 $Y2=0
cc_269 N_A3_M1022_g N_A2_M1010_g 0.00900058f $X=4.34 $Y=0.945 $X2=0 $Y2=0
cc_270 N_A3_M1012_g N_VPWR_c_491_n 0.00967855f $X=3.865 $Y=2.46 $X2=0 $Y2=0
cc_271 N_A3_M1012_g N_VPWR_c_497_n 0.005209f $X=3.865 $Y=2.46 $X2=0 $Y2=0
cc_272 N_A3_M1013_g N_VPWR_c_497_n 0.005209f $X=4.315 $Y=2.46 $X2=0 $Y2=0
cc_273 N_A3_M1012_g N_VPWR_c_486_n 0.0052541f $X=3.865 $Y=2.46 $X2=0 $Y2=0
cc_274 N_A3_M1013_g N_VPWR_c_486_n 0.00983474f $X=4.315 $Y=2.46 $X2=0 $Y2=0
cc_275 N_A3_M1012_g N_A_699_392#_c_640_n 0.0119936f $X=3.865 $Y=2.46 $X2=0 $Y2=0
cc_276 N_A3_M1013_g N_A_699_392#_c_640_n 0.0168287f $X=4.315 $Y=2.46 $X2=0 $Y2=0
cc_277 A3 N_A_699_392#_c_640_n 0.0732544f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_278 N_A3_c_324_n N_A_699_392#_c_640_n 0.00310615f $X=4.315 $Y=1.62 $X2=0
+ $Y2=0
cc_279 A3 N_A_699_392#_c_642_n 0.0387446f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_280 A3 N_A_699_392#_c_645_n 0.0185769f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_281 N_A3_M1021_g N_VGND_c_716_n 0.0068292f $X=3.91 $Y=0.945 $X2=0 $Y2=0
cc_282 N_A3_M1022_g N_VGND_c_716_n 0.00159705f $X=4.34 $Y=0.945 $X2=0 $Y2=0
cc_283 N_A3_M1022_g N_VGND_c_717_n 4.44968e-19 $X=4.34 $Y=0.945 $X2=0 $Y2=0
cc_284 N_A3_M1021_g N_VGND_c_724_n 0.00345209f $X=3.91 $Y=0.945 $X2=0 $Y2=0
cc_285 N_A3_M1022_g N_VGND_c_725_n 0.00399929f $X=4.34 $Y=0.945 $X2=0 $Y2=0
cc_286 N_A3_M1021_g N_VGND_c_727_n 0.00394323f $X=3.91 $Y=0.945 $X2=0 $Y2=0
cc_287 N_A3_M1022_g N_VGND_c_727_n 0.00469432f $X=4.34 $Y=0.945 $X2=0 $Y2=0
cc_288 N_A3_M1021_g N_A_492_125#_c_811_n 0.00427413f $X=3.91 $Y=0.945 $X2=0
+ $Y2=0
cc_289 N_A3_M1021_g N_A_492_125#_c_812_n 0.0146144f $X=3.91 $Y=0.945 $X2=0 $Y2=0
cc_290 N_A3_M1022_g N_A_492_125#_c_812_n 0.0109468f $X=4.34 $Y=0.945 $X2=0 $Y2=0
cc_291 A3 N_A_492_125#_c_812_n 0.0447473f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_292 N_A3_c_324_n N_A_492_125#_c_812_n 0.00384728f $X=4.315 $Y=1.62 $X2=0
+ $Y2=0
cc_293 A3 N_A_492_125#_c_813_n 0.0259104f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_294 N_A3_c_324_n N_A_492_125#_c_813_n 0.00106803f $X=4.315 $Y=1.62 $X2=0
+ $Y2=0
cc_295 N_A3_M1021_g N_A_492_125#_c_814_n 5.74244e-19 $X=3.91 $Y=0.945 $X2=0
+ $Y2=0
cc_296 N_A3_M1022_g N_A_492_125#_c_814_n 0.00722889f $X=4.34 $Y=0.945 $X2=0
+ $Y2=0
cc_297 A3 N_A_492_125#_c_815_n 0.0392531f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_298 N_A3_M1022_g N_A_492_125#_c_819_n 9.55648e-19 $X=4.34 $Y=0.945 $X2=0
+ $Y2=0
cc_299 A3 N_A_492_125#_c_819_n 0.0218995f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_300 N_A1_M1016_g N_A2_c_426_n 0.0250543f $X=5.2 $Y=0.945 $X2=-0.19 $Y2=-0.245
cc_301 N_A1_c_378_n N_A2_M1005_g 0.0250543f $X=5.715 $Y=1.62 $X2=0 $Y2=0
cc_302 N_A1_M1016_g N_A2_M1010_g 0.0223502f $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_303 N_A1_M1016_g N_A2_c_429_n 0.00894529f $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_304 N_A1_M1019_g N_A2_c_429_n 0.00894529f $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_305 N_A1_M1001_g N_A2_M1015_g 0.0243685f $X=5.715 $Y=2.46 $X2=0 $Y2=0
cc_306 N_A1_M1019_g N_A2_M1017_g 0.0255707f $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_307 N_A1_c_377_n A2 0.0199019f $X=5.71 $Y=1.62 $X2=0 $Y2=0
cc_308 N_A1_c_378_n A2 4.14111e-19 $X=5.715 $Y=1.62 $X2=0 $Y2=0
cc_309 N_A1_c_377_n N_A2_c_433_n 4.18284e-19 $X=5.71 $Y=1.62 $X2=0 $Y2=0
cc_310 N_A1_c_378_n N_A2_c_433_n 0.0182538f $X=5.715 $Y=1.62 $X2=0 $Y2=0
cc_311 N_A1_M1000_g N_VPWR_c_492_n 0.00868187f $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_312 N_A1_M1001_g N_VPWR_c_492_n 0.00334717f $X=5.715 $Y=2.46 $X2=0 $Y2=0
cc_313 N_A1_M1000_g N_VPWR_c_497_n 0.00460063f $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_314 N_A1_M1001_g N_VPWR_c_498_n 0.005209f $X=5.715 $Y=2.46 $X2=0 $Y2=0
cc_315 N_A1_M1000_g N_VPWR_c_486_n 0.00908665f $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_316 N_A1_M1001_g N_VPWR_c_486_n 0.0098256f $X=5.715 $Y=2.46 $X2=0 $Y2=0
cc_317 N_A1_M1000_g N_A_699_392#_c_642_n 0.0141255f $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_318 N_A1_M1001_g N_A_699_392#_c_642_n 0.0120733f $X=5.715 $Y=2.46 $X2=0 $Y2=0
cc_319 N_A1_c_377_n N_A_699_392#_c_642_n 0.0346511f $X=5.71 $Y=1.62 $X2=0 $Y2=0
cc_320 N_A1_c_378_n N_A_699_392#_c_642_n 0.00475748f $X=5.715 $Y=1.62 $X2=0
+ $Y2=0
cc_321 N_A1_M1001_g N_A_699_392#_c_644_n 7.29338e-19 $X=5.715 $Y=2.46 $X2=0
+ $Y2=0
cc_322 N_A1_M1000_g N_A_971_392#_c_687_n 3.4665e-19 $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_323 N_A1_M1000_g N_A_971_392#_c_690_n 0.0143112f $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_324 N_A1_M1001_g N_A_971_392#_c_690_n 0.0129876f $X=5.715 $Y=2.46 $X2=0 $Y2=0
cc_325 N_A1_M1000_g N_A_971_392#_c_688_n 8.1541e-19 $X=5.215 $Y=2.46 $X2=0 $Y2=0
cc_326 N_A1_M1001_g N_A_971_392#_c_688_n 0.00910977f $X=5.715 $Y=2.46 $X2=0
+ $Y2=0
cc_327 N_A1_M1016_g N_VGND_c_717_n 0.0076579f $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_328 N_A1_M1019_g N_VGND_c_717_n 4.18015e-19 $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_329 N_A1_M1016_g N_VGND_c_718_n 4.22423e-19 $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_330 N_A1_M1019_g N_VGND_c_718_n 0.00778124f $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_331 N_A1_M1016_g N_VGND_c_727_n 7.97988e-19 $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_332 N_A1_M1019_g N_VGND_c_727_n 7.97988e-19 $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_333 N_A1_M1016_g N_A_492_125#_c_815_n 0.0163028f $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_334 N_A1_M1016_g N_A_492_125#_c_816_n 0.00271758f $X=5.2 $Y=0.945 $X2=0 $Y2=0
cc_335 N_A1_M1019_g N_A_492_125#_c_817_n 0.0126598f $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_336 N_A1_c_377_n N_A_492_125#_c_817_n 0.0223244f $X=5.71 $Y=1.62 $X2=0 $Y2=0
cc_337 N_A1_c_378_n N_A_492_125#_c_817_n 0.00236025f $X=5.715 $Y=1.62 $X2=0
+ $Y2=0
cc_338 N_A1_M1019_g N_A_492_125#_c_818_n 8.31855e-19 $X=5.7 $Y=0.945 $X2=0 $Y2=0
cc_339 N_A1_c_377_n N_A_492_125#_c_820_n 0.0139157f $X=5.71 $Y=1.62 $X2=0 $Y2=0
cc_340 N_A1_c_378_n N_A_492_125#_c_820_n 0.00434354f $X=5.715 $Y=1.62 $X2=0
+ $Y2=0
cc_341 N_A2_M1005_g N_VPWR_c_492_n 6.54677e-19 $X=4.765 $Y=2.46 $X2=0 $Y2=0
cc_342 N_A2_M1005_g N_VPWR_c_497_n 0.005209f $X=4.765 $Y=2.46 $X2=0 $Y2=0
cc_343 N_A2_M1015_g N_VPWR_c_498_n 0.0053223f $X=6.205 $Y=2.46 $X2=0 $Y2=0
cc_344 N_A2_M1005_g N_VPWR_c_486_n 0.00983585f $X=4.765 $Y=2.46 $X2=0 $Y2=0
cc_345 N_A2_M1015_g N_VPWR_c_486_n 0.010243f $X=6.205 $Y=2.46 $X2=0 $Y2=0
cc_346 N_A2_M1005_g N_A_699_392#_c_642_n 0.014167f $X=4.765 $Y=2.46 $X2=0 $Y2=0
cc_347 N_A2_M1015_g N_A_699_392#_c_642_n 0.0138232f $X=6.205 $Y=2.46 $X2=0 $Y2=0
cc_348 A2 N_A_699_392#_c_642_n 0.0113921f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_349 N_A2_M1015_g N_A_699_392#_c_643_n 5.94541e-19 $X=6.205 $Y=2.46 $X2=0
+ $Y2=0
cc_350 A2 N_A_699_392#_c_643_n 0.0275157f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_351 N_A2_c_433_n N_A_699_392#_c_643_n 0.00349435f $X=6.28 $Y=1.62 $X2=0 $Y2=0
cc_352 N_A2_M1015_g N_A_699_392#_c_644_n 0.0109992f $X=6.205 $Y=2.46 $X2=0 $Y2=0
cc_353 N_A2_M1005_g N_A_971_392#_c_694_n 0.00235419f $X=4.765 $Y=2.46 $X2=0
+ $Y2=0
cc_354 N_A2_M1005_g N_A_971_392#_c_687_n 0.00671613f $X=4.765 $Y=2.46 $X2=0
+ $Y2=0
cc_355 N_A2_M1015_g N_A_971_392#_c_688_n 4.101e-19 $X=6.205 $Y=2.46 $X2=0 $Y2=0
cc_356 N_A2_c_430_n N_VGND_c_716_n 0.00599508f $X=4.845 $Y=0.18 $X2=0 $Y2=0
cc_357 N_A2_M1010_g N_VGND_c_717_n 0.0173258f $X=4.77 $Y=0.945 $X2=0 $Y2=0
cc_358 N_A2_c_429_n N_VGND_c_717_n 0.0175091f $X=6.125 $Y=0.18 $X2=0 $Y2=0
cc_359 N_A2_c_430_n N_VGND_c_717_n 0.00264835f $X=4.845 $Y=0.18 $X2=0 $Y2=0
cc_360 N_A2_c_429_n N_VGND_c_718_n 0.0232515f $X=6.125 $Y=0.18 $X2=0 $Y2=0
cc_361 N_A2_M1017_g N_VGND_c_718_n 0.0151404f $X=6.2 $Y=0.945 $X2=0 $Y2=0
cc_362 N_A2_c_429_n N_VGND_c_721_n 0.0184168f $X=6.125 $Y=0.18 $X2=0 $Y2=0
cc_363 N_A2_c_430_n N_VGND_c_725_n 0.00486043f $X=4.845 $Y=0.18 $X2=0 $Y2=0
cc_364 N_A2_c_429_n N_VGND_c_726_n 0.00730708f $X=6.125 $Y=0.18 $X2=0 $Y2=0
cc_365 N_A2_c_429_n N_VGND_c_727_n 0.032651f $X=6.125 $Y=0.18 $X2=0 $Y2=0
cc_366 N_A2_c_430_n N_VGND_c_727_n 0.00983503f $X=4.845 $Y=0.18 $X2=0 $Y2=0
cc_367 N_A2_c_426_n N_A_492_125#_c_815_n 9.05238e-19 $X=4.765 $Y=1.43 $X2=0
+ $Y2=0
cc_368 N_A2_M1010_g N_A_492_125#_c_815_n 0.0124384f $X=4.77 $Y=0.945 $X2=0 $Y2=0
cc_369 N_A2_c_429_n N_A_492_125#_c_816_n 0.00490374f $X=6.125 $Y=0.18 $X2=0
+ $Y2=0
cc_370 N_A2_M1017_g N_A_492_125#_c_817_n 0.0126004f $X=6.2 $Y=0.945 $X2=0 $Y2=0
cc_371 A2 N_A_492_125#_c_817_n 0.0379188f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_372 N_A2_c_433_n N_A_492_125#_c_817_n 0.00429604f $X=6.28 $Y=1.62 $X2=0 $Y2=0
cc_373 N_A2_M1017_g N_A_492_125#_c_818_n 0.00764782f $X=6.2 $Y=0.945 $X2=0 $Y2=0
cc_374 N_VPWR_M1008_d N_X_c_581_n 0.00165831f $X=1.06 $Y=1.84 $X2=0 $Y2=0
cc_375 N_VPWR_c_489_n N_X_c_581_n 0.0148589f $X=1.195 $Y=2.305 $X2=0 $Y2=0
cc_376 N_VPWR_c_490_n N_X_c_581_n 0.0062222f $X=2.095 $Y=1.985 $X2=0 $Y2=0
cc_377 N_VPWR_c_489_n N_X_c_582_n 0.0283501f $X=1.195 $Y=2.305 $X2=0 $Y2=0
cc_378 N_VPWR_c_490_n N_X_c_582_n 0.0339179f $X=2.095 $Y=1.985 $X2=0 $Y2=0
cc_379 N_VPWR_c_495_n N_X_c_582_n 0.0144623f $X=2.01 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_c_486_n N_X_c_582_n 0.0118344f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_488_n X 0.00634826f $X=0.295 $Y=1.985 $X2=0 $Y2=0
cc_382 N_VPWR_c_488_n X 0.0333923f $X=0.295 $Y=1.985 $X2=0 $Y2=0
cc_383 N_VPWR_c_489_n X 0.0277554f $X=1.195 $Y=2.305 $X2=0 $Y2=0
cc_384 N_VPWR_c_493_n X 0.0114106f $X=1.03 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_486_n X 0.00936481f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_c_497_n N_A_699_392#_c_641_n 0.00928115f $X=5.275 $Y=3.33 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_486_n N_A_699_392#_c_641_n 0.00768213f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_388 N_VPWR_M1000_d N_A_699_392#_c_642_n 0.00219516f $X=5.305 $Y=1.96 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_498_n N_A_699_392#_c_644_n 0.0145789f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_486_n N_A_699_392#_c_644_n 0.0120225f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_492_n N_A_971_392#_c_687_n 0.0120422f $X=5.44 $Y=2.8 $X2=0 $Y2=0
cc_392 N_VPWR_c_497_n N_A_971_392#_c_687_n 0.0109851f $X=5.275 $Y=3.33 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_486_n N_A_971_392#_c_687_n 0.00902188f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_394 N_VPWR_M1000_d N_A_971_392#_c_690_n 0.00422314f $X=5.305 $Y=1.96 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_492_n N_A_971_392#_c_690_n 0.0189268f $X=5.44 $Y=2.8 $X2=0 $Y2=0
cc_396 N_VPWR_c_492_n N_A_971_392#_c_688_n 0.0137357f $X=5.44 $Y=2.8 $X2=0 $Y2=0
cc_397 N_VPWR_c_498_n N_A_971_392#_c_688_n 0.0145567f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_486_n N_A_971_392#_c_688_n 0.0119773f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_X_c_576_n N_VGND_M1006_d 0.00230942f $X=1.45 $Y=1.045 $X2=0 $Y2=0
cc_400 X N_VGND_c_713_n 0.0225553f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_401 X N_VGND_c_713_n 0.00756924f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_402 N_X_c_576_n N_VGND_c_714_n 0.0135869f $X=1.45 $Y=1.045 $X2=0 $Y2=0
cc_403 N_X_c_577_n N_VGND_c_714_n 0.0286348f $X=1.615 $Y=0.515 $X2=0 $Y2=0
cc_404 X N_VGND_c_714_n 0.0164567f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_405 N_X_c_576_n N_VGND_c_715_n 0.00697079f $X=1.45 $Y=1.045 $X2=0 $Y2=0
cc_406 N_X_c_577_n N_VGND_c_715_n 0.0225912f $X=1.615 $Y=0.515 $X2=0 $Y2=0
cc_407 X N_VGND_c_719_n 0.0144922f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_408 N_X_c_577_n N_VGND_c_723_n 0.0109942f $X=1.615 $Y=0.515 $X2=0 $Y2=0
cc_409 N_X_c_577_n N_VGND_c_727_n 0.00904371f $X=1.615 $Y=0.515 $X2=0 $Y2=0
cc_410 X N_VGND_c_727_n 0.0118826f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_411 N_A_699_392#_c_642_n N_A_971_392#_M1005_s 0.00165831f $X=6.275 $Y=2.04
+ $X2=-0.19 $Y2=1.66
cc_412 N_A_699_392#_c_642_n N_A_971_392#_M1001_s 0.00208352f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_413 N_A_699_392#_c_642_n N_A_971_392#_c_694_n 0.014944f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_414 N_A_699_392#_c_641_n N_A_971_392#_c_687_n 0.018364f $X=4.54 $Y=2.475
+ $X2=0 $Y2=0
cc_415 N_A_699_392#_c_642_n N_A_971_392#_c_690_n 0.0372622f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_416 N_A_699_392#_c_642_n N_A_971_392#_c_688_n 0.0182003f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_417 N_A_699_392#_c_644_n N_A_971_392#_c_688_n 0.0201145f $X=6.44 $Y=2.815
+ $X2=0 $Y2=0
cc_418 N_A_699_392#_c_640_n N_A_492_125#_c_813_n 3.31765e-19 $X=4.435 $Y=2.08
+ $X2=0 $Y2=0
cc_419 N_A_699_392#_c_642_n N_A_492_125#_c_815_n 0.00375987f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_420 N_A_699_392#_c_642_n N_A_492_125#_c_817_n 0.00693341f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_421 N_A_699_392#_c_642_n N_A_492_125#_c_820_n 0.00273162f $X=6.275 $Y=2.04
+ $X2=0 $Y2=0
cc_422 N_VGND_c_715_n N_A_492_125#_c_808_n 0.0353611f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
cc_423 N_VGND_c_716_n N_A_492_125#_c_809_n 0.0141601f $X=4.125 $Y=0.775 $X2=0
+ $Y2=0
cc_424 N_VGND_c_724_n N_A_492_125#_c_809_n 0.063427f $X=3.96 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_727_n N_A_492_125#_c_809_n 0.0381741f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_715_n N_A_492_125#_c_810_n 0.0121618f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
cc_427 N_VGND_c_724_n N_A_492_125#_c_810_n 0.0222866f $X=3.96 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_727_n N_A_492_125#_c_810_n 0.0127763f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_716_n N_A_492_125#_c_811_n 0.0252717f $X=4.125 $Y=0.775 $X2=0
+ $Y2=0
cc_430 N_VGND_M1021_d N_A_492_125#_c_812_n 0.00176461f $X=3.985 $Y=0.625 $X2=0
+ $Y2=0
cc_431 N_VGND_c_716_n N_A_492_125#_c_812_n 0.0152916f $X=4.125 $Y=0.775 $X2=0
+ $Y2=0
cc_432 N_VGND_c_716_n N_A_492_125#_c_814_n 0.0124064f $X=4.125 $Y=0.775 $X2=0
+ $Y2=0
cc_433 N_VGND_c_717_n N_A_492_125#_c_814_n 0.012914f $X=4.985 $Y=0.775 $X2=0
+ $Y2=0
cc_434 N_VGND_c_725_n N_A_492_125#_c_814_n 0.00529503f $X=4.82 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_727_n N_A_492_125#_c_814_n 0.00766513f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_M1010_d N_A_492_125#_c_815_n 0.00176461f $X=4.845 $Y=0.625 $X2=0
+ $Y2=0
cc_437 N_VGND_c_717_n N_A_492_125#_c_815_n 0.0170777f $X=4.985 $Y=0.775 $X2=0
+ $Y2=0
cc_438 N_VGND_c_717_n N_A_492_125#_c_816_n 0.0135156f $X=4.985 $Y=0.775 $X2=0
+ $Y2=0
cc_439 N_VGND_c_718_n N_A_492_125#_c_816_n 0.012914f $X=5.915 $Y=0.775 $X2=0
+ $Y2=0
cc_440 N_VGND_c_721_n N_A_492_125#_c_816_n 0.00534275f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_c_727_n N_A_492_125#_c_816_n 0.00671416f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_M1019_d N_A_492_125#_c_817_n 0.00250873f $X=5.775 $Y=0.625 $X2=0
+ $Y2=0
cc_443 N_VGND_c_718_n N_A_492_125#_c_817_n 0.0209867f $X=5.915 $Y=0.775 $X2=0
+ $Y2=0
cc_444 N_VGND_c_718_n N_A_492_125#_c_818_n 0.0135481f $X=5.915 $Y=0.775 $X2=0
+ $Y2=0
cc_445 N_VGND_c_726_n N_A_492_125#_c_818_n 0.00702137f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_727_n N_A_492_125#_c_818_n 0.0100521f $X=6.48 $Y=0 $X2=0 $Y2=0

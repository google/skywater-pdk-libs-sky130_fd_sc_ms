* File: sky130_fd_sc_ms__o221ai_2.spice
* Created: Fri Aug 28 17:57:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o221ai_2.pex.spice"
.subckt sky130_fd_sc_ms__o221ai_2  VNB VPB C1 B1 B2 A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1017 N_Y_M1017_d N_C1_M1017_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1017_d N_C1_M1018_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_B1_M1012_g N_A_311_85#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1000 N_A_311_85#_M1000_d N_B2_M1000_g N_A_27_74#_M1012_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_311_85#_M1000_d N_B2_M1004_g N_A_27_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.14985 PD=1.02 PS=1.145 NRD=0 NRS=15.804 M=1 R=4.93333
+ SA=75001.1 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1016 N_A_27_74#_M1004_s N_B1_M1016_g N_A_311_85#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.14985 AS=0.1036 PD=1.145 PS=1.02 NRD=4.452 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_311_85#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1406 AS=0.1036 PD=1.12 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1001 N_A_311_85#_M1001_d N_A2_M1001_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.1406 PD=1.07 PS=1.12 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75002.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_311_85#_M1001_d N_A2_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.1258 PD=1.07 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75003.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1011_s N_A1_M1019_g N_A_311_85#_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2146 PD=1.08 PS=2.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_C1_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1013_d N_C1_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3528 PD=1.39 PS=1.75 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1008 N_A_379_368#_M1008_d N_B1_M1008_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1708 AS=0.3528 PD=1.425 PS=1.75 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.4
+ SB=90003.6 A=0.2016 P=2.6 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g N_A_379_368#_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.1708 PD=1.405 PS=1.425 NRD=1.7533 NRS=5.2599 M=1 R=6.22222
+ SA=90001.9 SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1002_d N_B2_M1009_g N_A_379_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.1792 PD=1.405 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.4
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1010 N_A_379_368#_M1009_s N_B1_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2072 PD=1.44 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.9
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1006 N_A_779_368#_M1006_d N_A1_M1006_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2072 PD=1.44 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.4
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_A2_M1005_g N_A_779_368#_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.9
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1005_d N_A2_M1007_g N_A_779_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.4
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1015 N_A_779_368#_M1007_s N_A1_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__o221ai_2.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ebufn_1 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_27_404# VPB pshort w=840000u l=180000u
+  ad=7.441e+11p pd=5.78e+06u as=2.352e+11p ps=2.24e+06u
M1001 a_569_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1002 a_229_74# A VGND VNB nlowvt w=550000u l=150000u
+  ad=1.4575e+11p pd=1.63e+06u as=3.759e+11p ps=3.75e+06u
M1003 a_229_74# A VPWR VPB pshort w=840000u l=180000u
+  ad=2.436e+11p pd=2.26e+06u as=0p ps=0u
M1004 Z a_229_74# a_569_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 a_569_74# a_27_404# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1006 Z a_229_74# a_569_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VGND TE_B a_27_404# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
.ends

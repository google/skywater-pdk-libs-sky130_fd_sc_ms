* File: sky130_fd_sc_ms__sdlclkp_1.pex.spice
* Created: Wed Sep  2 12:32:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%SCE 2 5 9 11 12 15 16
r35 15 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.455
+ $X2=0.407 $Y2=1.29
r36 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.455 $X2=0.385 $Y2=1.455
r37 12 16 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.625
+ $X2=0.385 $Y2=1.625
r38 9 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=1.29
r39 5 11 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.505 $Y=2.54
+ $X2=0.505 $Y2=1.96
r40 2 11 42.8297 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.407 $Y=1.773
+ $X2=0.407 $Y2=1.96
r41 1 15 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.477
+ $X2=0.407 $Y2=1.455
r42 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.407 $Y=1.477
+ $X2=0.407 $Y2=1.773
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%GATE 3 7 9 12 13
r43 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.795
+ $X2=0.97 $Y2=1.96
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.795
+ $X2=0.97 $Y2=1.63
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.795 $X2=0.97 $Y2=1.795
r46 9 13 5.98039 $w=4.78e-07 $l=2.4e-07 $layer=LI1_cond $X=1.045 $Y=2.035
+ $X2=1.045 $Y2=1.795
r47 7 14 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.925 $Y=0.835
+ $X2=0.925 $Y2=1.63
r48 3 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.895 $Y=2.54
+ $X2=0.895 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%A_318_74# 1 2 9 13 16 17 20 26 28 36
c74 28 0 8.55408e-20 $X=2.79 $Y=1.55
c75 9 0 1.79884e-19 $X=3 $Y=2.315
r76 35 36 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3 $Y=1.55 $X2=3.26
+ $Y2=1.55
r77 29 35 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.79 $Y=1.55 $X2=3
+ $Y2=1.55
r78 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.55 $X2=2.79 $Y2=1.55
r79 25 26 10.1887 $w=6.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=1.847
+ $X2=2.38 $Y2=1.847
r80 20 21 8.06167 $w=2.27e-07 $l=1.5e-07 $layer=LI1_cond $X=1.73 $Y=1 $X2=1.88
+ $Y2=1
r81 17 28 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=2.762 $Y=1.63
+ $X2=2.762 $Y2=1.55
r82 17 26 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.625 $Y=1.63
+ $X2=2.38 $Y2=1.63
r83 16 25 6.62291 $w=6.03e-07 $l=3.35e-07 $layer=LI1_cond $X=1.88 $Y=1.847
+ $X2=2.215 $Y2=1.847
r84 15 21 2.43258 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.88 $Y=1.12 $X2=1.88
+ $Y2=1
r85 15 16 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.88 $Y=1.12
+ $X2=1.88 $Y2=1.545
r86 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.385
+ $X2=3.26 $Y2=1.55
r87 11 13 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=3.26 $Y=1.385
+ $X2=3.26 $Y2=0.61
r88 7 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.715 $X2=3
+ $Y2=1.55
r89 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=3 $Y=1.715 $X2=3
+ $Y2=2.315
r90 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.215 $Y2=1.985
r91 1 20 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.37 $X2=1.73 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%A_288_48# 1 2 7 9 10 11 15 16 17 18 19 20
+ 22 25 28 29 30 32 33 34 36 37 38 42 44 46 49 53
c159 32 0 1.99229e-19 $X=3.495 $Y=0.88
c160 25 0 1.91872e-19 $X=3.535 $Y=2.67
c161 20 0 3.05753e-20 $X=2.755 $Y=0.995
r162 50 53 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.075 $Y=2.16
+ $X2=5.215 $Y2=2.16
r163 46 48 18.7692 $w=2.47e-07 $l=3.8e-07 $layer=LI1_cond $X=2.25 $Y=1.195
+ $X2=2.63 $Y2=1.195
r164 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.195 $X2=2.25 $Y2=1.195
r165 44 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=1.995
+ $X2=5.075 $Y2=2.16
r166 44 49 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.075 $Y=1.995
+ $X2=5.075 $Y2=1.13
r167 40 49 7.20219 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=0.965
+ $X2=5.065 $Y2=1.13
r168 40 42 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.065 $Y=0.965
+ $X2=5.065 $Y2=0.515
r169 39 42 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.065 $Y=0.425
+ $X2=5.065 $Y2=0.515
r170 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.9 $Y=0.34
+ $X2=5.065 $Y2=0.425
r171 37 38 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.9 $Y=0.34 $X2=4.26
+ $Y2=0.34
r172 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.175 $Y=0.425
+ $X2=4.26 $Y2=0.34
r173 35 36 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.175 $Y=0.425
+ $X2=4.175 $Y2=0.88
r174 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.09 $Y=0.965
+ $X2=4.175 $Y2=0.88
r175 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.09 $Y=0.965
+ $X2=3.58 $Y2=0.965
r176 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.495 $Y=0.88
+ $X2=3.58 $Y2=0.965
r177 31 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.495 $Y=0.425
+ $X2=3.495 $Y2=0.88
r178 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=0.34
+ $X2=3.495 $Y2=0.425
r179 29 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.41 $Y=0.34
+ $X2=2.715 $Y2=0.34
r180 28 48 2.92482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.03
+ $X2=2.63 $Y2=1.195
r181 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.715 $Y2=0.34
r182 27 28 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.63 $Y2=1.03
r183 23 25 157.427 $w=1.8e-07 $l=4.05e-07 $layer=POLY_cond $X=3.535 $Y=3.075
+ $X2=3.535 $Y2=2.67
r184 20 22 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.755 $Y=0.995
+ $X2=2.755 $Y2=0.645
r185 19 47 38.6443 $w=2.87e-07 $l=2.11849e-07 $layer=POLY_cond $X=2.415 $Y=1.07
+ $X2=2.25 $Y2=1.177
r186 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.68 $Y=1.07
+ $X2=2.755 $Y2=0.995
r187 18 19 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.68 $Y=1.07
+ $X2=2.415 $Y2=1.07
r188 16 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.445 $Y=3.15
+ $X2=3.535 $Y2=3.075
r189 16 17 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=3.445 $Y=3.15
+ $X2=2.08 $Y2=3.15
r190 13 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.99 $Y=3.075
+ $X2=2.08 $Y2=3.15
r191 13 15 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=1.99 $Y=3.075
+ $X2=1.99 $Y2=2.26
r192 12 47 43.6655 $w=2.87e-07 $l=3.39382e-07 $layer=POLY_cond $X=1.99 $Y=1.36
+ $X2=2.25 $Y2=1.177
r193 12 15 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=1.99 $Y=1.36 $X2=1.99
+ $Y2=2.26
r194 10 12 26.0485 $w=2.87e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.9 $Y=1.285
+ $X2=1.99 $Y2=1.36
r195 10 11 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.9 $Y=1.285
+ $X2=1.59 $Y2=1.285
r196 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.59 $Y2=1.285
r197 7 9 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.515 $Y2=0.74
r198 2 53 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=2.015 $X2=5.215 $Y2=2.16
r199 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.925
+ $Y=0.37 $X2=5.065 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%A_709_54# 1 2 9 13 15 17 20 22 29 32 34 35
+ 38 39 41 42 49 50 55
c124 50 0 1.28225e-19 $X=6.205 $Y=1.385
c125 49 0 1.17701e-19 $X=6.205 $Y=1.385
c126 35 0 8.87911e-20 $X=5.83 $Y=2.58
c127 22 0 3.71756e-19 $X=4.49 $Y=1.93
c128 9 0 8.55408e-20 $X=3.62 $Y=0.61
r129 50 59 57.0592 $w=3.21e-07 $l=3.8e-07 $layer=POLY_cond $X=6.205 $Y=1.385
+ $X2=6.585 $Y2=1.385
r130 50 57 13.514 $w=3.21e-07 $l=9e-08 $layer=POLY_cond $X=6.205 $Y=1.385
+ $X2=6.115 $Y2=1.385
r131 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.205
+ $Y=1.385 $X2=6.205 $Y2=1.385
r132 46 49 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=5.915 $Y=1.385
+ $X2=6.205 $Y2=1.385
r133 42 44 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.655 $Y=2.58
+ $X2=4.655 $Y2=2.735
r134 37 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.915 $Y=1.55
+ $X2=5.915 $Y2=1.385
r135 37 38 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.915 $Y=1.55
+ $X2=5.915 $Y2=2.495
r136 36 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=2.58
+ $X2=4.655 $Y2=2.58
r137 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.83 $Y=2.58
+ $X2=5.915 $Y2=2.495
r138 35 36 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=5.83 $Y=2.58
+ $X2=4.82 $Y2=2.58
r139 34 42 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=2.495
+ $X2=4.655 $Y2=2.58
r140 33 41 6.99524 $w=2.6e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=2.12
+ $X2=4.655 $Y2=1.93
r141 33 34 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.655 $Y=2.12
+ $X2=4.655 $Y2=2.495
r142 32 41 6.99524 $w=2.6e-07 $l=2.22261e-07 $layer=LI1_cond $X=4.585 $Y=1.74
+ $X2=4.655 $Y2=1.93
r143 32 39 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=4.585 $Y=1.74
+ $X2=4.585 $Y2=1.05
r144 27 39 6.45386 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.555 $Y=0.925
+ $X2=4.555 $Y2=1.05
r145 27 29 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=4.555 $Y=0.925
+ $X2=4.555 $Y2=0.82
r146 25 55 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.765 $Y=1.955
+ $X2=3.925 $Y2=1.955
r147 25 52 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.765 $Y=1.955
+ $X2=3.62 $Y2=1.955
r148 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.765
+ $Y=1.955 $X2=3.765 $Y2=1.955
r149 22 41 0.0189998 $w=3.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=1.93
+ $X2=4.655 $Y2=1.93
r150 22 24 21.9874 $w=3.78e-07 $l=7.25e-07 $layer=LI1_cond $X=4.49 $Y=1.93
+ $X2=3.765 $Y2=1.93
r151 18 59 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.585 $Y=1.55
+ $X2=6.585 $Y2=1.385
r152 18 20 344.008 $w=1.8e-07 $l=8.85e-07 $layer=POLY_cond $X=6.585 $Y=1.55
+ $X2=6.585 $Y2=2.435
r153 15 57 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.22
+ $X2=6.115 $Y2=1.385
r154 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.115 $Y=1.22
+ $X2=6.115 $Y2=0.79
r155 11 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=1.955
r156 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=2.67
r157 7 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.62 $Y=1.79
+ $X2=3.62 $Y2=1.955
r158 7 9 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=3.62 $Y=1.79
+ $X2=3.62 $Y2=0.61
r159 2 44 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.76 $X2=4.655 $Y2=2.735
r160 2 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.76 $X2=4.655 $Y2=1.905
r161 1 29 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.515 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%A_566_74# 1 2 7 9 12 15 19 22 28 31 34 38
c82 28 0 3.05753e-20 $X=3.155 $Y=0.76
c83 12 0 8.87911e-20 $X=4.43 $Y=2.32
c84 7 0 1.99229e-19 $X=4.3 $Y=1.22
r85 37 38 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=4.3 $Y=1.385 $X2=4.43
+ $Y2=1.385
r86 31 32 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=2.59
+ $X2=3.225 $Y2=2.425
r87 26 28 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.97 $Y=0.76
+ $X2=3.155 $Y2=0.76
r88 23 37 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.155 $Y=1.385
+ $X2=4.3 $Y2=1.385
r89 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=1.385 $X2=4.155 $Y2=1.385
r90 20 34 0.295496 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=3.39 $Y=1.385
+ $X2=3.23 $Y2=1.385
r91 20 22 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.39 $Y=1.385
+ $X2=4.155 $Y2=1.385
r92 19 32 13.5052 $w=3.18e-07 $l=3.75e-07 $layer=LI1_cond $X=3.23 $Y=2.05
+ $X2=3.23 $Y2=2.425
r93 16 34 6.56857 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=1.55
+ $X2=3.23 $Y2=1.385
r94 16 19 18.0069 $w=3.18e-07 $l=5e-07 $layer=LI1_cond $X=3.23 $Y=1.55 $X2=3.23
+ $Y2=2.05
r95 15 34 6.56857 $w=2.45e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.155 $Y=1.22
+ $X2=3.23 $Y2=1.385
r96 14 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0.925
+ $X2=3.155 $Y2=0.76
r97 14 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.155 $Y=0.925
+ $X2=3.155 $Y2=1.22
r98 10 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.43 $Y=1.55
+ $X2=4.43 $Y2=1.385
r99 10 12 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.43 $Y=1.55
+ $X2=4.43 $Y2=2.32
r100 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=1.22 $X2=4.3
+ $Y2=1.385
r101 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.3 $Y=1.22 $X2=4.3
+ $Y2=0.74
r102 2 31 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.895 $X2=3.225 $Y2=2.59
r103 2 19 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.895 $X2=3.225 $Y2=2.05
r104 1 26 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.37 $X2=2.97 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%CLK 3 5 7 10 12 13 14 16 17 23
c59 23 0 1.28225e-19 $X=5.495 $Y=1.52
c60 10 0 1.13508e-19 $X=5.755 $Y=0.79
r61 22 24 23.8705 $w=5.25e-07 $l=2.6e-07 $layer=POLY_cond $X=5.495 $Y=1.647
+ $X2=5.755 $Y2=1.647
r62 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=1.52 $X2=5.495 $Y2=1.52
r63 20 22 5.04952 $w=5.25e-07 $l=5.5e-08 $layer=POLY_cond $X=5.44 $Y=1.647
+ $X2=5.495 $Y2=1.647
r64 19 20 14.6895 $w=5.25e-07 $l=1.6e-07 $layer=POLY_cond $X=5.28 $Y=1.647
+ $X2=5.44 $Y2=1.647
r65 17 23 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.495 $Y=1.665
+ $X2=5.495 $Y2=1.52
r66 14 16 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=6.135 $Y=1.94
+ $X2=6.135 $Y2=2.435
r67 13 24 34.3153 $w=5.25e-07 $l=2.52733e-07 $layer=POLY_cond $X=5.83 $Y=1.865
+ $X2=5.755 $Y2=1.647
r68 12 14 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.045 $Y=1.865
+ $X2=6.135 $Y2=1.94
r69 12 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.045 $Y=1.865
+ $X2=5.83 $Y2=1.865
r70 8 24 32.6451 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=5.755 $Y=1.355
+ $X2=5.755 $Y2=1.647
r71 8 10 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=5.755 $Y=1.355
+ $X2=5.755 $Y2=0.79
r72 5 20 28.0673 $w=1.8e-07 $l=2.93e-07 $layer=POLY_cond $X=5.44 $Y=1.94
+ $X2=5.44 $Y2=1.647
r73 5 7 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.44 $Y=1.94 $X2=5.44
+ $Y2=2.435
r74 1 19 32.6451 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=5.28 $Y=1.355
+ $X2=5.28 $Y2=1.647
r75 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=5.28 $Y=1.355
+ $X2=5.28 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%A_1238_94# 1 2 7 9 12 13 14 16 18 21 24 25
+ 28
c58 21 0 2.79353e-20 $X=6.56 $Y=1.3
c59 16 0 8.55731e-20 $X=6.36 $Y=1.89
c60 13 0 1.17701e-19 $X=7.09 $Y=1.36
r61 28 30 16.1243 $w=4.78e-07 $l=4.35e-07 $layer=LI1_cond $X=6.405 $Y=0.615
+ $X2=6.405 $Y2=1.05
r62 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.08
+ $Y=1.465 $X2=7.08 $Y2=1.465
r63 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.645 $Y=1.465
+ $X2=7.08 $Y2=1.465
r64 21 22 9.30874 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.56 $Y=1.3
+ $X2=6.475 $Y2=1.465
r65 21 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.56 $Y=1.3 $X2=6.56
+ $Y2=1.05
r66 16 22 16.4581 $w=3.3e-07 $l=4.79062e-07 $layer=LI1_cond $X=6.36 $Y=1.89
+ $X2=6.475 $Y2=1.465
r67 16 18 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.36 $Y=1.89
+ $X2=6.36 $Y2=2.16
r68 15 25 14.0139 $w=3.5e-07 $l=8.5e-08 $layer=POLY_cond $X=7.09 $Y=1.55
+ $X2=7.09 $Y2=1.465
r69 13 25 17.3113 $w=3.5e-07 $l=1.05e-07 $layer=POLY_cond $X=7.09 $Y=1.36
+ $X2=7.09 $Y2=1.465
r70 13 14 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.09 $Y=1.36
+ $X2=7.09 $Y2=1.185
r71 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.19 $Y=0.74
+ $X2=7.19 $Y2=1.185
r72 7 15 35.6367 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.09 $Y=1.725
+ $X2=7.09 $Y2=1.55
r73 7 9 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=7.09 $Y=1.725 $X2=7.09
+ $Y2=2.4
r74 2 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=2.015 $X2=6.36 $Y2=2.16
r75 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.19
+ $Y=0.47 $X2=6.33 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 40
+ 41 42 44 49 68 69 75 78
r85 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r89 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r90 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r94 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r96 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.15 $Y2=3.33
r98 57 59 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r100 53 56 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r101 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 52 55 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r103 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 50 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r105 50 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 49 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.15 $Y2=3.33
r107 49 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 48 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 48 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r110 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 45 72 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r112 45 47 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r113 44 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 44 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 42 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 42 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 40 65 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.48 $Y2=3.33
r118 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.86 $Y2=3.33
r119 39 68 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=6.86 $Y2=3.33
r121 37 62 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.585 $Y=3.33
+ $X2=5.52 $Y2=3.33
r122 37 38 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.585 $Y=3.33
+ $X2=5.787 $Y2=3.33
r123 36 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 36 38 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=5.787 $Y2=3.33
r125 32 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=3.33
r126 32 34 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=2.225
r127 28 38 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.787 $Y=3.245
+ $X2=5.787 $Y2=3.33
r128 28 30 6.97157 $w=4.03e-07 $l=2.45e-07 $layer=LI1_cond $X=5.787 $Y=3.245
+ $X2=5.787 $Y2=3
r129 24 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=3.33
r130 24 26 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=2.67
r131 20 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r132 20 22 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.825
r133 16 72 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r134 16 18 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.295
r135 5 34 300 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=2 $X=6.675
+ $Y=2.015 $X2=6.86 $Y2=2.225
r136 4 30 600 $w=1.7e-07 $l=1.10517e-06 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=2.015 $X2=5.785 $Y2=3
r137 3 26 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=2.46 $X2=4.15 $Y2=2.67
r138 2 22 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.84 $X2=1.68 $Y2=2.825
r139 1 18 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%A_114_112# 1 2 3 4 16 18 20 21 22 26 27 28
+ 31 33 35 39 40
r103 39 40 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0.565
+ $X2=2.125 $Y2=0.565
r104 35 37 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.12 $Y=2.405
+ $X2=1.54 $Y2=2.405
r105 29 31 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.735 $Y=2.32
+ $X2=2.735 $Y2=2.05
r106 28 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.405
+ $X2=1.54 $Y2=2.405
r107 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=2.735 $Y2=2.32
r108 27 28 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=1.625 $Y2=2.405
r109 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.32
+ $X2=1.54 $Y2=2.405
r110 25 26 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.54 $Y=1.46
+ $X2=1.54 $Y2=2.32
r111 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=1.375
+ $X2=1.54 $Y2=1.46
r112 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.455 $Y=1.375
+ $X2=0.885 $Y2=1.375
r113 20 40 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=0.885 $Y=0.625
+ $X2=2.125 $Y2=0.625
r114 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.29
+ $X2=0.885 $Y2=1.375
r115 18 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.8 $Y=1.29 $X2=0.8
+ $Y2=1.12
r116 14 33 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.715 $Y=0.95
+ $X2=0.715 $Y2=1.12
r117 14 16 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=0.95
+ $X2=0.715 $Y2=0.83
r118 13 20 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.715 $Y=0.71
+ $X2=0.885 $Y2=0.625
r119 13 16 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=0.71
+ $X2=0.715 $Y2=0.83
r120 4 31 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=1.895 $X2=2.775 $Y2=2.05
r121 3 35 300 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=2.12 $X2=1.12 $Y2=2.405
r122 2 39 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.37 $X2=2.29 $Y2=0.565
r123 1 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.71 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%GCLK 1 2 9 13 14 15 16 23 32
r20 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=7.41 $Y=1.995 $X2=7.41
+ $Y2=2.035
r21 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.41 $Y=2.405
+ $X2=7.41 $Y2=2.775
r22 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=7.41 $Y=1.972
+ $X2=7.41 $Y2=1.995
r23 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=7.41 $Y=1.972
+ $X2=7.41 $Y2=1.82
r24 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=7.41 $Y=2.057
+ $X2=7.41 $Y2=2.405
r25 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=7.41 $Y=2.057
+ $X2=7.41 $Y2=2.035
r26 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.5 $Y=1.13 $X2=7.5
+ $Y2=1.82
r27 7 13 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=7.412 $Y=0.958
+ $X2=7.412 $Y2=1.13
r28 7 9 14.798 $w=3.43e-07 $l=4.43e-07 $layer=LI1_cond $X=7.412 $Y=0.958
+ $X2=7.412 $Y2=0.515
r29 2 14 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=7.18
+ $Y=1.84 $X2=7.4 $Y2=1.985
r30 2 16 400 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=7.18
+ $Y=1.84 $X2=7.4 $Y2=2.815
r31 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.37 $X2=7.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_1%VGND 1 2 3 4 5 16 18 22 26 30 33 34 35 37
+ 49 56 63 64 71 77 80
r85 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r86 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r87 71 74 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.22
+ $Y2=0.285
r88 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r89 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r90 64 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r91 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r92 61 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.065 $Y=0 $X2=6.94
+ $Y2=0
r93 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.065 $Y=0 $X2=7.44
+ $Y2=0
r94 60 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r95 60 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r96 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 57 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.66 $Y=0 $X2=5.535
+ $Y2=0
r98 57 59 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.66 $Y=0 $X2=6.48
+ $Y2=0
r99 56 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.815 $Y=0 $X2=6.94
+ $Y2=0
r100 56 59 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=6.48 $Y2=0
r101 55 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r102 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r103 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r104 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r105 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r106 49 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.535
+ $Y2=0
r107 49 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.04
+ $Y2=0
r108 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r109 45 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r110 45 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r111 44 47 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r112 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r113 42 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r114 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r115 41 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r116 41 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r117 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r118 38 67 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r119 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r120 37 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r121 37 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r122 35 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r123 35 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r124 33 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.6
+ $Y2=0
r125 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.835
+ $Y2=0
r126 32 51 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=4.08
+ $Y2=0
r127 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=0 $X2=3.835
+ $Y2=0
r128 28 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.94 $Y=0.085
+ $X2=6.94 $Y2=0
r129 28 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.94 $Y=0.085
+ $X2=6.94 $Y2=0.515
r130 24 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=0.085
+ $X2=5.535 $Y2=0
r131 24 26 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=5.535 $Y=0.085
+ $X2=5.535 $Y2=0.615
r132 20 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0
r133 20 22 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0.545
r134 16 67 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r135 16 18 34.3428 $w=2.48e-07 $l=7.45e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.83
r136 5 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.37 $X2=6.9 $Y2=0.515
r137 4 26 91 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=2 $X=5.355
+ $Y=0.37 $X2=5.495 $Y2=0.615
r138 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.4 $X2=3.835 $Y2=0.545
r139 2 74 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.56 $X2=1.22 $Y2=0.285
r140 1 18 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.83
.ends


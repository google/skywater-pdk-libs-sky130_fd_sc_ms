* File: sky130_fd_sc_ms__a22o_2.pxi.spice
* Created: Wed Sep  2 11:53:12 2020
* 
x_PM_SKY130_FD_SC_MS__A22O_2%A_81_48# N_A_81_48#_M1008_d N_A_81_48#_M1003_d
+ N_A_81_48#_c_70_n N_A_81_48#_M1002_g N_A_81_48#_M1005_g N_A_81_48#_c_72_n
+ N_A_81_48#_M1009_g N_A_81_48#_M1007_g N_A_81_48#_c_82_p N_A_81_48#_c_74_n
+ N_A_81_48#_c_75_n N_A_81_48#_c_83_p N_A_81_48#_c_110_p N_A_81_48#_c_97_p
+ N_A_81_48#_c_76_n N_A_81_48#_c_77_n N_A_81_48#_c_100_p N_A_81_48#_c_78_n
+ PM_SKY130_FD_SC_MS__A22O_2%A_81_48#
x_PM_SKY130_FD_SC_MS__A22O_2%A1 N_A1_M1010_g N_A1_M1008_g A1 N_A1_c_153_n
+ N_A1_c_154_n PM_SKY130_FD_SC_MS__A22O_2%A1
x_PM_SKY130_FD_SC_MS__A22O_2%B1 N_B1_M1003_g N_B1_M1006_g B1 N_B1_c_190_n
+ N_B1_c_191_n PM_SKY130_FD_SC_MS__A22O_2%B1
x_PM_SKY130_FD_SC_MS__A22O_2%B2 N_B2_M1011_g N_B2_M1000_g B2 N_B2_c_230_n
+ PM_SKY130_FD_SC_MS__A22O_2%B2
x_PM_SKY130_FD_SC_MS__A22O_2%A2 N_A2_M1004_g N_A2_M1001_g A2 N_A2_c_264_n
+ N_A2_c_265_n PM_SKY130_FD_SC_MS__A22O_2%A2
x_PM_SKY130_FD_SC_MS__A22O_2%VPWR N_VPWR_M1005_s N_VPWR_M1007_s N_VPWR_M1001_d
+ N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n
+ N_VPWR_c_295_n VPWR N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n
+ N_VPWR_c_289_n PM_SKY130_FD_SC_MS__A22O_2%VPWR
x_PM_SKY130_FD_SC_MS__A22O_2%X N_X_M1002_s N_X_M1005_d N_X_c_340_n N_X_c_337_n
+ N_X_c_342_n X X X X X N_X_c_339_n PM_SKY130_FD_SC_MS__A22O_2%X
x_PM_SKY130_FD_SC_MS__A22O_2%A_391_368# N_A_391_368#_M1010_d
+ N_A_391_368#_M1000_d N_A_391_368#_c_372_n N_A_391_368#_c_368_n
+ N_A_391_368#_c_369_n N_A_391_368#_c_370_n
+ PM_SKY130_FD_SC_MS__A22O_2%A_391_368#
x_PM_SKY130_FD_SC_MS__A22O_2%VGND N_VGND_M1002_d N_VGND_M1009_d N_VGND_M1011_d
+ N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n
+ N_VGND_c_401_n VGND N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n
+ N_VGND_c_405_n PM_SKY130_FD_SC_MS__A22O_2%VGND
x_PM_SKY130_FD_SC_MS__A22O_2%A_304_74# N_A_304_74#_M1008_s N_A_304_74#_M1004_d
+ N_A_304_74#_c_442_n N_A_304_74#_c_443_n N_A_304_74#_c_444_n
+ N_A_304_74#_c_481_p N_A_304_74#_c_445_n N_A_304_74#_c_446_n
+ N_A_304_74#_c_447_n PM_SKY130_FD_SC_MS__A22O_2%A_304_74#
cc_1 VNB N_A_81_48#_c_70_n 0.0199307f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.22
cc_2 VNB N_A_81_48#_M1005_g 0.00704621f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_3 VNB N_A_81_48#_c_72_n 0.0176642f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.22
cc_4 VNB N_A_81_48#_M1007_g 0.00570843f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=2.4
cc_5 VNB N_A_81_48#_c_74_n 0.0167228f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.095
cc_6 VNB N_A_81_48#_c_75_n 0.00613798f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.095
cc_7 VNB N_A_81_48#_c_76_n 7.42537e-19 $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.385
cc_8 VNB N_A_81_48#_c_77_n 0.00233643f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.55
cc_9 VNB N_A_81_48#_c_78_n 0.0926783f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.385
cc_10 VNB N_A1_M1008_g 0.0275155f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.22
cc_11 VNB N_A1_c_153_n 0.0242693f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_12 VNB N_A1_c_154_n 0.00392334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1006_g 0.0237683f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.22
cc_14 VNB N_B1_c_190_n 0.0227283f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_15 VNB N_B1_c_191_n 0.00472951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B2_M1011_g 0.0251119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB B2 0.00585622f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_18 VNB N_B2_c_230_n 0.0215953f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_19 VNB N_A2_M1004_g 0.0345407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_264_n 0.047419f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_21 VNB N_A2_c_265_n 0.00404344f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_22 VNB N_VPWR_c_289_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.385
cc_23 VNB X 0.00650146f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.22
cc_24 VNB N_VGND_c_396_n 0.0101995f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.55
cc_25 VNB N_VGND_c_397_n 0.0511447f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_26 VNB N_VGND_c_398_n 0.0134317f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_27 VNB N_VGND_c_399_n 0.00941023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_400_n 0.0389074f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.55
cc_29 VNB N_VGND_c_401_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.95
cc_30 VNB N_VGND_c_402_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.035
cc_31 VNB N_VGND_c_403_n 0.0199471f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.115
cc_32 VNB N_VGND_c_404_n 0.237175f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.385
cc_33 VNB N_VGND_c_405_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_304_74#_c_442_n 0.00370491f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_35 VNB N_A_304_74#_c_443_n 0.0048983f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_36 VNB N_A_304_74#_c_444_n 0.00412286f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.4
cc_37 VNB N_A_304_74#_c_445_n 0.0137f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_38 VNB N_A_304_74#_c_446_n 0.00735846f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_39 VNB N_A_304_74#_c_447_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=2.4
cc_40 VPB N_A_81_48#_M1005_g 0.024634f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_41 VPB N_A_81_48#_M1007_g 0.0244082f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=2.4
cc_42 VPB N_A1_M1010_g 0.0209585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A1_c_153_n 0.00552325f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_44 VPB N_A1_c_154_n 0.0024898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B1_M1003_g 0.0197297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_B1_c_190_n 0.00539327f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_47 VPB N_B1_c_191_n 0.00374496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_B2_M1000_g 0.0204985f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.22
cc_49 VPB B2 0.00573291f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=0.74
cc_50 VPB N_B2_c_230_n 0.00539477f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_51 VPB N_A2_M1001_g 0.02605f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.22
cc_52 VPB N_A2_c_264_n 0.0112708f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_53 VPB N_A2_c_265_n 0.00689237f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_54 VPB N_VPWR_c_290_n 0.0458603f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_55 VPB N_VPWR_c_291_n 0.00715805f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_56 VPB N_VPWR_c_292_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=2.4
cc_57 VPB N_VPWR_c_293_n 0.0517798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_294_n 0.017577f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=1.55
cc_59 VPB N_VPWR_c_295_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=1.95
cc_60 VPB N_VPWR_c_296_n 0.0182909f $X=-0.19 $Y=1.66 $X2=2.165 $Y2=0.76
cc_61 VPB N_VPWR_c_297_n 0.0411787f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.385
cc_62 VPB N_VPWR_c_298_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.385
cc_63 VPB N_VPWR_c_289_n 0.0856496f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.385
cc_64 VPB N_X_c_337_n 0.00202402f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_65 VPB X 0.00296132f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=1.22
cc_66 VPB N_X_c_339_n 0.00952367f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.55
cc_67 VPB N_A_391_368#_c_368_n 0.0138881f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_68 VPB N_A_391_368#_c_369_n 0.00322986f $X=-0.19 $Y=1.66 $X2=0.875 $Y2=2.4
cc_69 VPB N_A_391_368#_c_370_n 6.76734e-19 $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_70 N_A_81_48#_M1007_g N_A1_M1010_g 0.028559f $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_71 N_A_81_48#_c_82_p N_A1_M1010_g 0.00112695f $X=1.33 $Y=1.95 $X2=0 $Y2=0
cc_72 N_A_81_48#_c_83_p N_A1_M1010_g 0.0182384f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_73 N_A_81_48#_c_74_n N_A1_M1008_g 0.0160603f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_74 N_A_81_48#_c_76_n N_A1_M1008_g 0.0019081f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_75 N_A_81_48#_c_78_n N_A1_M1008_g 0.00473768f $X=1.325 $Y=1.385 $X2=0 $Y2=0
cc_76 N_A_81_48#_c_74_n N_A1_c_153_n 0.00126608f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_77 N_A_81_48#_c_83_p N_A1_c_153_n 7.14077e-19 $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A_81_48#_c_76_n N_A1_c_153_n 3.80775e-19 $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_79 N_A_81_48#_c_78_n N_A1_c_153_n 0.0210127f $X=1.325 $Y=1.385 $X2=0 $Y2=0
cc_80 N_A_81_48#_c_74_n N_A1_c_154_n 0.0243073f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_81 N_A_81_48#_c_83_p N_A1_c_154_n 0.0225056f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_82 N_A_81_48#_c_76_n N_A1_c_154_n 0.03304f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_83 N_A_81_48#_c_78_n N_A1_c_154_n 0.00260729f $X=1.325 $Y=1.385 $X2=0 $Y2=0
cc_84 N_A_81_48#_c_83_p N_B1_M1003_g 0.0142175f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_81_48#_c_74_n N_B1_M1006_g 0.00442568f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_86 N_A_81_48#_c_97_p N_B1_M1006_g 0.00514063f $X=2.165 $Y=0.76 $X2=0 $Y2=0
cc_87 N_A_81_48#_c_74_n N_B1_c_190_n 0.00355719f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_88 N_A_81_48#_c_83_p N_B1_c_190_n 2.24228e-19 $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_89 N_A_81_48#_c_100_p N_B1_c_190_n 2.2901e-19 $X=2.54 $Y=2.115 $X2=0 $Y2=0
cc_90 N_A_81_48#_c_74_n N_B1_c_191_n 0.0219116f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_91 N_A_81_48#_c_83_p N_B1_c_191_n 0.0251439f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_81_48#_c_100_p N_B1_c_191_n 0.00322171f $X=2.54 $Y=2.115 $X2=0 $Y2=0
cc_93 N_A_81_48#_c_83_p N_VPWR_M1007_s 0.00814324f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_81_48#_M1005_g N_VPWR_c_290_n 0.00770724f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A_81_48#_c_78_n N_VPWR_c_290_n 0.00150952f $X=1.325 $Y=1.385 $X2=0 $Y2=0
cc_96 N_A_81_48#_M1005_g N_VPWR_c_291_n 5.60169e-19 $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_81_48#_M1007_g N_VPWR_c_291_n 0.0145637f $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_81_48#_c_83_p N_VPWR_c_291_n 0.0196888f $X=2.455 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_81_48#_c_110_p N_VPWR_c_291_n 0.00237022f $X=1.415 $Y=2.035 $X2=0
+ $Y2=0
cc_100 N_A_81_48#_M1005_g N_VPWR_c_296_n 0.0048691f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_81_48#_M1007_g N_VPWR_c_296_n 0.00460063f $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_81_48#_M1005_g N_VPWR_c_289_n 0.00877338f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_81_48#_M1007_g N_VPWR_c_289_n 0.00908554f $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_81_48#_M1005_g N_X_c_340_n 0.00193479f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_81_48#_M1005_g N_X_c_337_n 0.008336f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_81_48#_M1005_g N_X_c_342_n 0.0130445f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_81_48#_M1007_g N_X_c_342_n 0.00474657f $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_81_48#_c_82_p N_X_c_342_n 0.00417842f $X=1.33 $Y=1.95 $X2=0 $Y2=0
cc_109 N_A_81_48#_c_110_p N_X_c_342_n 0.0133619f $X=1.415 $Y=2.035 $X2=0 $Y2=0
cc_110 N_A_81_48#_c_70_n X 0.0148558f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_111 N_A_81_48#_M1005_g X 0.0067259f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_81_48#_c_72_n X 0.0177235f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A_81_48#_M1007_g X 4.97449e-19 $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_81_48#_c_82_p X 0.0062516f $X=1.33 $Y=1.95 $X2=0 $Y2=0
cc_115 N_A_81_48#_c_75_n X 0.011439f $X=1.415 $Y=1.095 $X2=0 $Y2=0
cc_116 N_A_81_48#_c_76_n X 0.0222666f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A_81_48#_c_78_n X 0.0361511f $X=1.325 $Y=1.385 $X2=0 $Y2=0
cc_118 N_A_81_48#_M1005_g N_X_c_339_n 0.0175969f $X=0.875 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_81_48#_M1007_g N_X_c_339_n 0.00106863f $X=1.325 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_81_48#_c_82_p N_X_c_339_n 0.0132162f $X=1.33 $Y=1.95 $X2=0 $Y2=0
cc_121 N_A_81_48#_c_78_n N_X_c_339_n 0.00197664f $X=1.325 $Y=1.385 $X2=0 $Y2=0
cc_122 N_A_81_48#_c_83_p N_A_391_368#_M1010_d 0.00502116f $X=2.455 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_123 N_A_81_48#_c_83_p N_A_391_368#_c_372_n 0.0170259f $X=2.455 $Y=2.035 $X2=0
+ $Y2=0
cc_124 N_A_81_48#_c_100_p N_A_391_368#_c_368_n 0.0175414f $X=2.54 $Y=2.115 $X2=0
+ $Y2=0
cc_125 N_A_81_48#_M1007_g N_A_391_368#_c_369_n 4.90595e-19 $X=1.325 $Y=2.4 $X2=0
+ $Y2=0
cc_126 N_A_81_48#_c_75_n N_VGND_M1009_d 0.0030302f $X=1.415 $Y=1.095 $X2=0 $Y2=0
cc_127 N_A_81_48#_c_70_n N_VGND_c_397_n 0.00647412f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_128 N_A_81_48#_c_72_n N_VGND_c_398_n 0.00698798f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_129 N_A_81_48#_c_75_n N_VGND_c_398_n 0.0182898f $X=1.415 $Y=1.095 $X2=0 $Y2=0
cc_130 N_A_81_48#_c_78_n N_VGND_c_398_n 0.00259348f $X=1.325 $Y=1.385 $X2=0
+ $Y2=0
cc_131 N_A_81_48#_c_70_n N_VGND_c_402_n 0.00434272f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_132 N_A_81_48#_c_72_n N_VGND_c_402_n 0.00434272f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_81_48#_c_70_n N_VGND_c_404_n 0.00823889f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A_81_48#_c_72_n N_VGND_c_404_n 0.00825283f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_135 N_A_81_48#_c_74_n N_A_304_74#_M1008_s 0.00271234f $X=2 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_81_48#_c_74_n N_A_304_74#_c_442_n 0.021673f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_137 N_A_81_48#_M1008_d N_A_304_74#_c_443_n 0.00250873f $X=1.955 $Y=0.37 $X2=0
+ $Y2=0
cc_138 N_A_81_48#_c_74_n N_A_304_74#_c_443_n 0.00304353f $X=2 $Y=1.095 $X2=0
+ $Y2=0
cc_139 N_A_81_48#_c_97_p N_A_304_74#_c_443_n 0.0194097f $X=2.165 $Y=0.76 $X2=0
+ $Y2=0
cc_140 N_A_81_48#_c_74_n N_A_304_74#_c_446_n 0.0104256f $X=2 $Y=1.095 $X2=0
+ $Y2=0
cc_141 N_A1_M1010_g N_B1_M1003_g 0.0305861f $X=1.865 $Y=2.34 $X2=0 $Y2=0
cc_142 N_A1_M1008_g N_B1_M1006_g 0.0301069f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_c_153_n N_B1_c_190_n 0.0205009f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A1_c_154_n N_B1_c_190_n 3.16506e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_153_n N_B1_c_191_n 0.00276344f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A1_c_154_n N_B1_c_191_n 0.034584f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A1_M1010_g N_VPWR_c_291_n 0.00630856f $X=1.865 $Y=2.34 $X2=0 $Y2=0
cc_148 N_A1_M1010_g N_VPWR_c_297_n 0.00508554f $X=1.865 $Y=2.34 $X2=0 $Y2=0
cc_149 N_A1_M1010_g N_VPWR_c_289_n 0.00508379f $X=1.865 $Y=2.34 $X2=0 $Y2=0
cc_150 N_A1_M1010_g N_A_391_368#_c_372_n 0.00866597f $X=1.865 $Y=2.34 $X2=0
+ $Y2=0
cc_151 N_A1_M1010_g N_A_391_368#_c_369_n 0.00203526f $X=1.865 $Y=2.34 $X2=0
+ $Y2=0
cc_152 N_A1_M1008_g N_VGND_c_398_n 0.00174891f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1008_g N_VGND_c_400_n 0.00278247f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_M1008_g N_VGND_c_404_n 0.00359137f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_M1008_g N_A_304_74#_c_442_n 0.00730569f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A1_M1008_g N_A_304_74#_c_443_n 0.008259f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_M1008_g N_A_304_74#_c_444_n 0.00395315f $X=1.88 $Y=0.74 $X2=0 $Y2=0
cc_158 N_B1_M1006_g N_B2_M1011_g 0.0500418f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_159 N_B1_M1003_g N_B2_M1000_g 0.0196708f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_160 N_B1_c_191_n N_B2_M1000_g 3.72642e-19 $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_161 N_B1_M1003_g B2 3.32938e-19 $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_162 N_B1_c_190_n B2 4.13747e-19 $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_163 N_B1_c_191_n B2 0.0297654f $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_164 N_B1_c_190_n N_B2_c_230_n 0.0214219f $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_165 N_B1_c_191_n N_B2_c_230_n 4.14948e-19 $X=2.33 $Y=1.515 $X2=0 $Y2=0
cc_166 N_B1_M1003_g N_VPWR_c_297_n 8.89343e-19 $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_167 N_B1_M1003_g N_A_391_368#_c_372_n 0.00986711f $X=2.315 $Y=2.34 $X2=0
+ $Y2=0
cc_168 N_B1_M1003_g N_A_391_368#_c_368_n 0.0107571f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_169 N_B1_M1003_g N_A_391_368#_c_369_n 0.00141162f $X=2.315 $Y=2.34 $X2=0
+ $Y2=0
cc_170 N_B1_M1003_g N_A_391_368#_c_370_n 5.9276e-19 $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_171 N_B1_M1006_g N_VGND_c_400_n 0.00278271f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B1_M1006_g N_VGND_c_404_n 0.00353949f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B1_M1006_g N_A_304_74#_c_442_n 4.62714e-19 $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B1_M1006_g N_A_304_74#_c_443_n 0.0127288f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B1_M1006_g N_A_304_74#_c_446_n 9.3266e-19 $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B2_M1011_g N_A2_M1004_g 0.024575f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B2_M1000_g N_A2_M1001_g 0.00972574f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_178 B2 N_A2_c_264_n 0.00380277f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B2_c_230_n N_A2_c_264_n 0.020946f $X=2.87 $Y=1.515 $X2=0 $Y2=0
cc_180 B2 N_A2_c_265_n 0.035317f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_181 N_B2_c_230_n N_A2_c_265_n 2.2561e-19 $X=2.87 $Y=1.515 $X2=0 $Y2=0
cc_182 N_B2_M1000_g N_VPWR_c_293_n 2.89901e-19 $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_183 N_B2_M1000_g N_VPWR_c_297_n 8.89343e-19 $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_184 N_B2_M1000_g N_A_391_368#_c_372_n 5.6976e-19 $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_185 N_B2_M1000_g N_A_391_368#_c_368_n 0.0122144f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_186 N_B2_M1000_g N_A_391_368#_c_370_n 0.0134078f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_187 B2 N_A_391_368#_c_370_n 0.0263427f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B2_c_230_n N_A_391_368#_c_370_n 6.58373e-19 $X=2.87 $Y=1.515 $X2=0
+ $Y2=0
cc_189 N_B2_M1011_g N_VGND_c_399_n 0.00225437f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B2_M1011_g N_VGND_c_400_n 0.00461464f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B2_M1011_g N_VGND_c_404_n 0.00908275f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_192 N_B2_M1011_g N_A_304_74#_c_443_n 0.00120883f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_193 N_B2_M1011_g N_A_304_74#_c_445_n 0.014921f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_194 B2 N_A_304_74#_c_445_n 0.0409488f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_195 N_B2_c_230_n N_A_304_74#_c_445_n 0.00423269f $X=2.87 $Y=1.515 $X2=0 $Y2=0
cc_196 N_B2_M1011_g N_A_304_74#_c_447_n 8.17877e-19 $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A2_M1001_g N_VPWR_c_293_n 0.0193639f $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_198 N_A2_c_264_n N_VPWR_c_293_n 0.00169678f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A2_c_265_n N_VPWR_c_293_n 0.0255649f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A2_M1001_g N_VPWR_c_297_n 0.00492916f $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_201 N_A2_M1001_g N_VPWR_c_289_n 0.00511769f $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_202 N_A2_M1001_g N_A_391_368#_c_368_n 6.34081e-19 $X=3.335 $Y=2.34 $X2=0
+ $Y2=0
cc_203 N_A2_M1001_g N_A_391_368#_c_370_n 5.8566e-19 $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_204 N_A2_M1004_g N_VGND_c_399_n 0.00600897f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A2_M1004_g N_VGND_c_403_n 0.00434272f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A2_M1004_g N_VGND_c_404_n 0.00824829f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A2_M1004_g N_A_304_74#_c_445_n 0.0185399f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A2_c_264_n N_A_304_74#_c_445_n 0.00285738f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_209 N_A2_c_265_n N_A_304_74#_c_445_n 0.0253731f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A2_M1004_g N_A_304_74#_c_447_n 0.0102372f $X=3.32 $Y=0.74 $X2=0 $Y2=0
cc_211 N_VPWR_c_291_n N_X_c_337_n 0.02342f $X=1.55 $Y=2.375 $X2=0 $Y2=0
cc_212 N_VPWR_c_296_n N_X_c_337_n 0.0122335f $X=1.385 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_289_n N_X_c_337_n 0.0099849f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_290_n N_X_c_342_n 0.0337292f $X=0.65 $Y=2.225 $X2=0 $Y2=0
cc_215 N_VPWR_M1005_s N_X_c_339_n 0.00446079f $X=0.525 $Y=1.84 $X2=0 $Y2=0
cc_216 N_VPWR_c_290_n N_X_c_339_n 0.016109f $X=0.65 $Y=2.225 $X2=0 $Y2=0
cc_217 N_VPWR_c_291_n N_A_391_368#_c_372_n 0.0406486f $X=1.55 $Y=2.375 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_293_n N_A_391_368#_c_368_n 0.0147692f $X=3.56 $Y=2.115 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_297_n N_A_391_368#_c_368_n 0.0649714f $X=3.395 $Y=3.33 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_289_n N_A_391_368#_c_368_n 0.0369098f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_291_n N_A_391_368#_c_369_n 0.0126523f $X=1.55 $Y=2.375 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_297_n N_A_391_368#_c_369_n 0.0236566f $X=3.395 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_289_n N_A_391_368#_c_369_n 0.0128296f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_293_n N_A_391_368#_c_370_n 0.0384784f $X=3.56 $Y=2.115 $X2=0
+ $Y2=0
cc_225 X N_VGND_c_397_n 0.0294122f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_226 X N_VGND_c_398_n 0.0182902f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_227 X N_VGND_c_402_n 0.0144922f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_228 X N_VGND_c_404_n 0.0118826f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_229 N_VGND_c_398_n N_A_304_74#_c_442_n 0.0291511f $X=1.125 $Y=0.675 $X2=0
+ $Y2=0
cc_230 N_VGND_c_399_n N_A_304_74#_c_443_n 0.00898192f $X=3.035 $Y=0.675 $X2=0
+ $Y2=0
cc_231 N_VGND_c_400_n N_A_304_74#_c_443_n 0.0544911f $X=2.87 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_404_n N_A_304_74#_c_443_n 0.0305408f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_398_n N_A_304_74#_c_444_n 0.0127054f $X=1.125 $Y=0.675 $X2=0
+ $Y2=0
cc_234 N_VGND_c_400_n N_A_304_74#_c_444_n 0.0233048f $X=2.87 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_404_n N_A_304_74#_c_444_n 0.0126653f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_M1011_d N_A_304_74#_c_445_n 0.00309832f $X=2.855 $Y=0.37 $X2=0
+ $Y2=0
cc_237 N_VGND_c_399_n N_A_304_74#_c_445_n 0.022455f $X=3.035 $Y=0.675 $X2=0
+ $Y2=0
cc_238 N_VGND_c_399_n N_A_304_74#_c_447_n 0.0191765f $X=3.035 $Y=0.675 $X2=0
+ $Y2=0
cc_239 N_VGND_c_403_n N_A_304_74#_c_447_n 0.0145639f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_404_n N_A_304_74#_c_447_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_241 N_A_304_74#_c_481_p A_491_74# 0.00196494f $X=2.585 $Y=1.01 $X2=-0.19
+ $Y2=-0.245

* File: sky130_fd_sc_ms__sdlclkp_1.pxi.spice
* Created: Wed Sep  2 12:32:03 2020
* 
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%SCE N_SCE_c_154_n N_SCE_M1008_g N_SCE_M1013_g
+ N_SCE_c_160_n SCE N_SCE_c_156_n N_SCE_c_157_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%SCE
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%GATE N_GATE_M1000_g N_GATE_M1012_g GATE
+ N_GATE_c_190_n N_GATE_c_191_n PM_SKY130_FD_SC_MS__SDLCLKP_1%GATE
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%A_318_74# N_A_318_74#_M1003_d
+ N_A_318_74#_M1021_d N_A_318_74#_M1011_g N_A_318_74#_M1015_g
+ N_A_318_74#_c_233_n N_A_318_74#_c_234_n N_A_318_74#_c_235_n
+ N_A_318_74#_c_236_n N_A_318_74#_c_237_n N_A_318_74#_c_238_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%A_318_74#
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%A_288_48# N_A_288_48#_M1005_s
+ N_A_288_48#_M1020_s N_A_288_48#_c_306_n N_A_288_48#_M1003_g
+ N_A_288_48#_c_307_n N_A_288_48#_c_308_n N_A_288_48#_M1021_g
+ N_A_288_48#_c_326_n N_A_288_48#_c_327_n N_A_288_48#_c_310_n
+ N_A_288_48#_c_311_n N_A_288_48#_c_312_n N_A_288_48#_M1017_g
+ N_A_288_48#_M1002_g N_A_288_48#_c_313_n N_A_288_48#_c_314_n
+ N_A_288_48#_c_315_n N_A_288_48#_c_316_n N_A_288_48#_c_317_n
+ N_A_288_48#_c_318_n N_A_288_48#_c_367_p N_A_288_48#_c_319_n
+ N_A_288_48#_c_320_n N_A_288_48#_c_321_n N_A_288_48#_c_322_n
+ N_A_288_48#_c_323_n N_A_288_48#_c_324_n N_A_288_48#_c_330_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%A_288_48#
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%A_709_54# N_A_709_54#_M1010_d
+ N_A_709_54#_M1001_d N_A_709_54#_M1016_g N_A_709_54#_M1018_g
+ N_A_709_54#_c_466_n N_A_709_54#_M1007_g N_A_709_54#_M1009_g
+ N_A_709_54#_c_477_n N_A_709_54#_c_468_n N_A_709_54#_c_469_n
+ N_A_709_54#_c_479_n N_A_709_54#_c_480_n N_A_709_54#_c_470_n
+ N_A_709_54#_c_471_n N_A_709_54#_c_482_n N_A_709_54#_c_483_n
+ N_A_709_54#_c_472_n N_A_709_54#_c_473_n N_A_709_54#_c_484_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%A_709_54#
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%A_566_74# N_A_566_74#_M1017_d
+ N_A_566_74#_M1011_d N_A_566_74#_c_589_n N_A_566_74#_M1010_g
+ N_A_566_74#_M1001_g N_A_566_74#_c_591_n N_A_566_74#_c_592_n
+ N_A_566_74#_c_593_n N_A_566_74#_c_594_n N_A_566_74#_c_599_n
+ N_A_566_74#_c_595_n N_A_566_74#_c_596_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%A_566_74#
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%CLK N_CLK_M1005_g N_CLK_c_675_n N_CLK_M1020_g
+ N_CLK_M1006_g N_CLK_c_676_n N_CLK_c_673_n N_CLK_c_678_n N_CLK_M1004_g CLK
+ N_CLK_c_674_n PM_SKY130_FD_SC_MS__SDLCLKP_1%CLK
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%A_1238_94# N_A_1238_94#_M1007_d
+ N_A_1238_94#_M1004_d N_A_1238_94#_c_730_n N_A_1238_94#_M1014_g
+ N_A_1238_94#_M1019_g N_A_1238_94#_c_731_n N_A_1238_94#_c_732_n
+ N_A_1238_94#_c_733_n N_A_1238_94#_c_740_n N_A_1238_94#_c_734_n
+ N_A_1238_94#_c_735_n N_A_1238_94#_c_736_n N_A_1238_94#_c_737_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%A_1238_94#
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%VPWR N_VPWR_M1008_s N_VPWR_M1021_s
+ N_VPWR_M1018_d N_VPWR_M1020_d N_VPWR_M1009_d N_VPWR_c_789_n N_VPWR_c_790_n
+ N_VPWR_c_791_n N_VPWR_c_792_n N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n
+ N_VPWR_c_796_n N_VPWR_c_797_n N_VPWR_c_798_n VPWR N_VPWR_c_799_n
+ N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_788_n N_VPWR_c_803_n N_VPWR_c_804_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%VPWR
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%A_114_112# N_A_114_112#_M1013_d
+ N_A_114_112#_M1017_s N_A_114_112#_M1000_d N_A_114_112#_M1011_s
+ N_A_114_112#_c_886_n N_A_114_112#_c_873_n N_A_114_112#_c_874_n
+ N_A_114_112#_c_875_n N_A_114_112#_c_876_n N_A_114_112#_c_877_n
+ N_A_114_112#_c_882_n N_A_114_112#_c_883_n N_A_114_112#_c_884_n
+ N_A_114_112#_c_878_n N_A_114_112#_c_885_n N_A_114_112#_c_879_n
+ N_A_114_112#_c_880_n PM_SKY130_FD_SC_MS__SDLCLKP_1%A_114_112#
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%GCLK N_GCLK_M1019_d N_GCLK_M1014_d
+ N_GCLK_c_976_n N_GCLK_c_977_n GCLK GCLK GCLK GCLK N_GCLK_c_978_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%GCLK
x_PM_SKY130_FD_SC_MS__SDLCLKP_1%VGND N_VGND_M1013_s N_VGND_M1012_d
+ N_VGND_M1016_d N_VGND_M1005_d N_VGND_M1019_s N_VGND_c_996_n N_VGND_c_997_n
+ N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n
+ VGND N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_1%VGND
cc_1 VNB N_SCE_c_154_n 0.0157839f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.773
cc_2 VNB N_SCE_M1013_g 0.0259568f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB N_SCE_c_156_n 0.0236738f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_4 VNB N_SCE_c_157_n 0.0150641f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_5 VNB N_GATE_M1012_g 0.0408954f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_6 VNB N_GATE_c_190_n 0.0075224f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_GATE_c_191_n 0.00329566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_318_74#_M1015_g 0.0389156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_318_74#_c_233_n 0.00339384f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_10 VNB N_A_318_74#_c_234_n 0.00231274f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.29
cc_11 VNB N_A_318_74#_c_235_n 0.00736224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_318_74#_c_236_n 0.00390824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_318_74#_c_237_n 0.00408366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_318_74#_c_238_n 0.044129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_48#_c_306_n 0.0220743f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_16 VNB N_A_288_48#_c_307_n 0.0226305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_288_48#_c_308_n 0.00998942f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.96
cc_18 VNB N_A_288_48#_M1021_g 0.0193086f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_19 VNB N_A_288_48#_c_310_n 0.0289975f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_20 VNB N_A_288_48#_c_311_n 0.0486968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_288_48#_c_312_n 0.0185017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_288_48#_c_313_n 0.00119764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_288_48#_c_314_n 0.00547716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_288_48#_c_315_n 0.00507066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_288_48#_c_316_n 3.42301e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_288_48#_c_317_n 0.00855195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_288_48#_c_318_n 0.00227124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_288_48#_c_319_n 0.0162494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_288_48#_c_320_n 0.0018167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_288_48#_c_321_n 0.00525123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_288_48#_c_322_n 0.0107853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_288_48#_c_323_n 0.0090122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_288_48#_c_324_n 0.00699471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_709_54#_M1016_g 0.0520948f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_35 VNB N_A_709_54#_c_466_n 0.0183947f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_36 VNB N_A_709_54#_M1009_g 0.00607584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_709_54#_c_468_n 0.00310352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_709_54#_c_469_n 0.00569356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_709_54#_c_470_n 0.00230943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_709_54#_c_471_n 0.00109471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_709_54#_c_472_n 0.00886798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_709_54#_c_473_n 0.0520876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_566_74#_c_589_n 0.0210688f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_44 VNB N_A_566_74#_M1001_g 0.002121f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_45 VNB N_A_566_74#_c_591_n 0.00288593f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_46 VNB N_A_566_74#_c_592_n 0.00111963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_566_74#_c_593_n 0.0123613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_566_74#_c_594_n 0.00271082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_566_74#_c_595_n 0.00512979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_566_74#_c_596_n 0.0506641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_CLK_M1005_g 0.0287493f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.96
cc_52 VNB N_CLK_M1006_g 0.0225156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_CLK_c_673_n 0.0389302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_CLK_c_674_n 0.00149199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1238_94#_c_730_n 0.00818435f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_56 VNB N_A_1238_94#_c_731_n 0.0203644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1238_94#_c_732_n 0.0216435f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.455
cc_58 VNB N_A_1238_94#_c_733_n 0.00126393f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.455
cc_59 VNB N_A_1238_94#_c_734_n 0.00338577f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.625
cc_60 VNB N_A_1238_94#_c_735_n 0.0110227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1238_94#_c_736_n 0.0137359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1238_94#_c_737_n 0.0126688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VPWR_c_788_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_114_112#_c_873_n 0.00158689f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_65 VNB N_A_114_112#_c_874_n 0.00325089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_114_112#_c_875_n 0.0152342f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.625
cc_67 VNB N_A_114_112#_c_876_n 0.00499122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_114_112#_c_877_n 0.0042758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_114_112#_c_878_n 0.00507239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_114_112#_c_879_n 0.0064939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_114_112#_c_880_n 0.00971962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_GCLK_c_976_n 0.0264315f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_73 VNB N_GCLK_c_977_n 0.0128764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_GCLK_c_978_n 0.0248543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_996_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_76 VNB N_VGND_c_997_n 0.0503666f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_77 VNB N_VGND_c_998_n 0.00818657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_999_n 0.0148257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1000_n 0.0138206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1001_n 0.0594191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1002_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1003_n 0.0191862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1004_n 0.0363448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1005_n 0.0336226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1006_n 0.0190343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1007_n 0.450913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1008_n 0.0174852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1009_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1010_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VPB N_SCE_c_154_n 0.00952442f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.773
cc_91 VPB N_SCE_M1008_g 0.0274725f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_92 VPB N_SCE_c_160_n 0.0209371f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.96
cc_93 VPB N_SCE_c_157_n 0.0123756f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_94 VPB N_GATE_M1000_g 0.0246442f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.96
cc_95 VPB N_GATE_c_190_n 0.0283429f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_96 VPB N_GATE_c_191_n 0.00393454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_318_74#_M1011_g 0.0259851f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_98 VPB N_A_318_74#_c_234_n 0.00391009f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_99 VPB N_A_318_74#_c_236_n 0.00739397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_318_74#_c_237_n 0.00364869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_318_74#_c_238_n 0.0212067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_288_48#_M1021_g 0.0428327f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_103 VPB N_A_288_48#_c_326_n 0.113012f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_104 VPB N_A_288_48#_c_327_n 0.0140012f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.29
cc_105 VPB N_A_288_48#_M1002_g 0.0311075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_288_48#_c_322_n 0.00786399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_288_48#_c_330_n 0.00791546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_709_54#_M1016_g 0.00830614f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_109 VPB N_A_709_54#_M1018_g 0.032817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_709_54#_M1009_g 0.0323645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_709_54#_c_477_n 0.0060628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_709_54#_c_469_n 0.00145732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_709_54#_c_479_n 0.00418248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_709_54#_c_480_n 0.0117992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_709_54#_c_470_n 0.00314059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_709_54#_c_482_n 0.00887083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_709_54#_c_483_n 0.00705426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_709_54#_c_484_n 0.0508441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_566_74#_M1001_g 0.0291734f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_120 VPB N_A_566_74#_c_592_n 0.00732788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_566_74#_c_599_n 0.00120182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_CLK_c_675_n 0.0211217f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_123 VPB N_CLK_c_676_n 0.0207408f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_124 VPB N_CLK_c_673_n 0.0376269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_CLK_c_678_n 0.0171835f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.455
cc_126 VPB N_CLK_c_674_n 0.00107524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_1238_94#_c_730_n 0.0372561f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.29
cc_128 VPB N_A_1238_94#_c_733_n 0.00336531f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_129 VPB N_A_1238_94#_c_740_n 0.00275677f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_130 VPB N_VPWR_c_789_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_131 VPB N_VPWR_c_790_n 0.0419079f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.625
cc_132 VPB N_VPWR_c_791_n 0.0160989f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_792_n 0.0118948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_793_n 0.016159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_794_n 0.0103958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_795_n 0.0349499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_796_n 0.0077576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_797_n 0.0202398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_798_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_799_n 0.0312656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_800_n 0.0651369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_801_n 0.0201101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_788_n 0.102449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_803_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_804_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_114_112#_c_877_n 0.00930031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_114_112#_c_882_n 0.0134128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_114_112#_c_883_n 0.0122028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_114_112#_c_884_n 0.00639338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_114_112#_c_885_n 0.0083372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB GCLK 0.0136079f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.455
cc_152 VPB GCLK 0.0416896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_GCLK_c_978_n 0.00778235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 N_SCE_c_160_n N_GATE_M1000_g 0.04427f $X=0.407 $Y=1.96 $X2=0 $Y2=0
cc_155 N_SCE_M1013_g N_GATE_M1012_g 0.0205103f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_156 N_SCE_c_156_n N_GATE_M1012_g 0.0173046f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_157 N_SCE_c_157_n N_GATE_M1012_g 0.00112397f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_158 N_SCE_c_154_n N_GATE_c_190_n 0.04427f $X=0.407 $Y=1.773 $X2=0 $Y2=0
cc_159 N_SCE_c_157_n N_GATE_c_190_n 0.00106303f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_160 N_SCE_c_154_n N_GATE_c_191_n 0.00242614f $X=0.407 $Y=1.773 $X2=0 $Y2=0
cc_161 N_SCE_c_157_n N_GATE_c_191_n 0.0184673f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_162 N_SCE_M1008_g N_VPWR_c_790_n 0.0234401f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_163 N_SCE_c_160_n N_VPWR_c_790_n 0.00506126f $X=0.407 $Y=1.96 $X2=0 $Y2=0
cc_164 N_SCE_c_157_n N_VPWR_c_790_n 0.0254849f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_165 N_SCE_M1008_g N_VPWR_c_799_n 0.00460063f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_166 N_SCE_M1008_g N_VPWR_c_788_n 0.00908061f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_167 N_SCE_M1013_g N_A_114_112#_c_886_n 0.00259685f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_168 N_SCE_M1013_g N_A_114_112#_c_873_n 0.00358583f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_169 N_SCE_M1013_g N_A_114_112#_c_874_n 0.00332504f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_170 N_SCE_c_156_n N_A_114_112#_c_876_n 0.00130413f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_171 N_SCE_c_157_n N_A_114_112#_c_876_n 0.0145604f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_172 N_SCE_M1008_g N_A_114_112#_c_883_n 4.56234e-19 $X=0.505 $Y=2.54 $X2=0
+ $Y2=0
cc_173 N_SCE_M1013_g N_A_114_112#_c_878_n 0.00419565f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_174 N_SCE_c_156_n N_A_114_112#_c_878_n 0.00118053f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_175 N_SCE_M1008_g N_A_114_112#_c_885_n 0.00133673f $X=0.505 $Y=2.54 $X2=0
+ $Y2=0
cc_176 N_SCE_M1013_g N_VGND_c_997_n 0.00819892f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_177 N_SCE_c_156_n N_VGND_c_997_n 0.00386581f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_178 N_SCE_c_157_n N_VGND_c_997_n 0.0216167f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_179 N_SCE_M1013_g N_VGND_c_1003_n 0.00432822f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_180 N_SCE_M1013_g N_VGND_c_1007_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_181 N_GATE_M1012_g N_A_318_74#_c_235_n 0.00108365f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_182 N_GATE_M1012_g N_A_288_48#_c_306_n 0.0251298f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_183 N_GATE_M1000_g N_VPWR_c_790_n 0.00322746f $X=0.895 $Y=2.54 $X2=0 $Y2=0
cc_184 N_GATE_c_191_n N_VPWR_c_790_n 8.45929e-19 $X=0.97 $Y=1.795 $X2=0 $Y2=0
cc_185 N_GATE_M1000_g N_VPWR_c_791_n 0.00340497f $X=0.895 $Y=2.54 $X2=0 $Y2=0
cc_186 N_GATE_M1000_g N_VPWR_c_799_n 0.005209f $X=0.895 $Y=2.54 $X2=0 $Y2=0
cc_187 N_GATE_M1000_g N_VPWR_c_788_n 0.00983388f $X=0.895 $Y=2.54 $X2=0 $Y2=0
cc_188 N_GATE_c_191_n N_A_114_112#_M1000_d 0.00250903f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_189 N_GATE_M1012_g N_A_114_112#_c_886_n 0.00510645f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_190 N_GATE_M1012_g N_A_114_112#_c_873_n 0.00455954f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_191 N_GATE_M1012_g N_A_114_112#_c_874_n 0.00216557f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_192 N_GATE_M1012_g N_A_114_112#_c_875_n 0.009786f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_193 N_GATE_c_190_n N_A_114_112#_c_875_n 9.51679e-19 $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_194 N_GATE_c_191_n N_A_114_112#_c_875_n 0.0314033f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_195 N_GATE_M1012_g N_A_114_112#_c_876_n 0.00215547f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_196 N_GATE_c_190_n N_A_114_112#_c_876_n 3.44092e-19 $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_197 N_GATE_c_191_n N_A_114_112#_c_876_n 0.00675183f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_198 N_GATE_M1000_g N_A_114_112#_c_877_n 0.00362102f $X=0.895 $Y=2.54 $X2=0
+ $Y2=0
cc_199 N_GATE_M1012_g N_A_114_112#_c_877_n 0.00428574f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_200 N_GATE_c_190_n N_A_114_112#_c_877_n 0.00161237f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_201 N_GATE_c_191_n N_A_114_112#_c_877_n 0.0424879f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_202 N_GATE_M1000_g N_A_114_112#_c_883_n 0.00357062f $X=0.895 $Y=2.54 $X2=0
+ $Y2=0
cc_203 N_GATE_c_190_n N_A_114_112#_c_883_n 5.86442e-19 $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_204 N_GATE_c_191_n N_A_114_112#_c_883_n 0.0215229f $X=0.97 $Y=1.795 $X2=0
+ $Y2=0
cc_205 N_GATE_M1012_g N_A_114_112#_c_878_n 0.00476476f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_206 N_GATE_M1000_g N_A_114_112#_c_885_n 0.00992115f $X=0.895 $Y=2.54 $X2=0
+ $Y2=0
cc_207 N_GATE_M1012_g N_A_114_112#_c_880_n 0.00917045f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_208 N_GATE_M1012_g N_VGND_c_1003_n 0.00340632f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_209 N_GATE_M1012_g N_VGND_c_1007_n 0.00487769f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_210 N_A_318_74#_c_233_n N_A_288_48#_c_306_n 0.00194041f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_211 N_A_318_74#_c_235_n N_A_288_48#_c_306_n 0.005869f $X=1.73 $Y=0.965 $X2=0
+ $Y2=0
cc_212 N_A_318_74#_c_233_n N_A_288_48#_c_307_n 0.00954194f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_213 N_A_318_74#_c_235_n N_A_288_48#_c_307_n 0.00448444f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_214 N_A_318_74#_c_236_n N_A_288_48#_c_307_n 4.8832e-19 $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_215 N_A_318_74#_c_233_n N_A_288_48#_M1021_g 0.008824f $X=1.88 $Y=1.545 $X2=0
+ $Y2=0
cc_216 N_A_318_74#_c_236_n N_A_288_48#_M1021_g 0.034245f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_217 N_A_318_74#_c_237_n N_A_288_48#_M1021_g 4.73542e-19 $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_218 N_A_318_74#_c_238_n N_A_288_48#_M1021_g 0.00476526f $X=3.26 $Y=1.55 $X2=0
+ $Y2=0
cc_219 N_A_318_74#_M1011_g N_A_288_48#_c_326_n 0.0123594f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_220 N_A_318_74#_c_234_n N_A_288_48#_c_310_n 0.00115318f $X=2.625 $Y=1.63
+ $X2=0 $Y2=0
cc_221 N_A_318_74#_c_237_n N_A_288_48#_c_310_n 9.741e-19 $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_222 N_A_318_74#_c_238_n N_A_288_48#_c_310_n 0.0114346f $X=3.26 $Y=1.55 $X2=0
+ $Y2=0
cc_223 N_A_318_74#_c_233_n N_A_288_48#_c_311_n 0.00509279f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_224 N_A_318_74#_c_235_n N_A_288_48#_c_311_n 0.00163563f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_225 N_A_318_74#_c_236_n N_A_288_48#_c_311_n 0.0045155f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_226 N_A_318_74#_M1015_g N_A_288_48#_c_312_n 0.0224891f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_227 N_A_318_74#_M1011_g N_A_288_48#_M1002_g 0.0114165f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_228 N_A_318_74#_M1015_g N_A_288_48#_c_313_n 0.00115934f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_229 N_A_318_74#_c_235_n N_A_288_48#_c_313_n 0.00472036f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_230 N_A_318_74#_M1015_g N_A_288_48#_c_314_n 0.0127767f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_231 N_A_318_74#_M1015_g N_A_288_48#_c_316_n 0.00543799f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_232 N_A_318_74#_M1015_g N_A_288_48#_c_318_n 0.00118267f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_233 N_A_318_74#_M1015_g N_A_288_48#_c_323_n 4.23122e-19 $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_234 N_A_318_74#_c_233_n N_A_288_48#_c_323_n 0.0176486f $X=1.88 $Y=1.545 $X2=0
+ $Y2=0
cc_235 N_A_318_74#_c_234_n N_A_288_48#_c_323_n 0.0101474f $X=2.625 $Y=1.63 $X2=0
+ $Y2=0
cc_236 N_A_318_74#_c_235_n N_A_288_48#_c_323_n 0.00760911f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_237 N_A_318_74#_c_236_n N_A_288_48#_c_323_n 0.0216474f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_238 N_A_318_74#_c_237_n N_A_288_48#_c_323_n 0.00707468f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_239 N_A_318_74#_c_238_n N_A_288_48#_c_323_n 3.53521e-19 $X=3.26 $Y=1.55 $X2=0
+ $Y2=0
cc_240 N_A_318_74#_M1011_g N_A_709_54#_M1016_g 0.0060669f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_241 N_A_318_74#_M1015_g N_A_709_54#_M1016_g 0.0878255f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_242 N_A_318_74#_M1015_g N_A_566_74#_c_591_n 0.00783189f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_243 N_A_318_74#_M1011_g N_A_566_74#_c_592_n 0.018786f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_244 N_A_318_74#_c_237_n N_A_566_74#_c_592_n 0.0121454f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_245 N_A_318_74#_c_238_n N_A_566_74#_c_592_n 0.0129634f $X=3.26 $Y=1.55 $X2=0
+ $Y2=0
cc_246 N_A_318_74#_M1015_g N_A_566_74#_c_594_n 0.00886883f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_247 N_A_318_74#_c_237_n N_A_566_74#_c_594_n 5.28074e-19 $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_248 N_A_318_74#_c_238_n N_A_566_74#_c_594_n 0.00594074f $X=3.26 $Y=1.55 $X2=0
+ $Y2=0
cc_249 N_A_318_74#_M1011_g N_A_566_74#_c_599_n 0.00515202f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_250 N_A_318_74#_M1015_g N_A_566_74#_c_595_n 0.0114381f $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_251 N_A_318_74#_c_237_n N_A_566_74#_c_595_n 0.0129997f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_252 N_A_318_74#_c_238_n N_A_566_74#_c_595_n 0.01049f $X=3.26 $Y=1.55 $X2=0
+ $Y2=0
cc_253 N_A_318_74#_c_236_n N_VPWR_M1021_s 0.00384768f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_254 N_A_318_74#_M1011_g N_VPWR_c_788_n 0.00112709f $X=3 $Y=2.315 $X2=0 $Y2=0
cc_255 N_A_318_74#_c_233_n N_A_114_112#_c_875_n 0.0137774f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_256 N_A_318_74#_c_235_n N_A_114_112#_c_875_n 0.0048023f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_257 N_A_318_74#_c_233_n N_A_114_112#_c_877_n 0.00636232f $X=1.88 $Y=1.545
+ $X2=0 $Y2=0
cc_258 N_A_318_74#_c_236_n N_A_114_112#_c_877_n 0.0495323f $X=2.38 $Y=1.847
+ $X2=0 $Y2=0
cc_259 N_A_318_74#_M1021_d N_A_114_112#_c_882_n 0.00562767f $X=2.08 $Y=1.84
+ $X2=0 $Y2=0
cc_260 N_A_318_74#_M1011_g N_A_114_112#_c_882_n 0.00197714f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_261 N_A_318_74#_c_234_n N_A_114_112#_c_882_n 0.00713243f $X=2.625 $Y=1.63
+ $X2=0 $Y2=0
cc_262 N_A_318_74#_c_236_n N_A_114_112#_c_882_n 0.0368719f $X=2.38 $Y=1.847
+ $X2=0 $Y2=0
cc_263 N_A_318_74#_M1011_g N_A_114_112#_c_884_n 0.00174016f $X=3 $Y=2.315 $X2=0
+ $Y2=0
cc_264 N_A_318_74#_c_234_n N_A_114_112#_c_884_n 0.00118245f $X=2.625 $Y=1.63
+ $X2=0 $Y2=0
cc_265 N_A_318_74#_c_236_n N_A_114_112#_c_884_n 0.018296f $X=2.38 $Y=1.847 $X2=0
+ $Y2=0
cc_266 N_A_318_74#_c_237_n N_A_114_112#_c_884_n 0.0197455f $X=2.79 $Y=1.55 $X2=0
+ $Y2=0
cc_267 N_A_318_74#_c_238_n N_A_114_112#_c_884_n 0.00184413f $X=3.26 $Y=1.55
+ $X2=0 $Y2=0
cc_268 N_A_318_74#_M1003_d N_A_114_112#_c_880_n 0.00669008f $X=1.59 $Y=0.37
+ $X2=0 $Y2=0
cc_269 N_A_318_74#_c_235_n N_A_114_112#_c_880_n 0.0255794f $X=1.73 $Y=0.965
+ $X2=0 $Y2=0
cc_270 N_A_318_74#_M1015_g N_VGND_c_1001_n 9.29978e-19 $X=3.26 $Y=0.61 $X2=0
+ $Y2=0
cc_271 N_A_288_48#_c_319_n N_A_709_54#_M1010_d 0.00266942f $X=4.9 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_288_48#_c_314_n N_A_709_54#_M1016_g 0.00362604f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_273 N_A_288_48#_c_316_n N_A_709_54#_M1016_g 0.00875253f $X=3.495 $Y=0.88
+ $X2=0 $Y2=0
cc_274 N_A_288_48#_c_317_n N_A_709_54#_M1016_g 0.0112599f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_275 N_A_288_48#_c_318_n N_A_709_54#_M1016_g 0.0019606f $X=3.58 $Y=0.965 $X2=0
+ $Y2=0
cc_276 N_A_288_48#_c_367_p N_A_709_54#_M1016_g 0.00159596f $X=4.175 $Y=0.88
+ $X2=0 $Y2=0
cc_277 N_A_288_48#_M1002_g N_A_709_54#_M1018_g 0.0419503f $X=3.535 $Y=2.67 $X2=0
+ $Y2=0
cc_278 N_A_288_48#_c_319_n N_A_709_54#_c_468_n 0.0187364f $X=4.9 $Y=0.34 $X2=0
+ $Y2=0
cc_279 N_A_288_48#_c_321_n N_A_709_54#_c_468_n 0.0181109f $X=5.065 $Y=0.515
+ $X2=0 $Y2=0
cc_280 N_A_288_48#_c_322_n N_A_709_54#_c_469_n 0.0304982f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_281 N_A_288_48#_c_330_n N_A_709_54#_c_479_n 0.0172409f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_282 N_A_288_48#_M1020_s N_A_709_54#_c_480_n 0.00732293f $X=5.07 $Y=2.015
+ $X2=0 $Y2=0
cc_283 N_A_288_48#_c_330_n N_A_709_54#_c_480_n 0.0254481f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_284 N_A_288_48#_c_322_n N_A_709_54#_c_470_n 0.00560081f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_285 N_A_288_48#_c_330_n N_A_709_54#_c_470_n 0.0115929f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_286 N_A_288_48#_c_324_n N_A_709_54#_c_471_n 0.0181109f $X=5.065 $Y=1.13 $X2=0
+ $Y2=0
cc_287 N_A_288_48#_c_322_n N_A_709_54#_c_482_n 0.0215371f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_288 N_A_288_48#_c_330_n N_A_709_54#_c_482_n 0.0111525f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_289 N_A_288_48#_c_322_n N_A_709_54#_c_472_n 0.00357445f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_290 N_A_288_48#_M1002_g N_A_709_54#_c_484_n 0.00650081f $X=3.535 $Y=2.67
+ $X2=0 $Y2=0
cc_291 N_A_288_48#_c_314_n N_A_566_74#_M1017_d 0.00256812f $X=3.41 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_292 N_A_288_48#_c_317_n N_A_566_74#_c_589_n 0.00554178f $X=4.09 $Y=0.965
+ $X2=0 $Y2=0
cc_293 N_A_288_48#_c_367_p N_A_566_74#_c_589_n 0.0123114f $X=4.175 $Y=0.88 $X2=0
+ $Y2=0
cc_294 N_A_288_48#_c_319_n N_A_566_74#_c_589_n 0.0114613f $X=4.9 $Y=0.34 $X2=0
+ $Y2=0
cc_295 N_A_288_48#_c_320_n N_A_566_74#_c_589_n 0.00278978f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_296 N_A_288_48#_c_321_n N_A_566_74#_c_589_n 0.00362229f $X=5.065 $Y=0.515
+ $X2=0 $Y2=0
cc_297 N_A_288_48#_c_330_n N_A_566_74#_M1001_g 5.6792e-19 $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_298 N_A_288_48#_c_311_n N_A_566_74#_c_591_n 2.9126e-19 $X=2.415 $Y=1.07 $X2=0
+ $Y2=0
cc_299 N_A_288_48#_c_312_n N_A_566_74#_c_591_n 0.00183864f $X=2.755 $Y=0.995
+ $X2=0 $Y2=0
cc_300 N_A_288_48#_c_313_n N_A_566_74#_c_591_n 0.00430473f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_301 N_A_288_48#_c_318_n N_A_566_74#_c_591_n 0.0100841f $X=3.58 $Y=0.965 $X2=0
+ $Y2=0
cc_302 N_A_288_48#_c_323_n N_A_566_74#_c_591_n 0.00848118f $X=2.25 $Y=1.195
+ $X2=0 $Y2=0
cc_303 N_A_288_48#_M1002_g N_A_566_74#_c_592_n 0.00494982f $X=3.535 $Y=2.67
+ $X2=0 $Y2=0
cc_304 N_A_288_48#_c_317_n N_A_566_74#_c_593_n 0.0502793f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_305 N_A_288_48#_c_318_n N_A_566_74#_c_593_n 0.0147362f $X=3.58 $Y=0.965 $X2=0
+ $Y2=0
cc_306 N_A_288_48#_c_313_n N_A_566_74#_c_594_n 0.0112956f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_307 N_A_288_48#_c_314_n N_A_566_74#_c_594_n 0.0209617f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_308 N_A_288_48#_c_316_n N_A_566_74#_c_594_n 0.021236f $X=3.495 $Y=0.88 $X2=0
+ $Y2=0
cc_309 N_A_288_48#_c_318_n N_A_566_74#_c_594_n 0.00374694f $X=3.58 $Y=0.965
+ $X2=0 $Y2=0
cc_310 N_A_288_48#_c_326_n N_A_566_74#_c_599_n 0.00546485f $X=3.445 $Y=3.15
+ $X2=0 $Y2=0
cc_311 N_A_288_48#_c_311_n N_A_566_74#_c_595_n 8.48984e-19 $X=2.415 $Y=1.07
+ $X2=0 $Y2=0
cc_312 N_A_288_48#_c_323_n N_A_566_74#_c_595_n 0.00421113f $X=2.25 $Y=1.195
+ $X2=0 $Y2=0
cc_313 N_A_288_48#_c_317_n N_A_566_74#_c_596_n 0.00521109f $X=4.09 $Y=0.965
+ $X2=0 $Y2=0
cc_314 N_A_288_48#_c_322_n N_A_566_74#_c_596_n 0.00202724f $X=5.075 $Y=1.995
+ $X2=0 $Y2=0
cc_315 N_A_288_48#_c_319_n N_CLK_M1005_g 0.0047004f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_316 N_A_288_48#_c_321_n N_CLK_M1005_g 0.00681907f $X=5.065 $Y=0.515 $X2=0
+ $Y2=0
cc_317 N_A_288_48#_c_322_n N_CLK_M1005_g 0.0109213f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_318 N_A_288_48#_c_324_n N_CLK_M1005_g 0.00328501f $X=5.065 $Y=1.13 $X2=0
+ $Y2=0
cc_319 N_A_288_48#_c_330_n N_CLK_c_675_n 0.00717552f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_320 N_A_288_48#_c_322_n N_CLK_c_673_n 0.00679921f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_321 N_A_288_48#_c_330_n N_CLK_c_673_n 0.0049217f $X=5.215 $Y=2.16 $X2=0 $Y2=0
cc_322 N_A_288_48#_c_322_n N_CLK_c_674_n 0.0323289f $X=5.075 $Y=1.995 $X2=0
+ $Y2=0
cc_323 N_A_288_48#_c_330_n N_CLK_c_674_n 0.00328366f $X=5.215 $Y=2.16 $X2=0
+ $Y2=0
cc_324 N_A_288_48#_M1021_g N_VPWR_c_791_n 0.02379f $X=1.99 $Y=2.26 $X2=0 $Y2=0
cc_325 N_A_288_48#_M1002_g N_VPWR_c_792_n 0.00760658f $X=3.535 $Y=2.67 $X2=0
+ $Y2=0
cc_326 N_A_288_48#_c_327_n N_VPWR_c_800_n 0.0563267f $X=2.08 $Y=3.15 $X2=0 $Y2=0
cc_327 N_A_288_48#_c_326_n N_VPWR_c_788_n 0.0554168f $X=3.445 $Y=3.15 $X2=0
+ $Y2=0
cc_328 N_A_288_48#_c_327_n N_VPWR_c_788_n 0.00800048f $X=2.08 $Y=3.15 $X2=0
+ $Y2=0
cc_329 N_A_288_48#_c_313_n N_A_114_112#_M1017_s 0.0084363f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_330 N_A_288_48#_c_315_n N_A_114_112#_M1017_s 6.08643e-19 $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_331 N_A_288_48#_c_306_n N_A_114_112#_c_886_n 0.00137149f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_332 N_A_288_48#_c_307_n N_A_114_112#_c_875_n 0.00258488f $X=1.9 $Y=1.285
+ $X2=0 $Y2=0
cc_333 N_A_288_48#_c_308_n N_A_114_112#_c_875_n 0.00935869f $X=1.59 $Y=1.285
+ $X2=0 $Y2=0
cc_334 N_A_288_48#_M1021_g N_A_114_112#_c_875_n 6.00271e-19 $X=1.99 $Y=2.26
+ $X2=0 $Y2=0
cc_335 N_A_288_48#_M1021_g N_A_114_112#_c_877_n 0.00908083f $X=1.99 $Y=2.26
+ $X2=0 $Y2=0
cc_336 N_A_288_48#_M1021_g N_A_114_112#_c_882_n 0.0244403f $X=1.99 $Y=2.26 $X2=0
+ $Y2=0
cc_337 N_A_288_48#_c_326_n N_A_114_112#_c_882_n 0.0148523f $X=3.445 $Y=3.15
+ $X2=0 $Y2=0
cc_338 N_A_288_48#_M1021_g N_A_114_112#_c_884_n 0.00390377f $X=1.99 $Y=2.26
+ $X2=0 $Y2=0
cc_339 N_A_288_48#_c_308_n N_A_114_112#_c_878_n 0.00137149f $X=1.59 $Y=1.285
+ $X2=0 $Y2=0
cc_340 N_A_288_48#_M1021_g N_A_114_112#_c_885_n 0.0045398f $X=1.99 $Y=2.26 $X2=0
+ $Y2=0
cc_341 N_A_288_48#_c_306_n N_A_114_112#_c_879_n 0.00622457f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_342 N_A_288_48#_c_311_n N_A_114_112#_c_879_n 0.00597962f $X=2.415 $Y=1.07
+ $X2=0 $Y2=0
cc_343 N_A_288_48#_c_312_n N_A_114_112#_c_879_n 0.00235306f $X=2.755 $Y=0.995
+ $X2=0 $Y2=0
cc_344 N_A_288_48#_c_313_n N_A_114_112#_c_879_n 0.0276253f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_345 N_A_288_48#_c_315_n N_A_114_112#_c_879_n 0.00627272f $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_346 N_A_288_48#_c_323_n N_A_114_112#_c_879_n 0.0142183f $X=2.25 $Y=1.195
+ $X2=0 $Y2=0
cc_347 N_A_288_48#_c_306_n N_A_114_112#_c_880_n 0.0154871f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_348 N_A_288_48#_c_307_n N_A_114_112#_c_880_n 7.62449e-19 $X=1.9 $Y=1.285
+ $X2=0 $Y2=0
cc_349 N_A_288_48#_c_311_n N_A_114_112#_c_880_n 0.00222971f $X=2.415 $Y=1.07
+ $X2=0 $Y2=0
cc_350 N_A_288_48#_c_317_n N_VGND_M1016_d 0.00663756f $X=4.09 $Y=0.965 $X2=0
+ $Y2=0
cc_351 N_A_288_48#_c_367_p N_VGND_M1016_d 0.00488787f $X=4.175 $Y=0.88 $X2=0
+ $Y2=0
cc_352 N_A_288_48#_c_320_n N_VGND_M1016_d 5.22721e-19 $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_353 N_A_288_48#_c_314_n N_VGND_c_998_n 0.01267f $X=3.41 $Y=0.34 $X2=0 $Y2=0
cc_354 N_A_288_48#_c_317_n N_VGND_c_998_n 0.013847f $X=4.09 $Y=0.965 $X2=0 $Y2=0
cc_355 N_A_288_48#_c_367_p N_VGND_c_998_n 0.020664f $X=4.175 $Y=0.88 $X2=0 $Y2=0
cc_356 N_A_288_48#_c_320_n N_VGND_c_998_n 0.0142265f $X=4.26 $Y=0.34 $X2=0 $Y2=0
cc_357 N_A_288_48#_c_319_n N_VGND_c_999_n 0.0112234f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_288_48#_c_321_n N_VGND_c_999_n 0.0259244f $X=5.065 $Y=0.515 $X2=0
+ $Y2=0
cc_359 N_A_288_48#_c_306_n N_VGND_c_1001_n 0.00315544f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_360 N_A_288_48#_c_312_n N_VGND_c_1001_n 0.00278237f $X=2.755 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_288_48#_c_314_n N_VGND_c_1001_n 0.0565673f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_362 N_A_288_48#_c_315_n N_VGND_c_1001_n 0.0120637f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_363 N_A_288_48#_c_319_n N_VGND_c_1004_n 0.0644063f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_364 N_A_288_48#_c_320_n N_VGND_c_1004_n 0.0120637f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_A_288_48#_c_306_n N_VGND_c_1007_n 0.00400711f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_366 N_A_288_48#_c_312_n N_VGND_c_1007_n 0.00363424f $X=2.755 $Y=0.995 $X2=0
+ $Y2=0
cc_367 N_A_288_48#_c_314_n N_VGND_c_1007_n 0.0322089f $X=3.41 $Y=0.34 $X2=0
+ $Y2=0
cc_368 N_A_288_48#_c_315_n N_VGND_c_1007_n 0.00644906f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_369 N_A_288_48#_c_319_n N_VGND_c_1007_n 0.036247f $X=4.9 $Y=0.34 $X2=0 $Y2=0
cc_370 N_A_288_48#_c_320_n N_VGND_c_1007_n 0.00644906f $X=4.26 $Y=0.34 $X2=0
+ $Y2=0
cc_371 N_A_288_48#_c_306_n N_VGND_c_1008_n 0.00542971f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_372 N_A_288_48#_c_314_n A_667_80# 6.48644e-19 $X=3.41 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_373 N_A_288_48#_c_316_n A_667_80# 0.00370274f $X=3.495 $Y=0.88 $X2=-0.19
+ $Y2=-0.245
cc_374 N_A_709_54#_M1016_g N_A_566_74#_c_589_n 0.0149957f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_375 N_A_709_54#_c_469_n N_A_566_74#_c_589_n 0.00622278f $X=4.585 $Y=1.74
+ $X2=0 $Y2=0
cc_376 N_A_709_54#_M1016_g N_A_566_74#_M1001_g 0.00510488f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_377 N_A_709_54#_c_477_n N_A_566_74#_M1001_g 0.0247865f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_378 N_A_709_54#_c_469_n N_A_566_74#_M1001_g 0.0106639f $X=4.585 $Y=1.74 $X2=0
+ $Y2=0
cc_379 N_A_709_54#_c_479_n N_A_566_74#_M1001_g 0.0069653f $X=4.655 $Y=2.495
+ $X2=0 $Y2=0
cc_380 N_A_709_54#_c_482_n N_A_566_74#_M1001_g 0.00182639f $X=4.655 $Y=1.905
+ $X2=0 $Y2=0
cc_381 N_A_709_54#_c_483_n N_A_566_74#_M1001_g 0.00584538f $X=4.655 $Y=2.58
+ $X2=0 $Y2=0
cc_382 N_A_709_54#_c_484_n N_A_566_74#_M1001_g 0.0312088f $X=3.925 $Y=1.955
+ $X2=0 $Y2=0
cc_383 N_A_709_54#_M1016_g N_A_566_74#_c_591_n 0.00101991f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_384 N_A_709_54#_M1016_g N_A_566_74#_c_592_n 0.0081516f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_385 N_A_709_54#_M1018_g N_A_566_74#_c_592_n 0.00659071f $X=3.925 $Y=2.67
+ $X2=0 $Y2=0
cc_386 N_A_709_54#_c_477_n N_A_566_74#_c_592_n 0.0269421f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_387 N_A_709_54#_M1016_g N_A_566_74#_c_593_n 0.0175999f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_388 N_A_709_54#_c_477_n N_A_566_74#_c_593_n 0.0538499f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_389 N_A_709_54#_c_469_n N_A_566_74#_c_593_n 0.0251783f $X=4.585 $Y=1.74 $X2=0
+ $Y2=0
cc_390 N_A_709_54#_c_484_n N_A_566_74#_c_593_n 0.00190784f $X=3.925 $Y=1.955
+ $X2=0 $Y2=0
cc_391 N_A_709_54#_M1016_g N_A_566_74#_c_594_n 2.77632e-19 $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_392 N_A_709_54#_M1016_g N_A_566_74#_c_596_n 0.0140122f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_393 N_A_709_54#_c_477_n N_A_566_74#_c_596_n 0.00829634f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_394 N_A_709_54#_c_469_n N_A_566_74#_c_596_n 0.0107273f $X=4.585 $Y=1.74 $X2=0
+ $Y2=0
cc_395 N_A_709_54#_c_471_n N_A_566_74#_c_596_n 0.00269107f $X=4.555 $Y=1.05
+ $X2=0 $Y2=0
cc_396 N_A_709_54#_c_484_n N_A_566_74#_c_596_n 0.00132739f $X=3.925 $Y=1.955
+ $X2=0 $Y2=0
cc_397 N_A_709_54#_c_468_n N_CLK_M1005_g 0.00101752f $X=4.515 $Y=0.82 $X2=0
+ $Y2=0
cc_398 N_A_709_54#_c_472_n N_CLK_M1005_g 3.97134e-19 $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_399 N_A_709_54#_c_479_n N_CLK_c_675_n 0.00407535f $X=4.655 $Y=2.495 $X2=0
+ $Y2=0
cc_400 N_A_709_54#_c_480_n N_CLK_c_675_n 0.0203723f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_401 N_A_709_54#_c_470_n N_CLK_c_675_n 0.00679172f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_402 N_A_709_54#_c_482_n N_CLK_c_675_n 6.02829e-19 $X=4.655 $Y=1.905 $X2=0
+ $Y2=0
cc_403 N_A_709_54#_c_483_n N_CLK_c_675_n 0.00649549f $X=4.655 $Y=2.58 $X2=0
+ $Y2=0
cc_404 N_A_709_54#_c_466_n N_CLK_M1006_g 0.0365055f $X=6.115 $Y=1.22 $X2=0 $Y2=0
cc_405 N_A_709_54#_c_472_n N_CLK_M1006_g 0.00389357f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_406 N_A_709_54#_M1009_g N_CLK_c_676_n 0.0241262f $X=6.585 $Y=2.435 $X2=0
+ $Y2=0
cc_407 N_A_709_54#_c_470_n N_CLK_c_676_n 0.0145221f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_408 N_A_709_54#_c_472_n N_CLK_c_676_n 0.00356073f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_409 N_A_709_54#_c_473_n N_CLK_c_676_n 0.0117901f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_410 N_A_709_54#_M1009_g N_CLK_c_673_n 0.0025851f $X=6.585 $Y=2.435 $X2=0
+ $Y2=0
cc_411 N_A_709_54#_c_480_n N_CLK_c_673_n 0.00582245f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_412 N_A_709_54#_c_470_n N_CLK_c_673_n 0.00388892f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_413 N_A_709_54#_c_473_n N_CLK_c_673_n 0.0365055f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_414 N_A_709_54#_c_470_n N_CLK_c_678_n 0.00437194f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_415 N_A_709_54#_c_470_n N_CLK_c_674_n 0.0172833f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_416 N_A_709_54#_c_472_n N_CLK_c_674_n 0.0150518f $X=6.205 $Y=1.385 $X2=0
+ $Y2=0
cc_417 N_A_709_54#_M1009_g N_A_1238_94#_c_730_n 0.0266952f $X=6.585 $Y=2.435
+ $X2=0 $Y2=0
cc_418 N_A_709_54#_c_473_n N_A_1238_94#_c_731_n 0.00914688f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_419 N_A_709_54#_M1009_g N_A_1238_94#_c_733_n 0.0186357f $X=6.585 $Y=2.435
+ $X2=0 $Y2=0
cc_420 N_A_709_54#_c_470_n N_A_1238_94#_c_733_n 0.0184253f $X=5.915 $Y=2.495
+ $X2=0 $Y2=0
cc_421 N_A_709_54#_c_472_n N_A_1238_94#_c_733_n 0.0297948f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_422 N_A_709_54#_c_473_n N_A_1238_94#_c_733_n 0.0163379f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_423 N_A_709_54#_M1009_g N_A_1238_94#_c_740_n 0.0163676f $X=6.585 $Y=2.435
+ $X2=0 $Y2=0
cc_424 N_A_709_54#_c_470_n N_A_1238_94#_c_740_n 0.0243177f $X=5.915 $Y=2.495
+ $X2=0 $Y2=0
cc_425 N_A_709_54#_c_466_n N_A_1238_94#_c_734_n 0.00421972f $X=6.115 $Y=1.22
+ $X2=0 $Y2=0
cc_426 N_A_709_54#_c_472_n N_A_1238_94#_c_734_n 0.00580698f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_427 N_A_709_54#_c_473_n N_A_1238_94#_c_734_n 0.00749726f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_428 N_A_709_54#_M1009_g N_A_1238_94#_c_735_n 0.00239413f $X=6.585 $Y=2.435
+ $X2=0 $Y2=0
cc_429 N_A_709_54#_c_473_n N_A_1238_94#_c_735_n 0.00244172f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_430 N_A_709_54#_c_473_n N_A_1238_94#_c_736_n 0.00899294f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_431 N_A_709_54#_c_466_n N_A_1238_94#_c_737_n 0.0110552f $X=6.115 $Y=1.22
+ $X2=0 $Y2=0
cc_432 N_A_709_54#_c_472_n N_A_1238_94#_c_737_n 0.00874612f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_433 N_A_709_54#_c_473_n N_A_1238_94#_c_737_n 0.0075575f $X=6.205 $Y=1.385
+ $X2=0 $Y2=0
cc_434 N_A_709_54#_c_477_n N_VPWR_M1018_d 0.00282686f $X=4.49 $Y=1.93 $X2=0
+ $Y2=0
cc_435 N_A_709_54#_c_480_n N_VPWR_M1020_d 0.011393f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_436 N_A_709_54#_c_470_n N_VPWR_M1020_d 0.00954303f $X=5.915 $Y=2.495 $X2=0
+ $Y2=0
cc_437 N_A_709_54#_M1018_g N_VPWR_c_792_n 0.0139769f $X=3.925 $Y=2.67 $X2=0
+ $Y2=0
cc_438 N_A_709_54#_c_477_n N_VPWR_c_792_n 0.0161306f $X=4.49 $Y=1.93 $X2=0 $Y2=0
cc_439 N_A_709_54#_c_479_n N_VPWR_c_792_n 0.0176013f $X=4.655 $Y=2.495 $X2=0
+ $Y2=0
cc_440 N_A_709_54#_c_480_n N_VPWR_c_793_n 0.0320496f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_441 N_A_709_54#_M1009_g N_VPWR_c_794_n 0.00389286f $X=6.585 $Y=2.435 $X2=0
+ $Y2=0
cc_442 N_A_709_54#_c_480_n N_VPWR_c_795_n 0.0116792f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_443 N_A_709_54#_c_483_n N_VPWR_c_795_n 0.0109794f $X=4.655 $Y=2.58 $X2=0
+ $Y2=0
cc_444 N_A_709_54#_M1009_g N_VPWR_c_797_n 0.00578748f $X=6.585 $Y=2.435 $X2=0
+ $Y2=0
cc_445 N_A_709_54#_M1018_g N_VPWR_c_800_n 0.00519349f $X=3.925 $Y=2.67 $X2=0
+ $Y2=0
cc_446 N_A_709_54#_M1018_g N_VPWR_c_788_n 0.00524044f $X=3.925 $Y=2.67 $X2=0
+ $Y2=0
cc_447 N_A_709_54#_M1009_g N_VPWR_c_788_n 0.00615499f $X=6.585 $Y=2.435 $X2=0
+ $Y2=0
cc_448 N_A_709_54#_c_480_n N_VPWR_c_788_n 0.0233324f $X=5.83 $Y=2.58 $X2=0 $Y2=0
cc_449 N_A_709_54#_c_483_n N_VPWR_c_788_n 0.0114852f $X=4.655 $Y=2.58 $X2=0
+ $Y2=0
cc_450 N_A_709_54#_M1016_g N_VGND_c_998_n 0.0012897f $X=3.62 $Y=0.61 $X2=0 $Y2=0
cc_451 N_A_709_54#_c_466_n N_VGND_c_1000_n 0.00313422f $X=6.115 $Y=1.22 $X2=0
+ $Y2=0
cc_452 N_A_709_54#_M1016_g N_VGND_c_1001_n 0.00447942f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_453 N_A_709_54#_c_466_n N_VGND_c_1005_n 0.00485498f $X=6.115 $Y=1.22 $X2=0
+ $Y2=0
cc_454 N_A_709_54#_M1016_g N_VGND_c_1007_n 0.0041113f $X=3.62 $Y=0.61 $X2=0
+ $Y2=0
cc_455 N_A_709_54#_c_466_n N_VGND_c_1007_n 0.00514438f $X=6.115 $Y=1.22 $X2=0
+ $Y2=0
cc_456 N_A_566_74#_c_596_n N_CLK_M1005_g 0.00232575f $X=4.43 $Y=1.385 $X2=0
+ $Y2=0
cc_457 N_A_566_74#_M1001_g N_CLK_c_673_n 0.00232575f $X=4.43 $Y=2.32 $X2=0 $Y2=0
cc_458 N_A_566_74#_M1001_g N_VPWR_c_792_n 0.00362771f $X=4.43 $Y=2.32 $X2=0
+ $Y2=0
cc_459 N_A_566_74#_c_599_n N_VPWR_c_792_n 0.00451843f $X=3.225 $Y=2.59 $X2=0
+ $Y2=0
cc_460 N_A_566_74#_M1001_g N_VPWR_c_795_n 0.00597358f $X=4.43 $Y=2.32 $X2=0
+ $Y2=0
cc_461 N_A_566_74#_c_599_n N_VPWR_c_800_n 0.00726695f $X=3.225 $Y=2.59 $X2=0
+ $Y2=0
cc_462 N_A_566_74#_M1001_g N_VPWR_c_788_n 0.00624688f $X=4.43 $Y=2.32 $X2=0
+ $Y2=0
cc_463 N_A_566_74#_c_599_n N_VPWR_c_788_n 0.00904504f $X=3.225 $Y=2.59 $X2=0
+ $Y2=0
cc_464 N_A_566_74#_c_599_n N_A_114_112#_c_882_n 0.0115948f $X=3.225 $Y=2.59
+ $X2=0 $Y2=0
cc_465 N_A_566_74#_c_592_n N_A_114_112#_c_884_n 0.0140286f $X=3.225 $Y=2.05
+ $X2=0 $Y2=0
cc_466 N_A_566_74#_c_589_n N_VGND_c_998_n 0.00168945f $X=4.3 $Y=1.22 $X2=0 $Y2=0
cc_467 N_A_566_74#_c_589_n N_VGND_c_1004_n 0.00278237f $X=4.3 $Y=1.22 $X2=0
+ $Y2=0
cc_468 N_A_566_74#_c_589_n N_VGND_c_1007_n 0.00363424f $X=4.3 $Y=1.22 $X2=0
+ $Y2=0
cc_469 N_CLK_c_676_n N_A_1238_94#_c_733_n 0.00309887f $X=6.045 $Y=1.865 $X2=0
+ $Y2=0
cc_470 N_CLK_c_675_n N_A_1238_94#_c_740_n 9.33565e-19 $X=5.44 $Y=1.94 $X2=0
+ $Y2=0
cc_471 N_CLK_c_676_n N_A_1238_94#_c_740_n 0.00144331f $X=6.045 $Y=1.865 $X2=0
+ $Y2=0
cc_472 N_CLK_c_678_n N_A_1238_94#_c_740_n 0.0163674f $X=6.135 $Y=1.94 $X2=0
+ $Y2=0
cc_473 N_CLK_M1006_g N_A_1238_94#_c_737_n 0.00166928f $X=5.755 $Y=0.79 $X2=0
+ $Y2=0
cc_474 N_CLK_c_675_n N_VPWR_c_793_n 0.00419332f $X=5.44 $Y=1.94 $X2=0 $Y2=0
cc_475 N_CLK_c_678_n N_VPWR_c_793_n 0.00381374f $X=6.135 $Y=1.94 $X2=0 $Y2=0
cc_476 N_CLK_c_675_n N_VPWR_c_795_n 0.00466962f $X=5.44 $Y=1.94 $X2=0 $Y2=0
cc_477 N_CLK_c_678_n N_VPWR_c_797_n 0.00578748f $X=6.135 $Y=1.94 $X2=0 $Y2=0
cc_478 N_CLK_c_675_n N_VPWR_c_788_n 0.00615499f $X=5.44 $Y=1.94 $X2=0 $Y2=0
cc_479 N_CLK_c_678_n N_VPWR_c_788_n 0.00615499f $X=6.135 $Y=1.94 $X2=0 $Y2=0
cc_480 N_CLK_M1005_g N_VGND_c_999_n 0.00310756f $X=5.28 $Y=0.74 $X2=0 $Y2=0
cc_481 N_CLK_M1006_g N_VGND_c_999_n 0.00381172f $X=5.755 $Y=0.79 $X2=0 $Y2=0
cc_482 N_CLK_c_673_n N_VGND_c_999_n 0.00109716f $X=5.83 $Y=1.865 $X2=0 $Y2=0
cc_483 N_CLK_c_674_n N_VGND_c_999_n 0.0173191f $X=5.495 $Y=1.52 $X2=0 $Y2=0
cc_484 N_CLK_M1005_g N_VGND_c_1004_n 0.00430908f $X=5.28 $Y=0.74 $X2=0 $Y2=0
cc_485 N_CLK_M1006_g N_VGND_c_1005_n 0.00507111f $X=5.755 $Y=0.79 $X2=0 $Y2=0
cc_486 N_CLK_M1005_g N_VGND_c_1007_n 0.0082568f $X=5.28 $Y=0.74 $X2=0 $Y2=0
cc_487 N_CLK_M1006_g N_VGND_c_1007_n 0.00514438f $X=5.755 $Y=0.79 $X2=0 $Y2=0
cc_488 N_A_1238_94#_c_740_n N_VPWR_c_793_n 0.00200687f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_489 N_A_1238_94#_c_730_n N_VPWR_c_794_n 0.0231026f $X=7.09 $Y=1.725 $X2=0
+ $Y2=0
cc_490 N_A_1238_94#_c_740_n N_VPWR_c_794_n 0.0313712f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_491 N_A_1238_94#_c_735_n N_VPWR_c_794_n 0.0119681f $X=7.08 $Y=1.465 $X2=0
+ $Y2=0
cc_492 N_A_1238_94#_c_740_n N_VPWR_c_797_n 0.0101104f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_493 N_A_1238_94#_c_730_n N_VPWR_c_801_n 0.00475445f $X=7.09 $Y=1.725 $X2=0
+ $Y2=0
cc_494 N_A_1238_94#_c_730_n N_VPWR_c_788_n 0.00942664f $X=7.09 $Y=1.725 $X2=0
+ $Y2=0
cc_495 N_A_1238_94#_c_740_n N_VPWR_c_788_n 0.0112627f $X=6.36 $Y=2.16 $X2=0
+ $Y2=0
cc_496 N_A_1238_94#_c_732_n N_GCLK_c_976_n 0.00840121f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_497 N_A_1238_94#_c_732_n N_GCLK_c_977_n 0.00343235f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_498 N_A_1238_94#_c_730_n GCLK 0.0247403f $X=7.09 $Y=1.725 $X2=0 $Y2=0
cc_499 N_A_1238_94#_c_733_n GCLK 0.00131809f $X=6.36 $Y=1.89 $X2=0 $Y2=0
cc_500 N_A_1238_94#_c_735_n GCLK 6.98006e-19 $X=7.08 $Y=1.465 $X2=0 $Y2=0
cc_501 N_A_1238_94#_c_730_n N_GCLK_c_978_n 0.0014504f $X=7.09 $Y=1.725 $X2=0
+ $Y2=0
cc_502 N_A_1238_94#_c_732_n N_GCLK_c_978_n 0.0159294f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_503 N_A_1238_94#_c_735_n N_GCLK_c_978_n 0.0261275f $X=7.08 $Y=1.465 $X2=0
+ $Y2=0
cc_504 N_A_1238_94#_c_737_n N_VGND_c_999_n 0.0101545f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_505 N_A_1238_94#_c_731_n N_VGND_c_1000_n 0.00451355f $X=7.09 $Y=1.36 $X2=0
+ $Y2=0
cc_506 N_A_1238_94#_c_732_n N_VGND_c_1000_n 0.0196053f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_507 N_A_1238_94#_c_735_n N_VGND_c_1000_n 0.0213215f $X=7.08 $Y=1.465 $X2=0
+ $Y2=0
cc_508 N_A_1238_94#_c_737_n N_VGND_c_1000_n 0.0556027f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_509 N_A_1238_94#_c_737_n N_VGND_c_1005_n 0.0150236f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_510 N_A_1238_94#_c_732_n N_VGND_c_1006_n 0.00434272f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_511 N_A_1238_94#_c_732_n N_VGND_c_1007_n 0.00828811f $X=7.09 $Y=1.185 $X2=0
+ $Y2=0
cc_512 N_A_1238_94#_c_737_n N_VGND_c_1007_n 0.0164774f $X=6.33 $Y=0.615 $X2=0
+ $Y2=0
cc_513 N_VPWR_M1021_s N_A_114_112#_c_877_n 0.00746412f $X=1.535 $Y=1.84 $X2=0
+ $Y2=0
cc_514 N_VPWR_M1021_s N_A_114_112#_c_882_n 0.0101094f $X=1.535 $Y=1.84 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_800_n N_A_114_112#_c_882_n 0.00575553f $X=3.985 $Y=3.33 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_788_n N_A_114_112#_c_882_n 0.030078f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_M1021_s N_A_114_112#_c_883_n 0.00203332f $X=1.535 $Y=1.84 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_790_n N_A_114_112#_c_883_n 0.00544977f $X=0.28 $Y=2.295 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_791_n N_A_114_112#_c_883_n 0.0260097f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_788_n N_A_114_112#_c_883_n 0.00909591f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_790_n N_A_114_112#_c_885_n 0.0149884f $X=0.28 $Y=2.295 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_791_n N_A_114_112#_c_885_n 0.0215741f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_799_n N_A_114_112#_c_885_n 0.0142106f $X=1.515 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_788_n N_A_114_112#_c_885_n 0.0118429f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_794_n GCLK 0.0298396f $X=6.86 $Y=2.225 $X2=0 $Y2=0
cc_526 N_VPWR_c_801_n GCLK 0.0155281f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_c_788_n GCLK 0.0128528f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_528 N_A_114_112#_c_880_n N_VGND_M1012_d 0.00979382f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_529 N_A_114_112#_c_886_n N_VGND_c_997_n 0.0150351f $X=0.71 $Y=0.83 $X2=0
+ $Y2=0
cc_530 N_A_114_112#_c_874_n N_VGND_c_997_n 0.00756924f $X=0.885 $Y=0.625 $X2=0
+ $Y2=0
cc_531 N_A_114_112#_c_879_n N_VGND_c_1001_n 0.0107474f $X=2.29 $Y=0.565 $X2=0
+ $Y2=0
cc_532 N_A_114_112#_c_880_n N_VGND_c_1001_n 0.0151341f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_533 N_A_114_112#_c_874_n N_VGND_c_1003_n 0.0083132f $X=0.885 $Y=0.625 $X2=0
+ $Y2=0
cc_534 N_A_114_112#_c_880_n N_VGND_c_1003_n 0.00360867f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_535 N_A_114_112#_c_874_n N_VGND_c_1007_n 0.0109521f $X=0.885 $Y=0.625 $X2=0
+ $Y2=0
cc_536 N_A_114_112#_c_879_n N_VGND_c_1007_n 0.00908767f $X=2.29 $Y=0.565 $X2=0
+ $Y2=0
cc_537 N_A_114_112#_c_880_n N_VGND_c_1007_n 0.0289707f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_538 N_A_114_112#_c_880_n N_VGND_c_1008_n 0.0242087f $X=2.125 $Y=0.565 $X2=0
+ $Y2=0
cc_539 N_GCLK_c_976_n N_VGND_c_1000_n 0.0302381f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_540 N_GCLK_c_976_n N_VGND_c_1006_n 0.0152332f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_541 N_GCLK_c_976_n N_VGND_c_1007_n 0.0125524f $X=7.405 $Y=0.515 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VGND a_1292_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=1.98545e+12p pd=1.63e+07u as=4.514e+11p ps=4.18e+06u
M1001 a_119_143# GATE a_119_395# VPB pshort w=840000u l=180000u
+  ad=4.704e+11p pd=4.48e+06u as=2.016e+11p ps=2.16e+06u
M1002 VPWR CLK a_324_79# VPB pshort w=840000u l=180000u
+  ad=2.4738e+12p pd=1.955e+07u as=2.394e+11p ps=2.25e+06u
M1003 VGND a_1292_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_354_105# a_324_79# VPWR VPB pshort w=840000u l=180000u
+  ad=3.907e+11p pd=2.99e+06u as=0p ps=0u
M1005 a_634_74# a_354_105# a_119_143# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=0p ps=0u
M1006 a_792_48# a_634_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VGND a_792_48# a_744_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 a_788_455# a_324_79# a_634_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 GCLK a_1292_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=8.008e+11p pd=5.91e+06u as=0p ps=0u
M1010 VPWR a_1292_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1292_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1012 a_1292_368# a_792_48# a_1292_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 VGND CLK a_324_79# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1014 VPWR a_792_48# a_788_455# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 GCLK a_1292_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_1292_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_744_74# a_354_105# a_634_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.1025e+11p ps=1.9e+06u
M1018 GCLK a_1292_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_792_48# a_1292_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.208e+11p ps=3.17e+06u
M1020 a_1292_368# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_354_105# a_324_79# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_792_48# a_634_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1023 a_119_143# SCE VGND VNB nlowvt w=550000u l=150000u
+  ad=5.61e+11p pd=4.24e+06u as=0p ps=0u
M1024 a_634_74# a_324_79# a_119_143# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_119_395# SCE VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND GATE a_119_143# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 GCLK a_1292_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

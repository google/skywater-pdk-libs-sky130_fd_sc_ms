* File: sky130_fd_sc_ms__fahcon_1.pxi.spice
* Created: Wed Sep  2 12:09:53 2020
* 
x_PM_SKY130_FD_SC_MS__FAHCON_1%A N_A_M1014_g N_A_M1020_g A N_A_c_223_n
+ N_A_c_224_n PM_SKY130_FD_SC_MS__FAHCON_1%A
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_27_100# N_A_27_100#_M1014_s N_A_27_100#_M1013_d
+ N_A_27_100#_M1020_s N_A_27_100#_M1008_d N_A_27_100#_M1021_g
+ N_A_27_100#_c_261_n N_A_27_100#_M1002_g N_A_27_100#_c_262_n
+ N_A_27_100#_c_273_n N_A_27_100#_c_284_n N_A_27_100#_c_263_n
+ N_A_27_100#_c_264_n N_A_27_100#_c_265_n N_A_27_100#_c_266_n
+ N_A_27_100#_c_267_n N_A_27_100#_c_275_n N_A_27_100#_c_268_n
+ N_A_27_100#_c_361_p N_A_27_100#_c_302_p N_A_27_100#_c_269_n
+ N_A_27_100#_c_309_p N_A_27_100#_c_270_n N_A_27_100#_c_271_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_27_100#
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_336_263# N_A_336_263#_M1024_s
+ N_A_336_263#_M1027_s N_A_336_263#_M1000_g N_A_336_263#_M1003_g
+ N_A_336_263#_c_387_n N_A_336_263#_c_388_n N_A_336_263#_M1011_g
+ N_A_336_263#_M1030_g N_A_336_263#_c_391_n N_A_336_263#_c_392_n
+ N_A_336_263#_c_393_n N_A_336_263#_c_398_n N_A_336_263#_c_394_n
+ N_A_336_263#_c_399_n N_A_336_263#_c_395_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_336_263#
x_PM_SKY130_FD_SC_MS__FAHCON_1%B N_B_M1008_g N_B_M1013_g N_B_c_507_n N_B_c_508_n
+ N_B_M1019_g N_B_M1015_g N_B_c_510_n N_B_c_493_n N_B_c_494_n N_B_c_495_n
+ N_B_M1027_g N_B_c_497_n N_B_c_498_n N_B_M1024_g N_B_M1001_g N_B_M1031_g
+ N_B_c_501_n N_B_c_502_n N_B_c_515_n N_B_c_503_n B N_B_c_504_n N_B_c_505_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%B
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_374_120# N_A_374_120#_M1003_d
+ N_A_374_120#_M1011_d N_A_374_120#_M1012_g N_A_374_120#_M1018_g
+ N_A_374_120#_M1022_g N_A_374_120#_M1010_g N_A_374_120#_c_631_n
+ N_A_374_120#_c_657_n N_A_374_120#_c_672_n N_A_374_120#_c_650_n
+ N_A_374_120#_c_632_n N_A_374_120#_c_633_n N_A_374_120#_c_652_n
+ N_A_374_120#_c_634_n N_A_374_120#_c_654_n N_A_374_120#_c_635_n
+ N_A_374_120#_c_636_n N_A_374_120#_c_637_n N_A_374_120#_c_638_n
+ N_A_374_120#_c_639_n N_A_374_120#_c_640_n N_A_374_120#_c_641_n
+ N_A_374_120#_c_666_n N_A_374_120#_c_716_p N_A_374_120#_c_642_n
+ N_A_374_120#_c_721_p N_A_374_120#_c_643_n N_A_374_120#_c_644_n
+ N_A_374_120#_c_645_n N_A_374_120#_c_776_p N_A_374_120#_c_646_n
+ N_A_374_120#_c_647_n N_A_374_120#_c_762_p
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_374_120#
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_372_365# N_A_372_365#_M1030_d
+ N_A_372_365#_M1000_d N_A_372_365#_M1016_g N_A_372_365#_M1023_g
+ N_A_372_365#_M1026_g N_A_372_365#_c_887_n N_A_372_365#_M1007_g
+ N_A_372_365#_c_907_n N_A_372_365#_c_912_n N_A_372_365#_c_889_n
+ N_A_372_365#_c_909_n N_A_372_365#_c_890_n N_A_372_365#_c_891_n
+ N_A_372_365#_c_892_n N_A_372_365#_c_903_n N_A_372_365#_c_893_n
+ N_A_372_365#_c_894_n N_A_372_365#_c_895_n N_A_372_365#_c_896_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_372_365#
x_PM_SKY130_FD_SC_MS__FAHCON_1%CI N_CI_c_1058_n N_CI_M1005_g N_CI_M1025_g
+ N_CI_M1006_g N_CI_c_1054_n N_CI_M1004_g N_CI_c_1055_n CI N_CI_c_1057_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%CI
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_1609_368# N_A_1609_368#_M1004_d
+ N_A_1609_368#_M1006_d N_A_1609_368#_M1010_d N_A_1609_368#_M1017_g
+ N_A_1609_368#_M1028_g N_A_1609_368#_c_1125_n N_A_1609_368#_c_1126_n
+ N_A_1609_368#_c_1127_n N_A_1609_368#_c_1118_n N_A_1609_368#_c_1128_n
+ N_A_1609_368#_c_1129_n N_A_1609_368#_c_1119_n N_A_1609_368#_c_1176_n
+ N_A_1609_368#_c_1120_n N_A_1609_368#_c_1131_n N_A_1609_368#_c_1121_n
+ N_A_1609_368#_c_1122_n N_A_1609_368#_c_1123_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_1609_368#
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_1744_94# N_A_1744_94#_M1026_d
+ N_A_1744_94#_M1007_d N_A_1744_94#_M1029_g N_A_1744_94#_M1009_g
+ N_A_1744_94#_c_1233_n N_A_1744_94#_c_1234_n N_A_1744_94#_c_1235_n
+ N_A_1744_94#_c_1236_n N_A_1744_94#_c_1237_n N_A_1744_94#_c_1288_n
+ N_A_1744_94#_c_1289_n N_A_1744_94#_c_1243_n N_A_1744_94#_c_1238_n
+ N_A_1744_94#_c_1239_n N_A_1744_94#_c_1240_n N_A_1744_94#_c_1241_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_1744_94#
x_PM_SKY130_FD_SC_MS__FAHCON_1%VPWR N_VPWR_M1020_d N_VPWR_M1027_d N_VPWR_M1005_d
+ N_VPWR_M1028_d N_VPWR_c_1341_n N_VPWR_c_1342_n N_VPWR_c_1343_n N_VPWR_c_1344_n
+ N_VPWR_c_1345_n N_VPWR_c_1346_n VPWR N_VPWR_c_1347_n N_VPWR_c_1348_n
+ N_VPWR_c_1349_n N_VPWR_c_1340_n N_VPWR_c_1351_n N_VPWR_c_1352_n
+ N_VPWR_c_1353_n PM_SKY130_FD_SC_MS__FAHCON_1%VPWR
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_244_368# N_A_244_368#_M1002_d
+ N_A_244_368#_M1015_d N_A_244_368#_M1021_d N_A_244_368#_M1019_d
+ N_A_244_368#_c_1443_n N_A_244_368#_c_1438_n N_A_244_368#_c_1434_n
+ N_A_244_368#_c_1439_n N_A_244_368#_c_1440_n N_A_244_368#_c_1435_n
+ N_A_244_368#_c_1436_n N_A_244_368#_c_1437_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_244_368#
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_1026_389# N_A_1026_389#_M1031_d
+ N_A_1026_389#_M1001_d N_A_1026_389#_c_1505_n N_A_1026_389#_c_1502_n
+ N_A_1026_389#_c_1512_n N_A_1026_389#_c_1528_n N_A_1026_389#_c_1506_n
+ N_A_1026_389#_c_1503_n N_A_1026_389#_c_1504_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_1026_389#
x_PM_SKY130_FD_SC_MS__FAHCON_1%COUT_N N_COUT_N_M1016_d N_COUT_N_M1012_d
+ N_COUT_N_c_1560_n N_COUT_N_c_1557_n N_COUT_N_c_1558_n COUT_N
+ PM_SKY130_FD_SC_MS__FAHCON_1%COUT_N
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_1264_421# N_A_1264_421#_M1018_d
+ N_A_1264_421#_M1023_d N_A_1264_421#_c_1614_n N_A_1264_421#_c_1612_n
+ N_A_1264_421#_c_1613_n N_A_1264_421#_c_1628_n
+ PM_SKY130_FD_SC_MS__FAHCON_1%A_1264_421#
x_PM_SKY130_FD_SC_MS__FAHCON_1%A_1719_368# N_A_1719_368#_M1022_d
+ N_A_1719_368#_M1007_s N_A_1719_368#_M1028_s N_A_1719_368#_c_1660_n
+ N_A_1719_368#_c_1668_n N_A_1719_368#_c_1682_n N_A_1719_368#_c_1671_n
+ N_A_1719_368#_c_1661_n N_A_1719_368#_c_1659_n N_A_1719_368#_c_1663_n
+ N_A_1719_368#_c_1664_n PM_SKY130_FD_SC_MS__FAHCON_1%A_1719_368#
x_PM_SKY130_FD_SC_MS__FAHCON_1%SUM N_SUM_M1009_d N_SUM_M1029_d N_SUM_c_1724_n
+ N_SUM_c_1725_n SUM SUM SUM SUM N_SUM_c_1726_n PM_SKY130_FD_SC_MS__FAHCON_1%SUM
x_PM_SKY130_FD_SC_MS__FAHCON_1%VGND N_VGND_M1014_d N_VGND_M1024_d N_VGND_M1025_d
+ N_VGND_M1017_d N_VGND_c_1752_n N_VGND_c_1753_n N_VGND_c_1754_n N_VGND_c_1755_n
+ N_VGND_c_1756_n N_VGND_c_1757_n VGND N_VGND_c_1758_n N_VGND_c_1759_n
+ N_VGND_c_1760_n N_VGND_c_1761_n N_VGND_c_1762_n N_VGND_c_1763_n
+ N_VGND_c_1764_n N_VGND_c_1765_n PM_SKY130_FD_SC_MS__FAHCON_1%VGND
cc_1 VNB A 0.00276866f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_2 VNB N_A_c_223_n 0.0257856f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_3 VNB N_A_c_224_n 0.0229732f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_4 VNB N_A_27_100#_c_261_n 0.0183307f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_5 VNB N_A_27_100#_c_262_n 0.0223604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_100#_c_263_n 0.00202176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_100#_c_264_n 0.00407438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_100#_c_265_n 0.0171513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_100#_c_266_n 0.00429524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_100#_c_267_n 0.00851536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_100#_c_268_n 0.0221956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_100#_c_269_n 2.23982e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_100#_c_270_n 0.00329264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_100#_c_271_n 0.0367782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_336_263#_M1000_g 0.0104452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_336_263#_M1003_g 0.024584f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.68
cc_17 VNB N_A_336_263#_c_387_n 0.11362f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.565
cc_18 VNB N_A_336_263#_c_388_n 0.0126136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_336_263#_M1011_g 0.00632706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_336_263#_M1030_g 0.0105446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_336_263#_c_391_n 0.00971789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_336_263#_c_392_n 0.0107696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_336_263#_c_393_n 0.0406512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_336_263#_c_394_n 0.00431118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_336_263#_c_395_n 0.00832616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_M1008_g 0.00174903f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.68
cc_27 VNB N_B_M1013_g 0.0179575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_M1015_g 0.0302102f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_29 VNB N_B_c_493_n 0.00481223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_494_n 0.0211049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_c_495_n 0.0113666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_M1027_g 0.00543189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_497_n 0.0120607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_498_n 0.0194078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_M1001_g 0.00618698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_M1031_g 0.0288972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_501_n 0.0113865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_c_502_n 0.00401217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_c_503_n 0.00820428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_c_504_n 0.00641946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_B_c_505_n 0.046151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_374_120#_M1022_g 0.0222867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_374_120#_M1010_g 0.00427439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_374_120#_c_631_n 0.0212883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_374_120#_c_632_n 0.00594268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_374_120#_c_633_n 7.31919e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_374_120#_c_634_n 0.0468432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_374_120#_c_635_n 0.00506327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_374_120#_c_636_n 0.00157626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_374_120#_c_637_n 0.0083239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_374_120#_c_638_n 0.00265861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_374_120#_c_639_n 0.0396421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_374_120#_c_640_n 0.00173497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_374_120#_c_641_n 0.00638116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_374_120#_c_642_n 0.00248282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_374_120#_c_643_n 6.63101e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_374_120#_c_644_n 0.00352111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_374_120#_c_645_n 0.0015849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_374_120#_c_646_n 0.0259068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_374_120#_c_647_n 0.00261967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_372_365#_M1016_g 0.0523454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_372_365#_M1026_g 0.0253605f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_63 VNB N_A_372_365#_c_887_n 0.0196747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_372_365#_M1007_g 0.00175936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_372_365#_c_889_n 0.0156978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_372_365#_c_890_n 0.0207932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_372_365#_c_891_n 0.00189243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_372_365#_c_892_n 8.9583e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_372_365#_c_893_n 0.0169664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_372_365#_c_894_n 0.0388652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_372_365#_c_895_n 0.0015507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_372_365#_c_896_n 0.00794384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_CI_M1025_g 0.0258645f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_74 VNB N_CI_c_1054_n 0.0191394f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.68
cc_75 VNB N_CI_c_1055_n 0.00480507f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_76 VNB CI 0.00375348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_CI_c_1057_n 0.0639096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1609_368#_M1017_g 0.0227718f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_79 VNB N_A_1609_368#_M1028_g 0.00399992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1609_368#_c_1118_n 0.00356954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1609_368#_c_1119_n 0.00649616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1609_368#_c_1120_n 0.00271406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1609_368#_c_1121_n 0.00160893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1609_368#_c_1122_n 0.00443794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1609_368#_c_1123_n 0.0546693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1744_94#_M1029_g 0.00181061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1744_94#_M1009_g 0.0291228f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_88 VNB N_A_1744_94#_c_1233_n 0.0111586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1744_94#_c_1234_n 0.00132064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1744_94#_c_1235_n 0.0249277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1744_94#_c_1236_n 0.00646303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1744_94#_c_1237_n 6.28752e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1744_94#_c_1238_n 0.00268638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1744_94#_c_1239_n 0.00233037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1744_94#_c_1240_n 0.0364143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1744_94#_c_1241_n 0.00144783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VPWR_c_1340_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_244_368#_c_1434_n 0.00232036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_244_368#_c_1435_n 0.0133774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_244_368#_c_1436_n 0.00124806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_244_368#_c_1437_n 0.00651639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1026_389#_c_1502_n 0.00127577f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.68
cc_103 VNB N_A_1026_389#_c_1503_n 0.00579039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1026_389#_c_1504_n 0.00279567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_COUT_N_c_1557_n 0.00214343f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_106 VNB N_COUT_N_c_1558_n 0.00787408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB COUT_N 0.008237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1264_421#_c_1612_n 0.00289742f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.565
cc_109 VNB N_A_1264_421#_c_1613_n 0.00744846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1719_368#_c_1659_n 0.0071406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_SUM_c_1724_n 0.0271795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_SUM_c_1725_n 0.0100432f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_113 VNB N_SUM_c_1726_n 0.0246985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1752_n 0.0125244f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.68
cc_115 VNB N_VGND_c_1753_n 0.0085717f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_116 VNB N_VGND_c_1754_n 0.00927156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1755_n 0.0178043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1756_n 0.00324082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1757_n 0.00299623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1758_n 0.0981815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1759_n 0.0712816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1760_n 0.0614777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1761_n 0.0194686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1762_n 0.62607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1763_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1764_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1765_n 0.0164819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VPB N_A_M1020_g 0.0276694f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_129 VPB A 0.00446856f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_130 VPB N_A_c_223_n 0.00553287f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_131 VPB N_A_27_100#_M1021_g 0.0248478f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.565
cc_132 VPB N_A_27_100#_c_273_n 0.0376001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_27_100#_c_263_n 0.00237823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_27_100#_c_275_n 0.00828968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_27_100#_c_268_n 0.0129758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_27_100#_c_269_n 0.00117848f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_27_100#_c_271_n 0.011349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_336_263#_M1000_g 0.023596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_336_263#_M1011_g 0.0204953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_336_263#_c_398_n 0.0100177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_336_263#_c_399_n 0.00254863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_336_263#_c_395_n 0.00252733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_B_M1008_g 0.0403356f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.68
cc_144 VPB N_B_c_507_n 0.0606695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_B_c_508_n 0.0141117f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_146 VPB N_B_M1019_g 0.0293506f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.68
cc_147 VPB N_B_c_510_n 0.0342594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_B_c_493_n 0.0764837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_B_M1027_g 0.0229719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_B_M1001_g 0.0305356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_B_c_502_n 0.00628871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_B_c_515_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_374_120#_M1012_g 0.0330029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_374_120#_M1010_g 0.0245836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_374_120#_c_650_n 0.00608987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_374_120#_c_632_n 7.41961e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_374_120#_c_652_n 0.00358359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_374_120#_c_634_n 0.0180647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_374_120#_c_654_n 0.00410022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_374_120#_c_636_n 0.00561954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_374_120#_c_646_n 0.0178807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_372_365#_M1023_g 0.0350185f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.35
cc_163 VPB N_A_372_365#_M1007_g 0.0232932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_372_365#_c_889_n 0.0145411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_372_365#_c_890_n 0.0131464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_372_365#_c_891_n 4.67518e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_372_365#_c_892_n 0.00260542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_372_365#_c_903_n 0.00253628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_372_365#_c_893_n 0.0274729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_372_365#_c_895_n 0.00582875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_372_365#_c_896_n 0.00405122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_CI_c_1058_n 0.0292191f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.87
cc_173 VPB N_CI_M1006_g 0.0245337f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_174 VPB N_CI_c_1055_n 0.00569459f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_175 VPB N_CI_c_1057_n 0.00276949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_1609_368#_M1028_g 0.0345713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1609_368#_c_1125_n 0.00535398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_1609_368#_c_1126_n 0.0032918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_1609_368#_c_1127_n 0.00860927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1609_368#_c_1128_n 0.0176956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1609_368#_c_1129_n 0.00335711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1609_368#_c_1119_n 0.00350838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1609_368#_c_1131_n 0.00910417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1609_368#_c_1121_n 0.0031916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1744_94#_M1029_g 0.0295659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1744_94#_c_1243_n 0.00215868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1744_94#_c_1238_n 0.00142549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1341_n 0.0109142f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_189 VPB N_VPWR_c_1342_n 0.0141473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1343_n 0.00796272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1344_n 0.00867824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1345_n 0.0744604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1346_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1347_n 0.0854831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1348_n 0.0710953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1349_n 0.0190763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1340_n 0.138899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1351_n 0.0261991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1352_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1353_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_244_368#_c_1438_n 0.00543079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_244_368#_c_1439_n 0.0281187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_244_368#_c_1440_n 0.0039844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_244_368#_c_1435_n 0.0110866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_244_368#_c_1436_n 0.00256092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1026_389#_c_1505_n 0.00286305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1026_389#_c_1506_n 0.00144881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1026_389#_c_1503_n 0.00584417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_COUT_N_c_1560_n 0.00595983f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_210 VPB N_COUT_N_c_1557_n 0.00357929f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.35
cc_211 VPB N_A_1264_421#_c_1614_n 0.0171205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1264_421#_c_1613_n 0.00456651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1719_368#_c_1660_n 0.0344337f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_214 VPB N_A_1719_368#_c_1661_n 7.33272e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1719_368#_c_1659_n 0.00111753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1719_368#_c_1663_n 0.0114364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1719_368#_c_1664_n 0.00646305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB SUM 0.0126749f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.68
cc_219 VPB SUM 0.0415472f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_SUM_c_1726_n 0.00770625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 N_A_M1020_g N_A_27_100#_M1021_g 0.0185506f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_222 A N_A_27_100#_M1021_g 0.00105919f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A_c_224_n N_A_27_100#_c_261_n 0.00599956f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_224 N_A_c_224_n N_A_27_100#_c_262_n 4.63962e-19 $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_225 N_A_M1020_g N_A_27_100#_c_273_n 0.0101365f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_226 A N_A_27_100#_c_284_n 0.0269361f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A_c_223_n N_A_27_100#_c_284_n 0.00316435f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A_c_224_n N_A_27_100#_c_284_n 0.0145611f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_229 A N_A_27_100#_c_263_n 0.0255848f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_230 N_A_c_223_n N_A_27_100#_c_263_n 3.07635e-19 $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_231 N_A_c_224_n N_A_27_100#_c_263_n 0.00320785f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_232 N_A_c_224_n N_A_27_100#_c_264_n 0.00329314f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_233 N_A_c_224_n N_A_27_100#_c_266_n 3.07421e-19 $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_234 N_A_M1020_g N_A_27_100#_c_275_n 0.00268437f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_235 A N_A_27_100#_c_275_n 0.00362344f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_236 N_A_c_223_n N_A_27_100#_c_275_n 0.00142717f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_237 N_A_M1020_g N_A_27_100#_c_268_n 0.00473806f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_238 A N_A_27_100#_c_268_n 0.0330896f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_239 N_A_c_223_n N_A_27_100#_c_268_n 0.00785935f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A_c_224_n N_A_27_100#_c_268_n 0.00411368f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_241 A N_A_27_100#_c_271_n 0.00225172f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A_c_223_n N_A_27_100#_c_271_n 0.0211859f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_243 N_A_M1020_g N_VPWR_c_1341_n 0.00520277f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_244 A N_VPWR_c_1341_n 0.0115555f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A_c_223_n N_VPWR_c_1341_n 2.11748e-19 $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A_M1020_g N_VPWR_c_1340_n 0.009906f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_M1020_g N_VPWR_c_1351_n 0.005209f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_M1020_g N_A_244_368#_c_1443_n 5.98685e-19 $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_249 A N_A_244_368#_c_1436_n 0.00351446f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_250 N_A_c_224_n N_VGND_c_1752_n 0.00691015f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_251 N_A_c_224_n N_VGND_c_1755_n 0.00405273f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_252 N_A_c_224_n N_VGND_c_1757_n 0.0043102f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_253 N_A_c_224_n N_VGND_c_1762_n 0.00424518f $X=0.54 $Y=1.35 $X2=0 $Y2=0
cc_254 N_A_27_100#_M1021_g N_A_336_263#_M1000_g 0.0111671f $X=1.13 $Y=2.34 $X2=0
+ $Y2=0
cc_255 N_A_27_100#_c_302_p N_A_336_263#_M1000_g 5.43423e-19 $X=2.565 $Y=1.97
+ $X2=0 $Y2=0
cc_256 N_A_27_100#_c_271_n N_A_336_263#_M1000_g 0.00957794f $X=1.365 $Y=1.515
+ $X2=0 $Y2=0
cc_257 N_A_27_100#_c_261_n N_A_336_263#_M1003_g 0.0093625f $X=1.365 $Y=1.35
+ $X2=0 $Y2=0
cc_258 N_A_27_100#_c_264_n N_A_336_263#_M1003_g 0.00134468f $X=1.16 $Y=0.98
+ $X2=0 $Y2=0
cc_259 N_A_27_100#_c_265_n N_A_336_263#_M1003_g 0.0138038f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_260 N_A_27_100#_c_270_n N_A_336_263#_M1003_g 0.00294732f $X=2.61 $Y=0.725
+ $X2=0 $Y2=0
cc_261 N_A_27_100#_c_265_n N_A_336_263#_c_387_n 0.0228054f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_262 N_A_27_100#_c_309_p N_A_336_263#_c_387_n 8.5248e-19 $X=2.61 $Y=0.81 $X2=0
+ $Y2=0
cc_263 N_A_27_100#_c_270_n N_A_336_263#_c_387_n 0.00621886f $X=2.61 $Y=0.725
+ $X2=0 $Y2=0
cc_264 N_A_27_100#_c_265_n N_A_336_263#_c_388_n 0.00261705f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_265 N_A_27_100#_c_302_p N_A_336_263#_M1011_g 0.00490249f $X=2.565 $Y=1.97
+ $X2=0 $Y2=0
cc_266 N_A_27_100#_c_269_n N_A_336_263#_M1011_g 0.00655126f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_267 N_A_27_100#_c_269_n N_A_336_263#_M1030_g 0.00557596f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_268 N_A_27_100#_c_309_p N_A_336_263#_M1030_g 0.00216292f $X=2.61 $Y=0.81
+ $X2=0 $Y2=0
cc_269 N_A_27_100#_c_261_n N_A_336_263#_c_391_n 0.00957794f $X=1.365 $Y=1.35
+ $X2=0 $Y2=0
cc_270 N_A_27_100#_c_269_n N_A_336_263#_c_392_n 0.00498649f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_271 N_A_27_100#_c_265_n N_A_336_263#_c_394_n 0.0148909f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_272 N_A_27_100#_c_270_n N_A_336_263#_c_394_n 0.00970476f $X=2.61 $Y=0.725
+ $X2=0 $Y2=0
cc_273 N_A_27_100#_c_302_p N_B_M1008_g 0.00623718f $X=2.565 $Y=1.97 $X2=0 $Y2=0
cc_274 N_A_27_100#_c_269_n N_B_M1008_g 0.0021474f $X=2.587 $Y=1.805 $X2=0 $Y2=0
cc_275 N_A_27_100#_c_265_n N_B_M1013_g 0.00311259f $X=2.445 $Y=0.34 $X2=0 $Y2=0
cc_276 N_A_27_100#_c_269_n N_B_M1013_g 0.00750782f $X=2.587 $Y=1.805 $X2=0 $Y2=0
cc_277 N_A_27_100#_c_309_p N_B_M1013_g 0.00145757f $X=2.61 $Y=0.81 $X2=0 $Y2=0
cc_278 N_A_27_100#_c_270_n N_B_M1013_g 0.00351516f $X=2.61 $Y=0.725 $X2=0 $Y2=0
cc_279 N_A_27_100#_c_302_p N_B_c_501_n 6.34148e-19 $X=2.565 $Y=1.97 $X2=0 $Y2=0
cc_280 N_A_27_100#_c_269_n N_B_c_501_n 0.0041365f $X=2.587 $Y=1.805 $X2=0 $Y2=0
cc_281 N_A_27_100#_c_302_p N_A_374_120#_c_657_n 0.00475392f $X=2.565 $Y=1.97
+ $X2=0 $Y2=0
cc_282 N_A_27_100#_M1008_d N_A_374_120#_c_650_n 0.00166235f $X=2.43 $Y=1.825
+ $X2=0 $Y2=0
cc_283 N_A_27_100#_c_269_n N_A_374_120#_c_632_n 0.0148202f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_284 N_A_27_100#_c_302_p N_A_374_120#_c_654_n 0.00125813f $X=2.565 $Y=1.97
+ $X2=0 $Y2=0
cc_285 N_A_27_100#_c_269_n N_A_374_120#_c_654_n 0.00735732f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_286 N_A_27_100#_c_309_p N_A_374_120#_c_635_n 0.0166677f $X=2.61 $Y=0.81 $X2=0
+ $Y2=0
cc_287 N_A_27_100#_c_265_n N_A_374_120#_c_641_n 0.00443994f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_288 N_A_27_100#_c_269_n N_A_374_120#_c_641_n 0.0220099f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_289 N_A_27_100#_c_309_p N_A_374_120#_c_641_n 0.0129662f $X=2.61 $Y=0.81 $X2=0
+ $Y2=0
cc_290 N_A_27_100#_c_265_n N_A_374_120#_c_666_n 0.00236531f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_291 N_A_27_100#_c_269_n N_A_374_120#_c_666_n 0.00132788f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_292 N_A_27_100#_c_309_p N_A_374_120#_c_666_n 0.00132788f $X=2.61 $Y=0.81
+ $X2=0 $Y2=0
cc_293 N_A_27_100#_c_265_n N_A_374_120#_c_647_n 0.026474f $X=2.445 $Y=0.34 $X2=0
+ $Y2=0
cc_294 N_A_27_100#_c_270_n N_A_374_120#_c_647_n 0.0166677f $X=2.61 $Y=0.725
+ $X2=0 $Y2=0
cc_295 N_A_27_100#_M1008_d N_A_372_365#_c_907_n 0.00322007f $X=2.43 $Y=1.825
+ $X2=0 $Y2=0
cc_296 N_A_27_100#_c_302_p N_A_372_365#_c_907_n 0.0202871f $X=2.565 $Y=1.97
+ $X2=0 $Y2=0
cc_297 N_A_27_100#_c_269_n N_A_372_365#_c_909_n 0.00154391f $X=2.587 $Y=1.805
+ $X2=0 $Y2=0
cc_298 N_A_27_100#_c_309_p N_A_372_365#_c_896_n 0.0810636f $X=2.61 $Y=0.81 $X2=0
+ $Y2=0
cc_299 N_A_27_100#_M1021_g N_VPWR_c_1341_n 0.00663526f $X=1.13 $Y=2.34 $X2=0
+ $Y2=0
cc_300 N_A_27_100#_c_263_n N_VPWR_c_1341_n 4.57879e-19 $X=1.08 $Y=1.515 $X2=0
+ $Y2=0
cc_301 N_A_27_100#_c_275_n N_VPWR_c_1341_n 0.0405544f $X=0.32 $Y=2.115 $X2=0
+ $Y2=0
cc_302 N_A_27_100#_c_271_n N_VPWR_c_1341_n 0.0024915f $X=1.365 $Y=1.515 $X2=0
+ $Y2=0
cc_303 N_A_27_100#_M1021_g N_VPWR_c_1347_n 0.00508554f $X=1.13 $Y=2.34 $X2=0
+ $Y2=0
cc_304 N_A_27_100#_M1021_g N_VPWR_c_1340_n 0.00508379f $X=1.13 $Y=2.34 $X2=0
+ $Y2=0
cc_305 N_A_27_100#_c_273_n N_VPWR_c_1340_n 0.0145596f $X=0.32 $Y=2.815 $X2=0
+ $Y2=0
cc_306 N_A_27_100#_c_273_n N_VPWR_c_1351_n 0.0176724f $X=0.32 $Y=2.815 $X2=0
+ $Y2=0
cc_307 N_A_27_100#_M1021_g N_A_244_368#_c_1443_n 0.00427396f $X=1.13 $Y=2.34
+ $X2=0 $Y2=0
cc_308 N_A_27_100#_c_271_n N_A_244_368#_c_1443_n 0.00463503f $X=1.365 $Y=1.515
+ $X2=0 $Y2=0
cc_309 N_A_27_100#_M1021_g N_A_244_368#_c_1438_n 0.0121357f $X=1.13 $Y=2.34
+ $X2=0 $Y2=0
cc_310 N_A_27_100#_c_261_n N_A_244_368#_c_1434_n 0.00906427f $X=1.365 $Y=1.35
+ $X2=0 $Y2=0
cc_311 N_A_27_100#_c_263_n N_A_244_368#_c_1434_n 0.00823046f $X=1.08 $Y=1.515
+ $X2=0 $Y2=0
cc_312 N_A_27_100#_c_264_n N_A_244_368#_c_1434_n 0.0145966f $X=1.16 $Y=0.98
+ $X2=0 $Y2=0
cc_313 N_A_27_100#_c_265_n N_A_244_368#_c_1434_n 0.0256318f $X=2.445 $Y=0.34
+ $X2=0 $Y2=0
cc_314 N_A_27_100#_c_361_p N_A_244_368#_c_1434_n 0.00193071f $X=0.975 $Y=0.98
+ $X2=0 $Y2=0
cc_315 N_A_27_100#_M1021_g N_A_244_368#_c_1440_n 0.00286862f $X=1.13 $Y=2.34
+ $X2=0 $Y2=0
cc_316 N_A_27_100#_M1021_g N_A_244_368#_c_1436_n 0.00283126f $X=1.13 $Y=2.34
+ $X2=0 $Y2=0
cc_317 N_A_27_100#_c_271_n N_A_244_368#_c_1436_n 0.00718613f $X=1.365 $Y=1.515
+ $X2=0 $Y2=0
cc_318 N_A_27_100#_c_261_n N_A_244_368#_c_1437_n 0.00405483f $X=1.365 $Y=1.35
+ $X2=0 $Y2=0
cc_319 N_A_27_100#_c_263_n N_A_244_368#_c_1437_n 0.0255954f $X=1.08 $Y=1.515
+ $X2=0 $Y2=0
cc_320 N_A_27_100#_c_271_n N_A_244_368#_c_1437_n 0.00454619f $X=1.365 $Y=1.515
+ $X2=0 $Y2=0
cc_321 N_A_27_100#_c_284_n N_VGND_M1014_d 0.0147137f $X=0.975 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_322 N_A_27_100#_c_263_n N_VGND_M1014_d 0.00140773f $X=1.08 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_323 N_A_27_100#_c_264_n N_VGND_M1014_d 0.00790169f $X=1.16 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_324 N_A_27_100#_c_361_p N_VGND_M1014_d 0.00812545f $X=0.975 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_27_100#_c_264_n N_VGND_c_1752_n 0.00244281f $X=1.16 $Y=0.98 $X2=0
+ $Y2=0
cc_326 N_A_27_100#_c_266_n N_VGND_c_1752_n 0.00852809f $X=1.245 $Y=0.34 $X2=0
+ $Y2=0
cc_327 N_A_27_100#_c_262_n N_VGND_c_1755_n 0.00811546f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_328 N_A_27_100#_c_262_n N_VGND_c_1757_n 0.0126814f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_329 N_A_27_100#_c_284_n N_VGND_c_1757_n 0.023226f $X=0.975 $Y=1.08 $X2=0
+ $Y2=0
cc_330 N_A_27_100#_c_264_n N_VGND_c_1757_n 0.0257037f $X=1.16 $Y=0.98 $X2=0
+ $Y2=0
cc_331 N_A_27_100#_c_265_n N_VGND_c_1758_n 0.0866992f $X=2.445 $Y=0.34 $X2=0
+ $Y2=0
cc_332 N_A_27_100#_c_266_n N_VGND_c_1758_n 0.0121867f $X=1.245 $Y=0.34 $X2=0
+ $Y2=0
cc_333 N_A_27_100#_c_309_p N_VGND_c_1758_n 0.00203854f $X=2.61 $Y=0.81 $X2=0
+ $Y2=0
cc_334 N_A_27_100#_c_262_n N_VGND_c_1762_n 0.00943591f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_335 N_A_27_100#_c_265_n N_VGND_c_1762_n 0.047609f $X=2.445 $Y=0.34 $X2=0
+ $Y2=0
cc_336 N_A_27_100#_c_266_n N_VGND_c_1762_n 0.00660921f $X=1.245 $Y=0.34 $X2=0
+ $Y2=0
cc_337 N_A_27_100#_c_309_p N_VGND_c_1762_n 0.00383647f $X=2.61 $Y=0.81 $X2=0
+ $Y2=0
cc_338 N_A_336_263#_M1011_g N_B_M1008_g 0.0402126f $X=2.79 $Y=2.245 $X2=0 $Y2=0
cc_339 N_A_336_263#_M1003_g N_B_M1013_g 0.0180264f $X=1.795 $Y=0.92 $X2=0 $Y2=0
cc_340 N_A_336_263#_c_387_n N_B_M1013_g 0.0165115f $X=2.75 $Y=0.22 $X2=0 $Y2=0
cc_341 N_A_336_263#_c_392_n N_B_M1013_g 0.00639877f $X=2.8 $Y=1.53 $X2=0 $Y2=0
cc_342 N_A_336_263#_M1011_g N_B_c_507_n 0.00991747f $X=2.79 $Y=2.245 $X2=0 $Y2=0
cc_343 N_A_336_263#_c_387_n N_B_M1015_g 0.00102202f $X=2.75 $Y=0.22 $X2=0 $Y2=0
cc_344 N_A_336_263#_M1011_g N_B_M1015_g 0.00111876f $X=2.79 $Y=2.245 $X2=0 $Y2=0
cc_345 N_A_336_263#_M1030_g N_B_M1015_g 0.020317f $X=2.825 $Y=0.985 $X2=0 $Y2=0
cc_346 N_A_336_263#_c_393_n N_B_M1015_g 0.0105107f $X=4.04 $Y=0.34 $X2=0 $Y2=0
cc_347 N_A_336_263#_c_395_n N_B_c_493_n 0.0132167f $X=4.207 $Y=1.805 $X2=0 $Y2=0
cc_348 N_A_336_263#_c_393_n N_B_c_494_n 0.00872718f $X=4.04 $Y=0.34 $X2=0 $Y2=0
cc_349 N_A_336_263#_c_399_n N_B_c_494_n 0.00168863f $X=4.21 $Y=1.97 $X2=0 $Y2=0
cc_350 N_A_336_263#_c_395_n N_B_c_494_n 0.0136706f $X=4.207 $Y=1.805 $X2=0 $Y2=0
cc_351 N_A_336_263#_c_398_n N_B_M1027_g 0.0124641f $X=4.21 $Y=2.8 $X2=0 $Y2=0
cc_352 N_A_336_263#_c_399_n N_B_M1027_g 0.0025949f $X=4.21 $Y=1.97 $X2=0 $Y2=0
cc_353 N_A_336_263#_c_395_n N_B_M1027_g 0.00401079f $X=4.207 $Y=1.805 $X2=0
+ $Y2=0
cc_354 N_A_336_263#_c_393_n N_B_c_498_n 0.0028132f $X=4.04 $Y=0.34 $X2=0 $Y2=0
cc_355 N_A_336_263#_c_395_n N_B_c_498_n 0.00331719f $X=4.207 $Y=1.805 $X2=0
+ $Y2=0
cc_356 N_A_336_263#_M1000_g N_B_c_501_n 0.030708f $X=1.77 $Y=2.245 $X2=0 $Y2=0
cc_357 N_A_336_263#_M1011_g N_B_c_501_n 0.00639877f $X=2.79 $Y=2.245 $X2=0 $Y2=0
cc_358 N_A_336_263#_M1011_g N_B_c_502_n 0.0269757f $X=2.79 $Y=2.245 $X2=0 $Y2=0
cc_359 N_A_336_263#_c_393_n N_B_c_503_n 0.00127276f $X=4.04 $Y=0.34 $X2=0 $Y2=0
cc_360 N_A_336_263#_c_393_n N_B_c_504_n 0.0199834f $X=4.04 $Y=0.34 $X2=0 $Y2=0
cc_361 N_A_336_263#_c_395_n N_B_c_504_n 0.0232924f $X=4.207 $Y=1.805 $X2=0 $Y2=0
cc_362 N_A_336_263#_M1000_g N_A_374_120#_c_657_n 0.0219108f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_363 N_A_336_263#_M1000_g N_A_374_120#_c_672_n 0.00720952f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_364 N_A_336_263#_M1011_g N_A_374_120#_c_650_n 0.0107473f $X=2.79 $Y=2.245
+ $X2=0 $Y2=0
cc_365 N_A_336_263#_M1000_g N_A_374_120#_c_632_n 0.0021725f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_366 N_A_336_263#_M1000_g N_A_374_120#_c_654_n 0.0118301f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_367 N_A_336_263#_c_391_n N_A_374_120#_c_654_n 4.04023e-19 $X=1.775 $Y=1.465
+ $X2=0 $Y2=0
cc_368 N_A_336_263#_c_391_n N_A_374_120#_c_635_n 0.00306829f $X=1.775 $Y=1.465
+ $X2=0 $Y2=0
cc_369 N_A_336_263#_c_387_n N_A_374_120#_c_641_n 0.00104935f $X=2.75 $Y=0.22
+ $X2=0 $Y2=0
cc_370 N_A_336_263#_M1030_g N_A_374_120#_c_641_n 0.00803161f $X=2.825 $Y=0.985
+ $X2=0 $Y2=0
cc_371 N_A_336_263#_c_393_n N_A_374_120#_c_641_n 0.0815908f $X=4.04 $Y=0.34
+ $X2=0 $Y2=0
cc_372 N_A_336_263#_c_394_n N_A_374_120#_c_641_n 0.00667255f $X=3.115 $Y=0.405
+ $X2=0 $Y2=0
cc_373 N_A_336_263#_M1003_g N_A_374_120#_c_647_n 0.00306829f $X=1.795 $Y=0.92
+ $X2=0 $Y2=0
cc_374 N_A_336_263#_c_387_n N_A_374_120#_c_647_n 0.00183342f $X=2.75 $Y=0.22
+ $X2=0 $Y2=0
cc_375 N_A_336_263#_M1011_g N_A_372_365#_c_907_n 0.0153265f $X=2.79 $Y=2.245
+ $X2=0 $Y2=0
cc_376 N_A_336_263#_M1000_g N_A_372_365#_c_912_n 0.00270446f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_377 N_A_336_263#_c_393_n N_A_372_365#_c_889_n 0.00857875f $X=4.04 $Y=0.34
+ $X2=0 $Y2=0
cc_378 N_A_336_263#_c_399_n N_A_372_365#_c_889_n 0.0093448f $X=4.21 $Y=1.97
+ $X2=0 $Y2=0
cc_379 N_A_336_263#_c_395_n N_A_372_365#_c_889_n 0.0235991f $X=4.207 $Y=1.805
+ $X2=0 $Y2=0
cc_380 N_A_336_263#_c_387_n N_A_372_365#_c_896_n 0.00407716f $X=2.75 $Y=0.22
+ $X2=0 $Y2=0
cc_381 N_A_336_263#_M1011_g N_A_372_365#_c_896_n 0.00983096f $X=2.79 $Y=2.245
+ $X2=0 $Y2=0
cc_382 N_A_336_263#_M1030_g N_A_372_365#_c_896_n 0.00608247f $X=2.825 $Y=0.985
+ $X2=0 $Y2=0
cc_383 N_A_336_263#_c_393_n N_A_372_365#_c_896_n 0.00661426f $X=4.04 $Y=0.34
+ $X2=0 $Y2=0
cc_384 N_A_336_263#_c_394_n N_A_372_365#_c_896_n 0.0119852f $X=3.115 $Y=0.405
+ $X2=0 $Y2=0
cc_385 N_A_336_263#_c_399_n N_VPWR_c_1342_n 0.0451696f $X=4.21 $Y=1.97 $X2=0
+ $Y2=0
cc_386 N_A_336_263#_c_398_n N_VPWR_c_1347_n 0.0139297f $X=4.21 $Y=2.8 $X2=0
+ $Y2=0
cc_387 N_A_336_263#_c_398_n N_VPWR_c_1340_n 0.0121627f $X=4.21 $Y=2.8 $X2=0
+ $Y2=0
cc_388 N_A_336_263#_M1003_g N_A_244_368#_c_1434_n 0.00875874f $X=1.795 $Y=0.92
+ $X2=0 $Y2=0
cc_389 N_A_336_263#_c_391_n N_A_244_368#_c_1434_n 0.00102961f $X=1.775 $Y=1.465
+ $X2=0 $Y2=0
cc_390 N_A_336_263#_M1000_g N_A_244_368#_c_1439_n 0.00524675f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_391 N_A_336_263#_M1011_g N_A_244_368#_c_1439_n 0.00128944f $X=2.79 $Y=2.245
+ $X2=0 $Y2=0
cc_392 N_A_336_263#_c_398_n N_A_244_368#_c_1439_n 0.00429093f $X=4.21 $Y=2.8
+ $X2=0 $Y2=0
cc_393 N_A_336_263#_M1011_g N_A_244_368#_c_1435_n 0.00142796f $X=2.79 $Y=2.245
+ $X2=0 $Y2=0
cc_394 N_A_336_263#_M1030_g N_A_244_368#_c_1435_n 5.75539e-19 $X=2.825 $Y=0.985
+ $X2=0 $Y2=0
cc_395 N_A_336_263#_c_393_n N_A_244_368#_c_1435_n 0.168229f $X=4.04 $Y=0.34
+ $X2=0 $Y2=0
cc_396 N_A_336_263#_M1000_g N_A_244_368#_c_1436_n 0.0114606f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_397 N_A_336_263#_M1000_g N_A_244_368#_c_1437_n 0.00187115f $X=1.77 $Y=2.245
+ $X2=0 $Y2=0
cc_398 N_A_336_263#_c_391_n N_A_244_368#_c_1437_n 0.00357513f $X=1.775 $Y=1.465
+ $X2=0 $Y2=0
cc_399 N_A_336_263#_c_393_n N_A_1026_389#_c_1502_n 9.14388e-19 $X=4.04 $Y=0.34
+ $X2=0 $Y2=0
cc_400 N_A_336_263#_c_393_n N_VGND_c_1753_n 0.0384539f $X=4.04 $Y=0.34 $X2=0
+ $Y2=0
cc_401 N_A_336_263#_c_388_n N_VGND_c_1758_n 0.0290452f $X=1.87 $Y=0.22 $X2=0
+ $Y2=0
cc_402 N_A_336_263#_c_393_n N_VGND_c_1758_n 0.0496789f $X=4.04 $Y=0.34 $X2=0
+ $Y2=0
cc_403 N_A_336_263#_c_394_n N_VGND_c_1758_n 0.0806442f $X=3.115 $Y=0.405 $X2=0
+ $Y2=0
cc_404 N_A_336_263#_c_387_n N_VGND_c_1762_n 0.0328229f $X=2.75 $Y=0.22 $X2=0
+ $Y2=0
cc_405 N_A_336_263#_c_388_n N_VGND_c_1762_n 0.00542545f $X=1.87 $Y=0.22 $X2=0
+ $Y2=0
cc_406 N_A_336_263#_c_393_n N_VGND_c_1762_n 0.0269422f $X=4.04 $Y=0.34 $X2=0
+ $Y2=0
cc_407 N_A_336_263#_c_394_n N_VGND_c_1762_n 0.0458316f $X=3.115 $Y=0.405 $X2=0
+ $Y2=0
cc_408 N_B_M1008_g N_A_374_120#_c_657_n 0.00175329f $X=2.34 $Y=2.245 $X2=0 $Y2=0
cc_409 N_B_M1008_g N_A_374_120#_c_650_n 0.0121772f $X=2.34 $Y=2.245 $X2=0 $Y2=0
cc_410 N_B_c_507_n N_A_374_120#_c_650_n 0.00285336f $X=3.31 $Y=3.11 $X2=0 $Y2=0
cc_411 N_B_M1019_g N_A_374_120#_c_650_n 0.00138352f $X=3.4 $Y=2.245 $X2=0 $Y2=0
cc_412 N_B_M1013_g N_A_374_120#_c_632_n 0.00116618f $X=2.385 $Y=0.985 $X2=0
+ $Y2=0
cc_413 N_B_c_501_n N_A_374_120#_c_632_n 0.00179652f $X=2.355 $Y=1.615 $X2=0
+ $Y2=0
cc_414 N_B_M1008_g N_A_374_120#_c_654_n 0.00167773f $X=2.34 $Y=2.245 $X2=0 $Y2=0
cc_415 N_B_c_501_n N_A_374_120#_c_635_n 0.00119961f $X=2.355 $Y=1.615 $X2=0
+ $Y2=0
cc_416 N_B_M1031_g N_A_374_120#_c_637_n 0.00132931f $X=5.285 $Y=0.69 $X2=0 $Y2=0
cc_417 N_B_c_505_n N_A_374_120#_c_637_n 3.79762e-19 $X=5.04 $Y=1.385 $X2=0 $Y2=0
cc_418 N_B_M1013_g N_A_374_120#_c_641_n 0.00778522f $X=2.385 $Y=0.985 $X2=0
+ $Y2=0
cc_419 N_B_M1015_g N_A_374_120#_c_641_n 0.00678832f $X=3.43 $Y=0.985 $X2=0 $Y2=0
cc_420 N_B_c_495_n N_A_374_120#_c_641_n 0.0048712f $X=3.99 $Y=1.475 $X2=0 $Y2=0
cc_421 N_B_c_498_n N_A_374_120#_c_641_n 0.00835586f $X=4.81 $Y=1.22 $X2=0 $Y2=0
cc_422 N_B_M1031_g N_A_374_120#_c_641_n 0.00722002f $X=5.285 $Y=0.69 $X2=0 $Y2=0
cc_423 N_B_c_502_n N_A_374_120#_c_641_n 4.83406e-19 $X=3.407 $Y=1.75 $X2=0 $Y2=0
cc_424 N_B_c_504_n N_A_374_120#_c_641_n 0.0134657f $X=4.9 $Y=1.385 $X2=0 $Y2=0
cc_425 N_B_c_505_n N_A_374_120#_c_641_n 0.00161804f $X=5.04 $Y=1.385 $X2=0 $Y2=0
cc_426 N_B_M1013_g N_A_374_120#_c_666_n 0.00166189f $X=2.385 $Y=0.985 $X2=0
+ $Y2=0
cc_427 N_B_c_501_n N_A_374_120#_c_666_n 7.68744e-19 $X=2.355 $Y=1.615 $X2=0
+ $Y2=0
cc_428 N_B_M1031_g N_A_374_120#_c_644_n 0.00115827f $X=5.285 $Y=0.69 $X2=0 $Y2=0
cc_429 N_B_M1001_g N_A_374_120#_c_646_n 0.0260222f $X=5.04 $Y=2.445 $X2=0 $Y2=0
cc_430 N_B_c_505_n N_A_374_120#_c_646_n 0.00431096f $X=5.04 $Y=1.385 $X2=0 $Y2=0
cc_431 N_B_M1013_g N_A_374_120#_c_647_n 0.00519945f $X=2.385 $Y=0.985 $X2=0
+ $Y2=0
cc_432 N_B_M1008_g N_A_372_365#_c_907_n 0.0142316f $X=2.34 $Y=2.245 $X2=0 $Y2=0
cc_433 N_B_M1015_g N_A_372_365#_c_889_n 0.00435531f $X=3.43 $Y=0.985 $X2=0 $Y2=0
cc_434 N_B_c_493_n N_A_372_365#_c_889_n 0.0138354f $X=3.915 $Y=3.035 $X2=0 $Y2=0
cc_435 N_B_c_494_n N_A_372_365#_c_889_n 0.00104939f $X=4.345 $Y=1.475 $X2=0
+ $Y2=0
cc_436 N_B_M1027_g N_A_372_365#_c_889_n 0.011688f $X=4.435 $Y=2.385 $X2=0 $Y2=0
cc_437 N_B_c_497_n N_A_372_365#_c_889_n 0.00647571f $X=4.735 $Y=1.475 $X2=0
+ $Y2=0
cc_438 N_B_M1001_g N_A_372_365#_c_889_n 0.0134193f $X=5.04 $Y=2.445 $X2=0 $Y2=0
cc_439 N_B_c_502_n N_A_372_365#_c_889_n 0.0072953f $X=3.407 $Y=1.75 $X2=0 $Y2=0
cc_440 N_B_c_504_n N_A_372_365#_c_889_n 0.0242833f $X=4.9 $Y=1.385 $X2=0 $Y2=0
cc_441 N_B_c_505_n N_A_372_365#_c_889_n 0.00272371f $X=5.04 $Y=1.385 $X2=0 $Y2=0
cc_442 N_B_M1015_g N_A_372_365#_c_896_n 0.0079635f $X=3.43 $Y=0.985 $X2=0 $Y2=0
cc_443 N_B_c_502_n N_A_372_365#_c_896_n 0.00471064f $X=3.407 $Y=1.75 $X2=0 $Y2=0
cc_444 N_B_c_493_n N_VPWR_c_1342_n 0.0021388f $X=3.915 $Y=3.035 $X2=0 $Y2=0
cc_445 N_B_M1027_g N_VPWR_c_1342_n 0.00409571f $X=4.435 $Y=2.385 $X2=0 $Y2=0
cc_446 N_B_c_497_n N_VPWR_c_1342_n 0.00551661f $X=4.735 $Y=1.475 $X2=0 $Y2=0
cc_447 N_B_M1001_g N_VPWR_c_1342_n 0.0150854f $X=5.04 $Y=2.445 $X2=0 $Y2=0
cc_448 N_B_c_504_n N_VPWR_c_1342_n 0.0131178f $X=4.9 $Y=1.385 $X2=0 $Y2=0
cc_449 N_B_M1001_g N_VPWR_c_1345_n 0.00648879f $X=5.04 $Y=2.445 $X2=0 $Y2=0
cc_450 N_B_c_508_n N_VPWR_c_1347_n 0.037974f $X=2.43 $Y=3.11 $X2=0 $Y2=0
cc_451 N_B_M1027_g N_VPWR_c_1347_n 0.00648879f $X=4.435 $Y=2.385 $X2=0 $Y2=0
cc_452 N_B_c_507_n N_VPWR_c_1340_n 0.021021f $X=3.31 $Y=3.11 $X2=0 $Y2=0
cc_453 N_B_c_508_n N_VPWR_c_1340_n 0.00617673f $X=2.43 $Y=3.11 $X2=0 $Y2=0
cc_454 N_B_c_510_n N_VPWR_c_1340_n 0.020539f $X=3.84 $Y=3.11 $X2=0 $Y2=0
cc_455 N_B_M1027_g N_VPWR_c_1340_n 0.00649272f $X=4.435 $Y=2.385 $X2=0 $Y2=0
cc_456 N_B_M1001_g N_VPWR_c_1340_n 0.00649272f $X=5.04 $Y=2.445 $X2=0 $Y2=0
cc_457 N_B_c_515_n N_VPWR_c_1340_n 0.00450763f $X=3.4 $Y=3.11 $X2=0 $Y2=0
cc_458 N_B_M1008_g N_A_244_368#_c_1439_n 0.0108311f $X=2.34 $Y=2.245 $X2=0 $Y2=0
cc_459 N_B_c_507_n N_A_244_368#_c_1439_n 0.0198022f $X=3.31 $Y=3.11 $X2=0 $Y2=0
cc_460 N_B_c_508_n N_A_244_368#_c_1439_n 0.00301961f $X=2.43 $Y=3.11 $X2=0 $Y2=0
cc_461 N_B_M1019_g N_A_244_368#_c_1439_n 0.0134297f $X=3.4 $Y=2.245 $X2=0 $Y2=0
cc_462 N_B_c_510_n N_A_244_368#_c_1439_n 0.00852151f $X=3.84 $Y=3.11 $X2=0 $Y2=0
cc_463 N_B_c_493_n N_A_244_368#_c_1439_n 0.00298988f $X=3.915 $Y=3.035 $X2=0
+ $Y2=0
cc_464 N_B_c_515_n N_A_244_368#_c_1439_n 0.00202929f $X=3.4 $Y=3.11 $X2=0 $Y2=0
cc_465 N_B_M1019_g N_A_244_368#_c_1435_n 0.0252623f $X=3.4 $Y=2.245 $X2=0 $Y2=0
cc_466 N_B_M1015_g N_A_244_368#_c_1435_n 0.0168273f $X=3.43 $Y=0.985 $X2=0 $Y2=0
cc_467 N_B_c_495_n N_A_244_368#_c_1435_n 0.0149705f $X=3.99 $Y=1.475 $X2=0 $Y2=0
cc_468 N_B_c_502_n N_A_244_368#_c_1435_n 0.00366082f $X=3.407 $Y=1.75 $X2=0
+ $Y2=0
cc_469 N_B_M1001_g N_A_1026_389#_c_1505_n 0.0110275f $X=5.04 $Y=2.445 $X2=0
+ $Y2=0
cc_470 N_B_c_498_n N_A_1026_389#_c_1502_n 8.75563e-19 $X=4.81 $Y=1.22 $X2=0
+ $Y2=0
cc_471 N_B_M1031_g N_A_1026_389#_c_1502_n 0.0128414f $X=5.285 $Y=0.69 $X2=0
+ $Y2=0
cc_472 N_B_M1031_g N_A_1026_389#_c_1512_n 0.00312633f $X=5.285 $Y=0.69 $X2=0
+ $Y2=0
cc_473 N_B_M1001_g N_A_1026_389#_c_1506_n 0.00265349f $X=5.04 $Y=2.445 $X2=0
+ $Y2=0
cc_474 N_B_c_505_n N_A_1026_389#_c_1506_n 0.00220282f $X=5.04 $Y=1.385 $X2=0
+ $Y2=0
cc_475 N_B_c_504_n N_A_1026_389#_c_1503_n 0.0190992f $X=4.9 $Y=1.385 $X2=0 $Y2=0
cc_476 N_B_c_505_n N_A_1026_389#_c_1503_n 0.017036f $X=5.04 $Y=1.385 $X2=0 $Y2=0
cc_477 N_B_c_498_n N_A_1026_389#_c_1504_n 2.99244e-19 $X=4.81 $Y=1.22 $X2=0
+ $Y2=0
cc_478 N_B_M1031_g N_A_1026_389#_c_1504_n 0.00482748f $X=5.285 $Y=0.69 $X2=0
+ $Y2=0
cc_479 N_B_c_504_n N_A_1026_389#_c_1504_n 0.00977411f $X=4.9 $Y=1.385 $X2=0
+ $Y2=0
cc_480 N_B_c_505_n N_A_1026_389#_c_1504_n 0.00402809f $X=5.04 $Y=1.385 $X2=0
+ $Y2=0
cc_481 N_B_c_498_n N_VGND_c_1753_n 0.00249524f $X=4.81 $Y=1.22 $X2=0 $Y2=0
cc_482 N_B_M1031_g N_VGND_c_1753_n 0.0044164f $X=5.285 $Y=0.69 $X2=0 $Y2=0
cc_483 N_B_c_504_n N_VGND_c_1753_n 0.00792756f $X=4.9 $Y=1.385 $X2=0 $Y2=0
cc_484 N_B_c_505_n N_VGND_c_1753_n 0.00265976f $X=5.04 $Y=1.385 $X2=0 $Y2=0
cc_485 N_B_c_498_n N_VGND_c_1758_n 0.00461464f $X=4.81 $Y=1.22 $X2=0 $Y2=0
cc_486 N_B_M1031_g N_VGND_c_1759_n 0.00423055f $X=5.285 $Y=0.69 $X2=0 $Y2=0
cc_487 N_B_c_498_n N_VGND_c_1762_n 0.00912981f $X=4.81 $Y=1.22 $X2=0 $Y2=0
cc_488 N_B_M1031_g N_VGND_c_1762_n 0.00786497f $X=5.285 $Y=0.69 $X2=0 $Y2=0
cc_489 N_A_374_120#_c_641_n N_A_372_365#_M1030_d 0.00514299f $X=5.855 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_490 N_A_374_120#_c_650_n N_A_372_365#_M1000_d 0.00623621f $X=3.095 $Y=2.65
+ $X2=0 $Y2=0
cc_491 N_A_374_120#_c_654_n N_A_372_365#_M1000_d 0.00503007f $X=2.01 $Y=1.745
+ $X2=0 $Y2=0
cc_492 N_A_374_120#_c_631_n N_A_372_365#_M1016_g 0.00916477f $X=6.985 $Y=1.13
+ $X2=0 $Y2=0
cc_493 N_A_374_120#_c_652_n N_A_372_365#_M1016_g 6.40864e-19 $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_494 N_A_374_120#_c_634_n N_A_372_365#_M1016_g 0.007221f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_495 N_A_374_120#_c_636_n N_A_372_365#_M1016_g 3.57482e-19 $X=5.735 $Y=1.64
+ $X2=0 $Y2=0
cc_496 N_A_374_120#_c_637_n N_A_372_365#_M1016_g 0.0045902f $X=5.702 $Y=1.475
+ $X2=0 $Y2=0
cc_497 N_A_374_120#_c_716_p N_A_372_365#_M1016_g 0.00709291f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_498 N_A_374_120#_c_642_n N_A_372_365#_M1016_g 0.00418011f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_499 N_A_374_120#_c_644_n N_A_372_365#_M1016_g 0.00440701f $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_500 N_A_374_120#_c_646_n N_A_372_365#_M1016_g 0.0181029f $X=5.575 $Y=1.64
+ $X2=0 $Y2=0
cc_501 N_A_374_120#_M1022_g N_A_372_365#_M1026_g 0.00987226f $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_502 N_A_374_120#_c_721_p N_A_372_365#_M1026_g 0.0102405f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_503 N_A_374_120#_M1010_g N_A_372_365#_c_887_n 0.0411135f $X=9.5 $Y=2.26 $X2=0
+ $Y2=0
cc_504 N_A_374_120#_c_639_n N_A_372_365#_c_887_n 0.00578673f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_505 N_A_374_120#_M1011_d N_A_372_365#_c_907_n 0.0053241f $X=2.88 $Y=1.825
+ $X2=0 $Y2=0
cc_506 N_A_374_120#_c_650_n N_A_372_365#_c_907_n 0.06129f $X=3.095 $Y=2.65 $X2=0
+ $Y2=0
cc_507 N_A_374_120#_c_657_n N_A_372_365#_c_912_n 0.0277311f $X=1.775 $Y=2.565
+ $X2=0 $Y2=0
cc_508 N_A_374_120#_c_650_n N_A_372_365#_c_912_n 0.0126173f $X=3.095 $Y=2.65
+ $X2=0 $Y2=0
cc_509 N_A_374_120#_c_654_n N_A_372_365#_c_912_n 0.0049846f $X=2.01 $Y=1.745
+ $X2=0 $Y2=0
cc_510 N_A_374_120#_c_635_n N_A_372_365#_c_912_n 0.00328015f $X=2.1 $Y=1.325
+ $X2=0 $Y2=0
cc_511 N_A_374_120#_c_636_n N_A_372_365#_c_889_n 0.0241822f $X=5.735 $Y=1.64
+ $X2=0 $Y2=0
cc_512 N_A_374_120#_c_642_n N_A_372_365#_c_889_n 0.0134696f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_513 N_A_374_120#_c_644_n N_A_372_365#_c_889_n 0.00188072f $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_514 N_A_374_120#_c_646_n N_A_372_365#_c_889_n 0.00744324f $X=5.575 $Y=1.64
+ $X2=0 $Y2=0
cc_515 N_A_374_120#_c_641_n N_A_372_365#_c_909_n 0.0110709f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_516 N_A_374_120#_c_652_n N_A_372_365#_c_890_n 0.0215322f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_517 N_A_374_120#_c_634_n N_A_372_365#_c_890_n 0.00213765f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_518 N_A_374_120#_c_643_n N_A_372_365#_c_890_n 0.0112688f $X=7.105 $Y=0.925
+ $X2=0 $Y2=0
cc_519 N_A_374_120#_c_652_n N_A_372_365#_c_891_n 0.00254666f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_520 N_A_374_120#_c_634_n N_A_372_365#_c_891_n 0.00134421f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_521 N_A_374_120#_c_716_p N_A_372_365#_c_891_n 0.011115f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_522 N_A_374_120#_c_652_n N_A_372_365#_c_892_n 0.0129058f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_523 N_A_374_120#_c_634_n N_A_372_365#_c_892_n 9.12819e-19 $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_524 N_A_374_120#_c_721_p N_A_372_365#_c_903_n 0.0114531f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_525 N_A_374_120#_M1012_g N_A_372_365#_c_893_n 0.0179651f $X=5.575 $Y=2.525
+ $X2=0 $Y2=0
cc_526 N_A_374_120#_c_652_n N_A_372_365#_c_893_n 8.06489e-19 $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_527 N_A_374_120#_c_634_n N_A_372_365#_c_893_n 0.017203f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_528 N_A_374_120#_c_639_n N_A_372_365#_c_894_n 0.00245381f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_529 N_A_374_120#_c_721_p N_A_372_365#_c_895_n 0.00965476f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_530 N_A_374_120#_M1011_d N_A_372_365#_c_896_n 0.00948865f $X=2.88 $Y=1.825
+ $X2=0 $Y2=0
cc_531 N_A_374_120#_c_641_n N_A_372_365#_c_896_n 0.0230041f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_532 N_A_374_120#_c_631_n N_CI_M1025_g 0.00955653f $X=6.985 $Y=1.13 $X2=0
+ $Y2=0
cc_533 N_A_374_120#_c_634_n N_CI_M1025_g 0.00321559f $X=6.985 $Y=1.295 $X2=0
+ $Y2=0
cc_534 N_A_374_120#_c_721_p N_CI_M1025_g 0.0113056f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_535 N_A_374_120#_c_721_p N_CI_c_1054_n 0.00896038f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_536 N_A_374_120#_c_721_p CI 0.00563052f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_537 N_A_374_120#_c_652_n N_CI_c_1057_n 5.14735e-19 $X=6.985 $Y=1.295 $X2=0
+ $Y2=0
cc_538 N_A_374_120#_c_634_n N_CI_c_1057_n 0.0288449f $X=6.985 $Y=1.295 $X2=0
+ $Y2=0
cc_539 N_A_374_120#_c_721_p N_CI_c_1057_n 0.00208687f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_540 N_A_374_120#_c_721_p N_A_1609_368#_M1004_d 0.00255432f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_541 N_A_374_120#_M1022_g N_A_1609_368#_M1017_g 0.0139157f $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_542 N_A_374_120#_c_640_n N_A_1609_368#_M1017_g 0.00305336f $X=9.582 $Y=1.26
+ $X2=0 $Y2=0
cc_543 N_A_374_120#_c_762_p N_A_1609_368#_M1017_g 2.03926e-19 $X=9.56 $Y=0.925
+ $X2=0 $Y2=0
cc_544 N_A_374_120#_c_721_p N_A_1609_368#_c_1118_n 0.0231003f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_545 N_A_374_120#_M1010_g N_A_1609_368#_c_1128_n 0.0192317f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_546 N_A_374_120#_M1010_g N_A_1609_368#_c_1129_n 0.00752003f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_547 N_A_374_120#_c_721_p N_A_1609_368#_c_1120_n 0.0178279f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_548 N_A_374_120#_M1010_g N_A_1609_368#_c_1131_n 0.00370188f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_549 N_A_374_120#_c_638_n N_A_1609_368#_c_1131_n 0.00871051f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_550 N_A_374_120#_c_639_n N_A_1609_368#_c_1131_n 0.00308826f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_551 N_A_374_120#_M1010_g N_A_1609_368#_c_1121_n 0.00479784f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_552 N_A_374_120#_c_638_n N_A_1609_368#_c_1122_n 0.0258294f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_553 N_A_374_120#_c_639_n N_A_1609_368#_c_1122_n 0.00214701f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_554 N_A_374_120#_c_638_n N_A_1609_368#_c_1123_n 3.10403e-19 $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_555 N_A_374_120#_c_639_n N_A_1609_368#_c_1123_n 0.0206892f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_556 N_A_374_120#_c_721_p N_A_1744_94#_M1026_d 0.0046102f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_557 N_A_374_120#_c_776_p N_A_1744_94#_M1026_d 0.00334362f $X=9.36 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_558 N_A_374_120#_c_762_p N_A_1744_94#_M1026_d 0.00198141f $X=9.56 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_559 N_A_374_120#_M1022_g N_A_1744_94#_c_1233_n 0.00395783f $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_560 N_A_374_120#_c_640_n N_A_1744_94#_c_1233_n 0.0200673f $X=9.582 $Y=1.26
+ $X2=0 $Y2=0
cc_561 N_A_374_120#_c_721_p N_A_1744_94#_c_1233_n 0.0144192f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_562 N_A_374_120#_c_776_p N_A_1744_94#_c_1233_n 0.00557132f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_563 N_A_374_120#_c_762_p N_A_1744_94#_c_1233_n 0.00727454f $X=9.56 $Y=0.925
+ $X2=0 $Y2=0
cc_564 N_A_374_120#_M1022_g N_A_1744_94#_c_1234_n 0.00959577f $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_565 N_A_374_120#_c_721_p N_A_1744_94#_c_1234_n 0.0241653f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_566 N_A_374_120#_c_776_p N_A_1744_94#_c_1234_n 0.00142094f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_567 N_A_374_120#_c_762_p N_A_1744_94#_c_1234_n 0.0106426f $X=9.56 $Y=0.925
+ $X2=0 $Y2=0
cc_568 N_A_374_120#_M1022_g N_A_1744_94#_c_1235_n 0.0098518f $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_569 N_A_374_120#_c_721_p N_A_1744_94#_c_1235_n 0.00384885f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_570 N_A_374_120#_c_776_p N_A_1744_94#_c_1235_n 0.00730033f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_571 N_A_374_120#_c_762_p N_A_1744_94#_c_1235_n 0.00953934f $X=9.56 $Y=0.925
+ $X2=0 $Y2=0
cc_572 N_A_374_120#_M1022_g N_A_1744_94#_c_1237_n 6.84725e-19 $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_573 N_A_374_120#_M1010_g N_A_1744_94#_c_1238_n 0.00247031f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_574 N_A_374_120#_c_638_n N_A_1744_94#_c_1238_n 0.0151235f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_575 N_A_374_120#_c_639_n N_A_1744_94#_c_1238_n 0.00193209f $X=9.58 $Y=1.425
+ $X2=0 $Y2=0
cc_576 N_A_374_120#_M1012_g N_VPWR_c_1345_n 0.00680602f $X=5.575 $Y=2.525 $X2=0
+ $Y2=0
cc_577 N_A_374_120#_M1012_g N_VPWR_c_1340_n 0.00649272f $X=5.575 $Y=2.525 $X2=0
+ $Y2=0
cc_578 N_A_374_120#_c_672_n N_A_244_368#_c_1438_n 0.0141144f $X=1.86 $Y=2.65
+ $X2=0 $Y2=0
cc_579 N_A_374_120#_c_666_n N_A_244_368#_c_1434_n 0.00131974f $X=2.305 $Y=0.925
+ $X2=0 $Y2=0
cc_580 N_A_374_120#_c_647_n N_A_244_368#_c_1434_n 0.0201235f $X=2.09 $Y=0.76
+ $X2=0 $Y2=0
cc_581 N_A_374_120#_c_672_n N_A_244_368#_c_1439_n 0.0127477f $X=1.86 $Y=2.65
+ $X2=0 $Y2=0
cc_582 N_A_374_120#_c_650_n N_A_244_368#_c_1439_n 0.0969641f $X=3.095 $Y=2.65
+ $X2=0 $Y2=0
cc_583 N_A_374_120#_c_650_n N_A_244_368#_c_1435_n 0.00843289f $X=3.095 $Y=2.65
+ $X2=0 $Y2=0
cc_584 N_A_374_120#_c_641_n N_A_244_368#_c_1435_n 0.0327138f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_585 N_A_374_120#_c_657_n N_A_244_368#_c_1436_n 0.0541992f $X=1.775 $Y=2.565
+ $X2=0 $Y2=0
cc_586 N_A_374_120#_c_632_n N_A_244_368#_c_1436_n 0.0069711f $X=2.01 $Y=1.66
+ $X2=0 $Y2=0
cc_587 N_A_374_120#_c_654_n N_A_244_368#_c_1436_n 0.0128838f $X=2.01 $Y=1.745
+ $X2=0 $Y2=0
cc_588 N_A_374_120#_c_654_n N_A_244_368#_c_1437_n 0.00411346f $X=2.01 $Y=1.745
+ $X2=0 $Y2=0
cc_589 N_A_374_120#_c_635_n N_A_244_368#_c_1437_n 0.0201235f $X=2.1 $Y=1.325
+ $X2=0 $Y2=0
cc_590 N_A_374_120#_c_641_n N_A_1026_389#_M1031_d 0.00538208f $X=5.855 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_591 N_A_374_120#_c_642_n N_A_1026_389#_M1031_d 0.00208559f $X=6.145 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_592 N_A_374_120#_c_644_n N_A_1026_389#_M1031_d 0.00883869f $X=6 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_593 N_A_374_120#_c_637_n N_A_1026_389#_c_1502_n 0.00715307f $X=5.702 $Y=1.475
+ $X2=0 $Y2=0
cc_594 N_A_374_120#_c_641_n N_A_1026_389#_c_1502_n 0.0156475f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_595 N_A_374_120#_c_642_n N_A_1026_389#_c_1502_n 4.25711e-19 $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_596 N_A_374_120#_c_644_n N_A_1026_389#_c_1502_n 0.0164358f $X=6 $Y=0.925
+ $X2=0 $Y2=0
cc_597 N_A_374_120#_c_641_n N_A_1026_389#_c_1528_n 0.00899783f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_598 N_A_374_120#_c_642_n N_A_1026_389#_c_1528_n 0.00817197f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_599 N_A_374_120#_c_644_n N_A_1026_389#_c_1528_n 0.0284519f $X=6 $Y=0.925
+ $X2=0 $Y2=0
cc_600 N_A_374_120#_M1012_g N_A_1026_389#_c_1506_n 0.00658216f $X=5.575 $Y=2.525
+ $X2=0 $Y2=0
cc_601 N_A_374_120#_c_636_n N_A_1026_389#_c_1503_n 0.0235409f $X=5.735 $Y=1.64
+ $X2=0 $Y2=0
cc_602 N_A_374_120#_c_637_n N_A_1026_389#_c_1503_n 0.00937212f $X=5.702 $Y=1.475
+ $X2=0 $Y2=0
cc_603 N_A_374_120#_c_646_n N_A_1026_389#_c_1503_n 0.00465684f $X=5.575 $Y=1.64
+ $X2=0 $Y2=0
cc_604 N_A_374_120#_c_637_n N_A_1026_389#_c_1504_n 0.013153f $X=5.702 $Y=1.475
+ $X2=0 $Y2=0
cc_605 N_A_374_120#_c_641_n N_A_1026_389#_c_1504_n 0.00471784f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_606 N_A_374_120#_c_646_n N_A_1026_389#_c_1504_n 2.62009e-19 $X=5.575 $Y=1.64
+ $X2=0 $Y2=0
cc_607 N_A_374_120#_c_716_p N_COUT_N_M1016_d 0.013849f $X=6.815 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_608 N_A_374_120#_c_643_n N_COUT_N_M1016_d 5.04966e-19 $X=7.105 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_609 N_A_374_120#_M1012_g N_COUT_N_c_1560_n 0.0100995f $X=5.575 $Y=2.525 $X2=0
+ $Y2=0
cc_610 N_A_374_120#_c_636_n N_COUT_N_c_1560_n 0.0022531f $X=5.735 $Y=1.64 $X2=0
+ $Y2=0
cc_611 N_A_374_120#_c_646_n N_COUT_N_c_1560_n 0.00292755f $X=5.575 $Y=1.64 $X2=0
+ $Y2=0
cc_612 N_A_374_120#_M1012_g N_COUT_N_c_1557_n 0.00245884f $X=5.575 $Y=2.525
+ $X2=0 $Y2=0
cc_613 N_A_374_120#_c_652_n N_COUT_N_c_1557_n 0.00397215f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_614 N_A_374_120#_c_634_n N_COUT_N_c_1557_n 6.77617e-19 $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_615 N_A_374_120#_c_637_n N_COUT_N_c_1557_n 0.0304246f $X=5.702 $Y=1.475 $X2=0
+ $Y2=0
cc_616 N_A_374_120#_c_646_n N_COUT_N_c_1557_n 0.00196317f $X=5.575 $Y=1.64 $X2=0
+ $Y2=0
cc_617 N_A_374_120#_c_633_n N_COUT_N_c_1558_n 0.0139862f $X=6.977 $Y=1.287 $X2=0
+ $Y2=0
cc_618 N_A_374_120#_c_634_n N_COUT_N_c_1558_n 0.00165279f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_619 N_A_374_120#_c_637_n N_COUT_N_c_1558_n 0.0141264f $X=5.702 $Y=1.475 $X2=0
+ $Y2=0
cc_620 N_A_374_120#_c_716_p N_COUT_N_c_1558_n 0.00699693f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_621 N_A_374_120#_c_642_n N_COUT_N_c_1558_n 0.00177565f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_622 N_A_374_120#_c_644_n N_COUT_N_c_1558_n 0.00727468f $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_623 N_A_374_120#_c_631_n COUT_N 0.00709084f $X=6.985 $Y=1.13 $X2=0 $Y2=0
cc_624 N_A_374_120#_c_634_n COUT_N 7.56021e-19 $X=6.985 $Y=1.295 $X2=0 $Y2=0
cc_625 N_A_374_120#_c_637_n COUT_N 0.00648383f $X=5.702 $Y=1.475 $X2=0 $Y2=0
cc_626 N_A_374_120#_c_716_p COUT_N 0.0299539f $X=6.815 $Y=0.925 $X2=0 $Y2=0
cc_627 N_A_374_120#_c_642_n COUT_N 0.00234721f $X=6.145 $Y=0.925 $X2=0 $Y2=0
cc_628 N_A_374_120#_c_643_n COUT_N 0.00262708f $X=7.105 $Y=0.925 $X2=0 $Y2=0
cc_629 N_A_374_120#_c_644_n COUT_N 0.00676707f $X=6 $Y=0.925 $X2=0 $Y2=0
cc_630 N_A_374_120#_c_645_n COUT_N 0.0260829f $X=6.96 $Y=0.925 $X2=0 $Y2=0
cc_631 N_A_374_120#_c_721_p N_A_1264_421#_M1018_d 0.0129911f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_632 N_A_374_120#_c_643_n N_A_1264_421#_M1018_d 0.00241431f $X=7.105 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_633 N_A_374_120#_c_645_n N_A_1264_421#_M1018_d 0.00131937f $X=6.96 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_634 N_A_374_120#_c_652_n N_A_1264_421#_c_1614_n 0.0160329f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_635 N_A_374_120#_c_634_n N_A_1264_421#_c_1614_n 0.00298281f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_636 N_A_374_120#_c_631_n N_A_1264_421#_c_1612_n 0.00540965f $X=6.985 $Y=1.13
+ $X2=0 $Y2=0
cc_637 N_A_374_120#_c_631_n N_A_1264_421#_c_1613_n 5.39759e-19 $X=6.985 $Y=1.13
+ $X2=0 $Y2=0
cc_638 N_A_374_120#_c_633_n N_A_1264_421#_c_1613_n 0.0491204f $X=6.977 $Y=1.287
+ $X2=0 $Y2=0
cc_639 N_A_374_120#_c_634_n N_A_1264_421#_c_1613_n 0.00411498f $X=6.985 $Y=1.295
+ $X2=0 $Y2=0
cc_640 N_A_374_120#_c_721_p N_A_1264_421#_c_1613_n 0.00757493f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_641 N_A_374_120#_c_643_n N_A_1264_421#_c_1613_n 0.00128603f $X=7.105 $Y=0.925
+ $X2=0 $Y2=0
cc_642 N_A_374_120#_c_645_n N_A_1264_421#_c_1613_n 0.00952721f $X=6.96 $Y=0.925
+ $X2=0 $Y2=0
cc_643 N_A_374_120#_c_631_n N_A_1264_421#_c_1628_n 4.58038e-19 $X=6.985 $Y=1.13
+ $X2=0 $Y2=0
cc_644 N_A_374_120#_c_721_p N_A_1264_421#_c_1628_n 0.0247429f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_645 N_A_374_120#_c_643_n N_A_1264_421#_c_1628_n 0.00135086f $X=7.105 $Y=0.925
+ $X2=0 $Y2=0
cc_646 N_A_374_120#_c_645_n N_A_1264_421#_c_1628_n 0.0103098f $X=6.96 $Y=0.925
+ $X2=0 $Y2=0
cc_647 N_A_374_120#_c_640_n N_A_1719_368#_M1022_d 8.95266e-19 $X=9.582 $Y=1.26
+ $X2=-0.19 $Y2=-0.245
cc_648 N_A_374_120#_c_762_p N_A_1719_368#_M1022_d 0.0031492f $X=9.56 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_649 N_A_374_120#_M1010_g N_A_1719_368#_c_1660_n 0.00582438f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_650 N_A_374_120#_M1022_g N_A_1719_368#_c_1668_n 0.00459564f $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_651 N_A_374_120#_c_776_p N_A_1719_368#_c_1668_n 5.68711e-19 $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_652 N_A_374_120#_c_762_p N_A_1719_368#_c_1668_n 0.00789043f $X=9.56 $Y=0.925
+ $X2=0 $Y2=0
cc_653 N_A_374_120#_M1022_g N_A_1719_368#_c_1671_n 5.94451e-19 $X=9.455 $Y=0.79
+ $X2=0 $Y2=0
cc_654 N_A_374_120#_c_640_n N_A_1719_368#_c_1671_n 0.00406789f $X=9.582 $Y=1.26
+ $X2=0 $Y2=0
cc_655 N_A_374_120#_c_776_p N_A_1719_368#_c_1671_n 7.05632e-19 $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_656 N_A_374_120#_c_762_p N_A_1719_368#_c_1671_n 0.00956585f $X=9.56 $Y=0.925
+ $X2=0 $Y2=0
cc_657 N_A_374_120#_M1010_g N_A_1719_368#_c_1661_n 0.00374674f $X=9.5 $Y=2.26
+ $X2=0 $Y2=0
cc_658 N_A_374_120#_c_641_n N_VGND_M1024_d 0.00856848f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_659 N_A_374_120#_c_721_p N_VGND_M1025_d 0.00607567f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_660 N_A_374_120#_c_641_n N_VGND_c_1753_n 0.0205911f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_661 N_A_374_120#_c_721_p N_VGND_c_1754_n 0.0228047f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_662 N_A_374_120#_c_631_n N_VGND_c_1759_n 0.00461464f $X=6.985 $Y=1.13 $X2=0
+ $Y2=0
cc_663 N_A_374_120#_M1022_g N_VGND_c_1760_n 7.64118e-19 $X=9.455 $Y=0.79 $X2=0
+ $Y2=0
cc_664 N_A_374_120#_c_631_n N_VGND_c_1762_n 0.00461089f $X=6.985 $Y=1.13 $X2=0
+ $Y2=0
cc_665 N_A_374_120#_c_645_n N_VGND_c_1762_n 0.00598527f $X=6.96 $Y=0.925 $X2=0
+ $Y2=0
cc_666 N_A_372_365#_c_890_n N_CI_c_1058_n 8.94599e-19 $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_667 N_A_372_365#_c_890_n N_CI_M1006_g 0.00752551f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_668 N_A_372_365#_M1026_g N_CI_c_1054_n 0.0172282f $X=8.645 $Y=0.79 $X2=0
+ $Y2=0
cc_669 N_A_372_365#_c_890_n N_CI_c_1055_n 0.00383194f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_670 N_A_372_365#_c_890_n CI 0.0139637f $X=8.735 $Y=1.665 $X2=0 $Y2=0
cc_671 N_A_372_365#_c_890_n N_CI_c_1057_n 0.010759f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_672 N_A_372_365#_c_894_n N_CI_c_1057_n 0.00883838f $X=8.64 $Y=1.465 $X2=0
+ $Y2=0
cc_673 N_A_372_365#_c_890_n N_A_1609_368#_c_1126_n 0.00891013f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_674 N_A_372_365#_M1007_g N_A_1609_368#_c_1127_n 0.00426854f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_675 N_A_372_365#_M1026_g N_A_1609_368#_c_1118_n 0.00489776f $X=8.645 $Y=0.79
+ $X2=0 $Y2=0
cc_676 N_A_372_365#_M1007_g N_A_1609_368#_c_1128_n 0.0192574f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_677 N_A_372_365#_c_890_n N_A_1609_368#_c_1128_n 0.00653851f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_A_372_365#_c_903_n N_A_1609_368#_c_1128_n 0.0030665f $X=8.88 $Y=1.665
+ $X2=0 $Y2=0
cc_679 N_A_372_365#_c_894_n N_A_1609_368#_c_1128_n 0.0023552f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_680 N_A_372_365#_c_895_n N_A_1609_368#_c_1128_n 0.0103938f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_681 N_A_372_365#_M1007_g N_A_1609_368#_c_1129_n 7.38955e-19 $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_682 N_A_372_365#_M1026_g N_A_1609_368#_c_1119_n 0.00161935f $X=8.645 $Y=0.79
+ $X2=0 $Y2=0
cc_683 N_A_372_365#_M1007_g N_A_1609_368#_c_1119_n 0.0131535f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_684 N_A_372_365#_c_890_n N_A_1609_368#_c_1119_n 0.0258452f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_685 N_A_372_365#_c_903_n N_A_1609_368#_c_1119_n 4.11576e-19 $X=8.88 $Y=1.665
+ $X2=0 $Y2=0
cc_686 N_A_372_365#_c_894_n N_A_1609_368#_c_1119_n 0.00286059f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_687 N_A_372_365#_c_895_n N_A_1609_368#_c_1119_n 0.035259f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_688 N_A_372_365#_c_890_n N_A_1609_368#_c_1120_n 0.00656895f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_689 N_A_372_365#_c_894_n N_A_1609_368#_c_1120_n 0.00173321f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_690 N_A_372_365#_M1026_g N_A_1744_94#_c_1233_n 0.00369877f $X=8.645 $Y=0.79
+ $X2=0 $Y2=0
cc_691 N_A_372_365#_c_887_n N_A_1744_94#_c_1233_n 0.0117677f $X=8.96 $Y=1.555
+ $X2=0 $Y2=0
cc_692 N_A_372_365#_c_903_n N_A_1744_94#_c_1233_n 0.00343619f $X=8.88 $Y=1.665
+ $X2=0 $Y2=0
cc_693 N_A_372_365#_c_894_n N_A_1744_94#_c_1233_n 0.0016731f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_694 N_A_372_365#_c_895_n N_A_1744_94#_c_1233_n 0.0126247f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_695 N_A_372_365#_M1026_g N_A_1744_94#_c_1234_n 0.00485843f $X=8.645 $Y=0.79
+ $X2=0 $Y2=0
cc_696 N_A_372_365#_M1026_g N_A_1744_94#_c_1236_n 0.00142168f $X=8.645 $Y=0.79
+ $X2=0 $Y2=0
cc_697 N_A_372_365#_M1007_g N_A_1744_94#_c_1243_n 0.0134554f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_698 N_A_372_365#_c_887_n N_A_1744_94#_c_1238_n 0.00360836f $X=8.96 $Y=1.555
+ $X2=0 $Y2=0
cc_699 N_A_372_365#_M1007_g N_A_1744_94#_c_1238_n 0.00493291f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_700 N_A_372_365#_c_903_n N_A_1744_94#_c_1238_n 0.00665675f $X=8.88 $Y=1.665
+ $X2=0 $Y2=0
cc_701 N_A_372_365#_c_894_n N_A_1744_94#_c_1238_n 8.74882e-19 $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_702 N_A_372_365#_c_895_n N_A_1744_94#_c_1238_n 0.0204939f $X=8.64 $Y=1.465
+ $X2=0 $Y2=0
cc_703 N_A_372_365#_c_889_n N_VPWR_c_1342_n 0.0103196f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_704 N_A_372_365#_c_890_n N_VPWR_c_1343_n 0.00553999f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_705 N_A_372_365#_M1023_g N_VPWR_c_1345_n 0.00680602f $X=6.23 $Y=2.525 $X2=0
+ $Y2=0
cc_706 N_A_372_365#_M1023_g N_VPWR_c_1340_n 0.00649272f $X=6.23 $Y=2.525 $X2=0
+ $Y2=0
cc_707 N_A_372_365#_c_889_n N_A_244_368#_c_1435_n 0.0458738f $X=6.335 $Y=1.665
+ $X2=0 $Y2=0
cc_708 N_A_372_365#_c_909_n N_A_244_368#_c_1435_n 6.46573e-19 $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_709 N_A_372_365#_c_896_n N_A_244_368#_c_1435_n 0.0913345f $X=3.11 $Y=0.81
+ $X2=0 $Y2=0
cc_710 N_A_372_365#_M1016_g N_A_1026_389#_c_1502_n 0.00269094f $X=6.215 $Y=0.69
+ $X2=0 $Y2=0
cc_711 N_A_372_365#_M1016_g N_A_1026_389#_c_1528_n 0.00257634f $X=6.215 $Y=0.69
+ $X2=0 $Y2=0
cc_712 N_A_372_365#_c_889_n N_A_1026_389#_c_1506_n 0.00698626f $X=6.335 $Y=1.665
+ $X2=0 $Y2=0
cc_713 N_A_372_365#_c_889_n N_A_1026_389#_c_1503_n 0.0200487f $X=6.335 $Y=1.665
+ $X2=0 $Y2=0
cc_714 N_A_372_365#_c_889_n N_A_1026_389#_c_1504_n 0.00407768f $X=6.335 $Y=1.665
+ $X2=0 $Y2=0
cc_715 N_A_372_365#_M1023_g N_COUT_N_c_1560_n 0.00544982f $X=6.23 $Y=2.525 $X2=0
+ $Y2=0
cc_716 N_A_372_365#_c_889_n N_COUT_N_c_1560_n 0.00763395f $X=6.335 $Y=1.665
+ $X2=0 $Y2=0
cc_717 N_A_372_365#_M1016_g N_COUT_N_c_1557_n 0.00576186f $X=6.215 $Y=0.69 $X2=0
+ $Y2=0
cc_718 N_A_372_365#_M1023_g N_COUT_N_c_1557_n 0.0106219f $X=6.23 $Y=2.525 $X2=0
+ $Y2=0
cc_719 N_A_372_365#_c_889_n N_COUT_N_c_1557_n 0.0169335f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_720 N_A_372_365#_c_891_n N_COUT_N_c_1557_n 0.00221145f $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_721 N_A_372_365#_c_892_n N_COUT_N_c_1557_n 0.0215117f $X=6.48 $Y=1.665 $X2=0
+ $Y2=0
cc_722 N_A_372_365#_c_893_n N_COUT_N_c_1557_n 0.00697578f $X=6.445 $Y=1.715
+ $X2=0 $Y2=0
cc_723 N_A_372_365#_M1016_g N_COUT_N_c_1558_n 0.0124216f $X=6.215 $Y=0.69 $X2=0
+ $Y2=0
cc_724 N_A_372_365#_c_889_n N_COUT_N_c_1558_n 0.00627834f $X=6.335 $Y=1.665
+ $X2=0 $Y2=0
cc_725 N_A_372_365#_c_890_n N_COUT_N_c_1558_n 0.00106401f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_726 N_A_372_365#_c_891_n N_COUT_N_c_1558_n 0.00204168f $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_727 N_A_372_365#_c_892_n N_COUT_N_c_1558_n 0.016714f $X=6.48 $Y=1.665 $X2=0
+ $Y2=0
cc_728 N_A_372_365#_c_893_n N_COUT_N_c_1558_n 0.00401651f $X=6.445 $Y=1.715
+ $X2=0 $Y2=0
cc_729 N_A_372_365#_M1016_g COUT_N 0.00394959f $X=6.215 $Y=0.69 $X2=0 $Y2=0
cc_730 N_A_372_365#_M1023_g N_A_1264_421#_c_1614_n 0.00448296f $X=6.23 $Y=2.525
+ $X2=0 $Y2=0
cc_731 N_A_372_365#_c_890_n N_A_1264_421#_c_1614_n 0.0183685f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_732 N_A_372_365#_c_891_n N_A_1264_421#_c_1614_n 0.0025169f $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_733 N_A_372_365#_c_892_n N_A_1264_421#_c_1614_n 0.0172606f $X=6.48 $Y=1.665
+ $X2=0 $Y2=0
cc_734 N_A_372_365#_c_893_n N_A_1264_421#_c_1614_n 0.00203204f $X=6.445 $Y=1.715
+ $X2=0 $Y2=0
cc_735 N_A_372_365#_c_890_n N_A_1264_421#_c_1613_n 0.0257367f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_736 N_A_372_365#_c_893_n N_A_1264_421#_c_1613_n 0.0018314f $X=6.445 $Y=1.715
+ $X2=0 $Y2=0
cc_737 N_A_372_365#_M1007_g N_A_1719_368#_c_1660_n 0.00590997f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_738 N_A_372_365#_M1007_g N_A_1719_368#_c_1663_n 0.00570581f $X=9.05 $Y=2.26
+ $X2=0 $Y2=0
cc_739 N_A_372_365#_M1016_g N_VGND_c_1759_n 0.00450499f $X=6.215 $Y=0.69 $X2=0
+ $Y2=0
cc_740 N_A_372_365#_M1026_g N_VGND_c_1760_n 0.00507111f $X=8.645 $Y=0.79 $X2=0
+ $Y2=0
cc_741 N_A_372_365#_M1016_g N_VGND_c_1762_n 0.00880111f $X=6.215 $Y=0.69 $X2=0
+ $Y2=0
cc_742 N_A_372_365#_M1026_g N_VGND_c_1762_n 0.00514438f $X=8.645 $Y=0.79 $X2=0
+ $Y2=0
cc_743 N_CI_M1006_g N_A_1609_368#_c_1125_n 0.00449487f $X=7.955 $Y=2.4 $X2=0
+ $Y2=0
cc_744 N_CI_c_1058_n N_A_1609_368#_c_1126_n 4.55672e-19 $X=7.45 $Y=1.88 $X2=0
+ $Y2=0
cc_745 N_CI_M1006_g N_A_1609_368#_c_1126_n 0.00337674f $X=7.955 $Y=2.4 $X2=0
+ $Y2=0
cc_746 N_CI_c_1057_n N_A_1609_368#_c_1126_n 0.00482584f $X=7.955 $Y=1.46 $X2=0
+ $Y2=0
cc_747 N_CI_M1006_g N_A_1609_368#_c_1127_n 0.00703369f $X=7.955 $Y=2.4 $X2=0
+ $Y2=0
cc_748 N_CI_M1025_g N_A_1609_368#_c_1118_n 0.0010225f $X=7.625 $Y=0.69 $X2=0
+ $Y2=0
cc_749 N_CI_c_1054_n N_A_1609_368#_c_1118_n 0.0077333f $X=8.135 $Y=1.22 $X2=0
+ $Y2=0
cc_750 N_CI_c_1054_n N_A_1609_368#_c_1119_n 0.00212997f $X=8.135 $Y=1.22 $X2=0
+ $Y2=0
cc_751 CI N_A_1609_368#_c_1119_n 0.0272258f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_752 N_CI_c_1057_n N_A_1609_368#_c_1119_n 0.0140906f $X=7.955 $Y=1.46 $X2=0
+ $Y2=0
cc_753 N_CI_M1006_g N_A_1609_368#_c_1176_n 0.00204464f $X=7.955 $Y=2.4 $X2=0
+ $Y2=0
cc_754 N_CI_c_1054_n N_A_1609_368#_c_1120_n 0.00309864f $X=8.135 $Y=1.22 $X2=0
+ $Y2=0
cc_755 N_CI_c_1054_n N_A_1744_94#_c_1236_n 0.00233599f $X=8.135 $Y=1.22 $X2=0
+ $Y2=0
cc_756 N_CI_c_1058_n N_VPWR_c_1343_n 0.00545554f $X=7.45 $Y=1.88 $X2=0 $Y2=0
cc_757 N_CI_M1006_g N_VPWR_c_1343_n 0.00287385f $X=7.955 $Y=2.4 $X2=0 $Y2=0
cc_758 CI N_VPWR_c_1343_n 0.00303328f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_759 N_CI_c_1057_n N_VPWR_c_1343_n 0.00184526f $X=7.955 $Y=1.46 $X2=0 $Y2=0
cc_760 N_CI_c_1058_n N_VPWR_c_1345_n 0.00424497f $X=7.45 $Y=1.88 $X2=0 $Y2=0
cc_761 N_CI_M1006_g N_VPWR_c_1348_n 0.005209f $X=7.955 $Y=2.4 $X2=0 $Y2=0
cc_762 N_CI_c_1058_n N_VPWR_c_1340_n 0.00674361f $X=7.45 $Y=1.88 $X2=0 $Y2=0
cc_763 N_CI_M1006_g N_VPWR_c_1340_n 0.00987933f $X=7.955 $Y=2.4 $X2=0 $Y2=0
cc_764 N_CI_c_1058_n N_A_1264_421#_c_1614_n 0.0203825f $X=7.45 $Y=1.88 $X2=0
+ $Y2=0
cc_765 N_CI_M1025_g N_A_1264_421#_c_1612_n 0.0050722f $X=7.625 $Y=0.69 $X2=0
+ $Y2=0
cc_766 N_CI_c_1058_n N_A_1264_421#_c_1613_n 0.0100311f $X=7.45 $Y=1.88 $X2=0
+ $Y2=0
cc_767 N_CI_M1025_g N_A_1264_421#_c_1613_n 0.0068341f $X=7.625 $Y=0.69 $X2=0
+ $Y2=0
cc_768 N_CI_c_1055_n N_A_1264_421#_c_1613_n 0.00709366f $X=7.45 $Y=1.79 $X2=0
+ $Y2=0
cc_769 CI N_A_1264_421#_c_1613_n 0.0240032f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_770 N_CI_c_1057_n N_A_1264_421#_c_1613_n 0.00937321f $X=7.955 $Y=1.46 $X2=0
+ $Y2=0
cc_771 N_CI_M1025_g N_A_1264_421#_c_1628_n 0.00188502f $X=7.625 $Y=0.69 $X2=0
+ $Y2=0
cc_772 N_CI_c_1057_n N_A_1264_421#_c_1628_n 0.00183254f $X=7.955 $Y=1.46 $X2=0
+ $Y2=0
cc_773 N_CI_M1006_g N_A_1719_368#_c_1663_n 0.0021613f $X=7.955 $Y=2.4 $X2=0
+ $Y2=0
cc_774 N_CI_M1025_g N_VGND_c_1754_n 0.00663758f $X=7.625 $Y=0.69 $X2=0 $Y2=0
cc_775 N_CI_c_1054_n N_VGND_c_1754_n 0.00496435f $X=8.135 $Y=1.22 $X2=0 $Y2=0
cc_776 CI N_VGND_c_1754_n 0.0188393f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_777 N_CI_c_1057_n N_VGND_c_1754_n 0.00126314f $X=7.955 $Y=1.46 $X2=0 $Y2=0
cc_778 N_CI_M1025_g N_VGND_c_1759_n 0.00434272f $X=7.625 $Y=0.69 $X2=0 $Y2=0
cc_779 N_CI_c_1054_n N_VGND_c_1760_n 0.00422942f $X=8.135 $Y=1.22 $X2=0 $Y2=0
cc_780 N_CI_M1025_g N_VGND_c_1762_n 0.00822896f $X=7.625 $Y=0.69 $X2=0 $Y2=0
cc_781 N_CI_c_1054_n N_VGND_c_1762_n 0.00789565f $X=8.135 $Y=1.22 $X2=0 $Y2=0
cc_782 N_A_1609_368#_c_1128_n N_A_1744_94#_M1007_d 0.00403264f $X=9.56 $Y=2.405
+ $X2=0 $Y2=0
cc_783 N_A_1609_368#_M1028_g N_A_1744_94#_M1029_g 0.0237597f $X=10.51 $Y=2.46
+ $X2=0 $Y2=0
cc_784 N_A_1609_368#_c_1123_n N_A_1744_94#_M1009_g 4.37715e-19 $X=10.12 $Y=1.425
+ $X2=0 $Y2=0
cc_785 N_A_1609_368#_c_1119_n N_A_1744_94#_c_1233_n 0.00551123f $X=8.18 $Y=1.82
+ $X2=0 $Y2=0
cc_786 N_A_1609_368#_c_1120_n N_A_1744_94#_c_1233_n 0.00189708f $X=8.35 $Y=0.965
+ $X2=0 $Y2=0
cc_787 N_A_1609_368#_c_1118_n N_A_1744_94#_c_1234_n 0.00528681f $X=8.35 $Y=0.515
+ $X2=0 $Y2=0
cc_788 N_A_1609_368#_M1017_g N_A_1744_94#_c_1235_n 0.00929458f $X=10.115 $Y=0.79
+ $X2=0 $Y2=0
cc_789 N_A_1609_368#_c_1118_n N_A_1744_94#_c_1236_n 0.00493016f $X=8.35 $Y=0.515
+ $X2=0 $Y2=0
cc_790 N_A_1609_368#_M1017_g N_A_1744_94#_c_1237_n 0.00583112f $X=10.115 $Y=0.79
+ $X2=0 $Y2=0
cc_791 N_A_1609_368#_c_1123_n N_A_1744_94#_c_1288_n 4.88932e-19 $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_792 N_A_1609_368#_M1017_g N_A_1744_94#_c_1289_n 0.00670132f $X=10.115 $Y=0.79
+ $X2=0 $Y2=0
cc_793 N_A_1609_368#_c_1128_n N_A_1744_94#_c_1243_n 0.0127355f $X=9.56 $Y=2.405
+ $X2=0 $Y2=0
cc_794 N_A_1609_368#_c_1131_n N_A_1744_94#_c_1243_n 0.0121068f $X=9.725 $Y=1.985
+ $X2=0 $Y2=0
cc_795 N_A_1609_368#_c_1121_n N_A_1744_94#_c_1238_n 0.00751988f $X=9.795 $Y=1.82
+ $X2=0 $Y2=0
cc_796 N_A_1609_368#_c_1123_n N_A_1744_94#_c_1239_n 2.25827e-19 $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_797 N_A_1609_368#_c_1123_n N_A_1744_94#_c_1240_n 0.0142432f $X=10.12 $Y=1.425
+ $X2=0 $Y2=0
cc_798 N_A_1609_368#_M1017_g N_A_1744_94#_c_1241_n 0.00434028f $X=10.115 $Y=0.79
+ $X2=0 $Y2=0
cc_799 N_A_1609_368#_c_1127_n N_VPWR_c_1343_n 0.0167478f $X=8.18 $Y=2.815 $X2=0
+ $Y2=0
cc_800 N_A_1609_368#_M1028_g N_VPWR_c_1344_n 0.00279397f $X=10.51 $Y=2.46 $X2=0
+ $Y2=0
cc_801 N_A_1609_368#_M1028_g N_VPWR_c_1348_n 0.00512156f $X=10.51 $Y=2.46 $X2=0
+ $Y2=0
cc_802 N_A_1609_368#_c_1127_n N_VPWR_c_1348_n 0.014549f $X=8.18 $Y=2.815 $X2=0
+ $Y2=0
cc_803 N_A_1609_368#_M1028_g N_VPWR_c_1340_n 0.00964926f $X=10.51 $Y=2.46 $X2=0
+ $Y2=0
cc_804 N_A_1609_368#_c_1127_n N_VPWR_c_1340_n 0.0119743f $X=8.18 $Y=2.815 $X2=0
+ $Y2=0
cc_805 N_A_1609_368#_c_1128_n N_VPWR_c_1340_n 0.0101865f $X=9.56 $Y=2.405 $X2=0
+ $Y2=0
cc_806 N_A_1609_368#_c_1126_n N_A_1264_421#_c_1613_n 0.0033079f $X=8.18 $Y=1.985
+ $X2=0 $Y2=0
cc_807 N_A_1609_368#_c_1128_n N_A_1719_368#_M1007_s 0.00990766f $X=9.56 $Y=2.405
+ $X2=0 $Y2=0
cc_808 N_A_1609_368#_M1028_g N_A_1719_368#_c_1660_n 0.00424229f $X=10.51 $Y=2.46
+ $X2=0 $Y2=0
cc_809 N_A_1609_368#_c_1128_n N_A_1719_368#_c_1660_n 0.0580047f $X=9.56 $Y=2.405
+ $X2=0 $Y2=0
cc_810 N_A_1609_368#_M1017_g N_A_1719_368#_c_1682_n 0.0120317f $X=10.115 $Y=0.79
+ $X2=0 $Y2=0
cc_811 N_A_1609_368#_c_1122_n N_A_1719_368#_c_1682_n 0.0177202f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_812 N_A_1609_368#_c_1123_n N_A_1719_368#_c_1682_n 0.00546304f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_813 N_A_1609_368#_c_1122_n N_A_1719_368#_c_1671_n 0.0103693f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_814 N_A_1609_368#_c_1123_n N_A_1719_368#_c_1671_n 6.85786e-19 $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_815 N_A_1609_368#_M1028_g N_A_1719_368#_c_1661_n 0.0136432f $X=10.51 $Y=2.46
+ $X2=0 $Y2=0
cc_816 N_A_1609_368#_c_1128_n N_A_1719_368#_c_1661_n 0.0319267f $X=9.56 $Y=2.405
+ $X2=0 $Y2=0
cc_817 N_A_1609_368#_c_1131_n N_A_1719_368#_c_1661_n 0.0321339f $X=9.725
+ $Y=1.985 $X2=0 $Y2=0
cc_818 N_A_1609_368#_M1017_g N_A_1719_368#_c_1659_n 0.00522589f $X=10.115
+ $Y=0.79 $X2=0 $Y2=0
cc_819 N_A_1609_368#_M1028_g N_A_1719_368#_c_1659_n 0.00553535f $X=10.51 $Y=2.46
+ $X2=0 $Y2=0
cc_820 N_A_1609_368#_c_1121_n N_A_1719_368#_c_1659_n 0.00612666f $X=9.795
+ $Y=1.82 $X2=0 $Y2=0
cc_821 N_A_1609_368#_c_1122_n N_A_1719_368#_c_1659_n 0.0247014f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_822 N_A_1609_368#_c_1123_n N_A_1719_368#_c_1659_n 0.0083239f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_823 N_A_1609_368#_c_1127_n N_A_1719_368#_c_1663_n 0.0215742f $X=8.18 $Y=2.815
+ $X2=0 $Y2=0
cc_824 N_A_1609_368#_c_1128_n N_A_1719_368#_c_1663_n 0.0256793f $X=9.56 $Y=2.405
+ $X2=0 $Y2=0
cc_825 N_A_1609_368#_M1028_g N_A_1719_368#_c_1664_n 0.0145572f $X=10.51 $Y=2.46
+ $X2=0 $Y2=0
cc_826 N_A_1609_368#_c_1121_n N_A_1719_368#_c_1664_n 0.0143027f $X=9.795 $Y=1.82
+ $X2=0 $Y2=0
cc_827 N_A_1609_368#_c_1122_n N_A_1719_368#_c_1664_n 0.00638832f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_828 N_A_1609_368#_c_1123_n N_A_1719_368#_c_1664_n 0.00514781f $X=10.12
+ $Y=1.425 $X2=0 $Y2=0
cc_829 N_A_1609_368#_M1028_g SUM 7.72509e-19 $X=10.51 $Y=2.46 $X2=0 $Y2=0
cc_830 N_A_1609_368#_c_1118_n N_VGND_c_1754_n 0.046757f $X=8.35 $Y=0.515 $X2=0
+ $Y2=0
cc_831 N_A_1609_368#_M1017_g N_VGND_c_1760_n 7.822e-19 $X=10.115 $Y=0.79 $X2=0
+ $Y2=0
cc_832 N_A_1609_368#_c_1118_n N_VGND_c_1760_n 0.0149802f $X=8.35 $Y=0.515 $X2=0
+ $Y2=0
cc_833 N_A_1609_368#_c_1118_n N_VGND_c_1762_n 0.0123195f $X=8.35 $Y=0.515 $X2=0
+ $Y2=0
cc_834 N_A_1609_368#_M1017_g N_VGND_c_1765_n 3.82766e-19 $X=10.115 $Y=0.79 $X2=0
+ $Y2=0
cc_835 N_A_1744_94#_M1029_g N_VPWR_c_1344_n 0.00402511f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_836 N_A_1744_94#_c_1239_n N_VPWR_c_1344_n 0.00282622f $X=10.975 $Y=1.465
+ $X2=0 $Y2=0
cc_837 N_A_1744_94#_c_1240_n N_VPWR_c_1344_n 4.62134e-19 $X=10.975 $Y=1.465
+ $X2=0 $Y2=0
cc_838 N_A_1744_94#_M1029_g N_VPWR_c_1349_n 0.005209f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_839 N_A_1744_94#_M1029_g N_VPWR_c_1340_n 0.00986057f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_840 N_A_1744_94#_c_1235_n N_A_1719_368#_c_1668_n 0.0126665f $X=10.155 $Y=0.34
+ $X2=0 $Y2=0
cc_841 N_A_1744_94#_M1009_g N_A_1719_368#_c_1682_n 9.73318e-19 $X=11.025 $Y=0.74
+ $X2=0 $Y2=0
cc_842 N_A_1744_94#_c_1235_n N_A_1719_368#_c_1682_n 0.00422317f $X=10.155
+ $Y=0.34 $X2=0 $Y2=0
cc_843 N_A_1744_94#_c_1288_n N_A_1719_368#_c_1682_n 0.0232007f $X=10.81 $Y=0.665
+ $X2=0 $Y2=0
cc_844 N_A_1744_94#_c_1289_n N_A_1719_368#_c_1682_n 0.00873869f $X=10.325
+ $Y=0.665 $X2=0 $Y2=0
cc_845 N_A_1744_94#_c_1241_n N_A_1719_368#_c_1682_n 0.012984f $X=10.952 $Y=1.3
+ $X2=0 $Y2=0
cc_846 N_A_1744_94#_M1029_g N_A_1719_368#_c_1661_n 6.6228e-19 $X=11.015 $Y=2.4
+ $X2=0 $Y2=0
cc_847 N_A_1744_94#_M1029_g N_A_1719_368#_c_1659_n 0.0011097f $X=11.015 $Y=2.4
+ $X2=0 $Y2=0
cc_848 N_A_1744_94#_M1009_g N_A_1719_368#_c_1659_n 9.70728e-19 $X=11.025 $Y=0.74
+ $X2=0 $Y2=0
cc_849 N_A_1744_94#_c_1240_n N_A_1719_368#_c_1659_n 0.0022592f $X=10.975
+ $Y=1.465 $X2=0 $Y2=0
cc_850 N_A_1744_94#_c_1241_n N_A_1719_368#_c_1659_n 0.0377889f $X=10.952 $Y=1.3
+ $X2=0 $Y2=0
cc_851 N_A_1744_94#_M1029_g N_A_1719_368#_c_1664_n 0.00206752f $X=11.015 $Y=2.4
+ $X2=0 $Y2=0
cc_852 N_A_1744_94#_M1009_g N_SUM_c_1724_n 0.00206311f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_853 N_A_1744_94#_c_1241_n N_SUM_c_1725_n 0.0133045f $X=10.952 $Y=1.3 $X2=0
+ $Y2=0
cc_854 N_A_1744_94#_M1029_g SUM 0.00453261f $X=11.015 $Y=2.4 $X2=0 $Y2=0
cc_855 N_A_1744_94#_c_1239_n SUM 0.00131984f $X=10.975 $Y=1.465 $X2=0 $Y2=0
cc_856 N_A_1744_94#_c_1240_n SUM 0.00152224f $X=10.975 $Y=1.465 $X2=0 $Y2=0
cc_857 N_A_1744_94#_M1029_g SUM 0.0137399f $X=11.015 $Y=2.4 $X2=0 $Y2=0
cc_858 N_A_1744_94#_M1029_g N_SUM_c_1726_n 0.00346572f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_859 N_A_1744_94#_M1009_g N_SUM_c_1726_n 0.00244621f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_860 N_A_1744_94#_c_1239_n N_SUM_c_1726_n 0.0245253f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_861 N_A_1744_94#_c_1240_n N_SUM_c_1726_n 0.00780138f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_862 N_A_1744_94#_c_1241_n N_SUM_c_1726_n 0.0058197f $X=10.952 $Y=1.3 $X2=0
+ $Y2=0
cc_863 N_A_1744_94#_c_1237_n N_VGND_M1017_d 0.00186454f $X=10.24 $Y=0.58 $X2=0
+ $Y2=0
cc_864 N_A_1744_94#_c_1288_n N_VGND_M1017_d 0.0204921f $X=10.81 $Y=0.665 $X2=0
+ $Y2=0
cc_865 N_A_1744_94#_c_1289_n N_VGND_M1017_d 7.71978e-19 $X=10.325 $Y=0.665 $X2=0
+ $Y2=0
cc_866 N_A_1744_94#_c_1241_n N_VGND_M1017_d 0.00477971f $X=10.952 $Y=1.3 $X2=0
+ $Y2=0
cc_867 N_A_1744_94#_c_1235_n N_VGND_c_1760_n 0.0794807f $X=10.155 $Y=0.34 $X2=0
+ $Y2=0
cc_868 N_A_1744_94#_c_1236_n N_VGND_c_1760_n 0.0236566f $X=9.105 $Y=0.34 $X2=0
+ $Y2=0
cc_869 N_A_1744_94#_c_1288_n N_VGND_c_1760_n 0.00335833f $X=10.81 $Y=0.665 $X2=0
+ $Y2=0
cc_870 N_A_1744_94#_M1009_g N_VGND_c_1761_n 0.00433175f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_871 N_A_1744_94#_c_1288_n N_VGND_c_1761_n 0.00123713f $X=10.81 $Y=0.665 $X2=0
+ $Y2=0
cc_872 N_A_1744_94#_M1009_g N_VGND_c_1762_n 0.0081522f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_873 N_A_1744_94#_c_1235_n N_VGND_c_1762_n 0.0460251f $X=10.155 $Y=0.34 $X2=0
+ $Y2=0
cc_874 N_A_1744_94#_c_1236_n N_VGND_c_1762_n 0.0128296f $X=9.105 $Y=0.34 $X2=0
+ $Y2=0
cc_875 N_A_1744_94#_c_1288_n N_VGND_c_1762_n 0.00972205f $X=10.81 $Y=0.665 $X2=0
+ $Y2=0
cc_876 N_A_1744_94#_M1009_g N_VGND_c_1765_n 0.0059428f $X=11.025 $Y=0.74 $X2=0
+ $Y2=0
cc_877 N_A_1744_94#_c_1235_n N_VGND_c_1765_n 0.0139023f $X=10.155 $Y=0.34 $X2=0
+ $Y2=0
cc_878 N_A_1744_94#_c_1288_n N_VGND_c_1765_n 0.0303579f $X=10.81 $Y=0.665 $X2=0
+ $Y2=0
cc_879 N_VPWR_c_1341_n N_A_244_368#_c_1443_n 0.0331183f $X=0.82 $Y=2.115 $X2=0
+ $Y2=0
cc_880 N_VPWR_c_1347_n N_A_244_368#_c_1439_n 0.145169f $X=4.545 $Y=3.33 $X2=0
+ $Y2=0
cc_881 N_VPWR_c_1340_n N_A_244_368#_c_1439_n 0.0793314f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_882 N_VPWR_c_1341_n N_A_244_368#_c_1440_n 0.0128734f $X=0.82 $Y=2.115 $X2=0
+ $Y2=0
cc_883 N_VPWR_c_1347_n N_A_244_368#_c_1440_n 0.0236204f $X=4.545 $Y=3.33 $X2=0
+ $Y2=0
cc_884 N_VPWR_c_1340_n N_A_244_368#_c_1440_n 0.0128244f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_1345_n N_A_1026_389#_c_1505_n 0.0137192f $X=7.645 $Y=3.33 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_1340_n N_A_1026_389#_c_1505_n 0.0119797f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_887 N_VPWR_c_1342_n N_A_1026_389#_c_1506_n 0.0619636f $X=4.71 $Y=1.97 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1342_n N_A_1026_389#_c_1503_n 0.00795683f $X=4.71 $Y=1.97 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1345_n N_COUT_N_c_1560_n 0.0138039f $X=7.645 $Y=3.33 $X2=0 $Y2=0
cc_890 N_VPWR_c_1340_n N_COUT_N_c_1560_n 0.0120041f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_891 N_VPWR_c_1343_n N_A_1264_421#_c_1614_n 0.0695727f $X=7.73 $Y=2.105 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1345_n N_A_1264_421#_c_1614_n 0.047919f $X=7.645 $Y=3.33 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1340_n N_A_1264_421#_c_1614_n 0.0408851f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1343_n N_A_1264_421#_c_1613_n 0.0101458f $X=7.73 $Y=2.105 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1344_n N_A_1719_368#_c_1660_n 0.0092835f $X=10.735 $Y=2.265
+ $X2=0 $Y2=0
cc_896 N_VPWR_c_1348_n N_A_1719_368#_c_1660_n 0.0832659f $X=10.65 $Y=3.33 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1340_n N_A_1719_368#_c_1660_n 0.0572275f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1348_n N_A_1719_368#_c_1663_n 0.0184392f $X=10.65 $Y=3.33 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1340_n N_A_1719_368#_c_1663_n 0.0123276f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1344_n SUM 0.0334356f $X=10.735 $Y=2.265 $X2=0 $Y2=0
cc_901 N_VPWR_c_1349_n SUM 0.0158876f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_902 N_VPWR_c_1340_n SUM 0.0130823f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_903 N_A_1026_389#_c_1505_n N_COUT_N_c_1560_n 0.0106892f $X=5.265 $Y=2.46
+ $X2=0 $Y2=0
cc_904 N_A_1026_389#_c_1506_n N_COUT_N_c_1560_n 0.0106892f $X=5.265 $Y=2.12
+ $X2=0 $Y2=0
cc_905 N_A_1026_389#_c_1506_n N_COUT_N_c_1557_n 0.00368919f $X=5.265 $Y=2.12
+ $X2=0 $Y2=0
cc_906 N_A_1026_389#_c_1503_n N_COUT_N_c_1557_n 0.00518184f $X=5.265 $Y=1.975
+ $X2=0 $Y2=0
cc_907 N_A_1026_389#_c_1528_n N_COUT_N_c_1558_n 2.58673e-19 $X=5.985 $Y=0.555
+ $X2=0 $Y2=0
cc_908 N_A_1026_389#_c_1502_n N_VGND_c_1753_n 0.0127853f $X=5.41 $Y=1.135 $X2=0
+ $Y2=0
cc_909 N_A_1026_389#_c_1512_n N_VGND_c_1759_n 0.00527357f $X=5.495 $Y=0.515
+ $X2=0 $Y2=0
cc_910 N_A_1026_389#_c_1528_n N_VGND_c_1759_n 0.0218686f $X=5.985 $Y=0.555 $X2=0
+ $Y2=0
cc_911 N_A_1026_389#_c_1512_n N_VGND_c_1762_n 0.00594062f $X=5.495 $Y=0.515
+ $X2=0 $Y2=0
cc_912 N_A_1026_389#_c_1528_n N_VGND_c_1762_n 0.0227237f $X=5.985 $Y=0.555 $X2=0
+ $Y2=0
cc_913 N_COUT_N_c_1560_n N_A_1264_421#_c_1614_n 0.00874091f $X=5.955 $Y=2.25
+ $X2=0 $Y2=0
cc_914 COUT_N N_A_1264_421#_c_1612_n 0.0144484f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_915 COUT_N N_VGND_c_1759_n 0.0146357f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_916 COUT_N N_VGND_c_1762_n 0.0121141f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_917 N_A_1264_421#_c_1612_n N_VGND_c_1754_n 0.0249694f $X=7.41 $Y=0.515 $X2=0
+ $Y2=0
cc_918 N_A_1264_421#_c_1613_n N_VGND_c_1754_n 0.00150931f $X=7.39 $Y=2.085 $X2=0
+ $Y2=0
cc_919 N_A_1264_421#_c_1612_n N_VGND_c_1759_n 0.0145094f $X=7.41 $Y=0.515 $X2=0
+ $Y2=0
cc_920 N_A_1264_421#_c_1612_n N_VGND_c_1762_n 0.011977f $X=7.41 $Y=0.515 $X2=0
+ $Y2=0
cc_921 N_A_1719_368#_c_1661_n SUM 0.00429068f $X=10.285 $Y=2.105 $X2=0 $Y2=0
cc_922 N_A_1719_368#_c_1664_n SUM 0.00429206f $X=10.54 $Y=1.845 $X2=0 $Y2=0
cc_923 N_A_1719_368#_c_1659_n N_SUM_c_1726_n 0.00383953f $X=10.54 $Y=1.76 $X2=0
+ $Y2=0
cc_924 N_A_1719_368#_c_1664_n N_SUM_c_1726_n 2.86124e-19 $X=10.54 $Y=1.845 $X2=0
+ $Y2=0
cc_925 N_A_1719_368#_c_1682_n N_VGND_M1017_d 0.0109476f $X=10.455 $Y=1.005 $X2=0
+ $Y2=0
cc_926 N_A_1719_368#_c_1659_n N_VGND_M1017_d 5.78655e-19 $X=10.54 $Y=1.76 $X2=0
+ $Y2=0
cc_927 N_SUM_c_1724_n N_VGND_c_1761_n 0.0124046f $X=11.24 $Y=0.515 $X2=0 $Y2=0
cc_928 N_SUM_c_1724_n N_VGND_c_1762_n 0.0102675f $X=11.24 $Y=0.515 $X2=0 $Y2=0
cc_929 N_SUM_c_1724_n N_VGND_c_1765_n 0.00117784f $X=11.24 $Y=0.515 $X2=0 $Y2=0

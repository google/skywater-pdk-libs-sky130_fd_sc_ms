* File: sky130_fd_sc_ms__o21ba_2.pxi.spice
* Created: Fri Aug 28 17:55:27 2020
* 
x_PM_SKY130_FD_SC_MS__O21BA_2%B1_N N_B1_N_M1006_g N_B1_N_M1002_g B1_N
+ N_B1_N_c_75_n N_B1_N_c_76_n PM_SKY130_FD_SC_MS__O21BA_2%B1_N
x_PM_SKY130_FD_SC_MS__O21BA_2%A_177_48# N_A_177_48#_M1011_s N_A_177_48#_M1010_d
+ N_A_177_48#_M1001_g N_A_177_48#_M1004_g N_A_177_48#_M1007_g
+ N_A_177_48#_M1005_g N_A_177_48#_c_105_n N_A_177_48#_c_106_n
+ N_A_177_48#_c_113_n N_A_177_48#_c_107_n N_A_177_48#_c_108_n
+ N_A_177_48#_c_114_n N_A_177_48#_c_109_n N_A_177_48#_c_110_n
+ PM_SKY130_FD_SC_MS__O21BA_2%A_177_48#
x_PM_SKY130_FD_SC_MS__O21BA_2%A_27_74# N_A_27_74#_M1006_s N_A_27_74#_M1002_s
+ N_A_27_74#_M1011_g N_A_27_74#_M1010_g N_A_27_74#_c_204_n N_A_27_74#_c_205_n
+ N_A_27_74#_c_206_n N_A_27_74#_c_207_n N_A_27_74#_c_208_n N_A_27_74#_c_209_n
+ N_A_27_74#_c_247_n N_A_27_74#_c_210_n N_A_27_74#_c_216_n
+ PM_SKY130_FD_SC_MS__O21BA_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O21BA_2%A2 N_A2_M1003_g N_A2_M1000_g A2 N_A2_c_293_n
+ N_A2_c_294_n PM_SKY130_FD_SC_MS__O21BA_2%A2
x_PM_SKY130_FD_SC_MS__O21BA_2%A1 N_A1_c_326_n N_A1_M1009_g N_A1_c_328_n
+ N_A1_M1008_g A1 PM_SKY130_FD_SC_MS__O21BA_2%A1
x_PM_SKY130_FD_SC_MS__O21BA_2%VPWR N_VPWR_M1002_d N_VPWR_M1005_s N_VPWR_M1009_d
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n VPWR N_VPWR_c_355_n
+ N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_351_n
+ PM_SKY130_FD_SC_MS__O21BA_2%VPWR
x_PM_SKY130_FD_SC_MS__O21BA_2%X N_X_M1001_s N_X_M1004_d N_X_c_396_n N_X_c_400_n
+ X X X PM_SKY130_FD_SC_MS__O21BA_2%X
x_PM_SKY130_FD_SC_MS__O21BA_2%VGND N_VGND_M1006_d N_VGND_M1007_d N_VGND_M1003_d
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ VGND N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n PM_SKY130_FD_SC_MS__O21BA_2%VGND
x_PM_SKY130_FD_SC_MS__O21BA_2%A_487_74# N_A_487_74#_M1011_d N_A_487_74#_M1008_d
+ N_A_487_74#_c_493_n N_A_487_74#_c_487_n N_A_487_74#_c_488_n
+ PM_SKY130_FD_SC_MS__O21BA_2%A_487_74#
cc_1 VNB N_B1_N_M1006_g 0.0415411f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.645
cc_2 VNB N_B1_N_M1002_g 0.00201544f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_3 VNB N_B1_N_c_75_n 0.0037649f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_B1_N_c_76_n 0.0578343f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_5 VNB N_A_177_48#_M1001_g 0.0234736f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_177_48#_M1004_g 0.00309659f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_7 VNB N_A_177_48#_M1007_g 0.0223256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_177_48#_M1005_g 0.00161918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_177_48#_c_105_n 0.0164379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_177_48#_c_106_n 0.00911858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_177_48#_c_107_n 0.00963453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_177_48#_c_108_n 0.00364368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_177_48#_c_109_n 0.00360224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_177_48#_c_110_n 0.055852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_M1011_g 0.0270364f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A_27_74#_c_204_n 0.0292115f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.465
cc_17 VNB N_A_27_74#_c_205_n 0.0111152f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_18 VNB N_A_27_74#_c_206_n 0.0194899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_207_n 0.00436079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_208_n 0.00988676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_209_n 0.00937892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_210_n 0.00298618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1000_g 0.00641921f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_24 VNB A2 0.0138799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_c_293_n 0.0335506f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_26 VNB N_A2_c_294_n 0.0186845f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_27 VNB N_A1_c_326_n 0.0657219f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.3
cc_28 VNB N_A1_M1009_g 0.00167594f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.645
cc_29 VNB N_A1_c_328_n 0.024572f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_30 VNB A1 0.00756722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_351_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_396_n 0.00199855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.00419424f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.465
cc_35 VNB N_VGND_c_431_n 0.00562672f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_36 VNB N_VGND_c_432_n 0.0136548f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_37 VNB N_VGND_c_433_n 0.00790898f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_38 VNB N_VGND_c_434_n 0.0174338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_435_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_436_n 0.0207632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_437_n 0.0310006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_438_n 0.017961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_439_n 0.239258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_440_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_441_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_487_74#_c_487_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_487_74#_c_488_n 0.0284841f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.465
cc_48 VPB N_B1_N_M1002_g 0.0304732f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_49 VPB N_B1_N_c_75_n 0.00716464f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_50 VPB N_A_177_48#_M1004_g 0.0240047f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_51 VPB N_A_177_48#_M1005_g 0.0259305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_177_48#_c_113_n 0.0028233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_177_48#_c_114_n 0.00697016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_177_48#_c_109_n 0.0015533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_M1010_g 0.0234758f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_56 VPB N_A_27_74#_c_204_n 0.0141697f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.465
cc_57 VPB N_A_27_74#_c_205_n 0.00121388f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_58 VPB N_A_27_74#_c_209_n 0.00308003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_27_74#_c_210_n 0.00274289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_74#_c_216_n 0.0346333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A2_M1000_g 0.0230544f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_62 VPB N_A1_M1009_g 0.0294115f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.645
cc_63 VPB N_VPWR_c_352_n 0.0163777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_353_n 0.0118719f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_65 VPB N_VPWR_c_354_n 0.0614424f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_66 VPB N_VPWR_c_355_n 0.0182672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_356_n 0.0351759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_357_n 0.0274805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_358_n 0.0271519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_351_n 0.0913386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_X_c_396_n 0.00171753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_X_c_400_n 0.0022412f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_73 N_B1_N_M1006_g N_A_177_48#_M1001_g 0.0214791f $X=0.485 $Y=0.645 $X2=0
+ $Y2=0
cc_74 N_B1_N_c_76_n N_A_177_48#_M1001_g 0.0120528f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_75 N_B1_N_c_76_n N_A_177_48#_M1004_g 0.030753f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_76 N_B1_N_M1006_g N_A_27_74#_c_206_n 0.00265886f $X=0.485 $Y=0.645 $X2=0
+ $Y2=0
cc_77 N_B1_N_M1006_g N_A_27_74#_c_207_n 0.0186832f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_78 N_B1_N_c_75_n N_A_27_74#_c_207_n 0.00749401f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_79 N_B1_N_c_76_n N_A_27_74#_c_207_n 0.00183826f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_80 N_B1_N_c_75_n N_A_27_74#_c_208_n 0.0199042f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_81 N_B1_N_c_76_n N_A_27_74#_c_208_n 0.00180238f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_82 N_B1_N_M1006_g N_A_27_74#_c_209_n 0.00407925f $X=0.485 $Y=0.645 $X2=0
+ $Y2=0
cc_83 N_B1_N_c_75_n N_A_27_74#_c_209_n 0.0360322f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_84 N_B1_N_c_76_n N_A_27_74#_c_209_n 0.00644828f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_85 N_B1_N_M1002_g N_A_27_74#_c_216_n 0.0340259f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_86 N_B1_N_c_75_n N_A_27_74#_c_216_n 0.0264749f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_87 N_B1_N_c_76_n N_A_27_74#_c_216_n 0.00146545f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_88 N_B1_N_M1002_g N_VPWR_c_352_n 0.00386043f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_89 N_B1_N_M1002_g N_VPWR_c_357_n 0.0046462f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_90 N_B1_N_M1002_g N_VPWR_c_351_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_91 N_B1_N_M1006_g X 8.0174e-19 $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_92 N_B1_N_M1006_g N_VGND_c_431_n 0.0151909f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_93 N_B1_N_M1006_g N_VGND_c_434_n 0.00383152f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_94 N_B1_N_M1006_g N_VGND_c_439_n 0.00761163f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_95 N_A_177_48#_c_106_n N_A_27_74#_M1011_g 0.00159319f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_96 N_A_177_48#_c_107_n N_A_27_74#_M1011_g 0.00286806f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_97 N_A_177_48#_c_108_n N_A_27_74#_M1011_g 0.0153446f $X=2.465 $Y=1.095 $X2=0
+ $Y2=0
cc_98 N_A_177_48#_c_109_n N_A_27_74#_M1011_g 0.0084954f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_99 N_A_177_48#_c_110_n N_A_27_74#_M1011_g 7.05618e-19 $X=1.5 $Y=1.465 $X2=0
+ $Y2=0
cc_100 N_A_177_48#_M1005_g N_A_27_74#_M1010_g 0.011479f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_101 N_A_177_48#_c_113_n N_A_27_74#_M1010_g 0.0116245f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_102 N_A_177_48#_c_114_n N_A_27_74#_M1010_g 0.012907f $X=2.61 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_177_48#_c_109_n N_A_27_74#_M1010_g 0.00294828f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_104 N_A_177_48#_M1005_g N_A_27_74#_c_204_n 0.00234568f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_105 N_A_177_48#_c_105_n N_A_27_74#_c_204_n 0.00223955f $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_106 N_A_177_48#_c_107_n N_A_27_74#_c_204_n 0.00108808f $X=1.515 $Y=1.095
+ $X2=0 $Y2=0
cc_107 N_A_177_48#_c_108_n N_A_27_74#_c_204_n 0.00283481f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_108 N_A_177_48#_c_110_n N_A_27_74#_c_204_n 0.0184494f $X=1.5 $Y=1.465 $X2=0
+ $Y2=0
cc_109 N_A_177_48#_c_109_n N_A_27_74#_c_205_n 0.00968053f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_110 N_A_177_48#_M1001_g N_A_27_74#_c_207_n 0.00150892f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_111 N_A_177_48#_M1001_g N_A_27_74#_c_209_n 0.00390955f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_112 N_A_177_48#_M1004_g N_A_27_74#_c_209_n 0.00252098f $X=1.05 $Y=2.4 $X2=0
+ $Y2=0
cc_113 N_A_177_48#_M1004_g N_A_27_74#_c_247_n 0.0185679f $X=1.05 $Y=2.4 $X2=0
+ $Y2=0
cc_114 N_A_177_48#_M1005_g N_A_27_74#_c_247_n 0.0199539f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_115 N_A_177_48#_c_107_n N_A_27_74#_c_247_n 0.00558461f $X=1.515 $Y=1.095
+ $X2=0 $Y2=0
cc_116 N_A_177_48#_c_114_n N_A_27_74#_c_247_n 0.0142173f $X=2.61 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_177_48#_c_110_n N_A_27_74#_c_247_n 0.00158125f $X=1.5 $Y=1.465 $X2=0
+ $Y2=0
cc_118 N_A_177_48#_M1005_g N_A_27_74#_c_210_n 0.0102452f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_119 N_A_177_48#_c_105_n N_A_27_74#_c_210_n 0.0253755f $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_120 N_A_177_48#_c_107_n N_A_27_74#_c_210_n 0.0177787f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_121 N_A_177_48#_c_109_n N_A_27_74#_c_210_n 0.0669377f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_122 N_A_177_48#_c_110_n N_A_27_74#_c_210_n 3.50755e-19 $X=1.5 $Y=1.465 $X2=0
+ $Y2=0
cc_123 N_A_177_48#_M1004_g N_A_27_74#_c_216_n 0.00655255f $X=1.05 $Y=2.4 $X2=0
+ $Y2=0
cc_124 N_A_177_48#_c_113_n N_A2_M1000_g 0.00974686f $X=2.61 $Y=2.695 $X2=0 $Y2=0
cc_125 N_A_177_48#_c_114_n N_A2_M1000_g 0.0127939f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_177_48#_c_109_n N_A2_M1000_g 0.00540378f $X=2.577 $Y=1.82 $X2=0 $Y2=0
cc_127 N_A_177_48#_c_114_n A2 0.00311529f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_177_48#_c_109_n A2 0.0287265f $X=2.577 $Y=1.82 $X2=0 $Y2=0
cc_129 N_A_177_48#_c_114_n N_A2_c_293_n 8.5668e-19 $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_177_48#_c_108_n N_A2_c_294_n 0.00465411f $X=2.465 $Y=1.095 $X2=0
+ $Y2=0
cc_131 N_A_177_48#_c_109_n N_A2_c_294_n 0.00220497f $X=2.577 $Y=1.82 $X2=0 $Y2=0
cc_132 N_A_177_48#_c_114_n N_A1_M1009_g 0.00316501f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_177_48#_M1004_g N_VPWR_c_352_n 0.0132167f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A_177_48#_M1005_g N_VPWR_c_352_n 0.00147156f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_177_48#_c_114_n N_VPWR_c_354_n 0.0264659f $X=2.61 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_177_48#_M1004_g N_VPWR_c_355_n 0.00490827f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_177_48#_M1005_g N_VPWR_c_355_n 0.00476846f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_177_48#_c_113_n N_VPWR_c_356_n 0.00968502f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_139 N_A_177_48#_M1004_g N_VPWR_c_358_n 0.00147957f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_177_48#_M1005_g N_VPWR_c_358_n 0.0145768f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_177_48#_c_113_n N_VPWR_c_358_n 0.019579f $X=2.61 $Y=2.695 $X2=0 $Y2=0
cc_142 N_A_177_48#_M1004_g N_VPWR_c_351_n 0.00968767f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_177_48#_M1005_g N_VPWR_c_351_n 0.00938661f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_177_48#_c_113_n N_VPWR_c_351_n 0.0111457f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_145 N_A_177_48#_M1001_g N_X_c_396_n 0.00395829f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_177_48#_M1004_g N_X_c_396_n 0.00543455f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_177_48#_M1007_g N_X_c_396_n 0.00162644f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_177_48#_M1005_g N_X_c_396_n 0.00365601f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_177_48#_c_107_n N_X_c_396_n 0.0323092f $X=1.515 $Y=1.095 $X2=0 $Y2=0
cc_150 N_A_177_48#_c_110_n N_X_c_396_n 0.0119574f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_151 N_A_177_48#_M1004_g N_X_c_400_n 0.00714132f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_177_48#_M1005_g N_X_c_400_n 0.00571892f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_177_48#_c_107_n N_X_c_400_n 0.0063182f $X=1.515 $Y=1.095 $X2=0 $Y2=0
cc_154 N_A_177_48#_c_110_n N_X_c_400_n 0.0073494f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_155 N_A_177_48#_M1001_g X 0.00957449f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_177_48#_M1007_g X 0.00944938f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_177_48#_c_106_n X 0.00535741f $X=2.145 $Y=0.515 $X2=0 $Y2=0
cc_158 N_A_177_48#_M1001_g X 0.00206898f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_177_48#_M1007_g X 0.00364888f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_177_48#_c_107_n X 0.00540984f $X=1.515 $Y=1.095 $X2=0 $Y2=0
cc_161 N_A_177_48#_c_110_n X 0.0018557f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A_177_48#_c_105_n N_VGND_M1007_d 9.80805e-19 $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_163 N_A_177_48#_c_107_n N_VGND_M1007_d 0.00270316f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_164 N_A_177_48#_M1001_g N_VGND_c_431_n 0.00455916f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_165 N_A_177_48#_M1007_g N_VGND_c_432_n 0.00631755f $X=1.39 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_177_48#_c_105_n N_VGND_c_432_n 0.00672294f $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_167 N_A_177_48#_c_106_n N_VGND_c_432_n 0.0323605f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_168 N_A_177_48#_c_107_n N_VGND_c_432_n 0.0130147f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_169 N_A_177_48#_c_110_n N_VGND_c_432_n 6.72142e-19 $X=1.5 $Y=1.465 $X2=0
+ $Y2=0
cc_170 N_A_177_48#_M1001_g N_VGND_c_436_n 0.00434272f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_177_48#_M1007_g N_VGND_c_436_n 0.00434272f $X=1.39 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_177_48#_c_106_n N_VGND_c_437_n 0.0110419f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_173 N_A_177_48#_M1001_g N_VGND_c_439_n 0.00821771f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_177_48#_M1007_g N_VGND_c_439_n 0.00825283f $X=1.39 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_177_48#_c_106_n N_VGND_c_439_n 0.00915013f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_176 N_A_177_48#_c_108_n N_A_487_74#_M1011_d 0.00196876f $X=2.465 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_177 N_A_177_48#_c_106_n N_A_487_74#_c_487_n 0.0182902f $X=2.145 $Y=0.515
+ $X2=0 $Y2=0
cc_178 N_A_177_48#_c_108_n N_A_487_74#_c_487_n 0.00637434f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_179 N_A_27_74#_c_205_n N_A2_M1000_g 0.0190676f $X=2.38 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A_27_74#_c_205_n A2 2.1389e-19 $X=2.38 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A_27_74#_c_205_n N_A2_c_293_n 0.0105614f $X=2.38 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A_27_74#_M1011_g N_A2_c_294_n 0.0315537f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A_27_74#_c_209_n N_VPWR_M1002_d 0.00111052f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_27_74#_c_247_n N_VPWR_M1002_d 0.00484485f $X=1.89 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_27_74#_c_216_n N_VPWR_M1002_d 0.00525937f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_27_74#_c_247_n N_VPWR_M1005_s 0.0201185f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_187 N_A_27_74#_c_210_n N_VPWR_M1005_s 0.0152989f $X=2.055 $Y=1.515 $X2=0
+ $Y2=0
cc_188 N_A_27_74#_c_247_n N_VPWR_c_352_n 0.0101555f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_189 N_A_27_74#_c_216_n N_VPWR_c_352_n 0.0174384f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_190 N_A_27_74#_M1010_g N_VPWR_c_356_n 0.00567889f $X=2.385 $Y=2.34 $X2=0
+ $Y2=0
cc_191 N_A_27_74#_c_216_n N_VPWR_c_357_n 0.006683f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_192 N_A_27_74#_M1010_g N_VPWR_c_358_n 0.00780796f $X=2.385 $Y=2.34 $X2=0
+ $Y2=0
cc_193 N_A_27_74#_c_247_n N_VPWR_c_358_n 0.0502813f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_194 N_A_27_74#_M1010_g N_VPWR_c_351_n 0.00610055f $X=2.385 $Y=2.34 $X2=0
+ $Y2=0
cc_195 N_A_27_74#_c_216_n N_VPWR_c_351_n 0.010015f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_196 N_A_27_74#_c_247_n N_X_M1004_d 0.00745752f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_197 N_A_27_74#_c_209_n N_X_c_396_n 0.0412824f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_198 N_A_27_74#_c_209_n N_X_c_400_n 0.0081428f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_199 N_A_27_74#_c_247_n N_X_c_400_n 0.0227357f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_200 N_A_27_74#_c_210_n N_X_c_400_n 0.00927682f $X=2.055 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A_27_74#_c_216_n N_X_c_400_n 0.00838524f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_202 N_A_27_74#_c_206_n X 0.00264902f $X=0.27 $Y=0.645 $X2=0 $Y2=0
cc_203 N_A_27_74#_c_207_n X 0.0117316f $X=0.625 $Y=1.045 $X2=0 $Y2=0
cc_204 N_A_27_74#_c_207_n N_VGND_M1006_d 0.00400349f $X=0.625 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_27_74#_c_207_n N_VGND_c_431_n 0.0189182f $X=0.625 $Y=1.045 $X2=0
+ $Y2=0
cc_206 N_A_27_74#_M1011_g N_VGND_c_432_n 0.00342609f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_27_74#_c_206_n N_VGND_c_434_n 0.00750773f $X=0.27 $Y=0.645 $X2=0
+ $Y2=0
cc_208 N_A_27_74#_M1011_g N_VGND_c_437_n 0.00434272f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_27_74#_M1011_g N_VGND_c_439_n 0.00826366f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_27_74#_c_206_n N_VGND_c_439_n 0.00854988f $X=0.27 $Y=0.645 $X2=0
+ $Y2=0
cc_211 N_A_27_74#_M1011_g N_A_487_74#_c_487_n 0.0070904f $X=2.36 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A2_M1000_g N_A1_c_326_n 0.0525526f $X=2.835 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A2_c_293_n N_A1_c_326_n 0.0175387f $X=2.88 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_214 A2 N_A1_c_328_n 0.00312957f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_215 N_A2_c_294_n N_A1_c_328_n 0.0256009f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_216 A2 A1 0.0302901f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_217 N_A2_c_293_n A1 2.48878e-19 $X=2.88 $Y=1.385 $X2=0 $Y2=0
cc_218 N_A2_M1000_g N_VPWR_c_354_n 0.00368017f $X=2.835 $Y=2.34 $X2=0 $Y2=0
cc_219 N_A2_M1000_g N_VPWR_c_356_n 0.00567889f $X=2.835 $Y=2.34 $X2=0 $Y2=0
cc_220 N_A2_M1000_g N_VPWR_c_351_n 0.00610055f $X=2.835 $Y=2.34 $X2=0 $Y2=0
cc_221 N_A2_c_294_n N_VGND_c_433_n 0.00416106f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_222 N_A2_c_294_n N_VGND_c_437_n 0.00324657f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_223 N_A2_c_294_n N_VGND_c_439_n 0.00410881f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_224 A2 N_A_487_74#_c_493_n 0.0215496f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A2_c_293_n N_A_487_74#_c_493_n 8.51764e-19 $X=2.88 $Y=1.385 $X2=0 $Y2=0
cc_226 N_A2_c_294_n N_A_487_74#_c_493_n 0.0104597f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_227 A2 N_A_487_74#_c_487_n 8.53117e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A2_c_294_n N_A_487_74#_c_487_n 0.00797172f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_229 N_A2_c_294_n N_A_487_74#_c_488_n 0.00142177f $X=2.88 $Y=1.22 $X2=0 $Y2=0
cc_230 N_A1_c_326_n N_VPWR_c_354_n 0.00223706f $X=3.345 $Y=1.64 $X2=0 $Y2=0
cc_231 N_A1_M1009_g N_VPWR_c_354_n 0.0275819f $X=3.345 $Y=2.34 $X2=0 $Y2=0
cc_232 A1 N_VPWR_c_354_n 0.0196739f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_233 N_A1_M1009_g N_VPWR_c_356_n 0.00492916f $X=3.345 $Y=2.34 $X2=0 $Y2=0
cc_234 N_A1_M1009_g N_VPWR_c_351_n 0.00511769f $X=3.345 $Y=2.34 $X2=0 $Y2=0
cc_235 N_A1_c_328_n N_VGND_c_433_n 0.00416106f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_236 N_A1_c_328_n N_VGND_c_438_n 0.00324657f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_237 N_A1_c_328_n N_VGND_c_439_n 0.00414389f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_238 N_A1_c_328_n N_A_487_74#_c_493_n 0.0135231f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_239 N_A1_c_328_n N_A_487_74#_c_487_n 6.42889e-19 $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_240 N_A1_c_326_n N_A_487_74#_c_488_n 0.00195015f $X=3.345 $Y=1.64 $X2=0 $Y2=0
cc_241 N_A1_c_328_n N_A_487_74#_c_488_n 0.010732f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_242 A1 N_A_487_74#_c_488_n 0.0255896f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_243 X N_VGND_c_431_n 0.0269864f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_244 X N_VGND_c_432_n 0.0175734f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_245 X N_VGND_c_436_n 0.0144922f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_246 X N_VGND_c_439_n 0.0118826f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_247 N_VGND_M1003_d N_A_487_74#_c_493_n 0.00789873f $X=2.865 $Y=0.37 $X2=0
+ $Y2=0
cc_248 N_VGND_c_433_n N_A_487_74#_c_493_n 0.0235778f $X=3.075 $Y=0.335 $X2=0
+ $Y2=0
cc_249 N_VGND_c_437_n N_A_487_74#_c_493_n 0.00227739f $X=2.91 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_c_438_n N_A_487_74#_c_493_n 0.00227739f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_251 N_VGND_c_439_n N_A_487_74#_c_493_n 0.00966343f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_252 N_VGND_c_433_n N_A_487_74#_c_487_n 0.00641885f $X=3.075 $Y=0.335 $X2=0
+ $Y2=0
cc_253 N_VGND_c_437_n N_A_487_74#_c_487_n 0.0141563f $X=2.91 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_439_n N_A_487_74#_c_487_n 0.0117515f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_433_n N_A_487_74#_c_488_n 0.00641885f $X=3.075 $Y=0.335 $X2=0
+ $Y2=0
cc_256 N_VGND_c_438_n N_A_487_74#_c_488_n 0.0145323f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_439_n N_A_487_74#_c_488_n 0.0119861f $X=3.6 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a21oi_4.pxi.spice
* Created: Wed Sep  2 11:51:51 2020
* 
x_PM_SKY130_FD_SC_MS__A21OI_4%A2 N_A2_M1003_g N_A2_M1002_g N_A2_M1005_g
+ N_A2_M1014_g N_A2_M1007_g N_A2_M1015_g N_A2_M1008_g N_A2_M1017_g A2 A2 A2
+ N_A2_c_97_n PM_SKY130_FD_SC_MS__A21OI_4%A2
x_PM_SKY130_FD_SC_MS__A21OI_4%A1 N_A1_M1000_g N_A1_M1011_g N_A1_M1001_g
+ N_A1_M1013_g N_A1_M1010_g N_A1_M1016_g N_A1_M1012_g N_A1_M1018_g A1 A1
+ N_A1_c_182_n N_A1_c_183_n PM_SKY130_FD_SC_MS__A21OI_4%A1
x_PM_SKY130_FD_SC_MS__A21OI_4%B1 N_B1_c_269_n N_B1_M1004_g N_B1_M1006_g
+ N_B1_M1009_g N_B1_M1019_g N_B1_M1021_g N_B1_c_266_n N_B1_c_267_n N_B1_M1020_g
+ B1 B1 N_B1_c_268_n PM_SKY130_FD_SC_MS__A21OI_4%B1
x_PM_SKY130_FD_SC_MS__A21OI_4%A_69_368# N_A_69_368#_M1003_s N_A_69_368#_M1005_s
+ N_A_69_368#_M1008_s N_A_69_368#_M1013_s N_A_69_368#_M1018_s
+ N_A_69_368#_M1006_s N_A_69_368#_M1020_s N_A_69_368#_c_327_n
+ N_A_69_368#_c_328_n N_A_69_368#_c_339_n N_A_69_368#_c_329_n
+ N_A_69_368#_c_347_n N_A_69_368#_c_351_n N_A_69_368#_c_353_n
+ N_A_69_368#_c_330_n N_A_69_368#_c_361_n N_A_69_368#_c_364_n
+ N_A_69_368#_c_366_n N_A_69_368#_c_367_n N_A_69_368#_c_331_n
+ N_A_69_368#_c_332_n N_A_69_368#_c_421_p N_A_69_368#_c_333_n
+ N_A_69_368#_c_334_n N_A_69_368#_c_356_n N_A_69_368#_c_360_n
+ N_A_69_368#_c_335_n N_A_69_368#_c_336_n PM_SKY130_FD_SC_MS__A21OI_4%A_69_368#
x_PM_SKY130_FD_SC_MS__A21OI_4%VPWR N_VPWR_M1003_d N_VPWR_M1007_d N_VPWR_M1011_d
+ N_VPWR_M1016_d N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n
+ N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n
+ VPWR N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_425_n N_VPWR_c_438_n
+ N_VPWR_c_439_n PM_SKY130_FD_SC_MS__A21OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A21OI_4%Y N_Y_M1000_d N_Y_M1010_d N_Y_M1009_s N_Y_M1021_s
+ N_Y_M1004_d N_Y_M1019_d N_Y_c_521_n N_Y_c_526_n N_Y_c_509_n N_Y_c_510_n
+ N_Y_c_511_n N_Y_c_552_n N_Y_c_512_n N_Y_c_533_n N_Y_c_513_n N_Y_c_564_n Y Y Y
+ N_Y_c_541_n PM_SKY130_FD_SC_MS__A21OI_4%Y
x_PM_SKY130_FD_SC_MS__A21OI_4%A_84_74# N_A_84_74#_M1002_d N_A_84_74#_M1014_d
+ N_A_84_74#_M1017_d N_A_84_74#_M1001_s N_A_84_74#_M1012_s N_A_84_74#_c_604_n
+ N_A_84_74#_c_605_n N_A_84_74#_c_606_n N_A_84_74#_c_607_n N_A_84_74#_c_608_n
+ N_A_84_74#_c_609_n N_A_84_74#_c_610_n N_A_84_74#_c_611_n N_A_84_74#_c_612_n
+ N_A_84_74#_c_613_n N_A_84_74#_c_614_n PM_SKY130_FD_SC_MS__A21OI_4%A_84_74#
x_PM_SKY130_FD_SC_MS__A21OI_4%VGND N_VGND_M1002_s N_VGND_M1015_s N_VGND_M1009_d
+ N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n N_VGND_c_679_n N_VGND_c_680_n
+ N_VGND_c_681_n VGND N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n
+ N_VGND_c_685_n N_VGND_c_686_n PM_SKY130_FD_SC_MS__A21OI_4%VGND
cc_1 VNB N_A2_M1002_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.74
cc_2 VNB N_A2_M1014_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.74
cc_3 VNB N_A2_M1015_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=0.74
cc_4 VNB N_A2_M1017_g 0.0229394f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=0.74
cc_5 VNB A2 0.00342206f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_A2_c_97_n 0.0812974f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.515
cc_7 VNB N_A1_M1000_g 0.0222136f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.4
cc_8 VNB N_A1_M1001_g 0.0221267f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_9 VNB N_A1_M1010_g 0.022172f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.4
cc_10 VNB N_A1_M1012_g 0.030436f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.4
cc_11 VNB N_A1_c_182_n 0.0024641f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.515
cc_12 VNB N_A1_c_183_n 0.0709613f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.515
cc_13 VNB N_B1_M1009_g 0.0301827f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_14 VNB N_B1_M1021_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.4
cc_15 VNB N_B1_c_266_n 0.0299697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_267_n 0.0634446f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.35
cc_17 VNB N_B1_c_268_n 0.0024641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_425_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_509_n 0.0309489f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.35
cc_20 VNB N_Y_c_510_n 0.00857879f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.35
cc_21 VNB N_Y_c_511_n 0.0138829f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=0.74
cc_22 VNB N_Y_c_512_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.515
cc_23 VNB N_Y_c_513_n 0.00215725f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_24 VNB Y 9.59717e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.515
cc_25 VNB Y 0.00160528f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.515
cc_26 VNB N_A_84_74#_c_604_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.4
cc_27 VNB N_A_84_74#_c_605_n 0.00326872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_84_74#_c_606_n 0.0126777f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.35
cc_29 VNB N_A_84_74#_c_607_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_84_74#_c_608_n 0.00766679f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.4
cc_31 VNB N_A_84_74#_c_609_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_84_74#_c_610_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_33 VNB N_A_84_74#_c_611_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_34 VNB N_A_84_74#_c_612_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_84_74#_c_613_n 0.00202435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_84_74#_c_614_n 0.00757932f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_37 VNB N_VGND_c_676_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_677_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=0.74
cc_39 VNB N_VGND_c_678_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.4
cc_40 VNB N_VGND_c_679_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=0.74
cc_41 VNB N_VGND_c_680_n 0.0258237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_681_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.68
cc_43 VNB N_VGND_c_682_n 0.068654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_683_n 0.0344157f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_45 VNB N_VGND_c_684_n 0.383272f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_46 VNB N_VGND_c_685_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.515
cc_47 VNB N_VGND_c_686_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.515
cc_48 VPB N_A2_M1003_g 0.0281481f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.4
cc_49 VPB N_A2_M1005_g 0.0204973f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.4
cc_50 VPB N_A2_M1007_g 0.020498f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=2.4
cc_51 VPB N_A2_M1008_g 0.0208043f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=2.4
cc_52 VPB A2 0.00967578f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_53 VPB N_A2_c_97_n 0.0123252f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.515
cc_54 VPB N_A1_M1011_g 0.0205244f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.74
cc_55 VPB N_A1_M1013_g 0.0208653f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.74
cc_56 VPB N_A1_M1016_g 0.0204965f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_57 VPB N_A1_M1018_g 0.0202515f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=0.74
cc_58 VPB N_A1_c_182_n 0.00596833f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.515
cc_59 VPB N_A1_c_183_n 0.0115952f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.515
cc_60 VPB N_B1_c_269_n 0.0157927f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.68
cc_61 VPB N_B1_M1006_g 0.0196385f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.74
cc_62 VPB N_B1_M1019_g 0.0200484f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.74
cc_63 VPB N_B1_c_266_n 0.00419796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B1_c_267_n 0.0132117f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.35
cc_65 VPB N_B1_M1020_g 0.0270635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_B1_c_268_n 0.00519532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_69_368#_c_327_n 0.018312f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_68 VPB N_A_69_368#_c_328_n 0.0345796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_69_368#_c_329_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=0.74
cc_70 VPB N_A_69_368#_c_330_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_69_368#_c_331_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.515
cc_72 VPB N_A_69_368#_c_332_n 0.00160153f $X=-0.19 $Y=1.66 $X2=1.97 $Y2=1.515
cc_73 VPB N_A_69_368#_c_333_n 0.0119556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_69_368#_c_334_n 0.0510465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_69_368#_c_335_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_69_368#_c_336_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_426_n 0.00554449f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=0.74
cc_78 VPB N_VPWR_c_427_n 0.00732691f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=2.4
cc_79 VPB N_VPWR_c_428_n 0.0049754f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=0.74
cc_80 VPB N_VPWR_c_429_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.68
cc_81 VPB N_VPWR_c_430_n 0.00768031f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.35
cc_82 VPB N_VPWR_c_431_n 0.0240735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_432_n 0.00458862f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_84 VPB N_VPWR_c_433_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_85 VPB N_VPWR_c_434_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_435_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.515
cc_87 VPB N_VPWR_c_436_n 0.0621381f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.565
cc_88 VPB N_VPWR_c_425_n 0.0911957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_438_n 0.00458862f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_90 VPB N_VPWR_c_439_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.565
cc_91 VPB Y 0.00116532f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.515
cc_92 N_A2_M1017_g N_A1_M1000_g 0.0179032f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A2_M1008_g N_A1_M1011_g 0.0163093f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_94 A2 N_A1_c_183_n 0.00401772f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A2_c_97_n N_A1_c_183_n 0.0163093f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A2_M1003_g N_A_69_368#_c_327_n 8.13654e-19 $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A2_M1003_g N_A_69_368#_c_328_n 0.00147311f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A2_M1003_g N_A_69_368#_c_339_n 0.0195837f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A2_M1005_g N_A_69_368#_c_339_n 0.012931f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_100 A2 N_A_69_368#_c_339_n 0.0282763f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A2_c_97_n N_A_69_368#_c_339_n 4.8724e-19 $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A2_M1003_g N_A_69_368#_c_329_n 6.74232e-19 $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A2_M1005_g N_A_69_368#_c_329_n 0.0121366f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A2_M1007_g N_A_69_368#_c_329_n 0.0119382f $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A2_M1008_g N_A_69_368#_c_329_n 6.50516e-19 $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A2_M1007_g N_A_69_368#_c_347_n 0.0128923f $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A2_M1008_g N_A_69_368#_c_347_n 0.012931f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_108 A2 N_A_69_368#_c_347_n 0.0391869f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A2_c_97_n N_A_69_368#_c_347_n 4.90062e-19 $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A2_M1008_g N_A_69_368#_c_351_n 8.84614e-19 $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_111 A2 N_A_69_368#_c_351_n 0.0122167f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A2_M1007_g N_A_69_368#_c_353_n 4.32482e-19 $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A2_M1008_g N_A_69_368#_c_353_n 0.00321805f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A2_M1008_g N_A_69_368#_c_330_n 0.00661618f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A2_M1005_g N_A_69_368#_c_356_n 8.84614e-19 $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A2_M1007_g N_A_69_368#_c_356_n 8.84614e-19 $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_117 A2 N_A_69_368#_c_356_n 0.0235495f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A2_c_97_n N_A_69_368#_c_356_n 5.52655e-19 $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A2_M1008_g N_A_69_368#_c_360_n 0.0020266f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A2_M1003_g N_VPWR_c_426_n 0.0153844f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A2_M1005_g N_VPWR_c_426_n 0.002979f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A2_M1007_g N_VPWR_c_427_n 0.0027763f $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A2_M1008_g N_VPWR_c_427_n 0.00156821f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A2_M1008_g N_VPWR_c_428_n 4.53839e-19 $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A2_M1003_g N_VPWR_c_431_n 0.00460063f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A2_M1005_g N_VPWR_c_433_n 0.005209f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A2_M1007_g N_VPWR_c_433_n 0.005209f $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A2_M1008_g N_VPWR_c_435_n 0.005209f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A2_M1003_g N_VPWR_c_425_n 0.00912799f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A2_M1005_g N_VPWR_c_425_n 0.00982266f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A2_M1007_g N_VPWR_c_425_n 0.00982266f $X=1.595 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A2_M1008_g N_VPWR_c_425_n 0.00982376f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A2_M1008_g Y 7.95334e-19 $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A2_M1017_g Y 8.33311e-19 $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_135 A2 Y 0.026396f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A2_c_97_n Y 3.70081e-19 $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A2_M1002_g N_A_84_74#_c_604_n 0.00159319f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A2_M1002_g N_A_84_74#_c_605_n 0.0167076f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A2_M1014_g N_A_84_74#_c_605_n 0.0130918f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_140 A2 N_A_84_74#_c_605_n 0.0402557f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A2_c_97_n N_A_84_74#_c_605_n 0.00474395f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A2_c_97_n N_A_84_74#_c_606_n 0.00120964f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A2_M1014_g N_A_84_74#_c_607_n 3.92313e-19 $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A2_M1015_g N_A_84_74#_c_607_n 3.92313e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_M1015_g N_A_84_74#_c_608_n 0.0130453f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1017_g N_A_84_74#_c_608_n 0.0128967f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_147 A2 N_A_84_74#_c_608_n 0.0604918f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_97_n N_A_84_74#_c_608_n 0.00258446f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A2_M1017_g N_A_84_74#_c_610_n 9.48753e-19 $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_150 A2 N_A_84_74#_c_612_n 0.0146029f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A2_c_97_n N_A_84_74#_c_612_n 0.00248733f $X=2.05 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A2_M1002_g N_VGND_c_676_n 0.0133724f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A2_M1014_g N_VGND_c_676_n 0.0103289f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1015_g N_VGND_c_676_n 4.71636e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1014_g N_VGND_c_677_n 0.00383152f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1015_g N_VGND_c_677_n 0.00383152f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_M1014_g N_VGND_c_678_n 4.71636e-19 $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1015_g N_VGND_c_678_n 0.0103289f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1017_g N_VGND_c_678_n 0.00968343f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1002_g N_VGND_c_680_n 0.00383152f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A2_M1017_g N_VGND_c_682_n 0.00383152f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A2_M1002_g N_VGND_c_684_n 0.00761822f $X=0.76 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A2_M1014_g N_VGND_c_684_n 0.0075754f $X=1.19 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A2_M1015_g N_VGND_c_684_n 0.0075754f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A2_M1017_g N_VGND_c_684_n 0.00757637f $X=2.05 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1018_g N_B1_c_267_n 0.0346225f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A1_c_182_n N_B1_c_267_n 7.56125e-19 $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A1_c_183_n N_B1_c_267_n 0.0138408f $X=3.845 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A1_c_182_n N_B1_c_268_n 0.0228558f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A1_c_183_n N_B1_c_268_n 4.14832e-19 $X=3.845 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A1_M1011_g N_A_69_368#_c_361_n 0.0176379f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A1_M1013_g N_A_69_368#_c_361_n 0.012696f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_c_183_n N_A_69_368#_c_361_n 2.53686e-19 $X=3.845 $Y=1.515 $X2=0
+ $Y2=0
cc_174 N_A1_M1016_g N_A_69_368#_c_364_n 0.0126573f $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A1_M1018_g N_A_69_368#_c_364_n 0.012696f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A1_M1018_g N_A_69_368#_c_366_n 8.84614e-19 $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A1_M1016_g N_A_69_368#_c_367_n 5.41755e-19 $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A1_M1018_g N_A_69_368#_c_367_n 0.00649085f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A1_M1018_g N_A_69_368#_c_332_n 0.00347836f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A1_M1011_g N_A_69_368#_c_335_n 5.87944e-19 $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A1_M1013_g N_A_69_368#_c_335_n 0.0089696f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A1_M1016_g N_A_69_368#_c_335_n 0.00877121f $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A1_M1018_g N_A_69_368#_c_335_n 5.64228e-19 $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A1_M1011_g N_VPWR_c_428_n 0.00850642f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_M1013_g N_VPWR_c_428_n 0.002979f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1013_g N_VPWR_c_429_n 0.005209f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1016_g N_VPWR_c_429_n 0.005209f $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_M1016_g N_VPWR_c_430_n 0.0027763f $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A1_M1018_g N_VPWR_c_430_n 0.00120619f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A1_M1011_g N_VPWR_c_435_n 0.00460063f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A1_M1018_g N_VPWR_c_436_n 0.00517089f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A1_M1011_g N_VPWR_c_425_n 0.00908665f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A1_M1013_g N_VPWR_c_425_n 0.00982266f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A1_M1016_g N_VPWR_c_425_n 0.00982266f $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A1_M1018_g N_VPWR_c_425_n 0.00977588f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A1_M1013_g N_Y_c_521_n 0.0138002f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A1_M1016_g N_Y_c_521_n 0.0116623f $X=3.395 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A1_M1018_g N_Y_c_521_n 0.0116236f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A1_c_182_n N_Y_c_521_n 0.0690241f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A1_c_183_n N_Y_c_521_n 0.0013318f $X=3.845 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A1_M1011_g N_Y_c_526_n 0.00509562f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A1_M1001_g N_Y_c_509_n 0.0176537f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A1_M1010_g N_Y_c_509_n 0.0139916f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_M1012_g N_Y_c_509_n 0.0176112f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_c_182_n N_Y_c_509_n 0.0794462f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A1_c_183_n N_Y_c_509_n 0.00741821f $X=3.845 $Y=1.515 $X2=0 $Y2=0
cc_207 N_A1_M1012_g N_Y_c_510_n 0.00455139f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1018_g N_Y_c_533_n 7.42905e-19 $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_M1000_g Y 0.00466718f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A1_M1000_g Y 0.00447162f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A1_M1011_g Y 0.00706146f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_M1001_g Y 0.00414079f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A1_M1013_g Y 0.00471932f $X=2.945 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A1_c_182_n Y 0.0336392f $X=3.77 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A1_c_183_n Y 0.019001f $X=3.845 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A1_M1000_g N_Y_c_541_n 0.0040538f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_M1000_g N_A_84_74#_c_608_n 5.67309e-19 $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1000_g N_A_84_74#_c_609_n 0.0118512f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_M1001_g N_A_84_74#_c_609_n 0.00799819f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_M1010_g N_A_84_74#_c_611_n 0.00804476f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_M1012_g N_A_84_74#_c_611_n 0.00807644f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1000_g N_A_84_74#_c_613_n 6.64397e-19 $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1001_g N_A_84_74#_c_613_n 0.00704884f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1010_g N_A_84_74#_c_613_n 0.00766985f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_M1012_g N_A_84_74#_c_613_n 9.18514e-19 $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1010_g N_A_84_74#_c_614_n 9.18514e-19 $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1012_g N_A_84_74#_c_614_n 0.00862162f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1000_g N_VGND_c_682_n 0.00278271f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1001_g N_VGND_c_682_n 0.00279469f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1010_g N_VGND_c_682_n 0.00279469f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1012_g N_VGND_c_682_n 0.00279469f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_M1000_g N_VGND_c_684_n 0.00353526f $X=2.48 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1001_g N_VGND_c_684_n 0.00352518f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1010_g N_VGND_c_684_n 0.00352518f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1012_g N_VGND_c_684_n 0.00357517f $X=3.77 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B1_c_269_n N_A_69_368#_c_331_n 0.0139961f $X=4.295 $Y=1.77 $X2=0 $Y2=0
cc_237 N_B1_M1006_g N_A_69_368#_c_331_n 0.0140221f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B1_M1019_g N_A_69_368#_c_333_n 0.0140221f $X=5.195 $Y=2.4 $X2=0 $Y2=0
cc_239 N_B1_M1020_g N_A_69_368#_c_333_n 0.0149887f $X=5.645 $Y=2.4 $X2=0 $Y2=0
cc_240 N_B1_M1020_g N_A_69_368#_c_334_n 0.00181594f $X=5.645 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B1_c_269_n N_VPWR_c_436_n 0.00333926f $X=4.295 $Y=1.77 $X2=0 $Y2=0
cc_242 N_B1_M1006_g N_VPWR_c_436_n 0.00333926f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_243 N_B1_M1019_g N_VPWR_c_436_n 0.00333926f $X=5.195 $Y=2.4 $X2=0 $Y2=0
cc_244 N_B1_M1020_g N_VPWR_c_436_n 0.00333926f $X=5.645 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B1_c_269_n N_VPWR_c_425_n 0.00422798f $X=4.295 $Y=1.77 $X2=0 $Y2=0
cc_246 N_B1_M1006_g N_VPWR_c_425_n 0.00422687f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B1_M1019_g N_VPWR_c_425_n 0.00422687f $X=5.195 $Y=2.4 $X2=0 $Y2=0
cc_248 N_B1_M1020_g N_VPWR_c_425_n 0.00426704f $X=5.645 $Y=2.4 $X2=0 $Y2=0
cc_249 N_B1_c_269_n N_Y_c_521_n 0.0136739f $X=4.295 $Y=1.77 $X2=0 $Y2=0
cc_250 N_B1_c_268_n N_Y_c_521_n 0.00872169f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_251 N_B1_c_267_n N_Y_c_509_n 0.00532991f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_252 N_B1_c_268_n N_Y_c_509_n 0.0131745f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_253 N_B1_M1009_g N_Y_c_510_n 0.00159319f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B1_M1009_g N_Y_c_511_n 0.0139178f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B1_M1021_g N_Y_c_511_n 0.0148751f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B1_c_266_n N_Y_c_511_n 0.0112784f $X=5.555 $Y=1.605 $X2=0 $Y2=0
cc_257 N_B1_c_267_n N_Y_c_511_n 0.00380788f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_258 N_B1_c_268_n N_Y_c_511_n 0.0446327f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_259 N_B1_M1006_g N_Y_c_552_n 0.012931f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B1_M1019_g N_Y_c_552_n 0.0132059f $X=5.195 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B1_c_267_n N_Y_c_552_n 4.89356e-19 $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_262 N_B1_c_268_n N_Y_c_552_n 0.0384911f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_263 N_B1_M1021_g N_Y_c_512_n 0.00159319f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_264 N_B1_c_269_n N_Y_c_533_n 0.0105482f $X=4.295 $Y=1.77 $X2=0 $Y2=0
cc_265 N_B1_M1006_g N_Y_c_533_n 0.010564f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_266 N_B1_M1019_g N_Y_c_533_n 5.73047e-19 $X=5.195 $Y=2.4 $X2=0 $Y2=0
cc_267 N_B1_c_267_n N_Y_c_533_n 5.54777e-19 $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_268 N_B1_c_268_n N_Y_c_533_n 0.0235495f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_269 N_B1_c_267_n N_Y_c_513_n 0.00645498f $X=5.285 $Y=1.605 $X2=0 $Y2=0
cc_270 N_B1_c_268_n N_Y_c_513_n 0.0214728f $X=5.08 $Y=1.515 $X2=0 $Y2=0
cc_271 N_B1_M1006_g N_Y_c_564_n 5.73047e-19 $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_272 N_B1_M1019_g N_Y_c_564_n 0.0116492f $X=5.195 $Y=2.4 $X2=0 $Y2=0
cc_273 N_B1_c_266_n N_Y_c_564_n 0.00332381f $X=5.555 $Y=1.605 $X2=0 $Y2=0
cc_274 N_B1_M1020_g N_Y_c_564_n 0.0123791f $X=5.645 $Y=2.4 $X2=0 $Y2=0
cc_275 N_B1_M1009_g N_A_84_74#_c_614_n 0.00301154f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_276 N_B1_M1009_g N_VGND_c_679_n 0.0133724f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_277 N_B1_M1021_g N_VGND_c_679_n 0.0133724f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_278 N_B1_M1009_g N_VGND_c_682_n 0.00383152f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B1_M1021_g N_VGND_c_683_n 0.00383152f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_280 N_B1_M1009_g N_VGND_c_684_n 0.00762539f $X=4.78 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B1_M1021_g N_VGND_c_684_n 0.00762539f $X=5.21 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_69_368#_c_339_n N_VPWR_M1003_d 0.00314376f $X=1.205 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_283 N_A_69_368#_c_347_n N_VPWR_M1007_d 0.00314376f $X=2.105 $Y=2.035 $X2=0
+ $Y2=0
cc_284 N_A_69_368#_c_361_n N_VPWR_M1011_d 0.00322834f $X=3.005 $Y=2.375 $X2=0
+ $Y2=0
cc_285 N_A_69_368#_c_364_n N_VPWR_M1016_d 0.00324075f $X=3.905 $Y=2.375 $X2=0
+ $Y2=0
cc_286 N_A_69_368#_c_328_n N_VPWR_c_426_n 0.0224614f $X=0.47 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A_69_368#_c_339_n N_VPWR_c_426_n 0.0148589f $X=1.205 $Y=2.035 $X2=0
+ $Y2=0
cc_288 N_A_69_368#_c_329_n N_VPWR_c_426_n 0.0234083f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_289 N_A_69_368#_c_329_n N_VPWR_c_427_n 0.0233699f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_290 N_A_69_368#_c_347_n N_VPWR_c_427_n 0.0126919f $X=2.105 $Y=2.035 $X2=0
+ $Y2=0
cc_291 N_A_69_368#_c_330_n N_VPWR_c_427_n 0.017024f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A_69_368#_c_330_n N_VPWR_c_428_n 0.0117266f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_293 N_A_69_368#_c_361_n N_VPWR_c_428_n 0.0148589f $X=3.005 $Y=2.375 $X2=0
+ $Y2=0
cc_294 N_A_69_368#_c_335_n N_VPWR_c_428_n 0.0122069f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_295 N_A_69_368#_c_335_n N_VPWR_c_429_n 0.0144776f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_296 N_A_69_368#_c_364_n N_VPWR_c_430_n 0.0126919f $X=3.905 $Y=2.375 $X2=0
+ $Y2=0
cc_297 N_A_69_368#_c_332_n N_VPWR_c_430_n 0.0101219f $X=4.155 $Y=2.99 $X2=0
+ $Y2=0
cc_298 N_A_69_368#_c_335_n N_VPWR_c_430_n 0.0121684f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_299 N_A_69_368#_c_328_n N_VPWR_c_431_n 0.011066f $X=0.47 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A_69_368#_c_329_n N_VPWR_c_433_n 0.0144623f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_301 N_A_69_368#_c_330_n N_VPWR_c_435_n 0.0109793f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_69_368#_c_331_n N_VPWR_c_436_n 0.0459191f $X=4.885 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_69_368#_c_332_n N_VPWR_c_436_n 0.0178163f $X=4.155 $Y=2.99 $X2=0
+ $Y2=0
cc_304 N_A_69_368#_c_333_n N_VPWR_c_436_n 0.0638408f $X=5.785 $Y=2.99 $X2=0
+ $Y2=0
cc_305 N_A_69_368#_c_336_n N_VPWR_c_436_n 0.0121867f $X=4.97 $Y=2.99 $X2=0 $Y2=0
cc_306 N_A_69_368#_c_328_n N_VPWR_c_425_n 0.00915947f $X=0.47 $Y=2.4 $X2=0 $Y2=0
cc_307 N_A_69_368#_c_329_n N_VPWR_c_425_n 0.0118344f $X=1.37 $Y=2.815 $X2=0
+ $Y2=0
cc_308 N_A_69_368#_c_330_n N_VPWR_c_425_n 0.00901959f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_69_368#_c_331_n N_VPWR_c_425_n 0.0258001f $X=4.885 $Y=2.99 $X2=0
+ $Y2=0
cc_310 N_A_69_368#_c_332_n N_VPWR_c_425_n 0.00958215f $X=4.155 $Y=2.99 $X2=0
+ $Y2=0
cc_311 N_A_69_368#_c_333_n N_VPWR_c_425_n 0.0355196f $X=5.785 $Y=2.99 $X2=0
+ $Y2=0
cc_312 N_A_69_368#_c_335_n N_VPWR_c_425_n 0.0118404f $X=3.17 $Y=2.455 $X2=0
+ $Y2=0
cc_313 N_A_69_368#_c_336_n N_VPWR_c_425_n 0.00660921f $X=4.97 $Y=2.99 $X2=0
+ $Y2=0
cc_314 N_A_69_368#_c_331_n N_Y_M1004_d 0.00165831f $X=4.885 $Y=2.99 $X2=0 $Y2=0
cc_315 N_A_69_368#_c_333_n N_Y_M1019_d 0.00165831f $X=5.785 $Y=2.99 $X2=0 $Y2=0
cc_316 N_A_69_368#_M1013_s N_Y_c_521_n 0.00314376f $X=3.035 $Y=1.84 $X2=0 $Y2=0
cc_317 N_A_69_368#_M1018_s N_Y_c_521_n 0.00761058f $X=3.935 $Y=1.84 $X2=0 $Y2=0
cc_318 N_A_69_368#_c_361_n N_Y_c_521_n 0.0132201f $X=3.005 $Y=2.375 $X2=0 $Y2=0
cc_319 N_A_69_368#_c_364_n N_Y_c_521_n 0.0315971f $X=3.905 $Y=2.375 $X2=0 $Y2=0
cc_320 N_A_69_368#_c_366_n N_Y_c_521_n 0.0149351f $X=4.03 $Y=2.46 $X2=0 $Y2=0
cc_321 N_A_69_368#_c_335_n N_Y_c_521_n 0.0171986f $X=3.17 $Y=2.455 $X2=0 $Y2=0
cc_322 N_A_69_368#_c_361_n N_Y_c_526_n 0.013677f $X=3.005 $Y=2.375 $X2=0 $Y2=0
cc_323 N_A_69_368#_M1006_s N_Y_c_552_n 0.00314376f $X=4.835 $Y=1.84 $X2=0 $Y2=0
cc_324 N_A_69_368#_c_421_p N_Y_c_552_n 0.0126919f $X=4.97 $Y=2.455 $X2=0 $Y2=0
cc_325 N_A_69_368#_c_331_n N_Y_c_533_n 0.0159318f $X=4.885 $Y=2.99 $X2=0 $Y2=0
cc_326 N_A_69_368#_c_333_n N_Y_c_564_n 0.0159318f $X=5.785 $Y=2.99 $X2=0 $Y2=0
cc_327 N_A_69_368#_c_327_n N_A_84_74#_c_606_n 0.00646892f $X=0.43 $Y=2.12 $X2=0
+ $Y2=0
cc_328 N_VPWR_M1011_d N_Y_c_521_n 0.00181945f $X=2.585 $Y=1.84 $X2=0 $Y2=0
cc_329 N_VPWR_M1016_d N_Y_c_521_n 0.0031478f $X=3.485 $Y=1.84 $X2=0 $Y2=0
cc_330 N_VPWR_M1011_d N_Y_c_526_n 0.00124247f $X=2.585 $Y=1.84 $X2=0 $Y2=0
cc_331 N_VPWR_M1011_d Y 0.00126138f $X=2.585 $Y=1.84 $X2=0 $Y2=0
cc_332 N_Y_c_509_n N_A_84_74#_M1001_s 0.00179574f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_333 N_Y_c_509_n N_A_84_74#_M1012_s 0.00379734f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_334 Y N_A_84_74#_c_608_n 0.0101919f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_335 N_Y_M1000_d N_A_84_74#_c_609_n 0.00176461f $X=2.555 $Y=0.37 $X2=0 $Y2=0
cc_336 N_Y_c_509_n N_A_84_74#_c_609_n 0.00397126f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_337 N_Y_c_541_n N_A_84_74#_c_609_n 0.0146809f $X=2.652 $Y=0.88 $X2=0 $Y2=0
cc_338 N_Y_M1010_d N_A_84_74#_c_611_n 0.00285125f $X=3.415 $Y=0.37 $X2=0 $Y2=0
cc_339 N_Y_c_509_n N_A_84_74#_c_611_n 0.0140305f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_340 N_Y_c_509_n N_A_84_74#_c_613_n 0.0172179f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_341 N_Y_c_509_n N_A_84_74#_c_614_n 0.0221161f $X=4.4 $Y=1.03 $X2=0 $Y2=0
cc_342 N_Y_c_510_n N_A_84_74#_c_614_n 0.0224421f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_343 N_Y_c_511_n N_VGND_M1009_d 0.00176461f $X=5.34 $Y=1.095 $X2=0 $Y2=0
cc_344 N_Y_c_510_n N_VGND_c_679_n 0.0182902f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_345 N_Y_c_511_n N_VGND_c_679_n 0.0171619f $X=5.34 $Y=1.095 $X2=0 $Y2=0
cc_346 N_Y_c_512_n N_VGND_c_679_n 0.0182902f $X=5.425 $Y=0.515 $X2=0 $Y2=0
cc_347 N_Y_c_510_n N_VGND_c_682_n 0.011066f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_348 N_Y_c_512_n N_VGND_c_683_n 0.011066f $X=5.425 $Y=0.515 $X2=0 $Y2=0
cc_349 N_Y_c_510_n N_VGND_c_684_n 0.00915947f $X=4.565 $Y=0.515 $X2=0 $Y2=0
cc_350 N_Y_c_512_n N_VGND_c_684_n 0.00915947f $X=5.425 $Y=0.515 $X2=0 $Y2=0
cc_351 N_A_84_74#_c_605_n N_VGND_M1002_s 0.00176461f $X=1.32 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_352 N_A_84_74#_c_608_n N_VGND_M1015_s 0.00176461f $X=2.18 $Y=1.095 $X2=0
+ $Y2=0
cc_353 N_A_84_74#_c_604_n N_VGND_c_676_n 0.0182902f $X=0.545 $Y=0.515 $X2=0
+ $Y2=0
cc_354 N_A_84_74#_c_605_n N_VGND_c_676_n 0.0171619f $X=1.32 $Y=1.095 $X2=0 $Y2=0
cc_355 N_A_84_74#_c_607_n N_VGND_c_676_n 0.0182488f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_356 N_A_84_74#_c_607_n N_VGND_c_677_n 0.00749631f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_357 N_A_84_74#_c_607_n N_VGND_c_678_n 0.0182488f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_358 N_A_84_74#_c_608_n N_VGND_c_678_n 0.0171619f $X=2.18 $Y=1.095 $X2=0 $Y2=0
cc_359 N_A_84_74#_c_610_n N_VGND_c_678_n 0.0112234f $X=2.35 $Y=0.34 $X2=0 $Y2=0
cc_360 N_A_84_74#_c_604_n N_VGND_c_680_n 0.011066f $X=0.545 $Y=0.515 $X2=0 $Y2=0
cc_361 N_A_84_74#_c_609_n N_VGND_c_682_n 0.0384655f $X=2.96 $Y=0.34 $X2=0 $Y2=0
cc_362 N_A_84_74#_c_610_n N_VGND_c_682_n 0.0121867f $X=2.35 $Y=0.34 $X2=0 $Y2=0
cc_363 N_A_84_74#_c_611_n N_VGND_c_682_n 0.033414f $X=3.82 $Y=0.34 $X2=0 $Y2=0
cc_364 N_A_84_74#_c_613_n N_VGND_c_682_n 0.0226572f $X=3.125 $Y=0.34 $X2=0 $Y2=0
cc_365 N_A_84_74#_c_614_n N_VGND_c_682_n 0.0227371f $X=3.985 $Y=0.34 $X2=0 $Y2=0
cc_366 N_A_84_74#_c_604_n N_VGND_c_684_n 0.00915947f $X=0.545 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_84_74#_c_607_n N_VGND_c_684_n 0.0062048f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_368 N_A_84_74#_c_609_n N_VGND_c_684_n 0.0216792f $X=2.96 $Y=0.34 $X2=0 $Y2=0
cc_369 N_A_84_74#_c_610_n N_VGND_c_684_n 0.00660921f $X=2.35 $Y=0.34 $X2=0 $Y2=0
cc_370 N_A_84_74#_c_611_n N_VGND_c_684_n 0.0187892f $X=3.82 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_84_74#_c_613_n N_VGND_c_684_n 0.0124022f $X=3.125 $Y=0.34 $X2=0 $Y2=0
cc_372 N_A_84_74#_c_614_n N_VGND_c_684_n 0.0125119f $X=3.985 $Y=0.34 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o22a_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o22a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.300000 3.735000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.710000 1.430000 3.235000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.430000 1.875000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.430000 2.500000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.350000 0.790000 0.820000 ;
        RECT 0.535000 0.820000 0.865000 1.130000 ;
        RECT 0.635000 1.130000 0.805000 1.820000 ;
        RECT 0.635000 1.820000 0.965000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  0.085000 0.365000 1.130000 ;
      RECT 0.135000  1.820000 0.465000 3.245000 ;
      RECT 0.965000  0.085000 1.295000 0.640000 ;
      RECT 0.975000  1.300000 1.305000 1.630000 ;
      RECT 1.135000  0.880000 2.295000 1.130000 ;
      RECT 1.135000  1.130000 1.305000 1.300000 ;
      RECT 1.135000  1.630000 1.305000 1.950000 ;
      RECT 1.135000  1.950000 2.680000 2.120000 ;
      RECT 1.135000  2.290000 1.790000 3.245000 ;
      RECT 1.505000  0.350000 2.795000 0.520000 ;
      RECT 1.505000  0.520000 1.835000 0.710000 ;
      RECT 2.005000  0.800000 2.295000 0.880000 ;
      RECT 2.350000  2.120000 2.680000 2.940000 ;
      RECT 2.465000  0.520000 2.795000 0.960000 ;
      RECT 2.465000  0.960000 3.725000 1.130000 ;
      RECT 2.965000  0.085000 3.295000 0.790000 ;
      RECT 3.400000  1.950000 3.730000 3.245000 ;
      RECT 3.475000  0.350000 3.725000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_ms__o22a_2
END LIBRARY

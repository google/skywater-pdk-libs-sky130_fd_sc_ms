* File: sky130_fd_sc_ms__nand4_2.spice
* Created: Fri Aug 28 17:44:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4_2.pex.spice"
.subckt sky130_fd_sc_ms__nand4_2  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_74#_M1003_d N_D_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1369 PD=2.05 PS=1.11 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1011_d N_D_M1011_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1369 PD=1.02 PS=1.11 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_304_74#_M1008_d N_C_M1008_g N_A_27_74#_M1011_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1014 N_A_304_74#_M1008_d N_C_M1014_g N_A_27_74#_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.23225 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_515_74#_M1007_d N_B_M1007_g N_A_304_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1983 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1015 N_A_515_74#_M1015_d N_B_M1015_g N_A_304_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_515_74#_M1015_d N_A_M1001_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_A_515_74#_M1010_d N_A_M1010_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.22325 AS=0.111 PD=2.15 PS=1.04 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_D_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12 AD=0.1736
+ AS=0.3192 PD=1.43 PS=2.81 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90003.9
+ A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1002_d N_D_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.1736
+ AS=0.1736 PD=1.43 PS=1.43 NRD=6.1464 NRS=0.8668 M=1 R=6.22222 SA=90000.7
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1006_s N_C_M1000_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.1736
+ AS=0.1624 PD=1.43 PS=1.41 NRD=4.3931 NRS=2.6201 M=1 R=6.22222 SA=90001.2
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1012_d N_C_M1012_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.3528
+ AS=0.1624 PD=1.75 PS=1.41 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6 SB=90002.5
+ A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3528 PD=1.39 PS=1.75 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5 SB=90001.7
+ A=0.2016 P=2.6 MULT=1
MM1013 N_Y_M1009_d N_B_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2128 PD=1.39 PS=1.5 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.9 SB=90001.2
+ A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2128 PD=1.39 PS=1.5 NRD=0 NRS=9.6727 M=1 R=6.22222 SA=90003.5 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.336 PD=1.39 PS=2.84 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.9 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__nand4_2.pxi.spice"
*
.ends
*
*

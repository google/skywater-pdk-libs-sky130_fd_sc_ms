* File: sky130_fd_sc_ms__nand4b_1.pex.spice
* Created: Wed Sep  2 12:14:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4B_1%A_N 3 7 8 11 13
c29 13 0 1.3408e-19 $X=0.61 $Y=1.22
c30 8 0 9.94899e-20 $X=0.72 $Y=1.295
r31 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.385
+ $X2=0.61 $Y2=1.55
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.385
+ $X2=0.61 $Y2=1.22
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r34 8 12 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r35 7 13 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.7 $Y=0.835 $X2=0.7
+ $Y2=1.22
r36 3 14 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=0.64 $Y=2.26 $X2=0.64
+ $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%D 3 7 8 11 13
c33 13 0 9.94899e-20 $X=1.15 $Y=1.22
c34 8 0 1.81676e-19 $X=1.2 $Y=1.295
r35 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.385
+ $X2=1.15 $Y2=1.55
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.385
+ $X2=1.15 $Y2=1.22
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.385 $X2=1.15 $Y2=1.385
r38 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.15 $Y=1.295 $X2=1.15
+ $Y2=1.385
r39 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.24 $Y=0.74 $X2=1.24
+ $Y2=1.22
r40 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.225 $Y=2.4
+ $X2=1.225 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%C 3 6 8 11 13
c33 13 0 1.57197e-19 $X=1.69 $Y=1.22
c34 11 0 1.78939e-19 $X=1.69 $Y=1.385
c35 8 0 1.45352e-19 $X=1.68 $Y=1.295
r36 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.55
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.22
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.385 $X2=1.69 $Y2=1.385
r39 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.385
r40 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.675 $Y=2.4
+ $X2=1.675 $Y2=1.55
r41 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.63 $Y=0.74 $X2=1.63
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%B 3 6 8 11 13
c35 13 0 1.45352e-19 $X=2.23 $Y=1.22
c36 8 0 2.48945e-19 $X=2.16 $Y=1.295
r37 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.385
+ $X2=2.23 $Y2=1.55
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.385
+ $X2=2.23 $Y2=1.22
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.385 $X2=2.23 $Y2=1.385
r40 8 12 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=2.22 $Y=1.295 $X2=2.22
+ $Y2=1.385
r41 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.245 $Y=2.4
+ $X2=2.245 $Y2=1.55
r42 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.14 $Y=0.74 $X2=2.14
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%A_27_112# 1 2 9 12 19 20 23 25 26 28 29 33
+ 34 37
c73 37 0 1.39345e-19 $X=2.77 $Y=1.22
r74 34 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.385
+ $X2=2.77 $Y2=1.55
r75 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.385
+ $X2=2.77 $Y2=1.22
r76 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.385 $X2=2.77 $Y2=1.385
r77 30 33 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.65 $Y=1.385
+ $X2=2.77 $Y2=1.385
r78 28 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=0.845
+ $X2=0.65 $Y2=0.845
r79 25 26 9.3668 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.342 $Y=1.985
+ $X2=0.342 $Y2=1.82
r80 23 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=1.22
+ $X2=2.65 $Y2=1.385
r81 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.65 $Y=1.01
+ $X2=2.65 $Y2=1.22
r82 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.565 $Y=0.925
+ $X2=2.65 $Y2=1.01
r83 20 29 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=2.565 $Y=0.925
+ $X2=0.65 $Y2=0.925
r84 19 28 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.275 $Y=0.845
+ $X2=0.485 $Y2=0.845
r85 14 19 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.19 $Y=1.01
+ $X2=0.275 $Y2=0.845
r86 14 26 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.19 $Y=1.01
+ $X2=0.19 $Y2=1.82
r87 12 38 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.695 $Y=2.4
+ $X2=2.695 $Y2=1.55
r88 9 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.68 $Y=0.74 $X2=2.68
+ $Y2=1.22
r89 2 25 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.27
+ $Y=1.84 $X2=0.415 $Y2=1.985
r90 1 28 182 $w=1.7e-07 $l=4.71434e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.485 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%VPWR 1 2 3 12 18 20 22 27 28 30 31 32 41 47
c46 2 0 8.7301e-20 $X=1.765 $Y=1.84
r47 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 41 46 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=3.082 $Y2=3.33
r51 41 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 32 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 32 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 32 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 30 39 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.95 $Y2=3.33
r58 29 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.95 $Y2=3.33
r60 27 35 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.95 $Y2=3.33
r62 26 39 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.95 $Y2=3.33
r64 22 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.97 $Y=2.145
+ $X2=2.97 $Y2=2.825
r65 20 46 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=3.082 $Y2=3.33
r66 20 25 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=2.825
r67 16 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r68 16 18 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.405
r69 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.95 $Y=1.985
+ $X2=0.95 $Y2=2.815
r70 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=3.33
r71 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=2.815
r72 3 25 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=2.97 $Y2=2.825
r73 3 22 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=2.97 $Y2=2.145
r74 2 18 300 $w=1.7e-07 $l=6.50961e-07 $layer=licon1_PDIFF $count=2 $X=1.765
+ $Y=1.84 $X2=1.95 $Y2=2.405
r75 1 15 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.84 $X2=0.95 $Y2=2.815
r76 1 12 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.84 $X2=0.95 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%Y 1 2 3 10 12 16 18 22 25 29 31 32 33
c59 29 0 1.78939e-19 $X=2.285 $Y=1.935
c60 10 0 8.7301e-20 $X=1.45 $Y=2.15
r61 29 33 3.35013 $w=4.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=1.935
+ $X2=2.16 $Y2=1.935
r62 29 31 5.86152 $w=3e-07 $l=1.75e-07 $layer=LI1_cond $X=2.285 $Y=1.935
+ $X2=2.46 $Y2=1.935
r63 26 33 8.84433 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.83 $Y=1.935
+ $X2=2.16 $Y2=1.935
r64 26 28 3.19851 $w=4.3e-07 $l=2.73e-07 $layer=LI1_cond $X=1.83 $Y=1.935
+ $X2=1.557 $Y2=1.935
r65 25 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=1.72
+ $X2=3.19 $Y2=1.05
r66 20 32 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.09 $Y=0.865
+ $X2=3.09 $Y2=1.05
r67 20 22 10.9015 $w=3.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.09 $Y=0.865
+ $X2=3.09 $Y2=0.515
r68 19 31 5.86152 $w=3e-07 $l=2.3103e-07 $layer=LI1_cond $X=2.635 $Y=1.805
+ $X2=2.46 $Y2=1.935
r69 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=1.805
+ $X2=3.19 $Y2=1.72
r70 18 19 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.105 $Y=1.805
+ $X2=2.635 $Y2=1.805
r71 14 31 0.793806 $w=3.5e-07 $l=2.15e-07 $layer=LI1_cond $X=2.46 $Y=2.15
+ $X2=2.46 $Y2=1.935
r72 14 16 21.8964 $w=3.48e-07 $l=6.65e-07 $layer=LI1_cond $X=2.46 $Y=2.15
+ $X2=2.46 $Y2=2.815
r73 10 28 3.7726 $w=3.3e-07 $l=2.63116e-07 $layer=LI1_cond $X=1.45 $Y=2.15
+ $X2=1.557 $Y2=1.935
r74 10 12 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.45 $Y=2.15
+ $X2=1.45 $Y2=2.815
r75 3 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.84 $X2=2.47 $Y2=1.985
r76 3 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.84 $X2=2.47 $Y2=2.815
r77 2 28 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.45 $Y2=1.985
r78 2 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.45 $Y2=2.815
r79 1 22 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.37 $X2=2.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_1%VGND 1 6 9 10 11 21 22
r27 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r28 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r29 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r30 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r31 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r32 11 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r33 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r34 9 14 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.72
+ $Y2=0
r35 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.02
+ $Y2=0
r36 8 18 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.2
+ $Y2=0
r37 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.02
+ $Y2=0
r38 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=0.085 $X2=1.02
+ $Y2=0
r39 4 6 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.02 $Y=0.085 $X2=1.02
+ $Y2=0.55
r40 1 6 182 $w=1.7e-07 $l=2.4995e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.56 $X2=1.02 $Y2=0.55
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR D1 a_27_392# VPB pshort w=840000u l=180000u
+  ad=2.1934e+12p pd=1.825e+07u as=1.5046e+12p ps=1.239e+07u
M1001 a_287_74# C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=6.6465e+11p ps=6.59e+06u
M1002 a_27_392# A2 a_750_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1003 a_750_392# A2 a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_287_74# B1 a_477_198# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.5105e+11p ps=8.36e+06u
M1005 a_477_198# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.295e+12p ps=1.09e+07u
M1006 X a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_477_198# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# C1 a_287_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_392# D1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1011 a_27_74# D1 a_27_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_27_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B1 a_27_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A1 a_477_198# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_27_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.608e+11p ps=5.66e+06u
M1016 X a_27_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_27_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_750_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_27_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_392# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_27_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A1 a_750_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_392# D1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_392# C1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR C1 a_27_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_477_198# B1 a_287_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_477_198# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__mux2i_4.pex.spice
* Created: Wed Sep  2 12:12:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A1 3 7 11 15 19 23 27 31 33 34 35 51 53
r84 52 53 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.87 $Y2=1.515
r85 50 52 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.72 $Y=1.515
+ $X2=1.855 $Y2=1.515
r86 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.72
+ $Y=1.515 $X2=1.72 $Y2=1.515
r87 48 50 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.72 $Y2=1.515
r88 47 48 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.515
+ $X2=1.405 $Y2=1.515
r89 46 47 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=0.955 $Y=1.515
+ $X2=1.355 $Y2=1.515
r90 45 46 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.515
+ $X2=0.955 $Y2=1.515
r91 43 45 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.7 $Y=1.515
+ $X2=0.925 $Y2=1.515
r92 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.515 $X2=0.7 $Y2=1.515
r93 41 43 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.7 $Y2=1.515
r94 39 41 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.505 $Y2=1.515
r95 35 51 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.72
+ $Y2=1.565
r96 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r97 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r98 33 44 0.53602 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.7
+ $Y2=1.565
r99 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.515
r100 29 31 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.795
r101 25 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=1.515
r102 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=2.4
r103 21 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=1.515
r104 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=2.4
r105 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=1.515
r106 17 19 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=0.795
r107 13 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.515
r108 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r109 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.515
r110 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.795
r111 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r112 5 7 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.795
r113 1 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.515
r114 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A0 3 7 11 15 19 23 25 29 33 35 36 37 53
r83 52 53 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.305 $Y=1.515
+ $X2=3.395 $Y2=1.515
r84 51 52 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.275 $Y=1.515
+ $X2=3.305 $Y2=1.515
r85 49 51 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.07 $Y=1.515
+ $X2=3.275 $Y2=1.515
r86 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.515 $X2=3.07 $Y2=1.515
r87 47 49 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=2.805 $Y=1.515
+ $X2=3.07 $Y2=1.515
r88 46 47 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.8 $Y=1.515
+ $X2=2.805 $Y2=1.515
r89 45 50 10.37 $w=4e-07 $l=3.4e-07 $layer=LI1_cond $X=2.73 $Y=1.565 $X2=3.07
+ $Y2=1.565
r90 44 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.73 $Y=1.515 $X2=2.8
+ $Y2=1.515
r91 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=1.515 $X2=2.73 $Y2=1.515
r92 42 44 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.315 $Y=1.515
+ $X2=2.73 $Y2=1.515
r93 40 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.3 $Y=1.515
+ $X2=2.315 $Y2=1.515
r94 37 50 1.525 $w=4e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.07
+ $Y2=1.565
r95 36 45 2.745 $w=4e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.73
+ $Y2=1.565
r96 31 35 18.8402 $w=1.65e-07 $l=9.40744e-08 $layer=POLY_cond $X=3.805 $Y=1.5
+ $X2=3.762 $Y2=1.425
r97 31 33 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=3.805 $Y=1.5 $X2=3.805
+ $Y2=2.4
r98 27 35 18.8402 $w=1.65e-07 $l=9.94987e-08 $layer=POLY_cond $X=3.705 $Y=1.35
+ $X2=3.762 $Y2=1.425
r99 27 29 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.705 $Y=1.35
+ $X2=3.705 $Y2=0.795
r100 25 35 6.66866 $w=1.5e-07 $l=1.32e-07 $layer=POLY_cond $X=3.63 $Y=1.425
+ $X2=3.762 $Y2=1.425
r101 25 53 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.63 $Y=1.425
+ $X2=3.395 $Y2=1.425
r102 21 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.68
+ $X2=3.305 $Y2=1.515
r103 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.305 $Y=1.68
+ $X2=3.305 $Y2=2.4
r104 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.35
+ $X2=3.275 $Y2=1.515
r105 17 19 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.275 $Y=1.35
+ $X2=3.275 $Y2=0.795
r106 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.35
+ $X2=2.8 $Y2=1.515
r107 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.8 $Y=1.35
+ $X2=2.8 $Y2=0.795
r108 9 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.68
+ $X2=2.805 $Y2=1.515
r109 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.805 $Y=1.68
+ $X2=2.805 $Y2=2.4
r110 5 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.68
+ $X2=2.315 $Y2=1.515
r111 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.315 $Y=1.68
+ $X2=2.315 $Y2=2.4
r112 1 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=1.515
r113 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A_1030_268# 1 2 9 11 13 16 18 20 23 27 31 35
+ 37 42 46 48 52 55 62 63 73
r129 70 71 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=6.335 $Y=1.505
+ $X2=6.67 $Y2=1.505
r130 69 70 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.14 $Y=1.505
+ $X2=6.335 $Y2=1.505
r131 68 69 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=5.745 $Y=1.505
+ $X2=6.14 $Y2=1.505
r132 67 68 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=5.69 $Y=1.505
+ $X2=5.745 $Y2=1.505
r133 59 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.675 $Y=1.505
+ $X2=6.765 $Y2=1.505
r134 59 71 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.675 $Y=1.505
+ $X2=6.67 $Y2=1.505
r135 55 63 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.74 $Y=1.71 $X2=9.74
+ $Y2=1.01
r136 50 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.66 $Y=0.845
+ $X2=9.66 $Y2=1.01
r137 50 52 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.66 $Y=0.845
+ $X2=9.66 $Y2=0.555
r138 49 62 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.455 $Y=1.795
+ $X2=9.32 $Y2=1.795
r139 48 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.655 $Y=1.795
+ $X2=9.74 $Y2=1.71
r140 48 49 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.655 $Y=1.795
+ $X2=9.455 $Y2=1.795
r141 44 62 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.32 $Y=1.88
+ $X2=9.32 $Y2=1.795
r142 44 46 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.32 $Y=1.88
+ $X2=9.32 $Y2=1.985
r143 43 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=1.795
+ $X2=6.755 $Y2=1.795
r144 42 62 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.185 $Y=1.795
+ $X2=9.32 $Y2=1.795
r145 42 43 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=9.185 $Y=1.795
+ $X2=6.84 $Y2=1.795
r146 40 67 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.315 $Y=1.505
+ $X2=5.69 $Y2=1.505
r147 40 64 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.315 $Y=1.505
+ $X2=5.24 $Y2=1.505
r148 39 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.315
+ $Y=1.505 $X2=5.315 $Y2=1.505
r149 37 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.755 $Y=1.505
+ $X2=6.755 $Y2=1.795
r150 37 59 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.675
+ $Y=1.505 $X2=6.675 $Y2=1.505
r151 37 39 47.32 $w=3.28e-07 $l=1.355e-06 $layer=LI1_cond $X=6.67 $Y=1.505
+ $X2=5.315 $Y2=1.505
r152 33 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.34
+ $X2=6.765 $Y2=1.505
r153 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.765 $Y=1.34
+ $X2=6.765 $Y2=0.78
r154 29 71 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=1.67
+ $X2=6.67 $Y2=1.505
r155 29 31 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=6.67 $Y=1.67
+ $X2=6.67 $Y2=2.4
r156 25 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.34
+ $X2=6.335 $Y2=1.505
r157 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.335 $Y=1.34
+ $X2=6.335 $Y2=0.78
r158 21 69 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.67
+ $X2=6.14 $Y2=1.505
r159 21 23 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=6.14 $Y=1.67
+ $X2=6.14 $Y2=2.4
r160 18 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=1.505
r161 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.745 $Y=1.34
+ $X2=5.745 $Y2=0.86
r162 14 67 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.69 $Y=1.67
+ $X2=5.69 $Y2=1.505
r163 14 16 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.69 $Y=1.67
+ $X2=5.69 $Y2=2.4
r164 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.34
+ $X2=5.315 $Y2=1.505
r165 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.315 $Y=1.34
+ $X2=5.315 $Y2=0.86
r166 7 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.67
+ $X2=5.24 $Y2=1.505
r167 7 9 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.24 $Y=1.67 $X2=5.24
+ $Y2=2.4
r168 2 46 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.215
+ $Y=1.84 $X2=9.35 $Y2=1.985
r169 1 52 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.45
+ $Y=0.41 $X2=9.66 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%S 3 5 7 10 12 14 17 19 21 24 26 28 31 33 35
+ 38 40 41 42 43 44 71
c115 33 0 1.15153e-19 $X=9.375 $Y=1.26
r116 69 71 13.7714 $w=3.15e-07 $l=9e-08 $layer=POLY_cond $X=9.285 $Y=1.425
+ $X2=9.375 $Y2=1.425
r117 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.285
+ $Y=1.425 $X2=9.285 $Y2=1.425
r118 67 69 24.4825 $w=3.15e-07 $l=1.6e-07 $layer=POLY_cond $X=9.125 $Y=1.425
+ $X2=9.285 $Y2=1.425
r119 66 67 38.254 $w=3.15e-07 $l=2.5e-07 $layer=POLY_cond $X=8.875 $Y=1.425
+ $X2=9.125 $Y2=1.425
r120 65 66 39.019 $w=3.15e-07 $l=2.55e-07 $layer=POLY_cond $X=8.62 $Y=1.425
+ $X2=8.875 $Y2=1.425
r121 63 65 2.29524 $w=3.15e-07 $l=1.5e-08 $layer=POLY_cond $X=8.605 $Y=1.425
+ $X2=8.62 $Y2=1.425
r122 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.605
+ $Y=1.425 $X2=8.605 $Y2=1.425
r123 61 63 24.4825 $w=3.15e-07 $l=1.6e-07 $layer=POLY_cond $X=8.445 $Y=1.425
+ $X2=8.605 $Y2=1.425
r124 59 61 27.5429 $w=3.15e-07 $l=1.8e-07 $layer=POLY_cond $X=8.265 $Y=1.425
+ $X2=8.445 $Y2=1.425
r125 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.265
+ $Y=1.425 $X2=8.265 $Y2=1.425
r126 57 59 14.5365 $w=3.15e-07 $l=9.5e-08 $layer=POLY_cond $X=8.17 $Y=1.425
+ $X2=8.265 $Y2=1.425
r127 56 57 58.9111 $w=3.15e-07 $l=3.85e-07 $layer=POLY_cond $X=7.785 $Y=1.425
+ $X2=8.17 $Y2=1.425
r128 55 56 25.2476 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.62 $Y=1.425
+ $X2=7.785 $Y2=1.425
r129 53 55 5.35556 $w=3.15e-07 $l=3.5e-08 $layer=POLY_cond $X=7.585 $Y=1.425
+ $X2=7.62 $Y2=1.425
r130 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.585
+ $Y=1.425 $X2=7.585 $Y2=1.425
r131 51 53 35.1936 $w=3.15e-07 $l=2.3e-07 $layer=POLY_cond $X=7.355 $Y=1.425
+ $X2=7.585 $Y2=1.425
r132 50 51 28.3079 $w=3.15e-07 $l=1.85e-07 $layer=POLY_cond $X=7.17 $Y=1.425
+ $X2=7.355 $Y2=1.425
r133 44 70 2.40092 $w=3.58e-07 $l=7.5e-08 $layer=LI1_cond $X=9.36 $Y=1.36
+ $X2=9.285 $Y2=1.36
r134 43 70 12.965 $w=3.58e-07 $l=4.05e-07 $layer=LI1_cond $X=8.88 $Y=1.36
+ $X2=9.285 $Y2=1.36
r135 43 64 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=8.88 $Y=1.36
+ $X2=8.605 $Y2=1.36
r136 42 64 6.56252 $w=3.58e-07 $l=2.05e-07 $layer=LI1_cond $X=8.4 $Y=1.36
+ $X2=8.605 $Y2=1.36
r137 42 60 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=8.4 $Y=1.36
+ $X2=8.265 $Y2=1.36
r138 41 60 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=7.92 $Y=1.36
+ $X2=8.265 $Y2=1.36
r139 41 54 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=1.36
+ $X2=7.585 $Y2=1.36
r140 40 54 4.64178 $w=3.58e-07 $l=1.45e-07 $layer=LI1_cond $X=7.44 $Y=1.36
+ $X2=7.585 $Y2=1.36
r141 36 71 30.6032 $w=3.15e-07 $l=2.70185e-07 $layer=POLY_cond $X=9.575 $Y=1.59
+ $X2=9.375 $Y2=1.425
r142 36 38 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=9.575 $Y=1.59
+ $X2=9.575 $Y2=2.26
r143 33 71 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.375 $Y=1.26
+ $X2=9.375 $Y2=1.425
r144 33 35 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.375 $Y=1.26
+ $X2=9.375 $Y2=0.78
r145 29 67 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.59
+ $X2=9.125 $Y2=1.425
r146 29 31 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=9.125 $Y=1.59
+ $X2=9.125 $Y2=2.26
r147 26 66 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.875 $Y=1.26
+ $X2=8.875 $Y2=1.425
r148 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.875 $Y=1.26
+ $X2=8.875 $Y2=0.78
r149 22 65 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.62 $Y=1.59
+ $X2=8.62 $Y2=1.425
r150 22 24 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=8.62 $Y=1.59
+ $X2=8.62 $Y2=2.4
r151 19 61 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.445 $Y=1.26
+ $X2=8.445 $Y2=1.425
r152 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.445 $Y=1.26
+ $X2=8.445 $Y2=0.78
r153 15 57 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.17 $Y=1.59
+ $X2=8.17 $Y2=1.425
r154 15 17 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=8.17 $Y=1.59
+ $X2=8.17 $Y2=2.4
r155 12 56 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.785 $Y=1.26
+ $X2=7.785 $Y2=1.425
r156 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.785 $Y=1.26
+ $X2=7.785 $Y2=0.78
r157 8 55 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.62 $Y=1.59 $X2=7.62
+ $Y2=1.425
r158 8 10 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=7.62 $Y=1.59
+ $X2=7.62 $Y2=2.4
r159 5 51 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.355 $Y=1.26
+ $X2=7.355 $Y2=1.425
r160 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.355 $Y=1.26
+ $X2=7.355 $Y2=0.78
r161 1 50 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.17 $Y=1.59 $X2=7.17
+ $Y2=1.425
r162 1 3 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=7.17 $Y=1.59 $X2=7.17
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 37 39 40 41 45
+ 49 51 53 59 61 63 67 69 70 73 75 77 78 79 86 91
r121 91 92 1.37742 $w=6.2e-07 $l=7e-08 $layer=LI1_cond $X=3.865 $Y=1.965
+ $X2=3.865 $Y2=2.035
r122 86 91 5.90323 $w=6.2e-07 $l=3e-07 $layer=LI1_cond $X=3.865 $Y=1.665
+ $X2=3.865 $Y2=1.965
r123 79 82 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.08 $Y=2.035
+ $X2=3.08 $Y2=2.23
r124 70 86 9.50836 $w=6.2e-07 $l=1.83712e-07 $layer=LI1_cond $X=4 $Y=1.55
+ $X2=3.865 $Y2=1.665
r125 69 85 4.20453 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4 $Y=1.18 $X2=4
+ $Y2=1.057
r126 69 70 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4 $Y=1.18 $X2=4
+ $Y2=1.55
r127 68 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.035
+ $X2=3.08 $Y2=2.035
r128 67 92 8.52869 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.865 $Y2=2.035
r129 67 68 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.245 $Y2=2.035
r130 64 78 7.45506 $w=2.07e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=1.057
+ $X2=2.085 $Y2=1.057
r131 64 66 36.9252 $w=2.43e-07 $l=7.85e-07 $layer=LI1_cond $X=2.25 $Y=1.057
+ $X2=3.035 $Y2=1.057
r132 63 85 2.90557 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.915 $Y=1.057
+ $X2=4 $Y2=1.057
r133 63 66 41.3939 $w=2.43e-07 $l=8.8e-07 $layer=LI1_cond $X=3.915 $Y=1.057
+ $X2=3.035 $Y2=1.057
r134 62 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=2.035
+ $X2=2.08 $Y2=2.035
r135 61 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.035
+ $X2=3.08 $Y2=2.035
r136 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.915 $Y=2.035
+ $X2=2.245 $Y2=2.035
r137 57 78 0.261258 $w=3.3e-07 $l=1.22e-07 $layer=LI1_cond $X=2.085 $Y=0.935
+ $X2=2.085 $Y2=1.057
r138 57 59 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.085 $Y=0.935
+ $X2=2.085 $Y2=0.68
r139 54 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.035
+ $X2=1.18 $Y2=2.035
r140 53 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=2.035
+ $X2=2.08 $Y2=2.035
r141 53 54 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.915 $Y=2.035
+ $X2=1.265 $Y2=2.035
r142 52 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=1.095
+ $X2=1.14 $Y2=1.095
r143 51 78 7.45506 $w=2.07e-07 $l=1.83016e-07 $layer=LI1_cond $X=1.92 $Y=1.095
+ $X2=2.085 $Y2=1.057
r144 51 52 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.92 $Y=1.095
+ $X2=1.225 $Y2=1.095
r145 47 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.035
r146 47 49 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.57
r147 43 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.01
+ $X2=1.14 $Y2=1.095
r148 43 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.14 $Y=1.01
+ $X2=1.14 $Y2=0.82
r149 42 72 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=0.365 $Y=2.035
+ $X2=0.24 $Y2=1.97
r150 41 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=1.18 $Y2=2.035
r151 41 42 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=0.365 $Y2=2.035
r152 39 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=1.14 $Y2=1.095
r153 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=0.365 $Y2=1.095
r154 35 72 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=2.12 $X2=0.24
+ $Y2=1.97
r155 35 37 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=2.12
+ $X2=0.24 $Y2=2.4
r156 31 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r157 31 33 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.57
r158 10 91 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=1.84 $X2=4.08 $Y2=1.965
r159 9 82 600 $w=1.7e-07 $l=4.7355e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.84 $X2=3.08 $Y2=2.23
r160 8 77 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.035
r161 7 75 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.035
r162 7 49 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.57
r163 6 72 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r164 6 37 300 $w=1.7e-07 $l=6.28331e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.4
r165 5 85 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.425 $X2=3.92 $Y2=1.02
r166 4 66 182 $w=1.7e-07 $l=6.70242e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.425 $X2=3.035 $Y2=1.02
r167 3 59 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.425 $X2=2.085 $Y2=0.68
r168 2 45 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.425 $X2=1.14 $Y2=0.82
r169 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.425 $X2=0.28 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A_119_368# 1 2 3 4 15 17 18 21 25 27 29 32
r61 31 32 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=2.902
+ $X2=5.3 $Y2=2.902
r62 25 31 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=5.472 $Y=2.902
+ $X2=5.465 $Y2=2.902
r63 25 27 30.331 $w=3.43e-07 $l=9.08e-07 $layer=LI1_cond $X=5.472 $Y=2.902
+ $X2=6.38 $Y2=2.902
r64 24 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.715 $Y=2.99
+ $X2=1.59 $Y2=2.99
r65 24 32 233.888 $w=1.68e-07 $l=3.585e-06 $layer=LI1_cond $X=1.715 $Y=2.99
+ $X2=5.3 $Y2=2.99
r66 19 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.59 $Y2=2.99
r67 19 21 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.59 $Y2=2.455
r68 17 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=2.99
+ $X2=1.59 $Y2=2.99
r69 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.99
+ $X2=0.895 $Y2=2.99
r70 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r71 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.73 $Y2=2.415
r72 4 27 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=1.84 $X2=6.38 $Y2=2.815
r73 3 31 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.84 $X2=5.465 $Y2=2.815
r74 2 21 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.455
r75 1 15 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A_481_368# 1 2 3 4 13 15 17 21 26 31 35 40
+ 42
r73 35 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.045 $Y=2.475
+ $X2=5.045 $Y2=2.65
r74 31 33 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.58 $Y=2.455
+ $X2=3.58 $Y2=2.65
r75 26 28 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.58 $Y=2.455
+ $X2=2.58 $Y2=2.65
r76 22 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.56 $Y=2.475
+ $X2=7.395 $Y2=2.475
r77 21 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.23 $Y=2.475
+ $X2=8.395 $Y2=2.475
r78 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.23 $Y=2.475
+ $X2=7.56 $Y2=2.475
r79 18 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=2.475
+ $X2=5.045 $Y2=2.475
r80 17 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=2.475
+ $X2=7.395 $Y2=2.475
r81 17 18 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=7.23 $Y=2.475
+ $X2=5.13 $Y2=2.475
r82 16 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.65
+ $X2=3.58 $Y2=2.65
r83 15 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.65
+ $X2=5.045 $Y2=2.65
r84 15 16 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=4.96 $Y=2.65
+ $X2=3.745 $Y2=2.65
r85 14 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.65
+ $X2=2.58 $Y2=2.65
r86 13 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=2.65
+ $X2=3.58 $Y2=2.65
r87 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=2.65
+ $X2=2.745 $Y2=2.65
r88 4 42 300 $w=1.7e-07 $l=6.9925e-07 $layer=licon1_PDIFF $count=2 $X=8.26
+ $Y=1.84 $X2=8.395 $Y2=2.475
r89 3 40 300 $w=1.7e-07 $l=6.9925e-07 $layer=licon1_PDIFF $count=2 $X=7.26
+ $Y=1.84 $X2=7.395 $Y2=2.475
r90 2 31 600 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.84 $X2=3.58 $Y2=2.455
r91 1 26 600 $w=1.7e-07 $l=6.97029e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.84 $X2=2.58 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%VPWR 1 2 3 4 5 6 19 23 27 31 33 36 37 39 43
+ 46 48 56 61 66 72 75 78 82
r129 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r131 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r132 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r133 70 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r134 70 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r135 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r136 67 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.01 $Y=3.33
+ $X2=8.885 $Y2=3.33
r137 67 69 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.01 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 66 81 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.857 $Y2=3.33
r139 66 69 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.36 $Y2=3.33
r140 65 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r141 65 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r142 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r143 62 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=7.895 $Y2=3.33
r144 62 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=8.4 $Y2=3.33
r145 61 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.76 $Y=3.33
+ $X2=8.885 $Y2=3.33
r146 61 64 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.76 $Y=3.33
+ $X2=8.4 $Y2=3.33
r147 60 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 60 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r150 57 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.06 $Y=3.33
+ $X2=6.895 $Y2=3.33
r151 57 59 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.06 $Y=3.33
+ $X2=7.44 $Y2=3.33
r152 56 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=3.33
+ $X2=7.895 $Y2=3.33
r153 56 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.73 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 55 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r155 54 55 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r156 50 54 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r157 50 51 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r158 48 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.895 $Y2=3.33
r159 48 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.48 $Y2=3.33
r160 46 55 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 46 51 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r162 42 43 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.915 $Y=2.03
+ $X2=6.08 $Y2=2.03
r163 37 81 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.857 $Y2=3.33
r164 37 39 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.195
r165 34 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=3.245
+ $X2=8.885 $Y2=3.33
r166 34 36 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=8.885 $Y=3.245
+ $X2=8.885 $Y2=2.555
r167 33 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=2.22
+ $X2=8.885 $Y2=2.135
r168 33 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.885 $Y=2.22
+ $X2=8.885 $Y2=2.555
r169 29 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.895 $Y=3.245
+ $X2=7.895 $Y2=3.33
r170 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.895 $Y=3.245
+ $X2=7.895 $Y2=2.815
r171 25 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.895 $Y=3.245
+ $X2=6.895 $Y2=3.33
r172 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.895 $Y=3.245
+ $X2=6.895 $Y2=2.815
r173 23 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.76 $Y=2.135
+ $X2=8.885 $Y2=2.135
r174 23 43 174.845 $w=1.68e-07 $l=2.68e-06 $layer=LI1_cond $X=8.76 $Y=2.135
+ $X2=6.08 $Y2=2.135
r175 19 42 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=5.89 $Y=2.03
+ $X2=5.915 $Y2=2.03
r176 19 21 26.5365 $w=3.78e-07 $l=8.75e-07 $layer=LI1_cond $X=5.89 $Y=2.03
+ $X2=5.015 $Y2=2.03
r177 6 39 300 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_PDIFF $count=2 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=2.195
r178 5 45 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=8.71
+ $Y=1.84 $X2=8.845 $Y2=2.135
r179 5 36 600 $w=1.7e-07 $l=7.79583e-07 $layer=licon1_PDIFF $count=1 $X=8.71
+ $Y=1.84 $X2=8.845 $Y2=2.555
r180 4 31 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=7.71
+ $Y=1.84 $X2=7.895 $Y2=2.815
r181 3 27 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=1.84 $X2=6.895 $Y2=2.815
r182 2 42 600 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=1.84 $X2=5.915 $Y2=2.03
r183 1 21 300 $w=1.7e-07 $l=5.96825e-07 $layer=licon1_PDIFF $count=2 $X=4.495
+ $Y=1.84 $X2=5.015 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A_114_85# 1 2 3 4 15 17 18 21 23 26 28 29 31
+ 35 37 38 39 41
c109 35 0 1.15153e-19 $X=8.66 $Y=0.555
r110 43 44 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=7.57 $Y=0.665
+ $X2=7.57 $Y2=0.925
r111 41 43 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=7.57 $Y=0.555
+ $X2=7.57 $Y2=0.665
r112 38 39 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.355 $Y=0.705
+ $X2=5.525 $Y2=0.705
r113 33 35 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.66 $Y=0.84
+ $X2=8.66 $Y2=0.555
r114 32 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=0.925
+ $X2=7.57 $Y2=0.925
r115 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.495 $Y=0.925
+ $X2=8.66 $Y2=0.84
r116 31 32 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.495 $Y=0.925
+ $X2=7.735 $Y2=0.925
r117 29 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=0.665
+ $X2=7.57 $Y2=0.665
r118 29 39 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=7.405 $Y=0.665
+ $X2=5.525 $Y2=0.665
r119 28 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.765 $Y=0.745
+ $X2=5.355 $Y2=0.745
r120 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.68 $Y=0.66
+ $X2=4.765 $Y2=0.745
r121 25 26 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.68 $Y=0.425
+ $X2=4.68 $Y2=0.66
r122 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0.34
+ $X2=1.57 $Y2=0.34
r123 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.595 $Y=0.34
+ $X2=4.68 $Y2=0.425
r124 23 24 186.588 $w=1.68e-07 $l=2.86e-06 $layer=LI1_cond $X=4.595 $Y=0.34
+ $X2=1.735 $Y2=0.34
r125 19 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.425
+ $X2=1.57 $Y2=0.34
r126 19 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.57 $Y=0.425
+ $X2=1.57 $Y2=0.675
r127 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.34
+ $X2=1.57 $Y2=0.34
r128 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=0.34
+ $X2=0.875 $Y2=0.34
r129 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=0.425
+ $X2=0.875 $Y2=0.34
r130 13 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.71 $Y=0.425
+ $X2=0.71 $Y2=0.675
r131 4 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.52
+ $Y=0.41 $X2=8.66 $Y2=0.555
r132 3 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.43
+ $Y=0.41 $X2=7.57 $Y2=0.555
r133 2 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.425 $X2=1.57 $Y2=0.675
r134 1 15 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.425 $X2=0.71 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%A_475_85# 1 2 3 4 13 20 22 26 27
r44 26 27 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.55 $Y=1.045
+ $X2=6.385 $Y2=1.045
r45 24 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=5.53 $Y=1.085
+ $X2=6.385 $Y2=1.085
r46 22 24 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.425 $Y=1.085
+ $X2=5.53 $Y2=1.085
r47 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.34 $Y=1
+ $X2=4.425 $Y2=1.085
r48 19 20 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.34 $Y=0.765
+ $X2=4.34 $Y2=1
r49 15 18 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.585 $Y=0.68
+ $X2=3.49 $Y2=0.68
r50 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.255 $Y=0.68
+ $X2=4.34 $Y2=0.765
r51 13 18 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.255 $Y=0.68
+ $X2=3.49 $Y2=0.68
r52 4 26 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.41
+ $Y=0.41 $X2=6.55 $Y2=1.005
r53 3 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.49 $X2=5.53 $Y2=1.085
r54 2 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.425 $X2=3.49 $Y2=0.68
r55 1 15 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.425 $X2=2.585 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2I_4%VGND 1 2 3 4 5 18 20 22 26 30 33 34 35 37 45
+ 55 56 59 63 70 76
r95 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r96 71 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r97 70 73 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.06 $Y=0 $X2=7.06
+ $Y2=0.325
r98 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r99 64 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r100 63 66 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.04 $Y=0 $X2=6.04
+ $Y2=0.325
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r102 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r103 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r104 53 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r105 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r106 50 76 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.325 $Y=0 $X2=8.115
+ $Y2=0
r107 50 52 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.325 $Y=0
+ $X2=8.88 $Y2=0
r108 49 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r109 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r110 46 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.06
+ $Y2=0
r111 46 48 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=0
+ $X2=5.52 $Y2=0
r112 45 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=0 $X2=6.04
+ $Y2=0
r113 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.875 $Y=0
+ $X2=5.52 $Y2=0
r114 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r115 40 44 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.56
+ $Y2=0
r116 39 43 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.56
+ $Y2=0
r117 39 40 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 37 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=5.06
+ $Y2=0
r119 37 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.935 $Y=0
+ $X2=4.56 $Y2=0
r120 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r121 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r122 35 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r123 33 52 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.995 $Y=0
+ $X2=8.88 $Y2=0
r124 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.995 $Y=0 $X2=9.16
+ $Y2=0
r125 32 55 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=9.84 $Y2=0
r126 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.325 $Y=0 $X2=9.16
+ $Y2=0
r127 28 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.16 $Y=0.085
+ $X2=9.16 $Y2=0
r128 28 30 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=9.16 $Y=0.085
+ $X2=9.16 $Y2=0.555
r129 24 76 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0
r130 24 26 12.8964 $w=4.18e-07 $l=4.7e-07 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0.555
r131 23 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.225 $Y=0 $X2=7.06
+ $Y2=0
r132 22 76 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.905 $Y=0 $X2=8.115
+ $Y2=0
r133 22 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.905 $Y=0
+ $X2=7.225 $Y2=0
r134 21 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.04
+ $Y2=0
r135 20 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.895 $Y=0 $X2=7.06
+ $Y2=0
r136 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.205
+ $Y2=0
r137 16 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r138 16 18 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.325
r139 5 30 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.95
+ $Y=0.41 $X2=9.16 $Y2=0.555
r140 4 26 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=7.86
+ $Y=0.41 $X2=8.115 $Y2=0.555
r141 3 73 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=6.84
+ $Y=0.41 $X2=7.06 $Y2=0.325
r142 2 66 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=5.82
+ $Y=0.49 $X2=6.04 $Y2=0.325
r143 1 18 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.18 $X2=5.02 $Y2=0.325
.ends


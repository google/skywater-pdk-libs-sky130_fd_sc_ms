# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__nor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 0.935000 1.920000 ;
        RECT 0.605000 1.920000 1.795000 2.170000 ;
        RECT 1.625000 2.170000 6.135000 2.190000 ;
        RECT 1.625000 2.190000 4.020000 2.340000 ;
        RECT 3.850000 2.020000 6.135000 2.170000 ;
        RECT 5.805000 0.330000 6.135000 2.020000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.310000 1.350000 4.965000 1.510000 ;
        RECT 1.310000 1.510000 2.755000 1.520000 ;
        RECT 1.310000 1.520000 1.640000 1.680000 ;
        RECT 2.045000 1.180000 4.965000 1.350000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785000 0.340000 5.635000 0.670000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.674800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 1.875000 1.180000 ;
        RECT 1.545000 0.350000 1.875000 0.840000 ;
        RECT 1.545000 0.840000 5.305000 1.010000 ;
        RECT 2.140000 1.750000 5.305000 1.850000 ;
        RECT 2.140000 1.850000 3.680000 2.000000 ;
        RECT 2.545000 0.350000 2.875000 0.840000 ;
        RECT 3.350000 1.680000 5.305000 1.750000 ;
        RECT 5.135000 1.010000 5.305000 1.680000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.110000  1.820000 0.360000 2.340000 ;
      RECT 0.110000  2.340000 1.340000 2.510000 ;
      RECT 0.110000  2.510000 0.360000 2.980000 ;
      RECT 0.115000  0.085000 0.365000 1.130000 ;
      RECT 0.560000  2.680000 0.890000 3.245000 ;
      RECT 1.045000  0.085000 1.375000 0.840000 ;
      RECT 1.090000  2.510000 6.615000 2.530000 ;
      RECT 1.090000  2.530000 4.735000 2.680000 ;
      RECT 1.090000  2.680000 1.340000 2.980000 ;
      RECT 1.540000  2.850000 4.285000 2.905000 ;
      RECT 1.540000  2.905000 5.265000 3.075000 ;
      RECT 2.045000  0.085000 2.375000 0.670000 ;
      RECT 3.055000  0.085000 3.365000 0.670000 ;
      RECT 4.485000  2.360000 6.615000 2.510000 ;
      RECT 4.485000  2.680000 4.735000 2.735000 ;
      RECT 4.935000  2.700000 5.265000 2.905000 ;
      RECT 5.465000  2.530000 5.635000 3.000000 ;
      RECT 5.835000  2.700000 6.165000 3.245000 ;
      RECT 6.365000  1.820000 6.615000 2.360000 ;
      RECT 6.365000  2.530000 6.615000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ms__nor3_4

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__ha_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__ha_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.582000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.450000 1.390000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.582000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.550000 1.630000 ;
        RECT 0.125000 1.630000 0.295000 2.320000 ;
        RECT 0.125000 2.320000 2.120000 2.520000 ;
        RECT 1.790000 1.450000 2.120000 2.320000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.865000 1.820000 5.195000 2.170000 ;
        RECT 4.885000 0.350000 5.215000 1.130000 ;
        RECT 4.885000 1.130000 5.055000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.546600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.820000 4.675000 2.170000 ;
        RECT 3.975000 0.880000 4.675000 1.050000 ;
        RECT 4.505000 1.050000 4.675000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 0.890000 1.110000 ;
      RECT 0.115000  1.110000 2.460000 1.130000 ;
      RECT 0.115000  2.690000 0.445000 3.245000 ;
      RECT 0.565000  1.980000 0.895000 2.150000 ;
      RECT 0.720000  1.130000 2.460000 1.280000 ;
      RECT 0.720000  1.280000 0.890000 1.980000 ;
      RECT 0.935000  0.085000 1.265000 0.600000 ;
      RECT 1.015000  2.690000 1.400000 3.245000 ;
      RECT 1.365000  0.770000 2.465000 0.940000 ;
      RECT 1.795000  0.085000 2.125000 0.600000 ;
      RECT 2.290000  1.280000 3.035000 1.610000 ;
      RECT 2.290000  1.610000 2.460000 2.340000 ;
      RECT 2.290000  2.340000 5.555000 2.510000 ;
      RECT 2.295000  0.255000 3.315000 0.425000 ;
      RECT 2.295000  0.425000 2.465000 0.770000 ;
      RECT 2.630000  1.920000 3.490000 2.170000 ;
      RECT 2.635000  0.595000 2.805000 0.940000 ;
      RECT 2.635000  0.940000 3.490000 1.110000 ;
      RECT 2.985000  0.425000 3.315000 0.770000 ;
      RECT 3.080000  2.680000 3.845000 3.245000 ;
      RECT 3.320000  1.110000 3.490000 1.220000 ;
      RECT 3.320000  1.220000 4.330000 1.550000 ;
      RECT 3.320000  1.550000 3.490000 1.920000 ;
      RECT 3.545000  0.085000 3.875000 0.710000 ;
      RECT 4.415000  2.680000 4.745000 3.245000 ;
      RECT 4.455000  0.085000 4.705000 0.710000 ;
      RECT 5.225000  1.300000 5.555000 1.630000 ;
      RECT 5.315000  2.680000 5.645000 3.245000 ;
      RECT 5.385000  1.630000 5.555000 2.340000 ;
      RECT 5.395000  0.085000 5.645000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__ha_2
END LIBRARY

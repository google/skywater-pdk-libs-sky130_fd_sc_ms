* File: sky130_fd_sc_ms__o211a_2.pex.spice
* Created: Wed Sep  2 12:20:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O211A_2%C1 3 5 7 8 15
c25 8 0 1.40395e-19 $X=0.24 $Y=1.295
r26 14 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.51 $Y2=1.385
r27 11 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.385
+ $X2=0.495 $Y2=1.385
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r29 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r30 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.22
+ $X2=0.51 $Y2=1.385
r31 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=1.22 $X2=0.51
+ $Y2=0.74
r32 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=1.385
r33 1 3 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%B1 3 7 9 12 13
c38 13 0 1.11966e-19 $X=0.96 $Y=1.515
c39 12 0 1.40395e-19 $X=0.96 $Y=1.515
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.96 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.96 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.515 $X2=0.96 $Y2=1.515
r43 9 13 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.96 $Y2=1.565
r44 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.035 $Y=2.34
+ $X2=1.035 $Y2=1.68
r45 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.9 $Y=0.74 $X2=0.9
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%A2 3 7 9 12
c38 7 0 1.90452e-19 $X=1.495 $Y=2.34
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.515
+ $X2=1.5 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.515
+ $X2=1.5 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.515 $X2=1.5 $Y2=1.515
r42 9 13 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.5
+ $Y2=1.565
r43 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.495 $Y=2.34
+ $X2=1.495 $Y2=1.68
r44 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.41 $Y=0.74 $X2=1.41
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%A1 3 7 9 15 16
c39 16 0 7.84859e-20 $X=2.13 $Y=1.515
c40 15 0 1.82087e-19 $X=2.13 $Y=1.515
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r42 13 15 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.97 $Y=1.515
+ $X2=2.13 $Y2=1.515
r43 11 13 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.965 $Y=1.515
+ $X2=1.97 $Y2=1.515
r44 9 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r45 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.35
+ $X2=1.97 $Y2=1.515
r46 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.97 $Y=1.35 $X2=1.97
+ $Y2=0.74
r47 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.68
+ $X2=1.965 $Y2=1.515
r48 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.965 $Y=1.68
+ $X2=1.965 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%A_27_368# 1 2 3 10 12 13 15 16 18 20 22 23
+ 25 27 29 33 35 37 38 42 45
c120 42 0 7.65495e-20 $X=0.295 $Y=0.515
c121 38 0 1.82087e-19 $X=2.59 $Y=1.95
r122 51 52 10.3597 $w=4.42e-07 $l=9.5e-08 $layer=POLY_cond $X=2.835 $Y=1.455
+ $X2=2.93 $Y2=1.455
r123 49 51 17.9932 $w=4.42e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.455
+ $X2=2.835 $Y2=1.455
r124 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.465 $X2=2.67 $Y2=1.465
r125 46 48 17.702 $w=2.55e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.095
+ $X2=2.67 $Y2=1.465
r126 37 48 9.25285 $w=2.55e-07 $l=2.0106e-07 $layer=LI1_cond $X=2.59 $Y=1.63
+ $X2=2.67 $Y2=1.465
r127 37 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.59 $Y=1.63
+ $X2=2.59 $Y2=1.95
r128 36 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=2.035
+ $X2=1.27 $Y2=2.035
r129 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=2.59 $Y2=1.95
r130 35 36 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=1.435 $Y2=2.035
r131 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.12
+ $X2=1.27 $Y2=2.035
r132 31 33 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.27 $Y=2.12
+ $X2=1.27 $Y2=2.715
r133 30 42 12.936 $w=5.47e-07 $l=7.23699e-07 $layer=LI1_cond $X=0.775 $Y=1.095
+ $X2=0.452 $Y2=0.515
r134 29 46 3.11056 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.095
+ $X2=2.67 $Y2=1.095
r135 29 30 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=2.505 $Y=1.095
+ $X2=0.775 $Y2=1.095
r136 28 40 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.435 $Y=2.035
+ $X2=0.27 $Y2=1.97
r137 27 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=2.035
+ $X2=1.27 $Y2=2.035
r138 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=2.035
+ $X2=0.435 $Y2=2.035
r139 23 40 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.27 $Y=2.12 $X2=0.27
+ $Y2=1.97
r140 23 25 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=0.27 $Y=2.12
+ $X2=0.27 $Y2=2.695
r141 20 54 28.321 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.36 $Y=1.185
+ $X2=3.36 $Y2=1.455
r142 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.36 $Y=1.185
+ $X2=3.36 $Y2=0.74
r143 16 54 8.17873 $w=4.42e-07 $l=7.5e-08 $layer=POLY_cond $X=3.285 $Y=1.455
+ $X2=3.36 $Y2=1.455
r144 16 52 38.7127 $w=4.42e-07 $l=3.55e-07 $layer=POLY_cond $X=3.285 $Y=1.455
+ $X2=2.93 $Y2=1.455
r145 16 18 320.685 $w=1.8e-07 $l=8.25e-07 $layer=POLY_cond $X=3.285 $Y=1.575
+ $X2=3.285 $Y2=2.4
r146 13 52 28.321 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.93 $Y=1.185
+ $X2=2.93 $Y2=1.455
r147 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.93 $Y=1.185
+ $X2=2.93 $Y2=0.74
r148 10 51 23.8576 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.835 $Y=1.725
+ $X2=2.835 $Y2=1.455
r149 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.835 $Y=1.725
+ $X2=2.835 $Y2=2.4
r150 3 45 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.84 $X2=1.27 $Y2=2.035
r151 3 33 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.84 $X2=1.27 $Y2=2.715
r152 2 40 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
r153 2 25 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.695
r154 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%VPWR 1 2 3 12 16 18 20 24 26 31 36 42 45 49
r48 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 40 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 37 45 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.375 $Y2=3.33
r55 37 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 36 48 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.617 $Y2=3.33
r57 36 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 35 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.77 $Y2=3.33
r61 32 34 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 31 45 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.375 $Y2=3.33
r63 31 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 29 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 26 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.77 $Y2=3.33
r67 26 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 24 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 20 23 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.56 $Y=1.985
+ $X2=3.56 $Y2=2.815
r71 18 48 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.617 $Y2=3.33
r72 18 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.815
r73 14 45 2.86223 $w=7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=3.245
+ $X2=2.375 $Y2=3.33
r74 14 16 14.8655 $w=6.98e-07 $l=8.7e-07 $layer=LI1_cond $X=2.375 $Y=3.245
+ $X2=2.375 $Y2=2.375
r75 10 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r76 10 12 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.375
r77 3 23 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.84 $X2=3.56 $Y2=2.815
r78 3 20 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.84 $X2=3.56 $Y2=1.985
r79 2 16 150 $w=1.7e-07 $l=7.45922e-07 $layer=licon1_PDIFF $count=4 $X=2.055
+ $Y=1.84 $X2=2.56 $Y2=2.375
r80 1 12 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.77 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%X 1 2 9 11 15 16 17 18 31 36
c30 17 0 1.11614e-19 $X=3.035 $Y=0.84
r31 24 31 3.52512 $w=2.53e-07 $l=7.8e-08 $layer=LI1_cond $X=3.107 $Y=1.003
+ $X2=3.107 $Y2=0.925
r32 18 42 3.65775 $w=2.28e-07 $l=7.3e-08 $layer=LI1_cond $X=3.12 $Y=1.337
+ $X2=3.12 $Y2=1.41
r33 18 36 2.10446 $w=2.28e-07 $l=4.2e-08 $layer=LI1_cond $X=3.12 $Y=1.337
+ $X2=3.12 $Y2=1.295
r34 18 36 2.15457 $w=2.28e-07 $l=4.3e-08 $layer=LI1_cond $X=3.12 $Y=1.252
+ $X2=3.12 $Y2=1.295
r35 18 38 6.11296 $w=2.28e-07 $l=1.22e-07 $layer=LI1_cond $X=3.12 $Y=1.252
+ $X2=3.12 $Y2=1.13
r36 17 38 5.73947 $w=2.53e-07 $l=1.24e-07 $layer=LI1_cond $X=3.107 $Y=1.006
+ $X2=3.107 $Y2=1.13
r37 17 24 0.135582 $w=2.53e-07 $l=3e-09 $layer=LI1_cond $X=3.107 $Y=1.006
+ $X2=3.107 $Y2=1.003
r38 17 31 0.180775 $w=2.53e-07 $l=4e-09 $layer=LI1_cond $X=3.107 $Y=0.921
+ $X2=3.107 $Y2=0.925
r39 16 17 18.3487 $w=2.53e-07 $l=4.06e-07 $layer=LI1_cond $X=3.107 $Y=0.515
+ $X2=3.107 $Y2=0.921
r40 15 42 21.4773 $w=2.18e-07 $l=4.1e-07 $layer=LI1_cond $X=3.115 $Y=1.82
+ $X2=3.115 $Y2=1.41
r41 9 15 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=1.985
+ $X2=3.06 $Y2=1.82
r42 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.06 $Y=1.985
+ $X2=3.06 $Y2=2.815
r43 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.84 $X2=3.06 $Y2=2.815
r44 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.84 $X2=3.06 $Y2=1.985
r45 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.005
+ $Y=0.37 $X2=3.145 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%A_195_74# 1 2 7 10 15
r27 15 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.185 $Y=0.595
+ $X2=2.185 $Y2=0.755
r28 10 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.19 $Y=0.595
+ $X2=1.19 $Y2=0.755
r29 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.755
+ $X2=1.19 $Y2=0.755
r30 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=0.755
+ $X2=2.185 $Y2=0.755
r31 7 8 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.02 $Y=0.755
+ $X2=1.355 $Y2=0.755
r32 2 15 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.37 $X2=2.185 $Y2=0.595
r33 1 10 182 $w=1.7e-07 $l=3.14643e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.37 $X2=1.19 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_2%VGND 1 2 3 12 16 18 20 22 24 32 37 43 46 50
r50 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r52 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r54 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r55 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 38 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.675
+ $Y2=0
r57 38 40 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.12
+ $Y2=0
r58 37 49 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.625
+ $Y2=0
r59 37 40 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.12
+ $Y2=0
r60 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r61 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 33 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.65
+ $Y2=0
r63 33 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=2.16
+ $Y2=0
r64 32 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.675
+ $Y2=0
r65 32 35 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.16
+ $Y2=0
r66 31 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r67 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 27 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r69 26 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r70 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r71 24 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.65
+ $Y2=0
r72 24 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.2
+ $Y2=0
r73 22 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r74 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r75 18 49 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.625 $Y2=0
r76 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.515
r77 14 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.085
+ $X2=2.675 $Y2=0
r78 14 16 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=2.675 $Y=0.085
+ $X2=2.675 $Y2=0.595
r79 10 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0
r80 10 12 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0.335
r81 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.37 $X2=3.575 $Y2=0.515
r82 2 16 182 $w=1.7e-07 $l=2.82622e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.37 $X2=2.715 $Y2=0.595
r83 1 12 182 $w=1.7e-07 $l=2.21811e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.37 $X2=1.69 $Y2=0.335
.ends


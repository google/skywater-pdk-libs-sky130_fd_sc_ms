* File: sky130_fd_sc_ms__o32a_1.pxi.spice
* Created: Wed Sep  2 12:26:10 2020
* 
x_PM_SKY130_FD_SC_MS__O32A_1%A_83_264# N_A_83_264#_M1006_d N_A_83_264#_M1011_d
+ N_A_83_264#_M1003_g N_A_83_264#_M1007_g N_A_83_264#_c_74_n N_A_83_264#_c_85_p
+ N_A_83_264#_c_142_p N_A_83_264#_c_81_n N_A_83_264#_c_109_p N_A_83_264#_c_75_n
+ N_A_83_264#_c_76_n N_A_83_264#_c_77_n N_A_83_264#_c_78_n N_A_83_264#_c_104_p
+ PM_SKY130_FD_SC_MS__O32A_1%A_83_264#
x_PM_SKY130_FD_SC_MS__O32A_1%A1 N_A1_M1005_g N_A1_M1010_g A1 N_A1_c_166_n
+ N_A1_c_167_n PM_SKY130_FD_SC_MS__O32A_1%A1
x_PM_SKY130_FD_SC_MS__O32A_1%A2 N_A2_M1009_g N_A2_M1002_g A2 N_A2_c_207_n
+ N_A2_c_208_n PM_SKY130_FD_SC_MS__O32A_1%A2
x_PM_SKY130_FD_SC_MS__O32A_1%A3 N_A3_M1011_g N_A3_M1008_g A3 N_A3_c_243_n
+ N_A3_c_244_n PM_SKY130_FD_SC_MS__O32A_1%A3
x_PM_SKY130_FD_SC_MS__O32A_1%B2 N_B2_M1001_g N_B2_M1006_g B2 N_B2_c_281_n
+ N_B2_c_282_n PM_SKY130_FD_SC_MS__O32A_1%B2
x_PM_SKY130_FD_SC_MS__O32A_1%B1 N_B1_M1004_g N_B1_M1000_g B1 B1 N_B1_c_324_n
+ PM_SKY130_FD_SC_MS__O32A_1%B1
x_PM_SKY130_FD_SC_MS__O32A_1%X N_X_M1007_s N_X_M1003_s N_X_c_354_n N_X_c_355_n
+ N_X_c_351_n X X N_X_c_352_n X PM_SKY130_FD_SC_MS__O32A_1%X
x_PM_SKY130_FD_SC_MS__O32A_1%VPWR N_VPWR_M1003_d N_VPWR_M1004_d N_VPWR_c_379_n
+ N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n VPWR
+ N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_378_n
+ PM_SKY130_FD_SC_MS__O32A_1%VPWR
x_PM_SKY130_FD_SC_MS__O32A_1%VGND N_VGND_M1007_d N_VGND_M1002_d N_VGND_c_423_n
+ N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n
+ VGND N_VGND_c_429_n N_VGND_c_430_n PM_SKY130_FD_SC_MS__O32A_1%VGND
x_PM_SKY130_FD_SC_MS__O32A_1%A_251_74# N_A_251_74#_M1010_d N_A_251_74#_M1008_d
+ N_A_251_74#_M1000_d N_A_251_74#_c_467_n N_A_251_74#_c_468_n
+ N_A_251_74#_c_469_n N_A_251_74#_c_470_n N_A_251_74#_c_488_n
+ N_A_251_74#_c_471_n N_A_251_74#_c_472_n PM_SKY130_FD_SC_MS__O32A_1%A_251_74#
cc_1 VNB N_A_83_264#_M1003_g 5.69697e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_264#_M1007_g 0.03041f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_3 VNB N_A_83_264#_c_74_n 2.45937e-19 $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_4 VNB N_A_83_264#_c_75_n 0.00753812f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=1.18
cc_5 VNB N_A_83_264#_c_76_n 0.0036728f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=1.95
cc_6 VNB N_A_83_264#_c_77_n 0.0337383f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.485
cc_7 VNB N_A_83_264#_c_78_n 0.0027277f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.485
cc_8 VNB N_A1_M1010_g 0.0314409f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_9 VNB N_A1_c_166_n 0.0243048f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_10 VNB N_A1_c_167_n 0.00547709f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_11 VNB N_A2_M1002_g 0.0305392f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_12 VNB N_A2_c_207_n 0.0262307f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_13 VNB N_A2_c_208_n 0.00165774f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_14 VNB N_A3_M1008_g 0.0316956f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_15 VNB N_A3_c_243_n 0.0262274f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_16 VNB N_A3_c_244_n 0.00165645f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_17 VNB N_B2_M1006_g 0.0326134f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_18 VNB N_B2_c_281_n 0.0249231f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_19 VNB N_B2_c_282_n 0.0051357f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_20 VNB N_B1_M1004_g 0.00797545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_M1000_g 0.0294724f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_22 VNB B1 0.0119477f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB N_B1_c_324_n 0.0670728f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.035
cc_24 VNB N_X_c_351_n 0.0250947f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_25 VNB N_X_c_352_n 0.0283371f $X=-0.19 $Y=-0.245 $X2=3.065 $Y2=2.035
cc_26 VNB X 0.0180876f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.485
cc_27 VNB N_VPWR_c_378_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_423_n 0.0109103f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_29 VNB N_VGND_c_424_n 0.00895062f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_30 VNB N_VGND_c_425_n 0.0216783f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_31 VNB N_VGND_c_426_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.035
cc_32 VNB N_VGND_c_427_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=2.12
cc_33 VNB N_VGND_c_428_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.4 $Y2=2.715
cc_34 VNB N_VGND_c_429_n 0.0474473f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.035
cc_35 VNB N_VGND_c_430_n 0.23222f $X=-0.19 $Y=-0.245 $X2=2.982 $Y2=0.865
cc_36 VNB N_A_251_74#_c_467_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.74
cc_37 VNB N_A_251_74#_c_468_n 0.0247434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_251_74#_c_469_n 0.00810708f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_39 VNB N_A_251_74#_c_470_n 0.00257219f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_40 VNB N_A_251_74#_c_471_n 0.00456757f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_41 VNB N_A_251_74#_c_472_n 0.0049404f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=1.18
cc_42 VPB N_A_83_264#_M1003_g 0.0305464f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_43 VPB N_A_83_264#_c_74_n 0.00283485f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_44 VPB N_A_83_264#_c_81_n 0.00364632f $X=-0.19 $Y=1.66 $X2=2.395 $Y2=2.715
cc_45 VPB N_A_83_264#_c_76_n 0.00141192f $X=-0.19 $Y=1.66 $X2=3.15 $Y2=1.95
cc_46 VPB N_A1_M1005_g 0.0218345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A1_c_166_n 0.00560643f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_48 VPB N_A1_c_167_n 0.00307875f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_49 VPB N_A2_M1009_g 0.021491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A2_c_207_n 0.00562335f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_51 VPB N_A2_c_208_n 0.00205011f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_52 VPB N_A3_M1011_g 0.0225257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A3_c_243_n 0.00562174f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_54 VPB N_A3_c_244_n 0.00200497f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_55 VPB N_B2_M1001_g 0.0224682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_B2_c_281_n 0.00553695f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_57 VPB N_B2_c_282_n 0.00308059f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_58 VPB N_B1_M1004_g 0.0263641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB B1 0.0119607f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_60 VPB N_X_c_354_n 0.0415472f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.32
cc_61 VPB N_X_c_355_n 0.0136968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_X_c_351_n 0.00750262f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.65
cc_63 VPB N_VPWR_c_379_n 0.0143084f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_64 VPB N_VPWR_c_380_n 0.00626527f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.74
cc_65 VPB N_VPWR_c_381_n 0.0145833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_382_n 0.0345959f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_67 VPB N_VPWR_c_383_n 0.0117986f $X=-0.19 $Y=1.66 $X2=2.4 $Y2=2.12
cc_68 VPB N_VPWR_c_384_n 0.0189171f $X=-0.19 $Y=1.66 $X2=2.595 $Y2=2.035
cc_69 VPB N_VPWR_c_385_n 0.0730231f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.485
cc_70 VPB N_VPWR_c_386_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.32
cc_71 VPB N_VPWR_c_378_n 0.116326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_A_83_264#_M1003_g N_A1_M1005_g 0.0174581f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_83_264#_c_74_n N_A1_M1005_g 0.00360669f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_74 N_A_83_264#_c_85_p N_A1_M1005_g 0.0177183f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_75 N_A_83_264#_M1007_g N_A1_M1010_g 0.023959f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A_83_264#_c_77_n N_A1_M1010_g 8.96112e-19 $X=0.58 $Y=1.485 $X2=0 $Y2=0
cc_77 N_A_83_264#_c_78_n N_A1_M1010_g 5.98792e-19 $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_78 N_A_83_264#_M1003_g N_A1_c_166_n 7.81769e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_83_264#_c_74_n N_A1_c_166_n 2.15441e-19 $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_80 N_A_83_264#_c_85_p N_A1_c_166_n 5.45341e-19 $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_83_264#_c_77_n N_A1_c_166_n 0.018763f $X=0.58 $Y=1.485 $X2=0 $Y2=0
cc_82 N_A_83_264#_c_78_n N_A1_c_166_n 0.00170039f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_83 N_A_83_264#_c_74_n N_A1_c_167_n 0.0102525f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_84 N_A_83_264#_c_85_p N_A1_c_167_n 0.0232864f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_83_264#_c_77_n N_A1_c_167_n 3.43727e-19 $X=0.58 $Y=1.485 $X2=0 $Y2=0
cc_86 N_A_83_264#_c_78_n N_A1_c_167_n 0.0240952f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_87 N_A_83_264#_c_85_p N_A2_M1009_g 0.0173173f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_83_264#_c_81_n N_A2_M1009_g 0.00337214f $X=2.395 $Y=2.715 $X2=0 $Y2=0
cc_89 N_A_83_264#_c_85_p N_A2_c_207_n 7.07929e-19 $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A_83_264#_c_85_p N_A2_c_208_n 0.0229716f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_85_p N_A3_M1011_g 0.0147916f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_81_n N_A3_M1011_g 0.0153314f $X=2.395 $Y=2.715 $X2=0 $Y2=0
cc_93 N_A_83_264#_c_104_p N_A3_M1011_g 2.7414e-19 $X=2.395 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_83_264#_c_104_p N_A3_c_243_n 7.71396e-19 $X=2.395 $Y=2.035 $X2=0 $Y2=0
cc_95 N_A_83_264#_c_85_p N_A3_c_244_n 0.01236f $X=2.205 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_83_264#_c_104_p N_A3_c_244_n 0.0114387f $X=2.395 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A_83_264#_c_81_n N_B2_M1001_g 0.0166557f $X=2.395 $Y=2.715 $X2=0 $Y2=0
cc_98 N_A_83_264#_c_109_p N_B2_M1001_g 0.0143596f $X=3.065 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_76_n N_B2_M1001_g 0.0034179f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_104_p N_B2_M1001_g 5.7874e-19 $X=2.395 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_83_264#_c_75_n N_B2_M1006_g 0.0135416f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_76_n N_B2_M1006_g 0.00313735f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_103 N_A_83_264#_c_109_p N_B2_c_281_n 0.00102545f $X=3.065 $Y=2.035 $X2=0
+ $Y2=0
cc_104 N_A_83_264#_c_75_n N_B2_c_281_n 0.00152828f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_76_n N_B2_c_281_n 0.00201924f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_106 N_A_83_264#_c_109_p N_B2_c_282_n 0.0207439f $X=3.065 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_83_264#_c_75_n N_B2_c_282_n 0.0136544f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_76_n N_B2_c_282_n 0.0329497f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_109 N_A_83_264#_c_104_p N_B2_c_282_n 0.00329911f $X=2.395 $Y=2.035 $X2=0
+ $Y2=0
cc_110 N_A_83_264#_c_81_n N_B1_M1004_g 0.00334894f $X=2.395 $Y=2.715 $X2=0 $Y2=0
cc_111 N_A_83_264#_c_109_p N_B1_M1004_g 0.00917584f $X=3.065 $Y=2.035 $X2=0
+ $Y2=0
cc_112 N_A_83_264#_c_76_n N_B1_M1004_g 0.0147089f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_75_n N_B1_M1000_g 0.0197418f $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_76_n B1 0.0428502f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_75_n N_B1_c_324_n 6.70187e-19 $X=3.15 $Y=1.18 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_76_n N_B1_c_324_n 0.00900681f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_117 N_A_83_264#_M1003_g N_X_c_354_n 0.0148069f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_83_264#_M1003_g N_X_c_355_n 0.00321211f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_83_264#_c_74_n N_X_c_355_n 0.00565814f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_120 N_A_83_264#_c_78_n N_X_c_355_n 0.00151667f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_121 N_A_83_264#_M1007_g N_X_c_351_n 0.00424574f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_83_264#_c_74_n N_X_c_351_n 0.00535845f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_123 N_A_83_264#_c_77_n N_X_c_351_n 0.0101571f $X=0.58 $Y=1.485 $X2=0 $Y2=0
cc_124 N_A_83_264#_c_78_n N_X_c_351_n 0.0249376f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_125 N_A_83_264#_M1007_g N_X_c_352_n 0.0075748f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_83_264#_M1007_g X 0.00423703f $X=0.61 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_83_264#_c_77_n X 0.00343503f $X=0.58 $Y=1.485 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_78_n X 0.0102842f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_129 N_A_83_264#_c_74_n N_VPWR_M1003_d 0.00217698f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_83_264#_c_85_p N_VPWR_M1003_d 0.0125407f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_83_264#_c_142_p N_VPWR_M1003_d 0.00269585f $X=0.785 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_132 N_A_83_264#_M1003_g N_VPWR_c_379_n 0.00521232f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_133 N_A_83_264#_c_85_p N_VPWR_c_379_n 0.0128995f $X=2.205 $Y=2.035 $X2=0
+ $Y2=0
cc_134 N_A_83_264#_c_142_p N_VPWR_c_379_n 0.0116292f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_135 N_A_83_264#_c_77_n N_VPWR_c_379_n 3.5264e-19 $X=0.58 $Y=1.485 $X2=0 $Y2=0
cc_136 N_A_83_264#_c_109_p N_VPWR_c_383_n 0.0118099f $X=3.065 $Y=2.035 $X2=0
+ $Y2=0
cc_137 N_A_83_264#_M1003_g N_VPWR_c_384_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_83_264#_c_81_n N_VPWR_c_385_n 0.0122433f $X=2.395 $Y=2.715 $X2=0
+ $Y2=0
cc_139 N_A_83_264#_M1003_g N_VPWR_c_378_n 0.00990469f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_140 N_A_83_264#_c_81_n N_VPWR_c_378_n 0.0134094f $X=2.395 $Y=2.715 $X2=0
+ $Y2=0
cc_141 N_A_83_264#_c_85_p A_251_368# 0.00953889f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_83_264#_c_85_p A_335_368# 0.01606f $X=2.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_83_264#_c_109_p A_551_368# 0.0191624f $X=3.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_83_264#_c_76_n A_551_368# 0.00141422f $X=3.15 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_83_264#_M1007_g N_VGND_c_423_n 0.00737997f $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_83_264#_c_77_n N_VGND_c_423_n 2.61167e-19 $X=0.58 $Y=1.485 $X2=0
+ $Y2=0
cc_147 N_A_83_264#_c_78_n N_VGND_c_423_n 0.00279673f $X=0.7 $Y=1.485 $X2=0 $Y2=0
cc_148 N_A_83_264#_M1007_g N_VGND_c_425_n 0.00434272f $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_83_264#_M1007_g N_VGND_c_430_n 0.00825303f $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_83_264#_c_75_n N_A_251_74#_c_468_n 0.0147887f $X=3.15 $Y=1.18 $X2=0
+ $Y2=0
cc_151 N_A_83_264#_M1007_g N_A_251_74#_c_469_n 5.42515e-19 $X=0.61 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_83_264#_M1006_d N_A_251_74#_c_471_n 0.00431143f $X=2.755 $Y=0.37
+ $X2=0 $Y2=0
cc_153 N_A_83_264#_c_75_n N_A_251_74#_c_471_n 0.0277999f $X=3.15 $Y=1.18 $X2=0
+ $Y2=0
cc_154 N_A1_M1005_g N_A2_M1009_g 0.073253f $X=1.165 $Y=2.34 $X2=0 $Y2=0
cc_155 N_A1_M1010_g N_A2_M1002_g 0.0217728f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_156 N_A1_c_166_n N_A2_c_207_n 0.020661f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_157 N_A1_c_167_n N_A2_c_207_n 0.00244893f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A1_c_166_n N_A2_c_208_n 3.90049e-19 $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A1_c_167_n N_A2_c_208_n 0.0327917f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A1_M1005_g N_X_c_354_n 8.52238e-19 $X=1.165 $Y=2.34 $X2=0 $Y2=0
cc_161 N_A1_M1010_g N_X_c_352_n 4.46111e-19 $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_162 N_A1_M1005_g N_VPWR_c_379_n 0.0184077f $X=1.165 $Y=2.34 $X2=0 $Y2=0
cc_163 N_A1_M1005_g N_VPWR_c_385_n 0.0059286f $X=1.165 $Y=2.34 $X2=0 $Y2=0
cc_164 N_A1_M1005_g N_VPWR_c_378_n 0.00610055f $X=1.165 $Y=2.34 $X2=0 $Y2=0
cc_165 N_A1_M1010_g N_VGND_c_423_n 0.00606053f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_166 N_A1_c_166_n N_VGND_c_423_n 7.53427e-19 $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A1_c_167_n N_VGND_c_423_n 0.00553853f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A1_M1010_g N_VGND_c_427_n 0.00434272f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_169 N_A1_M1010_g N_VGND_c_430_n 0.0082141f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_170 N_A1_M1010_g N_A_251_74#_c_467_n 0.00725678f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_171 N_A1_M1010_g N_A_251_74#_c_469_n 0.0056999f $X=1.18 $Y=0.69 $X2=0 $Y2=0
cc_172 N_A1_c_166_n N_A_251_74#_c_469_n 2.37442e-19 $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A1_c_167_n N_A_251_74#_c_469_n 0.00726085f $X=1.12 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A2_M1009_g N_A3_M1011_g 0.0470587f $X=1.585 $Y=2.34 $X2=0 $Y2=0
cc_175 N_A2_c_208_n N_A3_M1011_g 6.85212e-19 $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A2_M1002_g N_A3_M1008_g 0.0261471f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_177 N_A2_c_207_n N_A3_c_243_n 0.0201104f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A2_c_208_n N_A3_c_243_n 0.00114936f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A2_c_207_n N_A3_c_244_n 0.00114936f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A2_c_208_n N_A3_c_244_n 0.0276388f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A2_M1009_g N_VPWR_c_385_n 0.0059286f $X=1.585 $Y=2.34 $X2=0 $Y2=0
cc_182 N_A2_M1009_g N_VPWR_c_378_n 0.00610055f $X=1.585 $Y=2.34 $X2=0 $Y2=0
cc_183 N_A2_M1002_g N_VGND_c_424_n 0.00472263f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_184 N_A2_M1002_g N_VGND_c_427_n 0.00434272f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_185 N_A2_M1002_g N_VGND_c_430_n 0.0082141f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_186 N_A2_M1002_g N_A_251_74#_c_467_n 0.00915605f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_187 N_A2_M1002_g N_A_251_74#_c_468_n 0.0117933f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_188 N_A2_c_207_n N_A_251_74#_c_468_n 9.79877e-19 $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A2_c_208_n N_A_251_74#_c_468_n 0.019847f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A2_M1002_g N_A_251_74#_c_469_n 0.0027332f $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_191 N_A2_c_207_n N_A_251_74#_c_469_n 3.0499e-19 $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_192 N_A2_c_208_n N_A_251_74#_c_469_n 0.00541082f $X=1.66 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A2_M1002_g N_A_251_74#_c_488_n 6.53479e-19 $X=1.61 $Y=0.69 $X2=0 $Y2=0
cc_194 N_A3_M1011_g N_B2_M1001_g 0.0107312f $X=2.125 $Y=2.34 $X2=0 $Y2=0
cc_195 N_A3_c_244_n N_B2_M1001_g 3.38956e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A3_M1008_g N_B2_M1006_g 0.0253778f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_197 N_A3_c_243_n N_B2_c_281_n 0.0206294f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A3_c_244_n N_B2_c_281_n 3.80681e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A3_M1011_g N_B2_c_282_n 2.66708e-19 $X=2.125 $Y=2.34 $X2=0 $Y2=0
cc_200 N_A3_c_243_n N_B2_c_282_n 0.00187654f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A3_c_244_n N_B2_c_282_n 0.0346782f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_202 N_A3_M1011_g N_VPWR_c_385_n 0.00584999f $X=2.125 $Y=2.34 $X2=0 $Y2=0
cc_203 N_A3_M1011_g N_VPWR_c_378_n 0.00610055f $X=2.125 $Y=2.34 $X2=0 $Y2=0
cc_204 N_A3_M1008_g N_VGND_c_424_n 0.00590558f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_205 N_A3_M1008_g N_VGND_c_429_n 0.00432912f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_206 N_A3_M1008_g N_VGND_c_430_n 0.00818188f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_207 N_A3_M1008_g N_A_251_74#_c_467_n 6.8749e-19 $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_208 N_A3_M1008_g N_A_251_74#_c_468_n 0.0145861f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_209 N_A3_c_243_n N_A_251_74#_c_468_n 0.00134262f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A3_c_244_n N_A_251_74#_c_468_n 0.0259036f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_211 N_A3_M1008_g N_A_251_74#_c_470_n 0.00250516f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_212 N_A3_M1008_g N_A_251_74#_c_488_n 0.00693236f $X=2.18 $Y=0.69 $X2=0 $Y2=0
cc_213 N_B2_M1001_g N_B1_M1004_g 0.0343415f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_214 N_B2_c_282_n N_B1_M1004_g 3.06315e-19 $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_215 N_B2_M1006_g N_B1_M1000_g 0.0231667f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_216 N_B2_M1006_g N_B1_c_324_n 0.00411837f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_217 N_B2_c_281_n N_B1_c_324_n 0.0152263f $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_218 N_B2_c_282_n N_B1_c_324_n 3.41341e-19 $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_219 N_B2_M1001_g N_VPWR_c_380_n 0.00305131f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_220 N_B2_M1001_g N_VPWR_c_385_n 0.00576265f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_221 N_B2_M1001_g N_VPWR_c_378_n 0.00610055f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_222 N_B2_M1006_g N_VGND_c_429_n 0.00290288f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_223 N_B2_M1006_g N_VGND_c_430_n 0.00360251f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_224 N_B2_M1006_g N_A_251_74#_c_468_n 0.00155078f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_225 N_B2_c_282_n N_A_251_74#_c_468_n 0.00217387f $X=2.74 $Y=1.515 $X2=0 $Y2=0
cc_226 N_B2_M1006_g N_A_251_74#_c_471_n 0.0152406f $X=2.68 $Y=0.69 $X2=0 $Y2=0
cc_227 N_B1_M1004_g N_VPWR_c_380_n 0.00748953f $X=3.26 $Y=2.34 $X2=0 $Y2=0
cc_228 N_B1_M1004_g N_VPWR_c_382_n 0.0150684f $X=3.26 $Y=2.34 $X2=0 $Y2=0
cc_229 B1 N_VPWR_c_383_n 0.020013f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_230 N_B1_c_324_n N_VPWR_c_383_n 0.00105029f $X=3.57 $Y=1.345 $X2=0 $Y2=0
cc_231 N_B1_M1004_g N_VPWR_c_385_n 0.00492916f $X=3.26 $Y=2.34 $X2=0 $Y2=0
cc_232 N_B1_M1004_g N_VPWR_c_378_n 0.00511769f $X=3.26 $Y=2.34 $X2=0 $Y2=0
cc_233 N_B1_M1000_g N_VGND_c_429_n 0.00290288f $X=3.275 $Y=0.69 $X2=0 $Y2=0
cc_234 N_B1_M1000_g N_VGND_c_430_n 0.00363413f $X=3.275 $Y=0.69 $X2=0 $Y2=0
cc_235 N_B1_M1000_g N_A_251_74#_c_471_n 0.0130694f $X=3.275 $Y=0.69 $X2=0 $Y2=0
cc_236 B1 N_A_251_74#_c_472_n 0.0210212f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_237 N_B1_c_324_n N_A_251_74#_c_472_n 0.00210773f $X=3.57 $Y=1.345 $X2=0 $Y2=0
cc_238 N_X_c_354_n N_VPWR_c_379_n 0.027028f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_239 N_X_c_354_n N_VPWR_c_384_n 0.0158876f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_240 N_X_c_354_n N_VPWR_c_378_n 0.0130823f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_241 N_X_c_352_n N_VGND_c_423_n 0.0277278f $X=0.395 $Y=0.515 $X2=0 $Y2=0
cc_242 N_X_c_352_n N_VGND_c_425_n 0.021034f $X=0.395 $Y=0.515 $X2=0 $Y2=0
cc_243 N_X_c_352_n N_VGND_c_430_n 0.0173537f $X=0.395 $Y=0.515 $X2=0 $Y2=0
cc_244 X N_A_251_74#_c_469_n 0.00259535f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_245 N_VGND_c_423_n N_A_251_74#_c_467_n 0.0255177f $X=0.895 $Y=0.515 $X2=0
+ $Y2=0
cc_246 N_VGND_c_424_n N_A_251_74#_c_467_n 0.018426f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_VGND_c_427_n N_A_251_74#_c_467_n 0.0144922f $X=1.73 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_430_n N_A_251_74#_c_467_n 0.0118826f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_424_n N_A_251_74#_c_468_n 0.0241019f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_250 N_VGND_c_423_n N_A_251_74#_c_469_n 0.00163629f $X=0.895 $Y=0.515 $X2=0
+ $Y2=0
cc_251 N_VGND_c_424_n N_A_251_74#_c_470_n 0.00879395f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_VGND_c_429_n N_A_251_74#_c_470_n 0.0152637f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_430_n N_A_251_74#_c_470_n 0.0121407f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_429_n N_A_251_74#_c_471_n 0.0348412f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_430_n N_A_251_74#_c_471_n 0.0286968f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_429_n N_A_251_74#_c_472_n 0.0116085f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_430_n N_A_251_74#_c_472_n 0.00928389f $X=3.6 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__xor3_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__xor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.180000 1.285000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.771000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.920000 1.350000 5.250000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.875000 1.180000 7.205000 1.685000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.755000 0.400000 9.005000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.120000 0.085000 ;
        RECT 0.625000  0.085000 1.195000 0.490000 ;
        RECT 5.315000  0.085000 5.565000 0.680000 ;
        RECT 8.245000  0.085000 8.575000 1.180000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.120000 3.415000 ;
        RECT 0.770000 2.260000 1.100000 3.245000 ;
        RECT 4.950000 1.950000 5.200000 3.245000 ;
        RECT 8.225000 1.950000 8.555000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.650000 0.445000 0.660000 ;
      RECT 0.085000 0.660000 1.965000 0.830000 ;
      RECT 0.085000 0.830000 0.445000 1.300000 ;
      RECT 0.085000 1.300000 0.255000 2.260000 ;
      RECT 0.085000 2.260000 0.600000 2.980000 ;
      RECT 0.425000 1.470000 0.750000 1.920000 ;
      RECT 0.425000 1.920000 1.625000 1.940000 ;
      RECT 0.425000 1.940000 1.700000 2.090000 ;
      RECT 1.370000 2.090000 1.700000 2.905000 ;
      RECT 1.370000 2.905000 3.895000 3.075000 ;
      RECT 1.455000 1.000000 1.625000 1.920000 ;
      RECT 1.795000 0.830000 1.965000 1.260000 ;
      RECT 1.795000 1.260000 2.760000 1.430000 ;
      RECT 1.930000 1.940000 2.260000 2.565000 ;
      RECT 1.930000 2.565000 3.555000 2.735000 ;
      RECT 2.135000 0.290000 3.215000 0.460000 ;
      RECT 2.135000 0.460000 2.385000 1.090000 ;
      RECT 2.430000 1.430000 2.760000 2.395000 ;
      RECT 2.590000 0.630000 2.850000 1.090000 ;
      RECT 2.590000 1.090000 2.760000 1.260000 ;
      RECT 2.965000 1.875000 3.215000 2.395000 ;
      RECT 3.020000 0.460000 3.215000 1.875000 ;
      RECT 3.385000 0.255000 5.145000 0.425000 ;
      RECT 3.385000 0.425000 3.555000 2.565000 ;
      RECT 3.725000 0.595000 4.805000 0.765000 ;
      RECT 3.725000 0.765000 3.895000 1.435000 ;
      RECT 3.725000 1.435000 4.055000 1.735000 ;
      RECT 3.725000 1.905000 4.395000 2.755000 ;
      RECT 3.725000 2.755000 3.895000 2.905000 ;
      RECT 4.065000 0.935000 4.395000 1.265000 ;
      RECT 4.225000 1.265000 4.395000 1.905000 ;
      RECT 4.580000 0.765000 4.805000 1.130000 ;
      RECT 4.580000 1.130000 4.750000 2.980000 ;
      RECT 4.975000 0.425000 5.145000 0.850000 ;
      RECT 4.975000 0.850000 6.025000 1.020000 ;
      RECT 5.405000 1.950000 5.625000 1.990000 ;
      RECT 5.405000 1.990000 5.855000 2.840000 ;
      RECT 5.420000 1.190000 6.365000 1.360000 ;
      RECT 5.420000 1.360000 5.625000 1.950000 ;
      RECT 5.775000 0.255000 7.645000 0.425000 ;
      RECT 5.775000 0.425000 6.025000 0.850000 ;
      RECT 5.805000 1.530000 6.195000 1.820000 ;
      RECT 6.025000 1.820000 6.195000 2.905000 ;
      RECT 6.025000 2.905000 7.605000 3.075000 ;
      RECT 6.195000 0.595000 7.305000 0.765000 ;
      RECT 6.195000 0.765000 6.365000 1.190000 ;
      RECT 6.365000 1.550000 6.705000 2.735000 ;
      RECT 6.535000 0.935000 6.705000 1.550000 ;
      RECT 6.875000 1.855000 7.645000 2.025000 ;
      RECT 6.875000 2.025000 7.205000 2.735000 ;
      RECT 6.885000 0.765000 7.305000 0.925000 ;
      RECT 7.435000 2.195000 7.985000 2.525000 ;
      RECT 7.435000 2.525000 7.605000 2.905000 ;
      RECT 7.475000 0.425000 7.645000 1.855000 ;
      RECT 7.815000 0.400000 8.065000 0.860000 ;
      RECT 7.815000 0.860000 7.985000 2.195000 ;
      RECT 8.255000 1.350000 8.585000 1.780000 ;
    LAYER mcon ;
      RECT 3.035000 1.580000 3.205000 1.750000 ;
      RECT 5.435000 1.580000 5.605000 1.750000 ;
      RECT 6.395000 1.580000 6.565000 1.750000 ;
      RECT 8.315000 1.580000 8.485000 1.750000 ;
    LAYER met1 ;
      RECT 2.975000 1.550000 3.265000 1.595000 ;
      RECT 2.975000 1.595000 5.665000 1.735000 ;
      RECT 2.975000 1.735000 3.265000 1.780000 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 6.335000 1.550000 6.625000 1.595000 ;
      RECT 6.335000 1.595000 8.545000 1.735000 ;
      RECT 6.335000 1.735000 6.625000 1.780000 ;
      RECT 8.255000 1.550000 8.545000 1.595000 ;
      RECT 8.255000 1.735000 8.545000 1.780000 ;
  END
END sky130_fd_sc_ms__xor3_1

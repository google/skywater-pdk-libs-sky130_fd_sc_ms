* File: sky130_fd_sc_ms__a21o_2.spice
* Created: Wed Sep  2 11:51:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21o_2.pex.spice"
.subckt sky130_fd_sc_ms__a21o_2  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_84_244#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1003_d N_A_84_244#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2442 PD=1.02 PS=1.4 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1004 N_A_84_244#_M1004_d N_B1_M1004_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2442 PD=1.02 PS=1.4 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 A_484_74# N_A1_M1008_g N_A_84_244#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_484_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75002.3 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_84_244#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1002 N_X_M1001_d N_A_84_244#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1007 N_A_404_392#_M1007_d N_B1_M1007_g N_A_84_244#_M1007_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_404_392#_M1007_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_404_392#_M1000_d N_A2_M1000_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__a21o_2.pxi.spice"
*
.ends
*
*

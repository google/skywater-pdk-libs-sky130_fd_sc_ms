* NGSPICE file created from sky130_fd_sc_ms__dfrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_1656_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.33593e+12p ps=1.182e+07u
M1001 a_493_387# a_299_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.262e+11p pd=2.14e+06u as=0p ps=0u
M1002 a_821_138# a_493_387# a_701_463# VNB nlowvt w=420000u l=150000u
+  ad=9.03e+10p pd=1.27e+06u as=1.407e+11p ps=1.51e+06u
M1003 VGND a_1867_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_1266_74# a_299_387# a_833_400# VPB pshort w=1e+06u l=180000u
+  ad=4.39e+11p pd=3.4e+06u as=3.5125e+11p ps=2.95e+06u
M1005 VPWR a_1867_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=1.82245e+12p pd=1.716e+07u as=3.64e+11p ps=2.89e+06u
M1006 VGND RESET_B a_894_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_701_463# a_299_387# a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.541e+11p ps=2.89e+06u
M1008 VPWR a_833_400# a_791_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 VGND RESET_B a_117_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_1471_493# a_493_387# a_1266_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_1867_409# a_1266_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 a_894_138# a_833_400# a_821_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_1518_203# a_1476_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1014 a_701_463# a_493_387# a_30_78# VPB pshort w=420000u l=180000u
+  ad=2.31e+11p pd=2.78e+06u as=2.31e+11p ps=2.78e+06u
M1015 VPWR a_1518_203# a_1471_493# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1476_81# a_299_387# a_1266_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.58e+11p ps=3.28e+06u
M1017 a_1518_203# a_1266_74# a_1656_81# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1018 a_30_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR RESET_B a_30_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1518_203# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1021 VPWR CLK a_299_387# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.1375e+11p ps=2.92e+06u
M1022 a_791_463# a_299_387# a_701_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_299_387# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.45475e+11p ps=2.15e+06u
M1024 VPWR a_1266_74# a_1518_203# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_493_387# a_299_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1026 a_117_78# D a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1266_74# a_493_387# a_833_400# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.921e+11p ps=2.81e+06u
M1028 a_1867_409# a_1266_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1029 a_833_400# a_701_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_701_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_833_400# a_701_463# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o32a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__o32a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 1.350000 2.315000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.855000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.180000 4.685000 2.890000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.350000 3.715000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.960000 1.050000 1.130000 ;
        RECT 0.535000 1.130000 0.705000 1.820000 ;
        RECT 0.535000 1.820000 0.895000 2.980000 ;
        RECT 0.720000 0.350000 1.050000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.085000 0.540000 0.790000 ;
      RECT 0.115000  0.790000 0.365000 1.140000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.875000  1.320000 1.235000 1.650000 ;
      RECT 1.065000  1.650000 1.235000 1.950000 ;
      RECT 1.065000  1.950000 4.185000 2.120000 ;
      RECT 1.065000  2.290000 1.600000 3.245000 ;
      RECT 1.220000  0.085000 1.550000 1.130000 ;
      RECT 1.720000  0.350000 2.050000 1.010000 ;
      RECT 1.720000  1.010000 3.050000 1.180000 ;
      RECT 2.220000  0.085000 2.550000 0.840000 ;
      RECT 2.675000  2.120000 3.110000 2.880000 ;
      RECT 2.720000  0.350000 4.615000 0.520000 ;
      RECT 2.720000  0.520000 3.050000 1.010000 ;
      RECT 3.220000  0.715000 4.185000 1.045000 ;
      RECT 3.815000  2.290000 4.145000 3.245000 ;
      RECT 4.015000  1.045000 4.185000 1.950000 ;
      RECT 4.355000  0.520000 4.615000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ms__o32a_2
END LIBRARY

* File: sky130_fd_sc_ms__o21bai_4.pex.spice
* Created: Wed Sep  2 12:22:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21BAI_4%A1 3 7 11 15 19 23 25 29 33 35 36 37 38 39
+ 57
r82 56 57 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.41 $Y=1.515 $X2=1.5
+ $Y2=1.515
r83 55 56 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.41 $Y2=1.515
r84 53 55 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.265 $Y=1.515
+ $X2=1.405 $Y2=1.515
r85 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r86 51 53 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=0.975 $Y=1.515
+ $X2=1.265 $Y2=1.515
r87 50 51 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.975 $Y2=1.515
r88 48 50 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.96 $Y2=1.515
r89 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r90 46 48 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.515
+ $X2=0.585 $Y2=1.515
r91 44 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.51 $Y2=1.515
r92 39 54 11.1224 $w=4.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.265 $Y2=1.565
r93 38 54 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r94 37 38 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r95 37 49 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r96 36 49 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r97 31 35 18.8402 $w=1.65e-07 $l=7.74597e-08 $layer=POLY_cond $X=1.86 $Y=1.5
+ $X2=1.855 $Y2=1.425
r98 31 33 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=1.86 $Y=1.5 $X2=1.86
+ $Y2=2.4
r99 27 35 18.8402 $w=1.65e-07 $l=8.44097e-08 $layer=POLY_cond $X=1.835 $Y=1.35
+ $X2=1.855 $Y2=1.425
r100 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.835 $Y=1.35
+ $X2=1.835 $Y2=0.74
r101 25 35 6.66866 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=1.76 $Y=1.425
+ $X2=1.855 $Y2=1.425
r102 25 57 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.76 $Y=1.425
+ $X2=1.5 $Y2=1.425
r103 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.405 $Y2=1.515
r104 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.405 $Y2=0.74
r105 17 56 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.68
+ $X2=1.41 $Y2=1.515
r106 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.41 $Y=1.68
+ $X2=1.41 $Y2=2.4
r107 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.35
+ $X2=0.975 $Y2=1.515
r108 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.975 $Y=1.35
+ $X2=0.975 $Y2=0.74
r109 9 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=1.515
r110 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=2.4
r111 5 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.68
+ $X2=0.51 $Y2=1.515
r112 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.51 $Y=1.68 $X2=0.51
+ $Y2=2.4
r113 1 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r114 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%A2 3 7 9 13 17 21 25 29 33 35 36 37 38 52
c97 13 0 1.44963e-19 $X=2.695 $Y=0.74
c98 7 0 1.88192e-19 $X=2.31 $Y=2.4
r99 52 53 0.734756 $w=3.28e-07 $l=5e-09 $layer=POLY_cond $X=3.71 $Y=1.515
+ $X2=3.715 $Y2=1.515
r100 50 52 36.003 $w=3.28e-07 $l=2.45e-07 $layer=POLY_cond $X=3.465 $Y=1.515
+ $X2=3.71 $Y2=1.515
r101 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.515 $X2=3.465 $Y2=1.515
r102 48 50 37.4726 $w=3.28e-07 $l=2.55e-07 $layer=POLY_cond $X=3.21 $Y=1.515
+ $X2=3.465 $Y2=1.515
r103 47 48 12.4909 $w=3.28e-07 $l=8.5e-08 $layer=POLY_cond $X=3.125 $Y=1.515
+ $X2=3.21 $Y2=1.515
r104 45 47 49.9634 $w=3.28e-07 $l=3.4e-07 $layer=POLY_cond $X=2.785 $Y=1.515
+ $X2=3.125 $Y2=1.515
r105 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.515 $X2=2.785 $Y2=1.515
r106 43 45 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=2.76 $Y=1.515
+ $X2=2.785 $Y2=1.515
r107 42 43 9.55183 $w=3.28e-07 $l=6.5e-08 $layer=POLY_cond $X=2.695 $Y=1.515
+ $X2=2.76 $Y2=1.515
r108 38 51 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.465 $Y2=1.565
r109 37 51 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.465 $Y2=1.565
r110 37 46 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.785 $Y2=1.565
r111 36 46 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.785 $Y2=1.565
r112 31 53 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.715 $Y=1.35
+ $X2=3.715 $Y2=1.515
r113 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.715 $Y=1.35
+ $X2=3.715 $Y2=0.74
r114 27 52 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.68
+ $X2=3.71 $Y2=1.515
r115 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.71 $Y=1.68
+ $X2=3.71 $Y2=2.4
r116 23 48 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.68
+ $X2=3.21 $Y2=1.515
r117 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.21 $Y=1.68
+ $X2=3.21 $Y2=2.4
r118 19 47 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.125 $Y2=1.515
r119 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.125 $Y2=0.74
r120 15 43 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.68
+ $X2=2.76 $Y2=1.515
r121 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.76 $Y=1.68
+ $X2=2.76 $Y2=2.4
r122 11 42 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=2.695 $Y2=1.515
r123 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=2.695 $Y2=0.74
r124 10 35 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=2.4 $Y=1.425
+ $X2=2.295 $Y2=1.425
r125 9 42 25.362 $w=3.28e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.62 $Y=1.425
+ $X2=2.695 $Y2=1.515
r126 9 10 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.62 $Y=1.425
+ $X2=2.4 $Y2=1.425
r127 5 35 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.31 $Y=1.5
+ $X2=2.295 $Y2=1.425
r128 5 7 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=2.31 $Y=1.5 $X2=2.31
+ $Y2=2.4
r129 1 35 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=2.265 $Y=1.35
+ $X2=2.295 $Y2=1.425
r130 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.265 $Y=1.35
+ $X2=2.265 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%A_828_48# 1 2 9 13 17 21 25 29 31 40 41 43
+ 44 47 51 53 64
c116 64 0 2.90942e-20 $X=5.645 $Y=1.515
r117 61 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.145 $Y=1.515
+ $X2=5.235 $Y2=1.515
r118 60 61 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.77 $Y=1.515
+ $X2=5.145 $Y2=1.515
r119 59 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=4.645 $Y=1.515
+ $X2=4.77 $Y2=1.515
r120 49 51 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=6.45 $Y=1.11
+ $X2=6.45 $Y2=0.665
r121 45 47 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=6.43 $Y=2.12
+ $X2=6.43 $Y2=2.265
r122 43 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.305 $Y=2.035
+ $X2=6.43 $Y2=2.12
r123 43 44 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.305 $Y=2.035
+ $X2=5.965 $Y2=2.035
r124 42 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=1.195
+ $X2=5.88 $Y2=1.195
r125 41 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.325 $Y=1.195
+ $X2=6.45 $Y2=1.11
r126 41 42 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.325 $Y=1.195
+ $X2=5.965 $Y2=1.195
r127 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.88 $Y=1.95
+ $X2=5.965 $Y2=2.035
r128 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.88 $Y=1.68
+ $X2=5.88 $Y2=1.95
r129 38 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.555 $Y=1.515
+ $X2=5.645 $Y2=1.515
r130 38 62 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=5.555 $Y=1.515
+ $X2=5.235 $Y2=1.515
r131 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.555
+ $Y=1.515 $X2=5.555 $Y2=1.515
r132 34 59 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.535 $Y=1.515
+ $X2=4.645 $Y2=1.515
r133 34 56 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=4.535 $Y=1.515
+ $X2=4.215 $Y2=1.515
r134 33 37 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=4.535 $Y=1.515
+ $X2=5.555 $Y2=1.515
r135 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.535
+ $Y=1.515 $X2=4.535 $Y2=1.515
r136 31 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=1.515
+ $X2=5.88 $Y2=1.68
r137 31 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.88 $Y=1.515
+ $X2=5.88 $Y2=1.195
r138 31 37 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.795 $Y=1.515
+ $X2=5.555 $Y2=1.515
r139 27 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.645 $Y=1.35
+ $X2=5.645 $Y2=1.515
r140 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.645 $Y=1.35
+ $X2=5.645 $Y2=0.74
r141 23 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=1.68
+ $X2=5.235 $Y2=1.515
r142 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.235 $Y=1.68
+ $X2=5.235 $Y2=2.4
r143 19 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.35
+ $X2=5.145 $Y2=1.515
r144 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.145 $Y=1.35
+ $X2=5.145 $Y2=0.74
r145 15 60 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.68
+ $X2=4.77 $Y2=1.515
r146 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.77 $Y=1.68
+ $X2=4.77 $Y2=2.4
r147 11 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.645 $Y=1.35
+ $X2=4.645 $Y2=1.515
r148 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.645 $Y=1.35
+ $X2=4.645 $Y2=0.74
r149 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.215 $Y=1.35
+ $X2=4.215 $Y2=1.515
r150 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.215 $Y=1.35
+ $X2=4.215 $Y2=0.74
r151 2 47 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.335
+ $Y=2.12 $X2=6.47 $Y2=2.265
r152 1 51 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.345
+ $Y=0.52 $X2=6.49 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%B1_N 3 5 7 11 13 14
c38 5 0 1.36199e-19 $X=6.695 $Y=1.78
r39 17 19 40.4029 $w=3.4e-07 $l=2.85e-07 $layer=POLY_cond $X=6.245 $Y=1.66
+ $X2=6.53 $Y2=1.66
r40 13 14 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.96 $Y2=1.615
r41 13 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.615 $X2=6.53 $Y2=1.615
r42 9 22 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.705 $Y=1.45
+ $X2=6.705 $Y2=1.66
r43 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.705 $Y=1.45
+ $X2=6.705 $Y2=0.89
r44 5 22 1.41765 $w=3.4e-07 $l=1e-08 $layer=POLY_cond $X=6.695 $Y=1.66 $X2=6.705
+ $Y2=1.66
r45 5 19 23.3912 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.66
+ $X2=6.53 $Y2=1.66
r46 5 7 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=6.695 $Y=1.78
+ $X2=6.695 $Y2=2.54
r47 1 17 17.6285 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=6.245 $Y=1.87
+ $X2=6.245 $Y2=1.66
r48 1 3 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=6.245 $Y=1.87
+ $X2=6.245 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%A_28_368# 1 2 3 4 5 16 18 20 24 26 28 32 33
+ 36 38 42 47 50
c75 42 0 2.90942e-20 $X=3.985 $Y=2.375
r76 40 42 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.985 $Y=2.905
+ $X2=3.985 $Y2=2.375
r77 39 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=2.99
+ $X2=2.985 $Y2=2.99
r78 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.82 $Y=2.99
+ $X2=3.985 $Y2=2.905
r79 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.82 $Y=2.99
+ $X2=3.15 $Y2=2.99
r80 34 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=2.905
+ $X2=2.985 $Y2=2.99
r81 34 36 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.985 $Y=2.905
+ $X2=2.985 $Y2=2.455
r82 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=2.99
+ $X2=2.985 $Y2=2.99
r83 32 33 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.82 $Y=2.99
+ $X2=2.17 $Y2=2.99
r84 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=2.905
+ $X2=2.17 $Y2=2.99
r85 29 31 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.085 $Y=2.905
+ $X2=2.085 $Y2=2.4
r86 28 49 3.40825 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.085 $Y=2.12
+ $X2=2.085 $Y2=1.97
r87 28 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.085 $Y=2.12
+ $X2=2.085 $Y2=2.4
r88 27 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.27 $Y=2.035
+ $X2=1.145 $Y2=2.035
r89 26 49 3.40825 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=2 $Y=2.035
+ $X2=2.085 $Y2=1.97
r90 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2 $Y=2.035 $X2=1.27
+ $Y2=2.035
r91 22 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.12
+ $X2=1.145 $Y2=2.035
r92 22 24 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=1.145 $Y=2.12
+ $X2=1.145 $Y2=2.44
r93 21 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.37 $Y=2.035
+ $X2=0.245 $Y2=2.035
r94 20 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.145 $Y2=2.035
r95 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.37 $Y2=2.035
r96 16 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.035
r97 16 18 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.44
r98 5 42 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=3.8
+ $Y=1.84 $X2=3.985 $Y2=2.375
r99 4 36 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=1.84 $X2=2.985 $Y2=2.455
r100 3 49 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.085 $Y2=1.985
r101 3 31 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=1.95
+ $Y=1.84 $X2=2.085 $Y2=2.4
r102 2 47 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.035
r103 2 24 300 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.44
r104 1 45 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.035
r105 1 18 300 $w=1.7e-07 $l=6.68581e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%VPWR 1 2 3 4 5 18 22 26 30 32 34 37 38 39
+ 41 46 58 62 68 71 74 78
c90 22 0 1.88192e-19 $X=1.635 $Y=2.455
r91 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r92 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r93 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 66 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r96 66 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r97 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 63 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.105 $Y=3.33
+ $X2=5.98 $Y2=3.33
r99 63 65 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=3.33
+ $X2=6.48 $Y2=3.33
r100 62 77 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.977 $Y2=3.33
r101 62 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.48 $Y2=3.33
r102 61 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r103 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r104 58 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.855 $Y=3.33
+ $X2=5.98 $Y2=3.33
r105 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.855 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r108 54 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 53 56 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r111 51 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=1.635 $Y2=3.33
r112 51 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 50 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r116 47 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.695 $Y2=3.33
r117 47 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 46 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=3.33
+ $X2=1.635 $Y2=3.33
r119 46 49 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.47 $Y=3.33 $X2=1.2
+ $Y2=3.33
r120 44 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r122 41 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.695 $Y2=3.33
r123 41 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 39 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 39 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 37 56 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.91 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=3.33
+ $X2=4.995 $Y2=3.33
r128 36 60 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r129 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=4.995 $Y2=3.33
r130 32 77 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.977 $Y2=3.33
r131 32 34 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.265
r132 28 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=3.245
+ $X2=5.98 $Y2=3.33
r133 28 30 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.98 $Y=3.245
+ $X2=5.98 $Y2=2.455
r134 24 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=3.245
+ $X2=4.995 $Y2=3.33
r135 24 26 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.995 $Y=3.245
+ $X2=4.995 $Y2=2.355
r136 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=3.33
r137 20 22 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=2.455
r138 16 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r139 16 18 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.455
r140 5 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.785
+ $Y=2.12 $X2=6.92 $Y2=2.265
r141 4 30 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=5.875
+ $Y=2.12 $X2=6.02 $Y2=2.455
r142 3 26 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.86
+ $Y=1.84 $X2=4.995 $Y2=2.355
r143 2 22 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=2.455
r144 1 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%Y 1 2 3 4 5 6 19 21 23 27 29 31 35 39 41 42
+ 43 47 49 51 56 62 64 67 68
r103 67 68 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.665
r104 61 68 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.08 $Y=1.95
+ $X2=4.08 $Y2=1.665
r105 61 62 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.95
+ $X2=4.08 $Y2=2.035
r106 58 67 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.18
+ $X2=4.08 $Y2=1.295
r107 49 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.46 $Y=2.02 $X2=5.46
+ $Y2=1.935
r108 49 51 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=5.46 $Y=2.02
+ $X2=5.46 $Y2=2.815
r109 45 47 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.43 $Y=1.01
+ $X2=5.43 $Y2=0.86
r110 44 64 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=4.71 $Y=1.935
+ $X2=4.545 $Y2=1.985
r111 43 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.295 $Y=1.935
+ $X2=5.46 $Y2=1.935
r112 43 44 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.295 $Y=1.935
+ $X2=4.71 $Y2=1.935
r113 41 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.265 $Y=1.095
+ $X2=5.43 $Y2=1.01
r114 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.265 $Y=1.095
+ $X2=4.595 $Y2=1.095
r115 37 64 0.89609 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=4.545 $Y=2.12
+ $X2=4.545 $Y2=1.985
r116 37 39 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.545 $Y=2.12
+ $X2=4.545 $Y2=2.815
r117 33 42 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=1.095
+ $X2=4.595 $Y2=1.095
r118 33 58 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=1.095
+ $X2=4.08 $Y2=1.095
r119 33 35 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.43 $Y=1.01
+ $X2=4.43 $Y2=0.82
r120 32 62 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.195 $Y=2.035
+ $X2=4.08 $Y2=2.035
r121 31 64 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=4.38 $Y=2.035
+ $X2=4.545 $Y2=1.985
r122 31 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.38 $Y=2.035
+ $X2=4.195 $Y2=2.035
r123 30 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.65 $Y=2.035
+ $X2=3.485 $Y2=2.035
r124 29 62 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.965 $Y=2.035
+ $X2=4.08 $Y2=2.035
r125 29 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.965 $Y=2.035
+ $X2=3.65 $Y2=2.035
r126 25 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=2.12
+ $X2=3.485 $Y2=2.035
r127 25 27 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.485 $Y=2.12
+ $X2=3.485 $Y2=2.57
r128 24 54 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.495 $Y2=2.035
r129 23 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=2.035
+ $X2=3.485 $Y2=2.035
r130 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.32 $Y=2.035
+ $X2=2.62 $Y2=2.035
r131 19 54 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=2.12
+ $X2=2.495 $Y2=2.035
r132 19 21 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.495 $Y=2.12
+ $X2=2.495 $Y2=2.57
r133 6 66 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.84 $X2=5.46 $Y2=2.015
r134 6 51 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.84 $X2=5.46 $Y2=2.815
r135 5 64 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.545 $Y2=2.015
r136 5 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.545 $Y2=2.815
r137 4 56 600 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.84 $X2=3.485 $Y2=2.035
r138 4 27 600 $w=1.7e-07 $l=8.17282e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.84 $X2=3.485 $Y2=2.57
r139 3 54 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.84 $X2=2.535 $Y2=2.035
r140 3 21 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.84 $X2=2.535 $Y2=2.57
r141 2 47 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.37 $X2=5.43 $Y2=0.86
r142 1 35 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=4.29
+ $Y=0.37 $X2=4.43 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%A_27_74# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 42 45 46 51 52 53 56 58 62 64 65 66 67
c114 42 0 1.44963e-19 $X=2.91 $Y=0.515
r115 60 62 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.93 $Y=0.425
+ $X2=5.93 $Y2=0.515
r116 59 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=0.34
+ $X2=4.93 $Y2=0.34
r117 58 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.765 $Y=0.34
+ $X2=5.93 $Y2=0.425
r118 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.765 $Y=0.34
+ $X2=5.095 $Y2=0.34
r119 54 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=0.425
+ $X2=4.93 $Y2=0.34
r120 54 56 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.93 $Y=0.425
+ $X2=4.93 $Y2=0.635
r121 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0.34
+ $X2=4.93 $Y2=0.34
r122 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.765 $Y=0.34
+ $X2=4.095 $Y2=0.34
r123 49 51 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=3.93 $Y=0.67
+ $X2=3.93 $Y2=0.595
r124 48 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.93 $Y=0.425
+ $X2=4.095 $Y2=0.34
r125 48 51 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.93 $Y=0.425
+ $X2=3.93 $Y2=0.595
r126 47 66 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.075 $Y=0.755
+ $X2=2.95 $Y2=0.755
r127 46 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.765 $Y=0.755
+ $X2=3.93 $Y2=0.67
r128 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.765 $Y=0.755
+ $X2=3.075 $Y2=0.755
r129 44 66 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.84
+ $X2=2.95 $Y2=0.755
r130 44 45 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.95 $Y=0.84
+ $X2=2.95 $Y2=1.01
r131 40 66 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.67
+ $X2=2.95 $Y2=0.755
r132 40 42 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.95 $Y=0.67
+ $X2=2.95 $Y2=0.515
r133 39 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=1.095
+ $X2=2.05 $Y2=1.095
r134 38 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.825 $Y=1.095
+ $X2=2.95 $Y2=1.01
r135 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.825 $Y=1.095
+ $X2=2.135 $Y2=1.095
r136 34 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.05 $Y2=1.095
r137 34 36 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.05 $Y2=0.515
r138 33 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=1.095
+ $X2=1.19 $Y2=1.095
r139 32 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=1.095
+ $X2=2.05 $Y2=1.095
r140 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.965 $Y=1.095
+ $X2=1.275 $Y2=1.095
r141 28 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=1.01
+ $X2=1.19 $Y2=1.095
r142 28 30 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.19 $Y=1.01
+ $X2=1.19 $Y2=0.515
r143 26 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=1.095
+ $X2=1.19 $Y2=1.095
r144 26 27 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.105 $Y=1.095
+ $X2=0.365 $Y2=1.095
r145 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r146 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r147 7 62 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.72
+ $Y=0.37 $X2=5.93 $Y2=0.515
r148 6 56 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.37 $X2=4.93 $Y2=0.635
r149 5 51 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.79
+ $Y=0.37 $X2=3.93 $Y2=0.595
r150 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.77
+ $Y=0.37 $X2=2.91 $Y2=0.515
r151 3 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.91
+ $Y=0.37 $X2=2.05 $Y2=0.515
r152 2 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.05
+ $Y=0.37 $X2=1.19 $Y2=0.515
r153 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_4%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 40
+ 41 42 44 49 61 69 72 76
c97 34 0 1.36199e-19 $X=6.92 $Y=0.665
r98 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r99 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r100 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 67 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r102 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r103 63 66 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r104 61 75 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.977 $Y2=0
r105 61 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.48 $Y2=0
r106 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r107 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r108 57 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r109 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 54 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r111 54 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.16 $Y2=0
r112 53 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r113 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r114 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r115 50 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r116 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r117 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r118 49 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.2
+ $Y2=0
r119 47 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r120 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r121 44 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r122 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r123 42 67 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r124 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r125 42 63 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r126 40 59 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0
+ $X2=3.12 $Y2=0
r127 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r128 39 63 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.6
+ $Y2=0
r129 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r130 37 56 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.16 $Y2=0
r131 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.48
+ $Y2=0
r132 36 59 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=3.12 $Y2=0
r133 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.48
+ $Y2=0
r134 32 75 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r135 32 34 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.665
r136 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r137 28 30 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.335
r138 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0
r139 24 26 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0.675
r140 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r141 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.675
r142 16 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r143 16 18 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.675
r144 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.78
+ $Y=0.52 $X2=6.92 $Y2=0.665
r145 4 30 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.37 $X2=3.42 $Y2=0.335
r146 3 26 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.37 $X2=2.48 $Y2=0.675
r147 2 22 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.62 $Y2=0.675
r148 1 18 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends


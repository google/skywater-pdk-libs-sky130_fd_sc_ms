* File: sky130_fd_sc_ms__xor3_1.spice
* Created: Wed Sep  2 12:34:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xor3_1.pex.spice"
.subckt sky130_fd_sc_ms__xor3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_A_84_108#_M1019_g N_A_27_134#_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.34745 AS=0.1824 PD=1.81 PS=1.85 NRD=91.476 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1000 N_A_84_108#_M1000_d N_A_M1000_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1702 AS=0.34745 PD=1.41 PS=1.81 NRD=0 NRS=91.476 M=1 R=4.26667 SA=75001
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1015 N_A_416_86#_M1015_d N_B_M1015_g N_A_84_108#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.125283 AS=0.1702 PD=1.19547 PS=1.41 NRD=0 NRS=39.54 M=1 R=4.26667
+ SA=75001.1 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1006 N_A_27_134#_M1006_d N_A_452_288#_M1006_g N_A_416_86#_M1015_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.125326 AS=0.082217 PD=0.919245 PS=0.784528 NRD=12.852
+ NRS=20.712 M=1 R=2.8 SA=75002.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_387_392#_M1014_d N_B_M1014_g N_A_27_134#_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.169075 AS=0.190974 PD=1.275 PS=1.40075 NRD=15.468 NRS=36.552 M=1
+ R=4.26667 SA=75002 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1020 N_A_84_108#_M1020_d N_A_452_288#_M1020_g N_A_387_392#_M1014_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2848 AS=0.169075 PD=2.17 PS=1.275 NRD=31.872 NRS=15.468 M=1
+ R=4.26667 SA=75002.4 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_452_288#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3885 AS=0.2035 PD=2.53 PS=2.03 NRD=40.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1016 N_A_1218_396#_M1016_d N_A_1157_298#_M1016_g N_A_387_392#_M1016_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1696 AS=0.176 PD=1.17 PS=1.83 NRD=46.872 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1007 N_A_416_86#_M1007_d N_C_M1007_g N_A_1218_396#_M1016_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.24 AS=0.1696 PD=2.03 PS=1.17 NRD=8.436 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_C_M1017_g N_A_1157_298#_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.1197 PD=0.796552 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_X_M1018_d N_A_1218_396#_M1018_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_84_108#_M1005_g N_A_27_134#_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.235 AS=0.28 PD=1.47 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1002 N_A_84_108#_M1002_d N_A_M1002_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.184674 AS=0.235 PD=1.47283 PS=1.47 NRD=0 NRS=28.565 M=1 R=5.55556
+ SA=90000.8 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1012 N_A_387_392#_M1012_d N_B_M1012_g N_A_84_108#_M1002_d VPB PSHORT L=0.18
+ W=0.84 AD=0.146432 AS=0.155126 PD=1.32243 PS=1.23717 NRD=4.6886 NRS=19.1484
+ M=1 R=4.66667 SA=90001.4 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1008 N_A_27_134#_M1008_d N_A_452_288#_M1008_g N_A_387_392#_M1012_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.0928 AS=0.111568 PD=0.93 PS=1.00757 NRD=4.6098 NRS=7.683
+ M=1 R=3.55556 SA=90001.9 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1009 N_A_416_86#_M1009_d N_B_M1009_g N_A_27_134#_M1008_d VPB PSHORT L=0.18
+ W=0.64 AD=0.120714 AS=0.0928 PD=1.03351 PS=0.93 NRD=24.6053 NRS=0 M=1
+ R=3.55556 SA=90002.3 SB=90001 A=0.1152 P=1.64 MULT=1
MM1010 N_A_84_108#_M1010_d N_A_452_288#_M1010_g N_A_416_86#_M1009_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.4956 AS=0.158436 PD=2.86 PS=1.35649 NRD=52.7566 NRS=0 M=1
+ R=4.66667 SA=90002.2 SB=90000.5 A=0.1512 P=2.04 MULT=1
MM1021 N_VPWR_M1021_d N_B_M1021_g N_A_452_288#_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_1218_396#_M1001_d N_A_1157_298#_M1001_g N_A_416_86#_M1001_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.2415 AS=0.3066 PD=1.415 PS=2.41 NRD=70.3487
+ NRS=18.7544 M=1 R=4.66667 SA=90000.3 SB=90001 A=0.1512 P=2.04 MULT=1
MM1003 N_A_387_392#_M1003_d N_C_M1003_g N_A_1218_396#_M1001_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2856 AS=0.2415 PD=2.36 PS=1.415 NRD=12.8838 NRS=0 M=1 R=4.66667
+ SA=90001 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1013 N_VPWR_M1013_d N_C_M1013_g N_A_1157_298#_M1013_s VPB PSHORT L=0.18 W=0.64
+ AD=0.167564 AS=0.2432 PD=1.18545 PS=2.04 NRD=73.087 NRS=13.8491 M=1 R=3.55556
+ SA=90000.3 SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1004 N_X_M1004_d N_A_1218_396#_M1004_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.293236 PD=2.8 PS=2.07455 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ms__xor3_1.pxi.spice"
*
.ends
*
*

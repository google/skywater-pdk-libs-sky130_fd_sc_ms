* File: sky130_fd_sc_ms__a32oi_4.pxi.spice
* Created: Wed Sep  2 11:56:13 2020
* 
x_PM_SKY130_FD_SC_MS__A32OI_4%B2 N_B2_M1008_g N_B2_M1000_g N_B2_M1007_g
+ N_B2_M1015_g N_B2_M1032_g N_B2_M1010_g N_B2_M1014_g N_B2_M1035_g B2 B2 B2 B2
+ N_B2_c_149_n PM_SKY130_FD_SC_MS__A32OI_4%B2
x_PM_SKY130_FD_SC_MS__A32OI_4%B1 N_B1_M1018_g N_B1_M1009_g N_B1_M1028_g
+ N_B1_M1011_g N_B1_M1033_g N_B1_M1012_g N_B1_M1038_g N_B1_M1013_g B1 B1 B1 B1
+ B1 N_B1_c_228_n PM_SKY130_FD_SC_MS__A32OI_4%B1
x_PM_SKY130_FD_SC_MS__A32OI_4%A1 N_A1_M1016_g N_A1_M1005_g N_A1_M1017_g
+ N_A1_M1029_g N_A1_M1025_g N_A1_M1034_g N_A1_M1031_g N_A1_M1036_g A1 A1 A1
+ N_A1_c_316_n N_A1_c_317_n PM_SKY130_FD_SC_MS__A32OI_4%A1
x_PM_SKY130_FD_SC_MS__A32OI_4%A2 N_A2_M1001_g N_A2_M1002_g N_A2_M1006_g
+ N_A2_M1020_g N_A2_M1022_g N_A2_M1026_g N_A2_M1023_g N_A2_M1030_g A2 A2 A2 A2
+ N_A2_c_397_n PM_SKY130_FD_SC_MS__A32OI_4%A2
x_PM_SKY130_FD_SC_MS__A32OI_4%A3 N_A3_M1003_g N_A3_M1004_g N_A3_M1019_g
+ N_A3_M1024_g N_A3_M1021_g N_A3_M1037_g N_A3_M1027_g N_A3_M1039_g A3 A3 A3 A3
+ N_A3_c_485_n PM_SKY130_FD_SC_MS__A32OI_4%A3
x_PM_SKY130_FD_SC_MS__A32OI_4%A_27_368# N_A_27_368#_M1000_s N_A_27_368#_M1007_s
+ N_A_27_368#_M1014_s N_A_27_368#_M1011_d N_A_27_368#_M1013_d
+ N_A_27_368#_M1017_s N_A_27_368#_M1031_s N_A_27_368#_M1020_s
+ N_A_27_368#_M1030_s N_A_27_368#_M1019_d N_A_27_368#_M1027_d
+ N_A_27_368#_c_563_n N_A_27_368#_c_564_n N_A_27_368#_c_565_n
+ N_A_27_368#_c_660_p N_A_27_368#_c_566_n N_A_27_368#_c_587_n
+ N_A_27_368#_c_567_n N_A_27_368#_c_591_n N_A_27_368#_c_568_n
+ N_A_27_368#_c_668_p N_A_27_368#_c_598_n N_A_27_368#_c_599_n
+ N_A_27_368#_c_601_n N_A_27_368#_c_609_n N_A_27_368#_c_613_n
+ N_A_27_368#_c_618_n N_A_27_368#_c_569_n N_A_27_368#_c_625_n
+ N_A_27_368#_c_570_n N_A_27_368#_c_629_n N_A_27_368#_c_571_n
+ N_A_27_368#_c_643_n N_A_27_368#_c_572_n N_A_27_368#_c_573_n
+ N_A_27_368#_c_574_n N_A_27_368#_c_575_n N_A_27_368#_c_576_n
+ N_A_27_368#_c_577_n N_A_27_368#_c_578_n N_A_27_368#_c_632_n
+ N_A_27_368#_c_634_n N_A_27_368#_c_652_n PM_SKY130_FD_SC_MS__A32OI_4%A_27_368#
x_PM_SKY130_FD_SC_MS__A32OI_4%Y N_Y_M1018_s N_Y_M1033_s N_Y_M1005_s N_Y_M1034_s
+ N_Y_M1000_d N_Y_M1010_d N_Y_M1009_s N_Y_M1012_s N_Y_c_739_n N_Y_c_743_n
+ N_Y_c_731_n N_Y_c_759_n N_Y_c_763_n N_Y_c_732_n N_Y_c_744_n N_Y_c_748_n
+ N_Y_c_733_n N_Y_c_771_n N_Y_c_734_n N_Y_c_776_n N_Y_c_735_n Y Y Y N_Y_c_736_n
+ N_Y_c_737_n PM_SKY130_FD_SC_MS__A32OI_4%Y
x_PM_SKY130_FD_SC_MS__A32OI_4%VPWR N_VPWR_M1016_d N_VPWR_M1025_d N_VPWR_M1002_d
+ N_VPWR_M1026_d N_VPWR_M1003_s N_VPWR_M1021_s N_VPWR_c_853_n N_VPWR_c_854_n
+ N_VPWR_c_855_n N_VPWR_c_856_n N_VPWR_c_857_n N_VPWR_c_858_n N_VPWR_c_859_n
+ N_VPWR_c_860_n N_VPWR_c_861_n N_VPWR_c_862_n N_VPWR_c_863_n N_VPWR_c_864_n
+ N_VPWR_c_865_n N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n VPWR
+ N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_852_n N_VPWR_c_872_n
+ PM_SKY130_FD_SC_MS__A32OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A32OI_4%A_27_74# N_A_27_74#_M1008_d N_A_27_74#_M1015_d
+ N_A_27_74#_M1035_d N_A_27_74#_M1028_d N_A_27_74#_M1038_d N_A_27_74#_c_982_n
+ N_A_27_74#_c_983_n N_A_27_74#_c_984_n N_A_27_74#_c_985_n N_A_27_74#_c_986_n
+ N_A_27_74#_c_987_n N_A_27_74#_c_988_n N_A_27_74#_c_989_n N_A_27_74#_c_990_n
+ N_A_27_74#_c_991_n N_A_27_74#_c_992_n PM_SKY130_FD_SC_MS__A32OI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__A32OI_4%VGND N_VGND_M1008_s N_VGND_M1032_s N_VGND_M1004_d
+ N_VGND_M1024_d N_VGND_M1039_d N_VGND_c_1056_n N_VGND_c_1057_n N_VGND_c_1058_n
+ N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n VGND N_VGND_c_1062_n
+ N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n
+ N_VGND_c_1067_n N_VGND_c_1068_n N_VGND_c_1069_n N_VGND_c_1070_n
+ N_VGND_c_1071_n PM_SKY130_FD_SC_MS__A32OI_4%VGND
x_PM_SKY130_FD_SC_MS__A32OI_4%A_868_74# N_A_868_74#_M1005_d N_A_868_74#_M1029_d
+ N_A_868_74#_M1036_d N_A_868_74#_M1006_d N_A_868_74#_M1023_d
+ N_A_868_74#_c_1168_n N_A_868_74#_c_1169_n N_A_868_74#_c_1170_n
+ PM_SKY130_FD_SC_MS__A32OI_4%A_868_74#
x_PM_SKY130_FD_SC_MS__A32OI_4%A_1313_74# N_A_1313_74#_M1001_s
+ N_A_1313_74#_M1022_s N_A_1313_74#_M1004_s N_A_1313_74#_M1037_s
+ N_A_1313_74#_c_1208_n N_A_1313_74#_c_1209_n N_A_1313_74#_c_1210_n
+ N_A_1313_74#_c_1211_n N_A_1313_74#_c_1212_n N_A_1313_74#_c_1213_n
+ N_A_1313_74#_c_1214_n N_A_1313_74#_c_1215_n
+ PM_SKY130_FD_SC_MS__A32OI_4%A_1313_74#
cc_1 VNB N_B2_M1008_g 0.0336211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1015_g 0.0234867f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_B2_M1032_g 0.0234201f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_4 VNB N_B2_M1035_g 0.0245585f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_5 VNB B2 0.0166475f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_B2_c_149_n 0.0775011f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_7 VNB N_B1_M1018_g 0.022921f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_B1_M1028_g 0.0232068f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_9 VNB N_B1_M1033_g 0.0231908f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_10 VNB N_B1_M1038_g 0.030436f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_11 VNB B1 0.0107199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_228_n 0.0816839f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_13 VNB N_A1_M1005_g 0.0318671f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_14 VNB N_A1_M1029_g 0.0242232f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_15 VNB N_A1_M1034_g 0.0233769f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_16 VNB N_A1_M1036_g 0.0238886f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_17 VNB N_A1_c_316_n 0.00260092f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_18 VNB N_A1_c_317_n 0.0814353f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_19 VNB N_A2_M1001_g 0.0238306f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_A2_M1006_g 0.0230765f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_21 VNB N_A2_M1022_g 0.0230833f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_22 VNB N_A2_M1023_g 0.0306791f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_23 VNB A2 0.00526789f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_24 VNB N_A2_c_397_n 0.0807073f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_25 VNB N_A3_M1004_g 0.0305493f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_26 VNB N_A3_M1024_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_27 VNB N_A3_M1037_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_28 VNB N_A3_M1039_g 0.031746f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_29 VNB A3 0.016914f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_30 VNB N_A3_c_485_n 0.0837259f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_31 VNB N_Y_c_731_n 0.00392452f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_32 VNB N_Y_c_732_n 0.0109512f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.515
cc_33 VNB N_Y_c_733_n 0.00229834f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.515
cc_34 VNB N_Y_c_734_n 0.00104729f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_35 VNB N_Y_c_735_n 0.0096783f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_36 VNB N_Y_c_736_n 0.0236767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_737_n 0.00229613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_852_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_982_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_40 VNB N_A_27_74#_c_983_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_984_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.68
cc_42 VNB N_A_27_74#_c_985_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_986_n 0.00822418f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_44 VNB N_A_27_74#_c_987_n 0.0029327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_74#_c_988_n 0.00218829f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_A_27_74#_c_989_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_47 VNB N_A_27_74#_c_990_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_48 VNB N_A_27_74#_c_991_n 0.00240889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_992_n 0.00747294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1056_n 0.00568581f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_51 VNB N_VGND_c_1057_n 0.00544084f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_52 VNB N_VGND_c_1058_n 0.0115972f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_53 VNB N_VGND_c_1059_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_54 VNB N_VGND_c_1060_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1061_n 0.0416027f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_56 VNB N_VGND_c_1062_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1063_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_58 VNB N_VGND_c_1064_n 0.159911f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.515
cc_59 VNB N_VGND_c_1065_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.515
cc_60 VNB N_VGND_c_1066_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1067_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1068_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1069_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1070_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1071_n 0.562946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_868_74#_c_1168_n 0.00799024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_868_74#_c_1169_n 0.00583627f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_68 VNB N_A_868_74#_c_1170_n 0.0171655f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_69 VNB N_A_1313_74#_c_1208_n 0.0180757f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_70 VNB N_A_1313_74#_c_1209_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.425
+ $Y2=0.74
cc_71 VNB N_A_1313_74#_c_1210_n 0.00527187f $X=-0.19 $Y=-0.245 $X2=1.455
+ $Y2=1.68
cc_72 VNB N_A_1313_74#_c_1211_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.905
+ $Y2=1.68
cc_73 VNB N_A_1313_74#_c_1212_n 0.00526132f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_74 VNB N_A_1313_74#_c_1213_n 0.0034448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1313_74#_c_1214_n 0.00114016f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_76 VNB N_A_1313_74#_c_1215_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_77 VPB N_B2_M1000_g 0.025802f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_78 VPB N_B2_M1007_g 0.0201646f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_79 VPB N_B2_M1010_g 0.0196385f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_80 VPB N_B2_M1014_g 0.0212611f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=2.4
cc_81 VPB B2 0.0169834f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_82 VPB N_B2_c_149_n 0.0133123f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_83 VPB N_B1_M1009_g 0.0209262f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_84 VPB N_B1_M1011_g 0.0208009f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_85 VPB N_B1_M1012_g 0.0207967f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_86 VPB N_B1_M1013_g 0.0222043f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=0.74
cc_87 VPB B1 0.0152947f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_B1_c_228_n 0.0174314f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_89 VPB N_A1_M1016_g 0.0226074f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_90 VPB N_A1_M1017_g 0.0210655f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_91 VPB N_A1_M1025_g 0.0215784f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_92 VPB N_A1_M1031_g 0.0229133f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=2.4
cc_93 VPB N_A1_c_316_n 0.00941617f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_94 VPB N_A1_c_317_n 0.0161665f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_95 VPB N_A2_M1002_g 0.0228146f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_96 VPB N_A2_M1020_g 0.0214797f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_97 VPB N_A2_M1026_g 0.0210655f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_98 VPB N_A2_M1030_g 0.0213755f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=0.74
cc_99 VPB A2 0.0125708f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_100 VPB N_A2_c_397_n 0.016157f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_101 VPB N_A3_M1003_g 0.0223126f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_102 VPB N_A3_M1019_g 0.0210572f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_103 VPB N_A3_M1021_g 0.0222099f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_104 VPB N_A3_M1027_g 0.028716f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=2.4
cc_105 VPB A3 0.016582f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_106 VPB N_A3_c_485_n 0.0179538f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_107 VPB N_A_27_368#_c_563_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_108 VPB N_A_27_368#_c_564_n 0.00259172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_368#_c_565_n 0.00971634f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_110 VPB N_A_27_368#_c_566_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_111 VPB N_A_27_368#_c_567_n 0.00241371f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_112 VPB N_A_27_368#_c_568_n 0.00633239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_368#_c_569_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_368#_c_570_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_368#_c_571_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_368#_c_572_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_368#_c_573_n 0.0352219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_368#_c_574_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_368#_c_575_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_368#_c_576_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_368#_c_577_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_27_368#_c_578_n 0.00240256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_Y_c_732_n 0.00369236f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_124 VPB N_VPWR_c_853_n 0.00565985f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.68
cc_125 VPB N_VPWR_c_854_n 0.0083004f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.68
cc_126 VPB N_VPWR_c_855_n 0.00829947f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.35
cc_127 VPB N_VPWR_c_856_n 0.00510895f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_128 VPB N_VPWR_c_857_n 0.00510895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_858_n 0.00903683f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_130 VPB N_VPWR_c_859_n 0.107574f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_131 VPB N_VPWR_c_860_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_132 VPB N_VPWR_c_861_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_133 VPB N_VPWR_c_862_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_134 VPB N_VPWR_c_863_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.515
cc_135 VPB N_VPWR_c_864_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_136 VPB N_VPWR_c_865_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=1.515
cc_137 VPB N_VPWR_c_866_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.515
cc_138 VPB N_VPWR_c_867_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_868_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_140 VPB N_VPWR_c_869_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_870_n 0.0194498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_852_n 0.0927044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_872_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 N_B2_M1035_g N_B1_M1018_g 0.0168335f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_145 N_B2_M1014_g N_B1_M1009_g 0.027833f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_146 B2 B1 0.0289875f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_147 N_B2_c_149_n B1 0.00485343f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_148 B2 N_B1_c_228_n 2.25699e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B2_c_149_n N_B1_c_228_n 0.0168335f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_150 N_B2_M1000_g N_A_27_368#_c_563_n 0.0121621f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_151 N_B2_M1007_g N_A_27_368#_c_563_n 9.34759e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_152 B2 N_A_27_368#_c_563_n 0.0254478f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B2_M1000_g N_A_27_368#_c_564_n 0.012228f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_154 N_B2_M1007_g N_A_27_368#_c_564_n 0.0142904f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_155 N_B2_M1000_g N_A_27_368#_c_565_n 0.00282152f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_156 N_B2_M1010_g N_A_27_368#_c_566_n 0.0140221f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_157 N_B2_M1014_g N_A_27_368#_c_566_n 0.0141884f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_158 N_B2_M1007_g N_Y_c_739_n 0.012931f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_159 N_B2_M1010_g N_Y_c_739_n 0.012931f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_160 B2 N_Y_c_739_n 0.0391869f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B2_c_149_n N_Y_c_739_n 4.89709e-19 $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_162 N_B2_M1014_g N_Y_c_743_n 0.017729f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B2_M1007_g N_Y_c_744_n 0.0105388f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_164 N_B2_M1010_g N_Y_c_744_n 5.73047e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_165 B2 N_Y_c_744_n 0.0244752f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_166 N_B2_c_149_n N_Y_c_744_n 8.32165e-19 $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_167 N_B2_M1007_g N_Y_c_748_n 5.73047e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_168 N_B2_M1010_g N_Y_c_748_n 0.010564f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_169 N_B2_M1014_g N_Y_c_748_n 0.0116773f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_170 B2 N_Y_c_748_n 0.0202798f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_171 N_B2_c_149_n N_Y_c_748_n 5.54777e-19 $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_172 N_B2_M1000_g N_VPWR_c_859_n 0.00333901f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B2_M1007_g N_VPWR_c_859_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B2_M1010_g N_VPWR_c_859_n 0.00333926f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B2_M1014_g N_VPWR_c_859_n 0.00333926f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_176 N_B2_M1000_g N_VPWR_c_852_n 0.00426886f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_177 N_B2_M1007_g N_VPWR_c_852_n 0.00423129f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B2_M1010_g N_VPWR_c_852_n 0.00422687f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B2_M1014_g N_VPWR_c_852_n 0.00423254f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_180 N_B2_M1008_g N_A_27_74#_c_982_n 0.0101077f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B2_M1015_g N_A_27_74#_c_982_n 9.62944e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B2_M1008_g N_A_27_74#_c_983_n 0.0115433f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B2_M1015_g N_A_27_74#_c_983_n 0.0134851f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_184 B2 N_A_27_74#_c_983_n 0.0510636f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_185 N_B2_c_149_n N_A_27_74#_c_983_n 0.00394939f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_186 N_B2_M1008_g N_A_27_74#_c_984_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_187 B2 N_A_27_74#_c_984_n 0.0286342f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B2_M1015_g N_A_27_74#_c_985_n 3.92313e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B2_M1032_g N_A_27_74#_c_985_n 3.92313e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B2_M1032_g N_A_27_74#_c_986_n 0.0134594f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B2_M1035_g N_A_27_74#_c_986_n 0.0185794f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_192 B2 N_A_27_74#_c_986_n 0.0377574f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B2_c_149_n N_A_27_74#_c_986_n 0.00399488f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_194 N_B2_M1035_g N_A_27_74#_c_988_n 0.00109794f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_195 B2 N_A_27_74#_c_990_n 0.0146029f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_B2_c_149_n N_A_27_74#_c_990_n 0.00242817f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_197 N_B2_M1008_g N_VGND_c_1056_n 0.00571035f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_198 N_B2_M1015_g N_VGND_c_1056_n 0.0103415f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_199 N_B2_M1032_g N_VGND_c_1056_n 4.71636e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B2_M1015_g N_VGND_c_1057_n 4.71636e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B2_M1032_g N_VGND_c_1057_n 0.01032f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B2_M1035_g N_VGND_c_1057_n 0.00397166f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B2_M1008_g N_VGND_c_1062_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B2_M1015_g N_VGND_c_1063_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B2_M1032_g N_VGND_c_1063_n 0.00383152f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B2_M1035_g N_VGND_c_1064_n 0.00461464f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B2_M1008_g N_VGND_c_1071_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B2_M1015_g N_VGND_c_1071_n 0.0075754f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B2_M1032_g N_VGND_c_1071_n 0.0075754f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B2_M1035_g N_VGND_c_1071_n 0.00908708f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B1_M1013_g N_A1_M1016_g 0.0161572f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_212 B1 N_A1_c_316_n 0.0305566f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B1_c_228_n N_A1_c_316_n 0.0013644f $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_214 B1 N_A1_c_317_n 0.00200382f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_215 N_B1_c_228_n N_A1_c_317_n 0.0161572f $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_216 N_B1_M1009_g N_A_27_368#_c_587_n 0.00895541f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_217 N_B1_M1011_g N_A_27_368#_c_587_n 5.88728e-19 $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_218 N_B1_M1009_g N_A_27_368#_c_567_n 0.0119307f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_219 N_B1_M1011_g N_A_27_368#_c_567_n 0.0145175f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_220 N_B1_M1012_g N_A_27_368#_c_591_n 0.00895541f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B1_M1013_g N_A_27_368#_c_591_n 5.88728e-19 $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B1_M1012_g N_A_27_368#_c_568_n 0.0119307f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_223 N_B1_M1013_g N_A_27_368#_c_568_n 0.014668f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_224 N_B1_M1009_g N_A_27_368#_c_575_n 0.00211007f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_225 N_B1_M1012_g N_A_27_368#_c_576_n 0.00214324f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_226 N_B1_M1009_g N_Y_c_743_n 0.0145035f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_227 B1 N_Y_c_743_n 0.0331478f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_M1028_g N_Y_c_731_n 0.014265f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_M1033_g N_Y_c_731_n 0.0146892f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_230 B1 N_Y_c_731_n 0.115026f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B1_c_228_n N_Y_c_731_n 0.00707936f $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B1_M1011_g N_Y_c_759_n 0.0132272f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_233 N_B1_M1012_g N_Y_c_759_n 0.0145524f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_234 B1 N_Y_c_759_n 0.046225f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_B1_c_228_n N_Y_c_759_n 7.55656e-19 $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_236 N_B1_M1013_g N_Y_c_763_n 0.0138062f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_237 B1 N_Y_c_763_n 0.0247708f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B1_M1009_g N_Y_c_748_n 4.54422e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_239 N_B1_M1018_g N_Y_c_733_n 0.00904704f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1028_g N_Y_c_733_n 0.00906556f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B1_M1033_g N_Y_c_733_n 9.11723e-19 $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_242 B1 N_Y_c_733_n 0.0276216f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B1_c_228_n N_Y_c_733_n 0.00259156f $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B1_M1011_g N_Y_c_771_n 0.010574f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B1_M1012_g N_Y_c_771_n 4.54422e-19 $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_246 B1 N_Y_c_771_n 0.0246996f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_247 N_B1_c_228_n N_Y_c_771_n 8.55208e-19 $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_248 N_B1_M1038_g N_Y_c_734_n 0.00820324f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B1_M1013_g N_Y_c_776_n 0.0108127f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_250 B1 N_Y_c_776_n 0.0246996f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B1_c_228_n N_Y_c_776_n 8.53086e-19 $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_252 N_B1_M1038_g N_Y_c_736_n 0.00954049f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B1_c_228_n N_Y_c_736_n 0.0055357f $X=3.905 $Y=1.515 $X2=0 $Y2=0
cc_254 N_B1_M1009_g N_VPWR_c_859_n 0.00333896f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_255 N_B1_M1011_g N_VPWR_c_859_n 0.00333926f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B1_M1012_g N_VPWR_c_859_n 0.00333896f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B1_M1013_g N_VPWR_c_859_n 0.00333926f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B1_M1009_g N_VPWR_c_852_n 0.0042374f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_259 N_B1_M1011_g N_VPWR_c_852_n 0.00423664f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B1_M1012_g N_VPWR_c_852_n 0.00423662f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B1_M1013_g N_VPWR_c_852_n 0.00424819f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B1_M1018_g N_A_27_74#_c_986_n 5.7591e-19 $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_263 B1 N_A_27_74#_c_986_n 0.0156959f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_264 N_B1_M1018_g N_A_27_74#_c_987_n 0.0119575f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_265 N_B1_M1028_g N_A_27_74#_c_987_n 0.00934417f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B1_M1033_g N_A_27_74#_c_989_n 0.00805131f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B1_M1038_g N_A_27_74#_c_989_n 0.0092831f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_268 N_B1_M1028_g N_A_27_74#_c_991_n 4.46617e-19 $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B1_M1033_g N_A_27_74#_c_991_n 0.00767662f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B1_M1038_g N_A_27_74#_c_991_n 9.18514e-19 $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_271 N_B1_M1033_g N_A_27_74#_c_992_n 9.18514e-19 $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_272 N_B1_M1038_g N_A_27_74#_c_992_n 0.0087405f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_273 N_B1_M1018_g N_VGND_c_1064_n 0.00278271f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_274 N_B1_M1028_g N_VGND_c_1064_n 0.00278271f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_275 N_B1_M1033_g N_VGND_c_1064_n 0.00279469f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_276 N_B1_M1038_g N_VGND_c_1064_n 0.00279469f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_277 N_B1_M1018_g N_VGND_c_1071_n 0.00353526f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_278 N_B1_M1028_g N_VGND_c_1071_n 0.00354087f $X=2.78 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B1_M1033_g N_VGND_c_1071_n 0.00353176f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_280 N_B1_M1038_g N_VGND_c_1071_n 0.00357517f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B1_M1038_g N_A_868_74#_c_1168_n 0.00378887f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A1_M1036_g N_A2_M1001_g 0.0252537f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A1_M1031_g N_A2_M1002_g 0.0252537f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A1_c_317_n N_A2_c_397_n 0.0252537f $X=6.06 $Y=1.515 $X2=0 $Y2=0
cc_285 N_A1_M1016_g N_A_27_368#_c_568_n 0.00188262f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A1_M1016_g N_A_27_368#_c_598_n 0.00747416f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A1_M1016_g N_A_27_368#_c_599_n 0.0170384f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_288 N_A1_M1017_g N_A_27_368#_c_599_n 0.0129921f $X=5.045 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A1_M1025_g N_A_27_368#_c_601_n 0.0132511f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A1_M1031_g N_A_27_368#_c_601_n 0.0132511f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A1_M1016_g N_A_27_368#_c_577_n 8.39327e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A1_M1017_g N_A_27_368#_c_577_n 0.00867318f $X=5.045 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A1_M1025_g N_A_27_368#_c_577_n 0.00893294f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A1_M1031_g N_A_27_368#_c_577_n 5.52103e-19 $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_295 N_A1_M1025_g N_A_27_368#_c_578_n 5.52103e-19 $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A1_M1031_g N_A_27_368#_c_578_n 0.00893538f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A1_M1016_g N_Y_c_763_n 0.0128349f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A1_M1017_g N_Y_c_763_n 0.0119585f $X=5.045 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A1_M1025_g N_Y_c_763_n 0.0122174f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A1_M1031_g N_Y_c_763_n 0.0172616f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_301 N_A1_c_316_n N_Y_c_763_n 0.0940005f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_302 N_A1_c_317_n N_Y_c_763_n 0.00396338f $X=6.06 $Y=1.515 $X2=0 $Y2=0
cc_303 N_A1_M1036_g N_Y_c_732_n 0.0121716f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A1_c_316_n N_Y_c_732_n 0.0192758f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_305 N_A1_M1016_g N_Y_c_776_n 8.98219e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A1_M1029_g N_Y_c_735_n 0.0122111f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A1_M1034_g N_Y_c_735_n 0.014039f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A1_M1036_g N_Y_c_735_n 0.0177493f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A1_c_316_n N_Y_c_735_n 0.0426866f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_310 N_A1_c_317_n N_Y_c_735_n 0.00640561f $X=6.06 $Y=1.515 $X2=0 $Y2=0
cc_311 N_A1_M1005_g N_Y_c_736_n 0.0138679f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A1_c_316_n N_Y_c_736_n 0.0556202f $X=5.64 $Y=1.515 $X2=0 $Y2=0
cc_313 N_A1_c_317_n N_Y_c_736_n 0.00448128f $X=6.06 $Y=1.515 $X2=0 $Y2=0
cc_314 N_A1_M1029_g N_Y_c_737_n 0.0034533f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A1_M1034_g N_Y_c_737_n 2.36785e-19 $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A1_c_317_n N_Y_c_737_n 0.00456495f $X=6.06 $Y=1.515 $X2=0 $Y2=0
cc_317 N_A1_M1016_g N_VPWR_c_853_n 0.00884319f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_318 N_A1_M1017_g N_VPWR_c_853_n 0.00194999f $X=5.045 $Y=2.4 $X2=0 $Y2=0
cc_319 N_A1_M1025_g N_VPWR_c_854_n 0.00203999f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_320 N_A1_M1031_g N_VPWR_c_854_n 0.00203999f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_321 N_A1_M1016_g N_VPWR_c_859_n 0.00460063f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_322 N_A1_M1017_g N_VPWR_c_861_n 0.005209f $X=5.045 $Y=2.4 $X2=0 $Y2=0
cc_323 N_A1_M1025_g N_VPWR_c_861_n 0.005209f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_324 N_A1_M1031_g N_VPWR_c_863_n 0.005209f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A1_M1016_g N_VPWR_c_852_n 0.00910197f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_326 N_A1_M1017_g N_VPWR_c_852_n 0.00982082f $X=5.045 $Y=2.4 $X2=0 $Y2=0
cc_327 N_A1_M1025_g N_VPWR_c_852_n 0.00982526f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_328 N_A1_M1031_g N_VPWR_c_852_n 0.00982731f $X=6.045 $Y=2.4 $X2=0 $Y2=0
cc_329 N_A1_M1005_g N_A_27_74#_c_992_n 0.00314096f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1005_g N_VGND_c_1064_n 0.00292759f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1029_g N_VGND_c_1064_n 0.00291649f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1034_g N_VGND_c_1064_n 0.00291649f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1036_g N_VGND_c_1064_n 0.00291649f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1005_g N_VGND_c_1071_n 0.00363814f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A1_M1029_g N_VGND_c_1071_n 0.00359779f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A1_M1034_g N_VGND_c_1071_n 0.00359121f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1036_g N_VGND_c_1071_n 0.00359219f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1005_g N_A_868_74#_c_1168_n 0.00792667f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1029_g N_A_868_74#_c_1168_n 8.9082e-19 $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1005_g N_A_868_74#_c_1170_n 0.0114225f $X=4.7 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A1_M1029_g N_A_868_74#_c_1170_n 0.0107985f $X=5.2 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A1_M1034_g N_A_868_74#_c_1170_n 0.010218f $X=5.63 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A1_M1036_g N_A_868_74#_c_1170_n 0.010213f $X=6.06 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A1_M1036_g N_A_1313_74#_c_1212_n 2.90368e-19 $X=6.06 $Y=0.74 $X2=0
+ $Y2=0
cc_345 N_A2_M1030_g N_A3_M1003_g 0.0103658f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_346 A2 N_A3_M1003_g 0.00467145f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_347 A2 A3 0.0278076f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_348 A2 N_A3_c_485_n 0.0105679f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_349 N_A2_c_397_n N_A3_c_485_n 0.0127853f $X=7.995 $Y=1.515 $X2=0 $Y2=0
cc_350 N_A2_M1002_g N_A_27_368#_c_609_n 0.0187797f $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A2_M1020_g N_A_27_368#_c_609_n 0.0148922f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_352 A2 N_A_27_368#_c_609_n 0.0115282f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A2_c_397_n N_A_27_368#_c_609_n 0.00178335f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_354 N_A2_M1002_g N_A_27_368#_c_613_n 7.76211e-19 $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_355 N_A2_M1020_g N_A_27_368#_c_613_n 0.00417445f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_356 N_A2_M1026_g N_A_27_368#_c_613_n 8.84614e-19 $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_357 A2 N_A_27_368#_c_613_n 0.0235495f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_358 N_A2_c_397_n N_A_27_368#_c_613_n 5.48413e-19 $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_359 N_A2_M1002_g N_A_27_368#_c_618_n 7.77834e-19 $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A2_M1020_g N_A_27_368#_c_618_n 0.00343312f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A2_M1026_g N_A_27_368#_c_618_n 0.00351396f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A2_M1030_g N_A_27_368#_c_618_n 4.53616e-19 $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_363 N_A2_M1002_g N_A_27_368#_c_569_n 5.53945e-19 $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_364 N_A2_M1020_g N_A_27_368#_c_569_n 0.00804796f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_365 N_A2_M1026_g N_A_27_368#_c_569_n 0.00635606f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_366 N_A2_M1026_g N_A_27_368#_c_625_n 0.0132272f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_367 N_A2_M1030_g N_A_27_368#_c_625_n 0.0145524f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_368 A2 N_A_27_368#_c_625_n 0.046225f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_369 N_A2_c_397_n N_A_27_368#_c_625_n 7.5354e-19 $X=7.995 $Y=1.515 $X2=0 $Y2=0
cc_370 A2 N_A_27_368#_c_629_n 0.00580317f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A2_M1002_g N_A_27_368#_c_578_n 0.00883034f $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A2_M1020_g N_A_27_368#_c_578_n 5.43435e-19 $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_373 N_A2_M1020_g N_A_27_368#_c_632_n 4.64231e-19 $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_374 N_A2_M1026_g N_A_27_368#_c_632_n 0.00192359f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_375 A2 N_A_27_368#_c_634_n 0.0246997f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_376 N_A2_M1002_g N_Y_c_763_n 0.00534356f $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_377 N_A2_M1001_g N_Y_c_732_n 0.0131859f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_378 A2 N_Y_c_732_n 0.0189002f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_379 N_A2_M1001_g N_Y_c_735_n 0.0030096f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_380 N_A2_M1002_g N_VPWR_c_855_n 0.00206359f $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_381 N_A2_M1020_g N_VPWR_c_855_n 0.00202232f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_382 N_A2_M1026_g N_VPWR_c_856_n 0.00194999f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_383 N_A2_M1030_g N_VPWR_c_856_n 0.0125212f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_384 N_A2_M1002_g N_VPWR_c_863_n 0.0053223f $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_385 N_A2_M1020_g N_VPWR_c_865_n 0.005209f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_386 N_A2_M1026_g N_VPWR_c_865_n 0.005209f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_387 N_A2_M1030_g N_VPWR_c_867_n 0.00460063f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_388 N_A2_M1002_g N_VPWR_c_852_n 0.0101911f $X=6.505 $Y=2.4 $X2=0 $Y2=0
cc_389 N_A2_M1020_g N_VPWR_c_852_n 0.0098244f $X=7.045 $Y=2.4 $X2=0 $Y2=0
cc_390 N_A2_M1026_g N_VPWR_c_852_n 0.00982082f $X=7.495 $Y=2.4 $X2=0 $Y2=0
cc_391 N_A2_M1030_g N_VPWR_c_852_n 0.00909121f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_392 N_A2_M1023_g N_VGND_c_1058_n 0.00708914f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A2_M1001_g N_VGND_c_1064_n 0.00291649f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A2_M1006_g N_VGND_c_1064_n 0.00291649f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A2_M1022_g N_VGND_c_1064_n 0.00291649f $X=7.355 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A2_M1023_g N_VGND_c_1064_n 0.00291649f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A2_M1001_g N_VGND_c_1071_n 0.00359219f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_398 N_A2_M1006_g N_VGND_c_1071_n 0.00359171f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A2_M1022_g N_VGND_c_1071_n 0.00359171f $X=7.355 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A2_M1023_g N_VGND_c_1071_n 0.0036412f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A2_M1022_g N_A_868_74#_c_1169_n 3.85913e-19 $X=7.355 $Y=0.74 $X2=0
+ $Y2=0
cc_402 N_A2_M1023_g N_A_868_74#_c_1169_n 0.00311138f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_403 N_A2_M1001_g N_A_868_74#_c_1170_n 0.0142216f $X=6.49 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A2_M1006_g N_A_868_74#_c_1170_n 0.0106163f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A2_M1022_g N_A_868_74#_c_1170_n 0.010696f $X=7.355 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A2_M1023_g N_A_868_74#_c_1170_n 0.00974906f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_407 N_A2_M1023_g N_A_1313_74#_c_1208_n 0.0103942f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A2_c_397_n N_A_1313_74#_c_1208_n 0.00593111f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_409 N_A2_M1001_g N_A_1313_74#_c_1212_n 0.00669488f $X=6.49 $Y=0.74 $X2=0
+ $Y2=0
cc_410 N_A2_M1006_g N_A_1313_74#_c_1212_n 0.0037133f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_411 N_A2_M1022_g N_A_1313_74#_c_1212_n 3.85091e-19 $X=7.355 $Y=0.74 $X2=0
+ $Y2=0
cc_412 A2 N_A_1313_74#_c_1212_n 0.140642f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_413 N_A2_c_397_n N_A_1313_74#_c_1212_n 0.00389297f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_414 N_A2_M1006_g N_A_1313_74#_c_1213_n 0.0116925f $X=6.92 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A2_M1022_g N_A_1313_74#_c_1213_n 0.0140807f $X=7.355 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A2_c_397_n N_A_1313_74#_c_1213_n 0.0054755f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_417 N_A2_M1023_g N_A_1313_74#_c_1214_n 0.00945167f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_418 N_A3_M1003_g N_A_27_368#_c_570_n 0.0118126f $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A3_M1019_g N_A_27_368#_c_570_n 6.27806e-19 $X=8.995 $Y=2.4 $X2=0 $Y2=0
cc_420 N_A3_M1003_g N_A_27_368#_c_629_n 0.0151488f $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_421 N_A3_M1019_g N_A_27_368#_c_629_n 0.0145524f $X=8.995 $Y=2.4 $X2=0 $Y2=0
cc_422 A3 N_A_27_368#_c_629_n 0.0230473f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_423 N_A3_c_485_n N_A_27_368#_c_629_n 0.00346191f $X=10.05 $Y=1.515 $X2=0
+ $Y2=0
cc_424 N_A3_M1021_g N_A_27_368#_c_571_n 0.0119363f $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_425 N_A3_M1027_g N_A_27_368#_c_571_n 5.9891e-19 $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_426 N_A3_M1021_g N_A_27_368#_c_643_n 0.0135102f $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_427 N_A3_M1027_g N_A_27_368#_c_643_n 0.0135102f $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_428 A3 N_A_27_368#_c_643_n 0.0475502f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_429 N_A3_c_485_n N_A_27_368#_c_643_n 0.00105451f $X=10.05 $Y=1.515 $X2=0
+ $Y2=0
cc_430 N_A3_M1027_g N_A_27_368#_c_572_n 8.84614e-19 $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_431 A3 N_A_27_368#_c_572_n 0.0259449f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_432 N_A3_M1021_g N_A_27_368#_c_573_n 6.02881e-19 $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_433 N_A3_M1027_g N_A_27_368#_c_573_n 0.0121858f $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_434 N_A3_M1003_g N_A_27_368#_c_634_n 8.84614e-19 $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_435 N_A3_M1021_g N_A_27_368#_c_652_n 8.84614e-19 $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_436 A3 N_A_27_368#_c_652_n 0.0246996f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_437 N_A3_c_485_n N_A_27_368#_c_652_n 8.53086e-19 $X=10.05 $Y=1.515 $X2=0
+ $Y2=0
cc_438 N_A3_M1003_g N_VPWR_c_856_n 5.13171e-19 $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_439 N_A3_M1003_g N_VPWR_c_857_n 0.00194999f $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_440 N_A3_M1019_g N_VPWR_c_857_n 0.0125212f $X=8.995 $Y=2.4 $X2=0 $Y2=0
cc_441 N_A3_M1021_g N_VPWR_c_857_n 5.13171e-19 $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_442 N_A3_M1021_g N_VPWR_c_858_n 0.00204877f $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_443 N_A3_M1027_g N_VPWR_c_858_n 0.00342423f $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_444 N_A3_M1003_g N_VPWR_c_867_n 0.005209f $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_445 N_A3_M1019_g N_VPWR_c_869_n 0.00460063f $X=8.995 $Y=2.4 $X2=0 $Y2=0
cc_446 N_A3_M1021_g N_VPWR_c_869_n 0.005209f $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_447 N_A3_M1027_g N_VPWR_c_870_n 0.005209f $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_448 N_A3_M1003_g N_VPWR_c_852_n 0.00982648f $X=8.495 $Y=2.4 $X2=0 $Y2=0
cc_449 N_A3_M1019_g N_VPWR_c_852_n 0.00909043f $X=8.995 $Y=2.4 $X2=0 $Y2=0
cc_450 N_A3_M1021_g N_VPWR_c_852_n 0.00983056f $X=9.495 $Y=2.4 $X2=0 $Y2=0
cc_451 N_A3_M1027_g N_VPWR_c_852_n 0.00986439f $X=10.05 $Y=2.4 $X2=0 $Y2=0
cc_452 N_A3_M1004_g N_VGND_c_1058_n 0.0120602f $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A3_M1024_g N_VGND_c_1058_n 4.71636e-19 $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_454 N_A3_M1004_g N_VGND_c_1059_n 4.71636e-19 $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_455 N_A3_M1024_g N_VGND_c_1059_n 0.0103289f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A3_M1037_g N_VGND_c_1059_n 0.0103289f $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_457 N_A3_M1039_g N_VGND_c_1059_n 4.71636e-19 $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A3_M1037_g N_VGND_c_1061_n 5.67074e-19 $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A3_M1039_g N_VGND_c_1061_n 0.015057f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_460 A3 N_VGND_c_1061_n 0.023775f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_461 N_A3_M1004_g N_VGND_c_1065_n 0.00383152f $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A3_M1024_g N_VGND_c_1065_n 0.00383152f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A3_M1037_g N_VGND_c_1066_n 0.00383152f $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_464 N_A3_M1039_g N_VGND_c_1066_n 0.00383152f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_465 N_A3_M1004_g N_VGND_c_1071_n 0.0075754f $X=8.775 $Y=0.74 $X2=0 $Y2=0
cc_466 N_A3_M1024_g N_VGND_c_1071_n 0.0075754f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A3_M1037_g N_VGND_c_1071_n 0.0075754f $X=9.635 $Y=0.74 $X2=0 $Y2=0
cc_468 N_A3_M1039_g N_VGND_c_1071_n 0.0075754f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A3_M1004_g N_A_868_74#_c_1169_n 7.60322e-19 $X=8.775 $Y=0.74 $X2=0
+ $Y2=0
cc_470 N_A3_M1004_g N_A_1313_74#_c_1208_n 0.0169578f $X=8.775 $Y=0.74 $X2=0
+ $Y2=0
cc_471 A3 N_A_1313_74#_c_1208_n 0.010384f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_472 N_A3_c_485_n N_A_1313_74#_c_1208_n 0.00668938f $X=10.05 $Y=1.515 $X2=0
+ $Y2=0
cc_473 N_A3_M1004_g N_A_1313_74#_c_1209_n 3.92313e-19 $X=8.775 $Y=0.74 $X2=0
+ $Y2=0
cc_474 N_A3_M1024_g N_A_1313_74#_c_1209_n 3.92313e-19 $X=9.205 $Y=0.74 $X2=0
+ $Y2=0
cc_475 N_A3_M1024_g N_A_1313_74#_c_1210_n 0.0130453f $X=9.205 $Y=0.74 $X2=0
+ $Y2=0
cc_476 N_A3_M1037_g N_A_1313_74#_c_1210_n 0.0128967f $X=9.635 $Y=0.74 $X2=0
+ $Y2=0
cc_477 N_A3_M1039_g N_A_1313_74#_c_1210_n 0.00174382f $X=10.065 $Y=0.74 $X2=0
+ $Y2=0
cc_478 A3 N_A_1313_74#_c_1210_n 0.0663371f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_479 N_A3_c_485_n N_A_1313_74#_c_1210_n 0.00508394f $X=10.05 $Y=1.515 $X2=0
+ $Y2=0
cc_480 N_A3_M1037_g N_A_1313_74#_c_1211_n 3.92313e-19 $X=9.635 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A3_M1039_g N_A_1313_74#_c_1211_n 3.92313e-19 $X=10.065 $Y=0.74 $X2=0
+ $Y2=0
cc_482 A3 N_A_1313_74#_c_1215_n 0.0146029f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_483 N_A3_c_485_n N_A_1313_74#_c_1215_n 0.00272398f $X=10.05 $Y=1.515 $X2=0
+ $Y2=0
cc_484 N_A_27_368#_c_564_n N_Y_M1000_d 0.00213667f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_485 N_A_27_368#_c_566_n N_Y_M1010_d 0.00165831f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_486 N_A_27_368#_c_567_n N_Y_M1009_s 0.00218982f $X=3.015 $Y=2.99 $X2=0 $Y2=0
cc_487 N_A_27_368#_c_568_n N_Y_M1012_s 0.00218982f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_488 N_A_27_368#_M1007_s N_Y_c_739_n 0.00314376f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_489 N_A_27_368#_c_660_p N_Y_c_739_n 0.0126919f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_490 N_A_27_368#_M1014_s N_Y_c_743_n 0.00438498f $X=1.995 $Y=1.84 $X2=0 $Y2=0
cc_491 N_A_27_368#_c_587_n N_Y_c_743_n 0.0189268f $X=2.18 $Y=2.455 $X2=0 $Y2=0
cc_492 N_A_27_368#_M1011_d N_Y_c_759_n 0.00410979f $X=2.995 $Y=1.84 $X2=0 $Y2=0
cc_493 N_A_27_368#_c_591_n N_Y_c_759_n 0.0189268f $X=3.18 $Y=2.455 $X2=0 $Y2=0
cc_494 N_A_27_368#_M1013_d N_Y_c_763_n 0.0138787f $X=3.995 $Y=1.84 $X2=0 $Y2=0
cc_495 N_A_27_368#_M1017_s N_Y_c_763_n 0.00314376f $X=5.135 $Y=1.84 $X2=0 $Y2=0
cc_496 N_A_27_368#_M1031_s N_Y_c_763_n 0.00426067f $X=6.135 $Y=1.84 $X2=0 $Y2=0
cc_497 N_A_27_368#_c_668_p N_Y_c_763_n 0.0238381f $X=4.18 $Y=2.46 $X2=0 $Y2=0
cc_498 N_A_27_368#_c_599_n N_Y_c_763_n 0.0411093f $X=5.105 $Y=2.375 $X2=0 $Y2=0
cc_499 N_A_27_368#_c_601_n N_Y_c_763_n 0.0388605f $X=6.105 $Y=2.375 $X2=0 $Y2=0
cc_500 N_A_27_368#_c_577_n N_Y_c_763_n 0.0171986f $X=5.27 $Y=2.455 $X2=0 $Y2=0
cc_501 N_A_27_368#_c_578_n N_Y_c_763_n 0.0164617f $X=6.27 $Y=2.455 $X2=0 $Y2=0
cc_502 N_A_27_368#_M1031_s N_Y_c_732_n 0.0014058f $X=6.135 $Y=1.84 $X2=0 $Y2=0
cc_503 N_A_27_368#_c_564_n N_Y_c_744_n 0.0173278f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_504 N_A_27_368#_c_566_n N_Y_c_748_n 0.0159318f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_505 N_A_27_368#_c_567_n N_Y_c_771_n 0.0177084f $X=3.015 $Y=2.99 $X2=0 $Y2=0
cc_506 N_A_27_368#_c_568_n N_Y_c_776_n 0.0177084f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_507 N_A_27_368#_c_599_n N_VPWR_M1016_d 0.00426066f $X=5.105 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_508 N_A_27_368#_c_601_n N_VPWR_M1025_d 0.00537357f $X=6.105 $Y=2.375 $X2=0
+ $Y2=0
cc_509 N_A_27_368#_c_609_n N_VPWR_M1002_d 0.00740097f $X=7.105 $Y=2.375 $X2=0
+ $Y2=0
cc_510 N_A_27_368#_c_625_n N_VPWR_M1026_d 0.00410979f $X=8.105 $Y=2.035 $X2=0
+ $Y2=0
cc_511 N_A_27_368#_c_629_n N_VPWR_M1003_s 0.00536271f $X=9.105 $Y=2.035 $X2=0
+ $Y2=0
cc_512 N_A_27_368#_c_643_n N_VPWR_M1021_s 0.00531191f $X=10.11 $Y=2.035 $X2=0
+ $Y2=0
cc_513 N_A_27_368#_c_568_n N_VPWR_c_853_n 0.0103379f $X=4.015 $Y=2.99 $X2=0
+ $Y2=0
cc_514 N_A_27_368#_c_598_n N_VPWR_c_853_n 0.015382f $X=4.18 $Y=2.905 $X2=0 $Y2=0
cc_515 N_A_27_368#_c_599_n N_VPWR_c_853_n 0.0189268f $X=5.105 $Y=2.375 $X2=0
+ $Y2=0
cc_516 N_A_27_368#_c_577_n N_VPWR_c_853_n 0.0139233f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_517 N_A_27_368#_c_601_n N_VPWR_c_854_n 0.0208278f $X=6.105 $Y=2.375 $X2=0
+ $Y2=0
cc_518 N_A_27_368#_c_577_n N_VPWR_c_854_n 0.0139233f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_519 N_A_27_368#_c_578_n N_VPWR_c_854_n 0.0139233f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_520 N_A_27_368#_c_609_n N_VPWR_c_855_n 0.0200142f $X=7.105 $Y=2.375 $X2=0
+ $Y2=0
cc_521 N_A_27_368#_c_569_n N_VPWR_c_855_n 0.0139233f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_522 N_A_27_368#_c_578_n N_VPWR_c_855_n 0.0139233f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_523 N_A_27_368#_c_569_n N_VPWR_c_856_n 0.0202646f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_524 N_A_27_368#_c_625_n N_VPWR_c_856_n 0.0189268f $X=8.105 $Y=2.035 $X2=0
+ $Y2=0
cc_525 N_A_27_368#_c_570_n N_VPWR_c_856_n 0.0266809f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_526 N_A_27_368#_c_570_n N_VPWR_c_857_n 0.0266809f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_527 N_A_27_368#_c_629_n N_VPWR_c_857_n 0.0189268f $X=9.105 $Y=2.035 $X2=0
+ $Y2=0
cc_528 N_A_27_368#_c_571_n N_VPWR_c_857_n 0.0266809f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_529 N_A_27_368#_c_571_n N_VPWR_c_858_n 0.0266809f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_530 N_A_27_368#_c_643_n N_VPWR_c_858_n 0.0212346f $X=10.11 $Y=2.035 $X2=0
+ $Y2=0
cc_531 N_A_27_368#_c_573_n N_VPWR_c_858_n 0.0260696f $X=10.275 $Y=2.815 $X2=0
+ $Y2=0
cc_532 N_A_27_368#_c_564_n N_VPWR_c_859_n 0.0440623f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_27_368#_c_565_n N_VPWR_c_859_n 0.0235688f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_534 N_A_27_368#_c_566_n N_VPWR_c_859_n 0.0439866f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_535 N_A_27_368#_c_567_n N_VPWR_c_859_n 0.0421443f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_536 N_A_27_368#_c_568_n N_VPWR_c_859_n 0.0658009f $X=4.015 $Y=2.99 $X2=0
+ $Y2=0
cc_537 N_A_27_368#_c_574_n N_VPWR_c_859_n 0.0121867f $X=1.23 $Y=2.99 $X2=0 $Y2=0
cc_538 N_A_27_368#_c_575_n N_VPWR_c_859_n 0.0235512f $X=2.18 $Y=2.99 $X2=0 $Y2=0
cc_539 N_A_27_368#_c_576_n N_VPWR_c_859_n 0.0235512f $X=3.18 $Y=2.99 $X2=0 $Y2=0
cc_540 N_A_27_368#_c_577_n N_VPWR_c_861_n 0.0144776f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_541 N_A_27_368#_c_578_n N_VPWR_c_863_n 0.0145075f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_542 N_A_27_368#_c_569_n N_VPWR_c_865_n 0.0144623f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_543 N_A_27_368#_c_570_n N_VPWR_c_867_n 0.014549f $X=8.27 $Y=2.815 $X2=0 $Y2=0
cc_544 N_A_27_368#_c_571_n N_VPWR_c_869_n 0.014549f $X=9.27 $Y=2.815 $X2=0 $Y2=0
cc_545 N_A_27_368#_c_573_n N_VPWR_c_870_n 0.014549f $X=10.275 $Y=2.815 $X2=0
+ $Y2=0
cc_546 N_A_27_368#_c_564_n N_VPWR_c_852_n 0.0247865f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_547 N_A_27_368#_c_565_n N_VPWR_c_852_n 0.0127152f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_548 N_A_27_368#_c_566_n N_VPWR_c_852_n 0.0246722f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_549 N_A_27_368#_c_567_n N_VPWR_c_852_n 0.0236813f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_550 N_A_27_368#_c_568_n N_VPWR_c_852_n 0.036511f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_551 N_A_27_368#_c_569_n N_VPWR_c_852_n 0.0118344f $X=7.27 $Y=2.815 $X2=0
+ $Y2=0
cc_552 N_A_27_368#_c_570_n N_VPWR_c_852_n 0.0119743f $X=8.27 $Y=2.815 $X2=0
+ $Y2=0
cc_553 N_A_27_368#_c_571_n N_VPWR_c_852_n 0.0119743f $X=9.27 $Y=2.815 $X2=0
+ $Y2=0
cc_554 N_A_27_368#_c_573_n N_VPWR_c_852_n 0.0119743f $X=10.275 $Y=2.815 $X2=0
+ $Y2=0
cc_555 N_A_27_368#_c_574_n N_VPWR_c_852_n 0.00660921f $X=1.23 $Y=2.99 $X2=0
+ $Y2=0
cc_556 N_A_27_368#_c_575_n N_VPWR_c_852_n 0.0126924f $X=2.18 $Y=2.99 $X2=0 $Y2=0
cc_557 N_A_27_368#_c_576_n N_VPWR_c_852_n 0.0126924f $X=3.18 $Y=2.99 $X2=0 $Y2=0
cc_558 N_A_27_368#_c_577_n N_VPWR_c_852_n 0.0118404f $X=5.27 $Y=2.455 $X2=0
+ $Y2=0
cc_559 N_A_27_368#_c_578_n N_VPWR_c_852_n 0.0118887f $X=6.27 $Y=2.455 $X2=0
+ $Y2=0
cc_560 N_Y_c_763_n N_VPWR_M1016_d 0.00411513f $X=6.18 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_561 N_Y_c_763_n N_VPWR_M1025_d 0.00631322f $X=6.18 $Y=2.035 $X2=0 $Y2=0
cc_562 N_Y_c_731_n N_A_27_74#_M1028_d 0.00255298f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_563 N_Y_c_736_n N_A_27_74#_M1038_d 0.00372475f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_564 N_Y_c_733_n N_A_27_74#_c_986_n 0.009209f $X=2.565 $Y=0.86 $X2=0 $Y2=0
cc_565 N_Y_M1018_s N_A_27_74#_c_987_n 0.00176461f $X=2.425 $Y=0.37 $X2=0 $Y2=0
cc_566 N_Y_c_731_n N_A_27_74#_c_987_n 0.0039879f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_567 N_Y_c_733_n N_A_27_74#_c_987_n 0.0158692f $X=2.565 $Y=0.86 $X2=0 $Y2=0
cc_568 N_Y_M1033_s N_A_27_74#_c_989_n 0.00285125f $X=3.355 $Y=0.37 $X2=0 $Y2=0
cc_569 N_Y_c_731_n N_A_27_74#_c_989_n 0.0108211f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_570 N_Y_c_736_n N_A_27_74#_c_989_n 0.0012223f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_571 N_Y_c_731_n N_A_27_74#_c_991_n 0.0211547f $X=3.51 $Y=1.03 $X2=0 $Y2=0
cc_572 N_Y_c_736_n N_A_27_74#_c_992_n 0.0139452f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_573 N_Y_c_736_n N_A_868_74#_M1005_d 0.00299905f $X=4.82 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_574 N_Y_c_735_n N_A_868_74#_M1029_d 0.00177442f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_575 N_Y_c_735_n N_A_868_74#_M1036_d 0.00535397f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_576 N_Y_c_736_n N_A_868_74#_c_1168_n 0.0214055f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_577 N_Y_M1005_s N_A_868_74#_c_1170_n 0.00254491f $X=4.775 $Y=0.37 $X2=0 $Y2=0
cc_578 N_Y_M1034_s N_A_868_74#_c_1170_n 0.00179007f $X=5.705 $Y=0.37 $X2=0 $Y2=0
cc_579 N_Y_c_735_n N_A_868_74#_c_1170_n 0.0127448f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_580 N_Y_c_736_n N_A_868_74#_c_1170_n 0.00412076f $X=4.82 $Y=0.975 $X2=0 $Y2=0
cc_581 N_Y_c_737_n N_A_868_74#_c_1170_n 0.0755709f $X=5.15 $Y=0.975 $X2=0 $Y2=0
cc_582 N_Y_c_732_n N_A_1313_74#_c_1212_n 0.00356311f $X=6.265 $Y=1.95 $X2=0
+ $Y2=0
cc_583 N_Y_c_735_n N_A_1313_74#_c_1212_n 0.0284876f $X=6.18 $Y=0.95 $X2=0 $Y2=0
cc_584 N_A_27_74#_c_983_n N_VGND_M1008_s 0.00250873f $X=1.125 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_585 N_A_27_74#_c_986_n N_VGND_M1032_s 0.00245557f $X=2.05 $Y=1.095 $X2=0
+ $Y2=0
cc_586 N_A_27_74#_c_982_n N_VGND_c_1056_n 0.0191765f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_587 N_A_27_74#_c_983_n N_VGND_c_1056_n 0.0210288f $X=1.125 $Y=1.095 $X2=0
+ $Y2=0
cc_588 N_A_27_74#_c_985_n N_VGND_c_1056_n 0.0182488f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_589 N_A_27_74#_c_985_n N_VGND_c_1057_n 0.0182488f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_590 N_A_27_74#_c_986_n N_VGND_c_1057_n 0.020622f $X=2.05 $Y=1.095 $X2=0 $Y2=0
cc_591 N_A_27_74#_c_988_n N_VGND_c_1057_n 0.00779323f $X=2.22 $Y=0.34 $X2=0
+ $Y2=0
cc_592 N_A_27_74#_c_982_n N_VGND_c_1062_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_593 N_A_27_74#_c_985_n N_VGND_c_1063_n 0.00749631f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_594 N_A_27_74#_c_987_n N_VGND_c_1064_n 0.042902f $X=2.9 $Y=0.34 $X2=0 $Y2=0
cc_595 N_A_27_74#_c_988_n N_VGND_c_1064_n 0.0121867f $X=2.22 $Y=0.34 $X2=0 $Y2=0
cc_596 N_A_27_74#_c_989_n N_VGND_c_1064_n 0.033414f $X=3.76 $Y=0.34 $X2=0 $Y2=0
cc_597 N_A_27_74#_c_991_n N_VGND_c_1064_n 0.0227371f $X=3.065 $Y=0.34 $X2=0
+ $Y2=0
cc_598 N_A_27_74#_c_992_n N_VGND_c_1064_n 0.0227371f $X=3.925 $Y=0.34 $X2=0
+ $Y2=0
cc_599 N_A_27_74#_c_982_n N_VGND_c_1071_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_600 N_A_27_74#_c_985_n N_VGND_c_1071_n 0.0062048f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_601 N_A_27_74#_c_987_n N_VGND_c_1071_n 0.0241973f $X=2.9 $Y=0.34 $X2=0 $Y2=0
cc_602 N_A_27_74#_c_988_n N_VGND_c_1071_n 0.00660921f $X=2.22 $Y=0.34 $X2=0
+ $Y2=0
cc_603 N_A_27_74#_c_989_n N_VGND_c_1071_n 0.0187892f $X=3.76 $Y=0.34 $X2=0 $Y2=0
cc_604 N_A_27_74#_c_991_n N_VGND_c_1071_n 0.0125119f $X=3.065 $Y=0.34 $X2=0
+ $Y2=0
cc_605 N_A_27_74#_c_992_n N_VGND_c_1071_n 0.0125119f $X=3.925 $Y=0.34 $X2=0
+ $Y2=0
cc_606 N_A_27_74#_c_992_n N_A_868_74#_c_1168_n 0.0242706f $X=3.925 $Y=0.34 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1064_n N_A_868_74#_c_1168_n 0.0142249f $X=8.395 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1071_n N_A_868_74#_c_1168_n 0.011867f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_c_1058_n N_A_868_74#_c_1169_n 0.0231578f $X=8.56 $Y=0.595 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1064_n N_A_868_74#_c_1170_n 0.142724f $X=8.395 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1071_n N_A_868_74#_c_1170_n 0.120136f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_M1004_d N_A_1313_74#_c_1208_n 0.00299905f $X=8.415 $Y=0.37 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1058_n N_A_1313_74#_c_1208_n 0.0219827f $X=8.56 $Y=0.595 $X2=0
+ $Y2=0
cc_614 N_VGND_c_1058_n N_A_1313_74#_c_1209_n 0.0182488f $X=8.56 $Y=0.595 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1059_n N_A_1313_74#_c_1209_n 0.0182488f $X=9.42 $Y=0.595 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1065_n N_A_1313_74#_c_1209_n 0.00749631f $X=9.255 $Y=0 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1071_n N_A_1313_74#_c_1209_n 0.0062048f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_618 N_VGND_M1024_d N_A_1313_74#_c_1210_n 0.00176461f $X=9.28 $Y=0.37 $X2=0
+ $Y2=0
cc_619 N_VGND_c_1059_n N_A_1313_74#_c_1210_n 0.0171619f $X=9.42 $Y=0.595 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1061_n N_A_1313_74#_c_1210_n 0.00517071f $X=10.28 $Y=0.515 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1059_n N_A_1313_74#_c_1211_n 0.0182488f $X=9.42 $Y=0.595 $X2=0
+ $Y2=0
cc_622 N_VGND_c_1061_n N_A_1313_74#_c_1211_n 0.0243418f $X=10.28 $Y=0.515 $X2=0
+ $Y2=0
cc_623 N_VGND_c_1066_n N_A_1313_74#_c_1211_n 0.00749631f $X=10.115 $Y=0 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1071_n N_A_1313_74#_c_1211_n 0.0062048f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_625 N_A_868_74#_c_1170_n N_A_1313_74#_M1001_s 0.00179007f $X=7.835 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_626 N_A_868_74#_c_1170_n N_A_1313_74#_M1022_s 0.00212678f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
cc_627 N_A_868_74#_M1023_d N_A_1313_74#_c_1208_n 0.00388574f $X=7.86 $Y=0.37
+ $X2=0 $Y2=0
cc_628 N_A_868_74#_c_1169_n N_A_1313_74#_c_1208_n 0.0127309f $X=8 $Y=0.515 $X2=0
+ $Y2=0
cc_629 N_A_868_74#_c_1170_n N_A_1313_74#_c_1208_n 0.00339963f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
cc_630 N_A_868_74#_c_1170_n N_A_1313_74#_c_1212_n 0.0163588f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0
cc_631 N_A_868_74#_M1006_d N_A_1313_74#_c_1213_n 0.00217299f $X=6.995 $Y=0.37
+ $X2=0 $Y2=0
cc_632 N_A_868_74#_c_1170_n N_A_1313_74#_c_1213_n 0.0336602f $X=7.835 $Y=0.515
+ $X2=0 $Y2=0

* File: sky130_fd_sc_ms__xnor3_4.pex.spice
* Created: Wed Sep  2 12:33:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_75_227# 1 2 3 4 15 19 21 22 24 25 26 29 33
+ 34 35 37 38 42 47 48 51 56
c131 33 0 1.89638e-19 $X=1.26 $Y=0.53
r132 51 53 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.515 $Y=2.795
+ $X2=3.515 $Y2=2.99
r133 47 48 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.35
+ $X2=3.2 $Y2=0.35
r134 42 57 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.3
+ $X2=0.54 $Y2=1.465
r135 42 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.3
+ $X2=0.54 $Y2=1.135
r136 41 43 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=1.3
+ $X2=0.58 $Y2=1.465
r137 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.3 $X2=0.54 $Y2=1.3
r138 38 41 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=0.58 $Y=1.12
+ $X2=0.58 $Y2=1.3
r139 37 48 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=1.425 $Y=0.34
+ $X2=3.2 $Y2=0.34
r140 34 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.35 $Y=2.99
+ $X2=3.515 $Y2=2.99
r141 34 35 127.545 $w=1.68e-07 $l=1.955e-06 $layer=LI1_cond $X=3.35 $Y=2.99
+ $X2=1.395 $Y2=2.99
r142 31 33 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=1.3 $Y=1.035
+ $X2=1.3 $Y2=0.53
r143 30 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.3 $Y=0.425
+ $X2=1.425 $Y2=0.34
r144 30 33 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=1.3 $Y=0.425
+ $X2=1.3 $Y2=0.53
r145 27 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.395 $Y2=2.99
r146 27 29 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.72
r147 26 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.12 $X2=1.23
+ $Y2=2.035
r148 26 29 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=1.23 $Y=2.12 $X2=1.23
+ $Y2=2.72
r149 24 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=1.23 $Y2=2.035
r150 24 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=0.705 $Y2=2.035
r151 23 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.705 $Y=1.12
+ $X2=0.58 $Y2=1.12
r152 22 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.175 $Y=1.12
+ $X2=1.3 $Y2=1.035
r153 22 23 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.175 $Y=1.12
+ $X2=0.705 $Y2=1.12
r154 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.705 $Y2=2.035
r155 21 43 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.62 $Y2=1.465
r156 19 56 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.545 $Y=0.705
+ $X2=0.545 $Y2=1.135
r157 15 57 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=0.505 $Y=2.365
+ $X2=0.505 $Y2=1.465
r158 4 51 600 $w=1.7e-07 $l=1.03417e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.865 $X2=3.515 $Y2=2.795
r159 3 45 300 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.865 $X2=1.23 $Y2=2.035
r160 3 29 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.865 $X2=1.23 $Y2=2.72
r161 2 47 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.605 $X2=3.365 $Y2=0.36
r162 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.12
+ $Y=0.385 $X2=1.26 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A 3 7 9 12 13
c44 12 0 9.56919e-20 $X=1.08 $Y=1.54
c45 7 0 1.6832e-19 $X=1.045 $Y=0.705
r46 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.54
+ $X2=1.08 $Y2=1.705
r47 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.54
+ $X2=1.08 $Y2=1.375
r48 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.54 $X2=1.08 $Y2=1.54
r49 9 13 3.60138 $w=3.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.115 $Y=1.665
+ $X2=1.115 $Y2=1.54
r50 7 14 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.045 $Y=0.705
+ $X2=1.045 $Y2=1.375
r51 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.005 $Y=2.365
+ $X2=1.005 $Y2=1.705
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_386_23# 1 2 10 11 12 13 15 20 23 29 32 35
+ 37 38 40 42 44 46
c125 46 0 1.70037e-20 $X=3.685 $Y=1.54
c126 32 0 1.9098e-19 $X=3.16 $Y=1.54
c127 15 0 8.8275e-20 $X=2.245 $Y=2.185
c128 11 0 1.46697e-19 $X=2.995 $Y=0.19
c129 10 0 7.08805e-20 $X=2.005 $Y=0.815
r130 42 44 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.77 $Y=2.075
+ $X2=4.105 $Y2=2.075
r131 38 40 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.77 $Y=1.04
+ $X2=3.925 $Y2=1.04
r132 37 42 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685 $Y=1.95
+ $X2=3.77 $Y2=2.075
r133 36 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=1.705
+ $X2=3.685 $Y2=1.54
r134 36 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.685 $Y=1.705
+ $X2=3.685 $Y2=1.95
r135 35 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=1.375
+ $X2=3.685 $Y2=1.54
r136 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.685 $Y=1.125
+ $X2=3.77 $Y2=1.04
r137 34 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.685 $Y=1.125
+ $X2=3.685 $Y2=1.375
r138 32 49 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.54
+ $X2=3.16 $Y2=1.705
r139 32 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.54
+ $X2=3.16 $Y2=1.375
r140 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.16
+ $Y=1.54 $X2=3.16 $Y2=1.54
r141 29 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.54
+ $X2=3.685 $Y2=1.54
r142 29 31 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.6 $Y=1.54
+ $X2=3.16 $Y2=1.54
r143 23 49 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.205 $Y=2.285
+ $X2=3.205 $Y2=1.705
r144 20 48 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.07 $Y=0.925
+ $X2=3.07 $Y2=1.375
r145 17 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.07 $Y=0.265
+ $X2=3.07 $Y2=0.925
r146 13 25 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.245 $Y=1.395
+ $X2=2.005 $Y2=1.395
r147 13 15 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=2.245 $Y=1.47
+ $X2=2.245 $Y2=2.185
r148 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.995 $Y=0.19
+ $X2=3.07 $Y2=0.265
r149 11 12 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.995 $Y=0.19
+ $X2=2.08 $Y2=0.19
r150 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.005 $Y=1.32
+ $X2=2.005 $Y2=1.395
r151 8 10 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.005 $Y=1.32
+ $X2=2.005 $Y2=0.815
r152 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.005 $Y=0.265
+ $X2=2.08 $Y2=0.19
r153 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.005 $Y=0.265
+ $X2=2.005 $Y2=0.815
r154 2 44 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.84 $X2=4.105 $Y2=2.115
r155 1 40 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.445 $X2=3.925 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%B 3 5 8 9 10 13 18 19 22 25 29 33 34 35 40
+ 41
c133 40 0 1.9098e-19 $X=4.105 $Y=1.515
c134 29 0 1.70037e-20 $X=4.33 $Y=2.4
c135 22 0 2.17801e-20 $X=3.81 $Y=3.075
c136 5 0 1.19763e-19 $X=1.545 $Y=1.73
c137 3 0 1.70469e-19 $X=1.53 $Y=0.705
r138 41 42 33.1812 $w=2.76e-07 $l=1.9e-07 $layer=POLY_cond $X=4.14 $Y=1.515
+ $X2=4.33 $Y2=1.515
r139 39 41 6.11232 $w=2.76e-07 $l=3.5e-08 $layer=POLY_cond $X=4.105 $Y=1.515
+ $X2=4.14 $Y2=1.515
r140 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.515 $X2=4.105 $Y2=1.515
r141 35 40 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.105 $Y=1.665
+ $X2=4.105 $Y2=1.515
r142 32 33 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.665 $Y=1.64
+ $X2=2.665 $Y2=1.79
r143 27 42 12.7955 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.33 $Y=1.68
+ $X2=4.33 $Y2=1.515
r144 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.33 $Y=1.68
+ $X2=4.33 $Y2=2.4
r145 23 41 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=1.515
r146 23 25 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=0.815
r147 21 39 51.5181 $w=2.76e-07 $l=3.68375e-07 $layer=POLY_cond $X=3.81 $Y=1.68
+ $X2=4.105 $Y2=1.515
r148 21 22 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=3.81 $Y=1.68
+ $X2=3.81 $Y2=3.075
r149 20 34 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.785 $Y=3.15
+ $X2=2.695 $Y2=3.15
r150 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.735 $Y=3.15
+ $X2=3.81 $Y2=3.075
r151 19 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.735 $Y=3.15
+ $X2=2.785 $Y2=3.15
r152 18 33 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.695 $Y=2.185
+ $X2=2.695 $Y2=1.79
r153 16 34 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=3.075
+ $X2=2.695 $Y2=3.15
r154 16 18 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.695 $Y=3.075
+ $X2=2.695 $Y2=2.185
r155 13 32 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.62 $Y=0.925
+ $X2=2.62 $Y2=1.64
r156 9 34 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.605 $Y=3.15
+ $X2=2.695 $Y2=3.15
r157 9 10 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.605 $Y=3.15
+ $X2=1.635 $Y2=3.15
r158 6 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.545 $Y=3.075
+ $X2=1.635 $Y2=3.15
r159 6 8 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.545 $Y=3.075
+ $X2=1.545 $Y2=2.285
r160 5 31 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.545 $Y=1.73
+ $X2=1.545 $Y2=1.64
r161 5 8 215.734 $w=1.8e-07 $l=5.55e-07 $layer=POLY_cond $X=1.545 $Y=1.73
+ $X2=1.545 $Y2=2.285
r162 3 31 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.53 $Y=0.705
+ $X2=1.53 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_1024_300# 1 2 9 13 15 18 20 23 25 27 30 34
r86 31 34 6.33218 $w=5.08e-07 $l=2.7e-07 $layer=LI1_cond $X=6.525 $Y=2.245
+ $X2=6.795 $Y2=2.245
r87 27 29 4.25191 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.085
+ $X2=6.555 $Y2=1.17
r88 23 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.665
+ $X2=5.285 $Y2=1.83
r89 23 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.665
+ $X2=5.285 $Y2=1.5
r90 22 25 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=1.665
+ $X2=5.45 $Y2=1.665
r91 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.285
+ $Y=1.665 $X2=5.285 $Y2=1.665
r92 20 31 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=6.525 $Y=1.99
+ $X2=6.525 $Y2=2.245
r93 19 30 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.525 $Y=1.72
+ $X2=6.5 $Y2=1.635
r94 19 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.525 $Y=1.72
+ $X2=6.525 $Y2=1.99
r95 18 30 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=1.55 $X2=6.5
+ $Y2=1.635
r96 18 29 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=6.5 $Y=1.55 $X2=6.5
+ $Y2=1.17
r97 15 30 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.39 $Y=1.635 $X2=6.5
+ $Y2=1.635
r98 15 25 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.39 $Y=1.635
+ $X2=5.45 $Y2=1.635
r99 13 38 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=5.34 $Y=2.41
+ $X2=5.34 $Y2=1.83
r100 9 37 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.21 $Y=0.69 $X2=5.21
+ $Y2=1.5
r101 2 34 600 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=1 $X=6.65
+ $Y=1.84 $X2=6.795 $Y2=2.235
r102 1 27 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.41
+ $Y=0.81 $X2=6.555 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%C 3 7 10 11 13 16 21 24 27 28
c76 11 0 2.47917e-19 $X=6.77 $Y=1.35
r77 26 28 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.945 $Y=1.515
+ $X2=7.02 $Y2=1.515
r78 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.945
+ $Y=1.515 $X2=6.945 $Y2=1.515
r79 23 26 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.77 $Y=1.515
+ $X2=6.945 $Y2=1.515
r80 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.77 $Y=1.515
+ $X2=6.695 $Y2=1.515
r81 21 27 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.945 $Y=1.665
+ $X2=6.945 $Y2=1.515
r82 14 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.02 $Y=1.68
+ $X2=7.02 $Y2=1.515
r83 14 16 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=7.02 $Y=1.68
+ $X2=7.02 $Y2=2.16
r84 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.35
+ $X2=6.77 $Y2=1.515
r85 11 13 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.77 $Y=1.35 $X2=6.77
+ $Y2=1.02
r86 10 24 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.05 $Y=1.425
+ $X2=6.695 $Y2=1.425
r87 5 10 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.96 $Y=1.425 $X2=6.05
+ $Y2=1.425
r88 5 18 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.96 $Y=1.425
+ $X2=5.765 $Y2=1.425
r89 5 7 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=5.96 $Y=1.5 $X2=5.96
+ $Y2=2.41
r90 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=1.425
r91 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_1057_74# 1 2 9 11 13 16 18 20 23 25 27 28
+ 30 32 34 37 39 40 41 44 45 46 48 49 50 52 54 56 59 63 69 72 74
c159 74 0 1.96868e-19 $X=8.13 $Y=1.505
c160 72 0 1.17951e-19 $X=7.485 $Y=1.505
r161 82 83 5.14329 $w=3.28e-07 $l=3.5e-08 $layer=POLY_cond $X=9.12 $Y=1.505
+ $X2=9.155 $Y2=1.505
r162 81 82 58.0457 $w=3.28e-07 $l=3.95e-07 $layer=POLY_cond $X=8.725 $Y=1.505
+ $X2=9.12 $Y2=1.505
r163 80 81 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=8.67 $Y=1.505
+ $X2=8.725 $Y2=1.505
r164 79 80 55.1067 $w=3.28e-07 $l=3.75e-07 $layer=POLY_cond $X=8.295 $Y=1.505
+ $X2=8.67 $Y2=1.505
r165 78 79 11.0213 $w=3.28e-07 $l=7.5e-08 $layer=POLY_cond $X=8.22 $Y=1.505
+ $X2=8.295 $Y2=1.505
r166 73 74 112.786 $w=3.3e-07 $l=6.45e-07 $layer=POLY_cond $X=7.485 $Y=1.505
+ $X2=8.13 $Y2=1.505
r167 72 73 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.485
+ $Y=1.505 $X2=7.485 $Y2=1.505
r168 67 69 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=7.222 $Y=2.035
+ $X2=7.405 $Y2=2.035
r169 63 65 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.65 $Y=2.895
+ $X2=5.65 $Y2=2.99
r170 60 78 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=8.165 $Y=1.505
+ $X2=8.22 $Y2=1.505
r171 60 74 5.11212 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.165 $Y=1.505
+ $X2=8.13 $Y2=1.505
r172 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.165
+ $Y=1.505 $X2=8.165 $Y2=1.505
r173 57 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.49 $Y=1.505
+ $X2=7.405 $Y2=1.505
r174 57 59 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.49 $Y=1.505
+ $X2=8.165 $Y2=1.505
r175 56 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=1.95
+ $X2=7.405 $Y2=2.035
r176 55 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=1.67
+ $X2=7.405 $Y2=1.505
r177 55 56 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.405 $Y=1.67
+ $X2=7.405 $Y2=1.95
r178 54 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=1.34
+ $X2=7.405 $Y2=1.505
r179 53 54 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.405 $Y=1.18
+ $X2=7.405 $Y2=1.34
r180 51 67 0.22998 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=7.222 $Y=2.12
+ $X2=7.222 $Y2=2.035
r181 51 52 47.0614 $w=1.83e-07 $l=7.85e-07 $layer=LI1_cond $X=7.222 $Y=2.12
+ $X2=7.222 $Y2=2.905
r182 49 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.32 $Y=1.095
+ $X2=7.405 $Y2=1.18
r183 49 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.32 $Y=1.095
+ $X2=7.06 $Y2=1.095
r184 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.975 $Y=1.01
+ $X2=7.06 $Y2=1.095
r185 47 48 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.975 $Y=0.83
+ $X2=6.975 $Y2=1.01
r186 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.975 $Y2=0.83
r187 45 46 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.5 $Y2=0.745
r188 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=0.66
+ $X2=6.5 $Y2=0.745
r189 43 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.415 $Y=0.425
+ $X2=6.415 $Y2=0.66
r190 42 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=2.99
+ $X2=5.65 $Y2=2.99
r191 41 52 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.13 $Y=2.99
+ $X2=7.222 $Y2=2.905
r192 41 42 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=7.13 $Y=2.99
+ $X2=5.815 $Y2=2.99
r193 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=6.415 $Y2=0.425
r194 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=5.66 $Y2=0.34
r195 35 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.66 $Y2=0.34
r196 35 37 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.495 $Y2=0.515
r197 32 85 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.585 $Y=1.34
+ $X2=9.585 $Y2=1.505
r198 32 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.585 $Y=1.34
+ $X2=9.585 $Y2=0.86
r199 28 85 2.20427 $w=3.28e-07 $l=1.5e-08 $layer=POLY_cond $X=9.57 $Y=1.505
+ $X2=9.585 $Y2=1.505
r200 28 83 60.9848 $w=3.28e-07 $l=4.15e-07 $layer=POLY_cond $X=9.57 $Y=1.505
+ $X2=9.155 $Y2=1.505
r201 28 30 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=9.57 $Y=1.665
+ $X2=9.57 $Y2=2.4
r202 25 83 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.155 $Y=1.34
+ $X2=9.155 $Y2=1.505
r203 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.155 $Y=1.34
+ $X2=9.155 $Y2=0.86
r204 21 82 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.12 $Y=1.67
+ $X2=9.12 $Y2=1.505
r205 21 23 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=9.12 $Y=1.67
+ $X2=9.12 $Y2=2.4
r206 18 81 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.725 $Y=1.34
+ $X2=8.725 $Y2=1.505
r207 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.725 $Y=1.34
+ $X2=8.725 $Y2=0.86
r208 14 80 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.67
+ $X2=8.67 $Y2=1.505
r209 14 16 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=8.67 $Y=1.67
+ $X2=8.67 $Y2=2.4
r210 11 79 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.295 $Y=1.34
+ $X2=8.295 $Y2=1.505
r211 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.295 $Y=1.34
+ $X2=8.295 $Y2=0.86
r212 7 78 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.22 $Y=1.67
+ $X2=8.22 $Y2=1.505
r213 7 9 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=8.22 $Y=1.67 $X2=8.22
+ $Y2=2.4
r214 2 63 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.99 $X2=5.65 $Y2=2.895
r215 1 37 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.495 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_27_373# 1 2 3 4 15 17 18 20 23 24 25 29 34
+ 38 39 45 46 49
c107 29 0 6.75216e-20 $X=2.3 $Y=1.1
c108 25 0 1.83967e-19 $X=1.665 $Y=1.475
c109 20 0 1.6832e-19 $X=0.33 $Y=0.615
r110 49 51 29.2227 $w=2.78e-07 $l=7.1e-07 $layer=LI1_cond $X=0.225 $Y=2.01
+ $X2=0.225 $Y2=2.72
r111 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.035
r112 41 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.035
r113 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=2.035
+ $X2=0.24 $Y2=2.035
r114 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.535 $Y=2.035
+ $X2=1.68 $Y2=2.035
r115 38 39 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=1.535 $Y=2.035
+ $X2=0.385 $Y2=2.035
r116 34 36 7.40856 $w=4.18e-07 $l=2.7e-07 $layer=LI1_cond $X=2.515 $Y=2.38
+ $X2=2.515 $Y2=2.65
r117 29 31 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.26 $Y=1.1
+ $X2=2.26 $Y2=1.25
r118 27 46 29.3909 $w=1.98e-07 $l=5.3e-07 $layer=LI1_cond $X=1.665 $Y=2.565
+ $X2=1.665 $Y2=2.035
r119 25 46 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=1.665 $Y=1.475
+ $X2=1.665 $Y2=2.035
r120 25 26 13.8873 $w=2e-07 $l=2.25e-07 $layer=LI1_cond $X=1.665 $Y=1.475
+ $X2=1.665 $Y2=1.25
r121 23 49 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.225 $Y=1.985
+ $X2=0.225 $Y2=2.01
r122 23 24 6.72007 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=1.985
+ $X2=0.225 $Y2=1.845
r123 22 24 54.3455 $w=1.98e-07 $l=9.8e-07 $layer=LI1_cond $X=0.185 $Y=0.865
+ $X2=0.185 $Y2=1.845
r124 20 22 10.0564 $w=4.08e-07 $l=2.5e-07 $layer=LI1_cond $X=0.29 $Y=0.615
+ $X2=0.29 $Y2=0.865
r125 18 27 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.765 $Y=2.65
+ $X2=1.665 $Y2=2.565
r126 17 36 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.305 $Y=2.65
+ $X2=2.515 $Y2=2.65
r127 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.305 $Y=2.65
+ $X2=1.765 $Y2=2.65
r128 16 26 1.02909 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.765 $Y=1.25
+ $X2=1.665 $Y2=1.25
r129 15 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.135 $Y=1.25
+ $X2=2.26 $Y2=1.25
r130 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.135 $Y=1.25
+ $X2=1.765 $Y2=1.25
r131 4 34 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.865 $X2=2.47 $Y2=2.38
r132 3 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.865 $X2=0.28 $Y2=2.72
r133 3 49 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.865 $X2=0.28 $Y2=2.01
r134 2 29 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.605 $X2=2.3 $Y2=1.1
r135 1 20 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.385 $X2=0.33 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%VPWR 1 2 3 4 5 18 22 25 28 30 34 38 40 45 47
+ 49 54 62 70 76 79 82 85 89
r107 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r108 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r109 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r110 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 74 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r114 74 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 71 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=8.895 $Y2=3.33
r117 71 73 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.98 $Y=3.33
+ $X2=9.36 $Y2=3.33
r118 70 88 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.895 $Y2=3.33
r119 70 73 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.36 $Y2=3.33
r120 69 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 65 68 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 63 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=4.555 $Y2=3.33
r124 63 65 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 62 82 12.8484 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.797 $Y2=3.33
r126 62 68 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.44 $Y2=3.33
r127 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 60 61 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 58 61 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 57 60 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 57 58 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 55 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r134 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 54 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=3.33
+ $X2=4.555 $Y2=3.33
r136 54 60 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.39 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 52 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 49 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r140 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 47 69 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r142 47 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 47 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 45 46 3.52857 $w=6.23e-07 $l=1.2e-07 $layer=LI1_cond $X=7.797 $Y=2.41
+ $X2=7.797 $Y2=2.29
r145 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.835 $Y=1.985
+ $X2=9.835 $Y2=2.815
r146 38 88 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.835 $Y=3.245
+ $X2=9.895 $Y2=3.33
r147 38 43 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.835 $Y=3.245
+ $X2=9.835 $Y2=2.815
r148 34 37 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.895 $Y=1.985
+ $X2=8.895 $Y2=2.815
r149 32 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=3.245
+ $X2=8.895 $Y2=3.33
r150 32 37 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.895 $Y=3.245
+ $X2=8.895 $Y2=2.815
r151 31 82 12.8484 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=8.11 $Y=3.33
+ $X2=7.797 $Y2=3.33
r152 30 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.895 $Y2=3.33
r153 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.81 $Y=3.33 $X2=8.11
+ $Y2=3.33
r154 28 46 7.72815 $w=4.23e-07 $l=2.85e-07 $layer=LI1_cond $X=7.897 $Y=2.005
+ $X2=7.897 $Y2=2.29
r155 25 82 2.61429 $w=6.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.797 $Y=3.245
+ $X2=7.797 $Y2=3.33
r156 24 45 3.67435 $w=6.23e-07 $l=1.92e-07 $layer=LI1_cond $X=7.797 $Y=2.602
+ $X2=7.797 $Y2=2.41
r157 24 25 12.3053 $w=6.23e-07 $l=6.43e-07 $layer=LI1_cond $X=7.797 $Y=2.602
+ $X2=7.797 $Y2=3.245
r158 20 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=3.33
r159 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=2.815
r160 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r161 16 18 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.375
r162 5 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.795 $Y2=2.815
r163 5 40 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.795 $Y2=1.985
r164 4 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.895 $Y2=2.815
r165 4 34 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.895 $Y2=1.985
r166 3 45 150 $w=1.7e-07 $l=1.13476e-06 $layer=licon1_PDIFF $count=4 $X=7.11
+ $Y=1.84 $X2=7.995 $Y2=2.41
r167 3 28 600 $w=1.7e-07 $l=7.37902e-07 $layer=licon1_PDIFF $count=1 $X=7.11
+ $Y=1.84 $X2=7.77 $Y2=2.005
r168 2 22 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.84 $X2=4.555 $Y2=2.815
r169 1 18 300 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.865 $X2=0.73 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_327_373# 1 2 3 4 14 15 16 18 20 22 23 25
+ 30 33 35 36 42 43 46
c128 16 0 2.40512e-19 $X=2.245 $Y=1.59
r129 43 47 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.04 $Y=2.085
+ $X2=4.865 $Y2=2.085
r130 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r131 38 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r132 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r133 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r134 35 36 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=2.305 $Y2=2.035
r135 27 30 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=2.655 $Y=1.08
+ $X2=2.845 $Y2=1.08
r136 23 33 32.9995 $w=1.98e-07 $l=5.9e-07 $layer=LI1_cond $X=5.995 $Y=1.28
+ $X2=5.405 $Y2=1.28
r137 23 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.995 $Y=1.18
+ $X2=5.995 $Y2=0.81
r138 22 33 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.95 $Y=1.295
+ $X2=5.405 $Y2=1.295
r139 20 47 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.865 $Y=1.95
+ $X2=4.865 $Y2=2.085
r140 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.865 $Y=1.38
+ $X2=4.95 $Y2=1.295
r141 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.865 $Y=1.38
+ $X2=4.865 $Y2=1.95
r142 17 27 2.04652 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=1.205
+ $X2=2.655 $Y2=1.08
r143 17 18 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=2.655 $Y=1.205
+ $X2=2.655 $Y2=1.505
r144 15 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.555 $Y=1.59
+ $X2=2.655 $Y2=1.505
r145 15 16 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.555 $Y=1.59
+ $X2=2.245 $Y2=1.59
r146 14 46 1.05747 $w=3.1e-07 $l=2.5e-08 $layer=LI1_cond $X=2.09 $Y=1.965
+ $X2=2.09 $Y2=1.99
r147 13 16 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.245 $Y2=1.59
r148 13 14 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.09 $Y2=1.965
r149 4 43 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=1.99 $X2=5.115 $Y2=2.135
r150 3 46 600 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=1.635
+ $Y=1.865 $X2=2.02 $Y2=1.99
r151 2 25 182 $w=1.7e-07 $l=5.11664e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.37 $X2=5.995 $Y2=0.81
r152 1 30 182 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.605 $X2=2.845 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%A_321_77# 1 2 3 4 15 19 21 22 24 25 29 31 36
+ 37 38 41
c130 37 0 2.17577e-19 $X=2.725 $Y=0.69
c131 22 0 2.17801e-20 $X=3.145 $Y=2.455
r132 38 40 10.6978 $w=5.36e-07 $l=4.7e-07 $layer=LI1_cond $X=4.525 $Y=0.69
+ $X2=4.995 $Y2=0.69
r133 36 37 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=0.69
+ $X2=2.725 $Y2=0.69
r134 31 34 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.79 $Y=0.68
+ $X2=1.79 $Y2=0.795
r135 27 29 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.145 $Y=2.39
+ $X2=6.145 $Y2=2.135
r136 26 41 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.61 $Y=2.475
+ $X2=4.525 $Y2=2.465
r137 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.02 $Y=2.475
+ $X2=6.145 $Y2=2.39
r138 25 26 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=6.02 $Y=2.475
+ $X2=4.61 $Y2=2.475
r139 24 41 1.34256 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.525 $Y=2.37
+ $X2=4.525 $Y2=2.465
r140 23 38 7.59541 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=4.525 $Y=1.03
+ $X2=4.525 $Y2=0.69
r141 23 24 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=4.525 $Y=1.03
+ $X2=4.525 $Y2=2.37
r142 21 41 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.44 $Y=2.455
+ $X2=4.525 $Y2=2.465
r143 21 22 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=4.44 $Y=2.455
+ $X2=3.145 $Y2=2.455
r144 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.02 $Y=2.37
+ $X2=3.145 $Y2=2.455
r145 17 19 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=3.02 $Y=2.37
+ $X2=3.02 $Y2=2.04
r146 15 38 8.11642 $w=5.36e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.44 $Y=0.7
+ $X2=4.525 $Y2=0.69
r147 15 37 111.888 $w=1.68e-07 $l=1.715e-06 $layer=LI1_cond $X=4.44 $Y=0.7
+ $X2=2.725 $Y2=0.7
r148 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=1.79 $Y2=0.68
r149 14 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=2.555 $Y2=0.68
r150 4 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.05
+ $Y=1.99 $X2=6.185 $Y2=2.135
r151 3 19 300 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=2 $X=2.785
+ $Y=1.865 $X2=2.98 $Y2=2.04
r152 2 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.37 $X2=4.995 $Y2=0.515
r153 1 34 182 $w=1.7e-07 $l=4.93913e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.385 $X2=1.79 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%X 1 2 3 4 15 19 22 25 28 29 30 31 32 33 34
+ 35 36 37 38 58
r58 56 58 1.29853 $w=3.53e-07 $l=4e-08 $layer=LI1_cond $X=9.357 $Y=1.625
+ $X2=9.357 $Y2=1.665
r59 37 38 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=9.357 $Y=2.405
+ $X2=9.357 $Y2=2.775
r60 36 37 13.6345 $w=3.53e-07 $l=4.2e-07 $layer=LI1_cond $X=9.357 $Y=1.985
+ $X2=9.357 $Y2=2.405
r61 35 47 3.3083 $w=3.42e-07 $l=1.08305e-07 $layer=LI1_cond $X=9.357 $Y=1.522
+ $X2=9.37 $Y2=1.42
r62 35 56 3.3083 $w=3.42e-07 $l=1.03e-07 $layer=LI1_cond $X=9.357 $Y=1.522
+ $X2=9.357 $Y2=1.625
r63 35 36 9.67403 $w=3.53e-07 $l=2.98e-07 $layer=LI1_cond $X=9.357 $Y=1.687
+ $X2=9.357 $Y2=1.985
r64 35 58 0.71419 $w=3.53e-07 $l=2.2e-08 $layer=LI1_cond $X=9.357 $Y=1.687
+ $X2=9.357 $Y2=1.665
r65 34 47 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.37 $Y=1.295
+ $X2=9.37 $Y2=1.42
r66 33 34 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=0.925
+ $X2=9.37 $Y2=1.295
r67 32 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=0.555
+ $X2=9.37 $Y2=0.925
r68 28 29 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.46 $Y=2.005
+ $X2=8.46 $Y2=1.84
r69 26 31 1.0233 $w=2.05e-07 $l=1.03e-07 $layer=LI1_cond $X=8.675 $Y=1.522
+ $X2=8.572 $Y2=1.522
r70 25 35 3.24129 $w=2.05e-07 $l=1.77e-07 $layer=LI1_cond $X=9.18 $Y=1.522
+ $X2=9.357 $Y2=1.522
r71 25 26 27.3215 $w=2.03e-07 $l=5.05e-07 $layer=LI1_cond $X=9.18 $Y=1.522
+ $X2=8.675 $Y2=1.522
r72 23 31 5.56063 $w=1.87e-07 $l=1.11176e-07 $layer=LI1_cond $X=8.555 $Y=1.625
+ $X2=8.572 $Y2=1.522
r73 23 29 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.555 $Y=1.625
+ $X2=8.555 $Y2=1.84
r74 22 31 5.56063 $w=1.87e-07 $l=1.02e-07 $layer=LI1_cond $X=8.572 $Y=1.42
+ $X2=8.572 $Y2=1.522
r75 22 30 13.5255 $w=2.03e-07 $l=2.5e-07 $layer=LI1_cond $X=8.572 $Y=1.42
+ $X2=8.572 $Y2=1.17
r76 17 30 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.51 $Y=1.005
+ $X2=8.51 $Y2=1.17
r77 17 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.51 $Y=1.005
+ $X2=8.51 $Y2=0.635
r78 13 28 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=8.46 $Y=2.02
+ $X2=8.46 $Y2=2.005
r79 13 15 25.4498 $w=3.58e-07 $l=7.95e-07 $layer=LI1_cond $X=8.46 $Y=2.02
+ $X2=8.46 $Y2=2.815
r80 4 38 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.21
+ $Y=1.84 $X2=9.345 $Y2=2.815
r81 4 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.21
+ $Y=1.84 $X2=9.345 $Y2=1.985
r82 3 28 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=8.31
+ $Y=1.84 $X2=8.445 $Y2=2.005
r83 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.31
+ $Y=1.84 $X2=8.445 $Y2=2.815
r84 2 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.23
+ $Y=0.49 $X2=9.37 $Y2=0.635
r85 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.37
+ $Y=0.49 $X2=8.51 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_4%VGND 1 2 3 4 5 20 24 26 30 32 33 36 38 40 42
+ 44 52 58 61 77 81
c100 20 0 1.02947e-19 $X=0.83 $Y=0.615
r101 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r102 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r103 74 75 0.585834 $w=8.33e-07 $l=4e-08 $layer=LI1_cond $X=8 $Y=0.377 $X2=8.04
+ $Y2=0.377
r104 72 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r105 71 74 1.17167 $w=8.33e-07 $l=8e-08 $layer=LI1_cond $X=7.92 $Y=0.377 $X2=8
+ $Y2=0.377
r106 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r107 69 71 5.71188 $w=8.33e-07 $l=3.9e-07 $layer=LI1_cond $X=7.53 $Y=0.377
+ $X2=7.92 $Y2=0.377
r108 67 69 6.81032 $w=8.33e-07 $l=4.65e-07 $layer=LI1_cond $X=7.065 $Y=0.377
+ $X2=7.53 $Y2=0.377
r109 65 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r110 64 67 1.53782 $w=8.33e-07 $l=1.05e-07 $layer=LI1_cond $X=6.96 $Y=0.377
+ $X2=7.065 $Y2=0.377
r111 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r112 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r113 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r114 56 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r115 56 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r116 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r117 53 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.025 $Y=0 $X2=8.94
+ $Y2=0
r118 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=9.36 $Y2=0
r119 52 80 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.715 $Y=0
+ $X2=9.897 $Y2=0
r120 52 55 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.715 $Y=0
+ $X2=9.36 $Y2=0
r121 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r122 50 51 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r123 48 51 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r124 48 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r125 47 50 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r126 47 48 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r127 45 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.83
+ $Y2=0
r128 45 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.2
+ $Y2=0
r129 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r130 44 50 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r131 42 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r132 42 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r133 38 80 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.84 $Y=0.085
+ $X2=9.897 $Y2=0
r134 38 40 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=9.84 $Y=0.085
+ $X2=9.84 $Y2=0.635
r135 34 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.94 $Y=0.085
+ $X2=8.94 $Y2=0
r136 34 36 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.94 $Y=0.085
+ $X2=8.94 $Y2=0.635
r137 33 75 11.282 $w=8.33e-07 $l=4.35033e-07 $layer=LI1_cond $X=8.165 $Y=0
+ $X2=8.04 $Y2=0.377
r138 32 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=0 $X2=8.94
+ $Y2=0
r139 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.855 $Y=0 $X2=8.165
+ $Y2=0
r140 28 75 7.9472 $w=2.5e-07 $l=4.63e-07 $layer=LI1_cond $X=8.04 $Y=0.84
+ $X2=8.04 $Y2=0.377
r141 28 30 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.04 $Y=0.84
+ $X2=8.04 $Y2=1.005
r142 27 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r143 26 64 10.33 $w=8.33e-07 $l=4.05893e-07 $layer=LI1_cond $X=6.9 $Y=0 $X2=6.96
+ $Y2=0.377
r144 26 27 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.9 $Y=0 $X2=4.6
+ $Y2=0
r145 22 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r146 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.36
r147 18 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0
r148 18 20 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0.615
r149 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.49 $X2=9.8 $Y2=0.635
r150 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.8
+ $Y=0.49 $X2=8.94 $Y2=0.635
r151 3 74 91 $w=1.7e-07 $l=1.3763e-06 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.81 $X2=8 $Y2=0.325
r152 3 69 91 $w=1.7e-07 $l=8.95237e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.81 $X2=7.53 $Y2=0.325
r153 3 67 91 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.81 $X2=7.065 $Y2=0.325
r154 3 30 182 $w=1.7e-07 $l=1.32893e-06 $layer=licon1_NDIFF $count=1 $X=6.845
+ $Y=0.81 $X2=8.08 $Y2=1.005
r155 2 24 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.445 $X2=4.435 $Y2=0.36
r156 1 20 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.385 $X2=0.83 $Y2=0.615
.ends


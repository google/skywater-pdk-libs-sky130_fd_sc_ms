* File: sky130_fd_sc_ms__o311a_1.pxi.spice
* Created: Wed Sep  2 12:24:49 2020
* 
x_PM_SKY130_FD_SC_MS__O311A_1%C1 N_C1_M1010_g N_C1_M1004_g C1 N_C1_c_81_n
+ PM_SKY130_FD_SC_MS__O311A_1%C1
x_PM_SKY130_FD_SC_MS__O311A_1%B1 N_B1_M1002_g N_B1_M1008_g B1 N_B1_c_108_n
+ PM_SKY130_FD_SC_MS__O311A_1%B1
x_PM_SKY130_FD_SC_MS__O311A_1%A2 N_A2_M1007_g N_A2_M1003_g N_A2_c_141_n
+ N_A2_c_159_p N_A2_c_188_p N_A2_c_142_n N_A2_c_143_n A2 N_A2_c_144_n
+ N_A2_c_145_n PM_SKY130_FD_SC_MS__O311A_1%A2
x_PM_SKY130_FD_SC_MS__O311A_1%A3 N_A3_c_214_n N_A3_M1009_g N_A3_c_215_n
+ N_A3_c_216_n N_A3_c_210_n N_A3_M1005_g A3 A3 A3 N_A3_c_212_n N_A3_c_213_n
+ PM_SKY130_FD_SC_MS__O311A_1%A3
x_PM_SKY130_FD_SC_MS__O311A_1%A1 N_A1_M1001_g N_A1_M1000_g A1 N_A1_c_256_n
+ N_A1_c_257_n N_A1_c_258_n PM_SKY130_FD_SC_MS__O311A_1%A1
x_PM_SKY130_FD_SC_MS__O311A_1%A_31_387# N_A_31_387#_M1004_s N_A_31_387#_M1010_s
+ N_A_31_387#_M1008_d N_A_31_387#_M1011_g N_A_31_387#_M1006_g
+ N_A_31_387#_c_304_n N_A_31_387#_c_294_n N_A_31_387#_c_295_n
+ N_A_31_387#_c_296_n N_A_31_387#_c_297_n N_A_31_387#_c_307_n
+ N_A_31_387#_c_323_n N_A_31_387#_c_308_n N_A_31_387#_c_309_n
+ N_A_31_387#_c_298_n N_A_31_387#_c_299_n N_A_31_387#_c_300_n
+ N_A_31_387#_c_301_n N_A_31_387#_c_302_n PM_SKY130_FD_SC_MS__O311A_1%A_31_387#
x_PM_SKY130_FD_SC_MS__O311A_1%VPWR N_VPWR_M1010_d N_VPWR_M1001_d N_VPWR_c_416_n
+ N_VPWR_c_417_n VPWR N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n
+ N_VPWR_c_415_n N_VPWR_c_422_n N_VPWR_c_423_n PM_SKY130_FD_SC_MS__O311A_1%VPWR
x_PM_SKY130_FD_SC_MS__O311A_1%X N_X_M1006_d N_X_M1011_d N_X_c_469_n N_X_c_470_n
+ N_X_c_466_n X X X PM_SKY130_FD_SC_MS__O311A_1%X
x_PM_SKY130_FD_SC_MS__O311A_1%A_209_74# N_A_209_74#_M1002_d N_A_209_74#_M1005_d
+ N_A_209_74#_c_493_n N_A_209_74#_c_496_n N_A_209_74#_c_494_n
+ PM_SKY130_FD_SC_MS__O311A_1%A_209_74#
x_PM_SKY130_FD_SC_MS__O311A_1%VGND N_VGND_M1007_d N_VGND_M1000_d N_VGND_c_521_n
+ N_VGND_c_512_n VGND N_VGND_c_513_n N_VGND_c_514_n N_VGND_c_515_n
+ N_VGND_c_516_n PM_SKY130_FD_SC_MS__O311A_1%VGND
cc_1 VNB N_C1_M1010_g 0.0154393f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.435
cc_2 VNB N_C1_M1004_g 0.02469f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_3 VNB C1 0.0121164f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_C1_c_81_n 0.0546617f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_5 VNB N_B1_M1002_g 0.0196196f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.435
cc_6 VNB N_B1_M1008_g 0.0130036f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_7 VNB B1 0.00308495f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_B1_c_108_n 0.0295848f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_9 VNB N_A2_M1007_g 0.0210444f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.435
cc_10 VNB N_A2_c_141_n 0.00351602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_142_n 0.00486902f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.305
cc_12 VNB N_A2_c_143_n 0.0257001f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_13 VNB N_A2_c_144_n 0.0298977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_145_n 0.00245544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_210_n 0.0114682f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_16 VNB A3 0.00138988f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_17 VNB N_A3_c_212_n 0.0473444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A3_c_213_n 0.0213502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1001_g 0.011579f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.435
cc_20 VNB N_A1_c_256_n 0.0340747f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_21 VNB N_A1_c_257_n 0.0166185f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_22 VNB N_A1_c_258_n 0.0221309f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_23 VNB N_A_31_387#_M1006_g 0.0312993f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_24 VNB N_A_31_387#_c_294_n 0.019793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_31_387#_c_295_n 0.00527983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_31_387#_c_296_n 0.0106214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_31_387#_c_297_n 0.00304476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_31_387#_c_298_n 0.00424542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_31_387#_c_299_n 7.98615e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_31_387#_c_300_n 0.00695823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_31_387#_c_301_n 0.00336822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_31_387#_c_302_n 0.0291511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_415_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_466_n 0.0250799f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.305
cc_35 VNB X 0.0267037f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.305
cc_36 VNB X 0.013364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_209_74#_c_493_n 0.00406087f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.69
cc_38 VNB N_A_209_74#_c_494_n 0.0147102f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.305
cc_39 VNB N_VGND_c_512_n 0.00647919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_513_n 0.0873829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_514_n 0.0193554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_515_n 0.261122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_516_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C1_M1010_g 0.034242f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.435
cc_45 VPB N_B1_M1008_g 0.0272449f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.69
cc_46 VPB N_A2_M1003_g 0.0253086f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.69
cc_47 VPB N_A2_c_141_n 0.00176822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A2_c_142_n 0.00100657f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.305
cc_49 VPB N_A2_c_143_n 0.0129975f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.305
cc_50 VPB N_A3_c_214_n 0.0193107f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.47
cc_51 VPB N_A3_c_215_n 0.0362831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A3_c_216_n 0.00787f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.14
cc_53 VPB N_A3_c_210_n 0.00271961f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.69
cc_54 VPB A3 0.00232472f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.305
cc_55 VPB N_A1_M1001_g 0.0284942f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.435
cc_56 VPB N_A_31_387#_M1011_g 0.0280254f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.305
cc_57 VPB N_A_31_387#_c_304_n 0.0473207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_31_387#_c_296_n 0.00309737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_31_387#_c_297_n 0.00935005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_31_387#_c_307_n 0.00241627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_31_387#_c_308_n 0.0116725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_31_387#_c_309_n 9.36467e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_31_387#_c_298_n 0.00552399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_31_387#_c_299_n 7.96937e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_31_387#_c_301_n 0.00296303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_31_387#_c_302_n 0.00563363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_416_n 0.0115806f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_68 VPB N_VPWR_c_417_n 0.0105221f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.305
cc_69 VPB N_VPWR_c_418_n 0.0198977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_419_n 0.0607653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_420_n 0.0193973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_415_n 0.081852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_422_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_423_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_X_c_469_n 0.0366174f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_76 VPB N_X_c_470_n 0.00768928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_X_c_466_n 0.0132127f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.305
cc_78 N_C1_M1004_g N_B1_M1002_g 0.0311169f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_79 N_C1_M1010_g N_B1_M1008_g 0.0169558f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_80 N_C1_c_81_n B1 3.30694e-19 $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_81 N_C1_c_81_n N_B1_c_108_n 0.0311169f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_82 N_C1_M1010_g N_A_31_387#_c_304_n 0.0180387f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_83 N_C1_M1004_g N_A_31_387#_c_294_n 0.00844889f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_84 N_C1_M1010_g N_A_31_387#_c_295_n 0.00863954f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_85 N_C1_M1004_g N_A_31_387#_c_295_n 0.00858018f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_86 C1 N_A_31_387#_c_295_n 0.0233985f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_C1_c_81_n N_A_31_387#_c_295_n 0.00911304f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_88 N_C1_M1010_g N_A_31_387#_c_297_n 0.0195228f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_89 C1 N_A_31_387#_c_297_n 0.0206681f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_C1_c_81_n N_A_31_387#_c_297_n 0.00704075f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_91 N_C1_M1010_g N_A_31_387#_c_323_n 5.88427e-19 $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_92 N_C1_M1004_g N_A_31_387#_c_300_n 0.00848905f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_93 C1 N_A_31_387#_c_300_n 0.0155323f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_C1_c_81_n N_A_31_387#_c_300_n 0.00717614f $X=0.58 $Y=1.305 $X2=0 $Y2=0
cc_95 N_C1_M1010_g N_VPWR_c_416_n 0.00346378f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_96 N_C1_M1010_g N_VPWR_c_418_n 0.00640648f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_97 N_C1_M1010_g N_VPWR_c_415_n 0.00645424f $X=0.525 $Y=2.435 $X2=0 $Y2=0
cc_98 N_C1_M1004_g N_VGND_c_513_n 0.00434272f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_99 N_C1_M1004_g N_VGND_c_515_n 0.00442932f $X=0.58 $Y=0.69 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_A2_M1007_g 0.0159664f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_101 N_B1_M1008_g N_A2_c_141_n 0.00467318f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_102 B1 N_A2_c_144_n 0.00193925f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_108_n N_A2_c_144_n 0.020587f $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_104 B1 N_A2_c_145_n 0.0265356f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B1_c_108_n N_A2_c_145_n 3.50521e-19 $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_106 N_B1_M1008_g N_A3_c_216_n 0.0170362f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_107 N_B1_M1008_g N_A_31_387#_c_304_n 6.25242e-19 $X=1.075 $Y=2.435 $X2=0
+ $Y2=0
cc_108 N_B1_M1002_g N_A_31_387#_c_294_n 0.00129834f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_A_31_387#_c_295_n 0.00553928f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_110 N_B1_M1008_g N_A_31_387#_c_295_n 0.00341339f $X=1.075 $Y=2.435 $X2=0
+ $Y2=0
cc_111 B1 N_A_31_387#_c_295_n 0.0249634f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B1_M1008_g N_A_31_387#_c_296_n 0.0168875f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_113 B1 N_A_31_387#_c_296_n 0.0283256f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B1_c_108_n N_A_31_387#_c_296_n 0.00414882f $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_115 N_B1_M1008_g N_A_31_387#_c_307_n 0.00246751f $X=1.075 $Y=2.435 $X2=0
+ $Y2=0
cc_116 N_B1_M1008_g N_A_31_387#_c_323_n 0.0141124f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_117 N_B1_M1002_g N_A_31_387#_c_300_n 0.00138573f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_118 N_B1_M1008_g N_VPWR_c_416_n 0.00346343f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_119 N_B1_M1008_g N_VPWR_c_419_n 0.00639579f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_120 N_B1_M1008_g N_VPWR_c_415_n 0.00645424f $X=1.075 $Y=2.435 $X2=0 $Y2=0
cc_121 N_B1_M1002_g N_A_209_74#_c_493_n 0.00276611f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_122 B1 N_A_209_74#_c_496_n 0.0169224f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B1_c_108_n N_A_209_74#_c_496_n 0.00410213f $X=1.06 $Y=1.305 $X2=0 $Y2=0
cc_124 N_B1_M1002_g N_VGND_c_513_n 0.00461464f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_125 N_B1_M1002_g N_VGND_c_515_n 0.00910057f $X=0.97 $Y=0.69 $X2=0 $Y2=0
cc_126 N_A2_c_141_n N_A3_c_214_n 0.00974807f $X=1.72 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A2_M1003_g N_A3_c_215_n 0.00551412f $X=2.605 $Y=2.435 $X2=0 $Y2=0
cc_128 N_A2_c_141_n N_A3_c_215_n 0.0123672f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_129 N_A2_c_159_p N_A3_c_215_n 0.00484151f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_130 N_A2_c_145_n N_A3_c_215_n 2.41637e-19 $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_131 N_A2_c_144_n N_A3_c_216_n 0.0196974f $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_132 N_A2_c_145_n N_A3_c_216_n 0.0012802f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_133 N_A2_c_141_n N_A3_c_210_n 0.00456493f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_134 N_A2_c_142_n N_A3_c_210_n 4.02794e-19 $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_135 N_A2_c_143_n N_A3_c_210_n 0.00551412f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_136 N_A2_c_141_n A3 0.0510888f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_137 N_A2_c_159_p A3 0.0266856f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_138 N_A2_c_142_n A3 0.0472442f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_139 N_A2_c_143_n A3 0.00888973f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_140 N_A2_c_144_n A3 3.76918e-19 $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_141 N_A2_c_145_n A3 0.02617f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_142 N_A2_M1007_g N_A3_c_212_n 0.00206579f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_143 N_A2_c_143_n N_A3_c_212_n 3.04703e-19 $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_144 N_A2_c_144_n N_A3_c_212_n 0.0205549f $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_145 N_A2_c_145_n N_A3_c_212_n 0.00184761f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_146 N_A2_M1007_g N_A3_c_213_n 0.0166563f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_147 N_A2_M1003_g N_A1_M1001_g 0.0371701f $X=2.605 $Y=2.435 $X2=0 $Y2=0
cc_148 N_A2_c_159_p N_A1_M1001_g 6.21929e-19 $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_149 N_A2_c_142_n N_A1_M1001_g 0.00304909f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_150 N_A2_c_143_n N_A1_M1001_g 0.0177236f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_151 N_A2_c_143_n N_A1_c_256_n 3.52691e-19 $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_152 N_A2_c_141_n N_A_31_387#_c_296_n 0.0135297f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_153 N_A2_c_144_n N_A_31_387#_c_296_n 6.39279e-19 $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_154 N_A2_c_145_n N_A_31_387#_c_296_n 8.43332e-19 $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_155 N_A2_c_141_n N_A_31_387#_c_323_n 0.02354f $X=1.72 $Y=2.32 $X2=0 $Y2=0
cc_156 N_A2_M1003_g N_A_31_387#_c_308_n 0.0146238f $X=2.605 $Y=2.435 $X2=0 $Y2=0
cc_157 N_A2_c_159_p N_A_31_387#_c_308_n 0.0412579f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_158 N_A2_c_188_p N_A_31_387#_c_308_n 0.00648054f $X=1.805 $Y=2.405 $X2=0
+ $Y2=0
cc_159 N_A2_M1003_g N_A_31_387#_c_309_n 0.00707496f $X=2.605 $Y=2.435 $X2=0
+ $Y2=0
cc_160 N_A2_c_159_p N_A_31_387#_c_309_n 0.0138307f $X=2.515 $Y=2.405 $X2=0 $Y2=0
cc_161 N_A2_c_142_n N_A_31_387#_c_309_n 0.0408384f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_162 N_A2_c_142_n N_A_31_387#_c_299_n 0.0142132f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_163 N_A2_c_143_n N_A_31_387#_c_299_n 9.90056e-19 $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_164 N_A2_M1003_g N_VPWR_c_419_n 0.00479416f $X=2.605 $Y=2.435 $X2=0 $Y2=0
cc_165 N_A2_M1003_g N_VPWR_c_415_n 0.00645424f $X=2.605 $Y=2.435 $X2=0 $Y2=0
cc_166 N_A2_c_141_n A_323_387# 0.0107778f $X=1.72 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_167 N_A2_c_159_p A_323_387# 0.0253796f $X=2.515 $Y=2.405 $X2=-0.19 $Y2=-0.245
cc_168 N_A2_c_188_p A_323_387# 0.00310345f $X=1.805 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A2_c_159_p A_539_387# 0.00281032f $X=2.515 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A2_c_142_n A_539_387# 0.00336566f $X=2.68 $Y=1.61 $X2=-0.19 $Y2=-0.245
cc_171 N_A2_M1007_g N_A_209_74#_c_494_n 0.0203628f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_172 N_A2_c_145_n N_A_209_74#_c_494_n 0.00310605f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_173 N_A2_M1007_g N_VGND_c_521_n 0.0056177f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_174 N_A2_c_142_n N_VGND_c_521_n 0.0111729f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_175 N_A2_c_143_n N_VGND_c_521_n 0.00178249f $X=2.68 $Y=1.61 $X2=0 $Y2=0
cc_176 N_A2_c_144_n N_VGND_c_521_n 0.00385043f $X=1.6 $Y=1.305 $X2=0 $Y2=0
cc_177 N_A2_c_145_n N_VGND_c_521_n 0.0148018f $X=1.72 $Y=1.305 $X2=0 $Y2=0
cc_178 N_A2_M1007_g N_VGND_c_513_n 0.00281891f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_179 N_A2_M1007_g N_VGND_c_515_n 0.00357277f $X=1.51 $Y=0.69 $X2=0 $Y2=0
cc_180 N_A3_c_216_n N_A_31_387#_c_296_n 0.00301767f $X=1.615 $Y=1.785 $X2=0
+ $Y2=0
cc_181 N_A3_c_214_n N_A_31_387#_c_307_n 9.84805e-19 $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_182 N_A3_c_214_n N_A_31_387#_c_323_n 0.0211914f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_183 N_A3_c_216_n N_A_31_387#_c_323_n 0.00139178f $X=1.615 $Y=1.785 $X2=0
+ $Y2=0
cc_184 N_A3_c_214_n N_A_31_387#_c_308_n 0.0145796f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_185 N_A3_c_214_n N_VPWR_c_419_n 0.00479391f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_186 N_A3_c_214_n N_VPWR_c_415_n 0.00645424f $X=1.525 $Y=1.86 $X2=0 $Y2=0
cc_187 A3 A_323_387# 0.0096356f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_188 N_A3_c_213_n N_A_209_74#_c_494_n 0.0159594f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_189 A3 N_VGND_c_521_n 0.0233403f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A3_c_212_n N_VGND_c_521_n 0.00471366f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_191 N_A3_c_213_n N_VGND_c_521_n 0.0136627f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_192 N_A3_c_213_n N_VGND_c_513_n 0.00281891f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_193 N_A3_c_213_n N_VGND_c_515_n 0.00361247f $X=2.14 $Y=1.085 $X2=0 $Y2=0
cc_194 N_A1_M1001_g N_A_31_387#_M1011_g 0.0182893f $X=3.175 $Y=2.435 $X2=0 $Y2=0
cc_195 N_A1_c_257_n N_A_31_387#_M1006_g 0.00133094f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_196 N_A1_c_258_n N_A_31_387#_M1006_g 0.022713f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_197 N_A1_M1001_g N_A_31_387#_c_308_n 0.00638395f $X=3.175 $Y=2.435 $X2=0
+ $Y2=0
cc_198 N_A1_M1001_g N_A_31_387#_c_309_n 0.0251614f $X=3.175 $Y=2.435 $X2=0 $Y2=0
cc_199 N_A1_M1001_g N_A_31_387#_c_298_n 0.00814558f $X=3.175 $Y=2.435 $X2=0
+ $Y2=0
cc_200 N_A1_c_256_n N_A_31_387#_c_298_n 0.00316326f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_201 N_A1_c_257_n N_A_31_387#_c_298_n 0.0146979f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_202 N_A1_M1001_g N_A_31_387#_c_299_n 0.00382034f $X=3.175 $Y=2.435 $X2=0
+ $Y2=0
cc_203 N_A1_c_256_n N_A_31_387#_c_299_n 6.9887e-19 $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_204 N_A1_c_257_n N_A_31_387#_c_299_n 0.0140509f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_205 N_A1_M1001_g N_A_31_387#_c_301_n 0.00118148f $X=3.175 $Y=2.435 $X2=0
+ $Y2=0
cc_206 N_A1_c_257_n N_A_31_387#_c_301_n 0.00631056f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_207 N_A1_M1001_g N_A_31_387#_c_302_n 0.00908926f $X=3.175 $Y=2.435 $X2=0
+ $Y2=0
cc_208 N_A1_c_256_n N_A_31_387#_c_302_n 0.0063017f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_209 N_A1_c_257_n N_A_31_387#_c_302_n 3.45132e-19 $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_210 N_A1_M1001_g N_VPWR_c_417_n 0.0120593f $X=3.175 $Y=2.435 $X2=0 $Y2=0
cc_211 N_A1_M1001_g N_VPWR_c_419_n 0.00564767f $X=3.175 $Y=2.435 $X2=0 $Y2=0
cc_212 N_A1_M1001_g N_VPWR_c_415_n 0.00645424f $X=3.175 $Y=2.435 $X2=0 $Y2=0
cc_213 N_A1_c_257_n X 2.93139e-19 $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_214 N_A1_c_258_n X 6.59557e-19 $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_215 N_A1_c_258_n N_A_209_74#_c_494_n 0.00664776f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_216 N_A1_c_256_n N_VGND_c_521_n 0.00450164f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_217 N_A1_c_257_n N_VGND_c_521_n 0.0251429f $X=3.22 $Y=1.285 $X2=0 $Y2=0
cc_218 N_A1_c_258_n N_VGND_c_521_n 0.0111167f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_219 N_A1_c_258_n N_VGND_c_512_n 0.0146844f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_220 N_A1_c_258_n N_VGND_c_513_n 0.00383152f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_221 N_A1_c_258_n N_VGND_c_515_n 0.00374822f $X=3.22 $Y=1.12 $X2=0 $Y2=0
cc_222 N_A_31_387#_c_304_n N_VPWR_c_416_n 0.0373748f $X=0.3 $Y=2.08 $X2=0 $Y2=0
cc_223 N_A_31_387#_c_297_n N_VPWR_c_416_n 0.0238529f $X=0.75 $Y=1.725 $X2=0
+ $Y2=0
cc_224 N_A_31_387#_c_307_n N_VPWR_c_416_n 0.0079549f $X=1.3 $Y=2.785 $X2=0 $Y2=0
cc_225 N_A_31_387#_M1011_g N_VPWR_c_417_n 0.00389287f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_226 N_A_31_387#_c_308_n N_VPWR_c_417_n 0.0140386f $X=3.015 $Y=2.87 $X2=0
+ $Y2=0
cc_227 N_A_31_387#_c_309_n N_VPWR_c_417_n 0.06101f $X=3.1 $Y=2.785 $X2=0 $Y2=0
cc_228 N_A_31_387#_c_298_n N_VPWR_c_417_n 0.0197628f $X=3.595 $Y=1.705 $X2=0
+ $Y2=0
cc_229 N_A_31_387#_c_301_n N_VPWR_c_417_n 0.00620567f $X=3.76 $Y=1.515 $X2=0
+ $Y2=0
cc_230 N_A_31_387#_c_302_n N_VPWR_c_417_n 4.41165e-19 $X=3.76 $Y=1.515 $X2=0
+ $Y2=0
cc_231 N_A_31_387#_c_304_n N_VPWR_c_418_n 0.0132154f $X=0.3 $Y=2.08 $X2=0 $Y2=0
cc_232 N_A_31_387#_c_307_n N_VPWR_c_419_n 0.0131906f $X=1.3 $Y=2.785 $X2=0 $Y2=0
cc_233 N_A_31_387#_c_308_n N_VPWR_c_419_n 0.0626603f $X=3.015 $Y=2.87 $X2=0
+ $Y2=0
cc_234 N_A_31_387#_M1011_g N_VPWR_c_420_n 0.005209f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_31_387#_M1011_g N_VPWR_c_415_n 0.00990536f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_236 N_A_31_387#_c_304_n N_VPWR_c_415_n 0.0119049f $X=0.3 $Y=2.08 $X2=0 $Y2=0
cc_237 N_A_31_387#_c_307_n N_VPWR_c_415_n 0.011945f $X=1.3 $Y=2.785 $X2=0 $Y2=0
cc_238 N_A_31_387#_c_308_n N_VPWR_c_415_n 0.0596823f $X=3.015 $Y=2.87 $X2=0
+ $Y2=0
cc_239 N_A_31_387#_c_308_n A_323_387# 0.015221f $X=3.015 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_31_387#_c_308_n A_539_387# 0.00795586f $X=3.015 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_241 N_A_31_387#_c_309_n A_539_387# 0.00876676f $X=3.1 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_242 N_A_31_387#_M1011_g N_X_c_469_n 0.0101633f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_31_387#_M1011_g N_X_c_470_n 0.00257732f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_31_387#_c_301_n N_X_c_470_n 0.0027288f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_245 N_A_31_387#_M1011_g N_X_c_466_n 0.00490693f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A_31_387#_M1006_g N_X_c_466_n 0.00580334f $X=3.82 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_31_387#_c_301_n N_X_c_466_n 0.0332754f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A_31_387#_c_302_n N_X_c_466_n 0.00766421f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A_31_387#_M1006_g X 0.00812529f $X=3.82 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_31_387#_M1006_g X 0.0042952f $X=3.82 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_31_387#_c_301_n X 0.00153012f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_252 N_A_31_387#_c_302_n X 0.0012634f $X=3.76 $Y=1.515 $X2=0 $Y2=0
cc_253 N_A_31_387#_c_295_n A_131_74# 5.66122e-19 $X=0.665 $Y=1.64 $X2=-0.19
+ $Y2=-0.245
cc_254 N_A_31_387#_c_300_n A_131_74# 0.00269364f $X=0.665 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_255 N_A_31_387#_c_294_n N_A_209_74#_c_493_n 0.00424699f $X=0.365 $Y=0.515
+ $X2=0 $Y2=0
cc_256 N_A_31_387#_c_296_n N_A_209_74#_c_496_n 0.00334383f $X=1.135 $Y=1.725
+ $X2=0 $Y2=0
cc_257 N_A_31_387#_c_298_n N_VGND_c_521_n 0.00547315f $X=3.595 $Y=1.705 $X2=0
+ $Y2=0
cc_258 N_A_31_387#_c_301_n N_VGND_c_521_n 0.00405649f $X=3.76 $Y=1.515 $X2=0
+ $Y2=0
cc_259 N_A_31_387#_c_302_n N_VGND_c_521_n 6.53733e-19 $X=3.76 $Y=1.515 $X2=0
+ $Y2=0
cc_260 N_A_31_387#_M1006_g N_VGND_c_512_n 0.00538108f $X=3.82 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_31_387#_c_294_n N_VGND_c_513_n 0.0141395f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_262 N_A_31_387#_M1006_g N_VGND_c_514_n 0.00434272f $X=3.82 $Y=0.74 $X2=0
+ $Y2=0
cc_263 N_A_31_387#_M1006_g N_VGND_c_515_n 0.00824752f $X=3.82 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_31_387#_c_294_n N_VGND_c_515_n 0.0118342f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_265 N_A_31_387#_c_300_n N_VGND_c_515_n 0.00703783f $X=0.665 $Y=0.885 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_420_n N_X_c_469_n 0.01678f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_415_n N_X_c_469_n 0.0138209f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_417_n N_X_c_470_n 0.0398603f $X=3.52 $Y=2.125 $X2=0 $Y2=0
cc_269 X N_VGND_c_512_n 0.0164106f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_270 X N_VGND_c_514_n 0.0161257f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_271 X N_VGND_c_515_n 0.013291f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_272 N_A_209_74#_c_494_n N_VGND_M1007_d 0.00743158f $X=3.015 $Y=0.525
+ $X2=-0.19 $Y2=-0.245
cc_273 N_A_209_74#_M1005_d N_VGND_c_521_n 0.0325693f $X=2.305 $Y=0.37 $X2=0
+ $Y2=0
cc_274 N_A_209_74#_c_494_n N_VGND_c_521_n 0.106422f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
cc_275 N_A_209_74#_c_494_n N_VGND_c_512_n 0.0157478f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
cc_276 N_A_209_74#_c_493_n N_VGND_c_513_n 0.0204446f $X=1.225 $Y=0.61 $X2=0
+ $Y2=0
cc_277 N_A_209_74#_c_494_n N_VGND_c_513_n 0.103511f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0
cc_278 N_A_209_74#_c_493_n N_VGND_c_515_n 0.0126791f $X=1.225 $Y=0.61 $X2=0
+ $Y2=0
cc_279 N_A_209_74#_c_494_n N_VGND_c_515_n 0.0659666f $X=3.015 $Y=0.525 $X2=0
+ $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__or2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__or2b_1 A B_N VGND VNB VPB VPWR X
M1000 a_264_368# a_27_112# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=7.357e+11p ps=5.01e+06u
M1001 VGND A a_264_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_264_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=7.218e+11p ps=5.39e+06u
M1003 VGND B_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.685e+11p ps=2.44e+06u
M1004 a_356_368# a_27_112# a_264_368# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1005 VPWR B_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1006 VPWR A a_356_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_264_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


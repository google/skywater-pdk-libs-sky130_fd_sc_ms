* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_119_392# A2 a_203_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VPWR a_203_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_27_74# a_281_244# a_203_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_281_244# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 VGND a_203_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_203_392# a_281_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 VPWR A1 a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_281_244# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__clkbuf_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__clkbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.058400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.360000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 0.350000 2.660000 2.120000 ;
        RECT 2.430000 2.120000 2.660000 2.980000 ;
        RECT 3.275000 0.350000 3.500000 1.690000 ;
        RECT 3.275000 1.690000 3.545000 1.860000 ;
        RECT 3.340000 1.860000 3.545000 2.980000 ;
        RECT 4.075000 0.350000 4.340000 0.745000 ;
        RECT 4.170000 0.745000 4.340000 1.690000 ;
        RECT 4.170000 1.690000 4.430000 1.860000 ;
        RECT 4.230000 1.860000 4.430000 2.980000 ;
        RECT 5.025000 0.350000 5.255000 1.690000 ;
        RECT 5.025000 1.690000 5.350000 1.860000 ;
        RECT 5.140000 1.860000 5.350000 2.980000 ;
        RECT 5.935000 0.350000 6.185000 1.690000 ;
        RECT 5.935000 1.690000 6.245000 1.860000 ;
        RECT 6.040000 1.860000 6.245000 2.980000 ;
        RECT 6.865000 0.350000 7.115000 1.690000 ;
        RECT 6.865000 1.690000 7.150000 1.860000 ;
        RECT 6.945000 1.860000 7.150000 2.980000 ;
        RECT 7.795000 0.350000 8.045000 1.690000 ;
        RECT 7.795000 1.690000 8.050000 1.860000 ;
        RECT 7.840000 1.860000 8.050000 2.980000 ;
        RECT 8.725000 0.350000 8.975000 1.830000 ;
        RECT 8.725000 1.830000 8.970000 1.860000 ;
        RECT 8.750000 1.860000 8.970000 2.980000 ;
      LAYER mcon ;
        RECT 2.460000 1.950000 2.630000 2.120000 ;
        RECT 3.360000 1.950000 3.530000 2.120000 ;
        RECT 4.245000 1.950000 4.415000 2.120000 ;
        RECT 5.160000 1.950000 5.330000 2.120000 ;
        RECT 6.060000 1.950000 6.230000 2.120000 ;
        RECT 6.960000 1.950000 7.130000 2.120000 ;
        RECT 7.860000 1.950000 8.030000 2.120000 ;
        RECT 8.780000 1.950000 8.950000 2.120000 ;
      LAYER met1 ;
        RECT 2.390000 1.920000 9.090000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 0.115000  0.085000 0.365000 0.810000 ;
        RECT 0.975000  0.085000 1.225000 0.810000 ;
        RECT 1.855000  0.085000 2.185000 0.810000 ;
        RECT 2.865000  0.085000 3.035000 0.680000 ;
        RECT 3.670000  0.085000 3.895000 0.725000 ;
        RECT 4.510000  0.085000 4.835000 0.740000 ;
        RECT 5.435000  0.085000 5.765000 0.680000 ;
        RECT 6.365000  0.085000 6.695000 0.680000 ;
        RECT 7.295000  0.085000 7.625000 0.680000 ;
        RECT 8.225000  0.085000 8.555000 0.680000 ;
        RECT 9.155000  0.085000 9.485000 0.745000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.120000 1.950000 0.370000 3.245000 ;
        RECT 1.100000 2.290000 1.270000 3.245000 ;
        RECT 2.000000 2.290000 2.250000 3.245000 ;
        RECT 2.830000 2.030000 3.160000 3.245000 ;
        RECT 3.730000 2.030000 4.060000 3.245000 ;
        RECT 4.630000 2.030000 4.960000 3.245000 ;
        RECT 5.530000 2.030000 5.860000 3.245000 ;
        RECT 6.430000 2.030000 6.760000 3.245000 ;
        RECT 7.330000 2.030000 7.660000 3.245000 ;
        RECT 8.230000 2.030000 8.560000 3.245000 ;
        RECT 9.150000 2.030000 9.480000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545000 0.350000 0.795000 0.980000 ;
      RECT 0.545000 0.980000 2.135000 1.150000 ;
      RECT 0.570000 1.950000 2.135000 2.120000 ;
      RECT 0.570000 2.120000 0.900000 2.980000 ;
      RECT 1.425000 0.350000 1.675000 0.980000 ;
      RECT 1.470000 2.120000 1.800000 2.980000 ;
      RECT 1.965000 1.150000 2.135000 1.180000 ;
      RECT 1.965000 1.180000 2.210000 1.410000 ;
      RECT 1.965000 1.410000 2.135000 1.950000 ;
      RECT 2.835000 1.190000 3.105000 1.520000 ;
      RECT 3.670000 1.190000 4.000000 1.520000 ;
      RECT 4.510000 1.190000 4.840000 1.520000 ;
      RECT 5.425000 1.190000 5.755000 1.520000 ;
      RECT 6.365000 1.190000 6.695000 1.520000 ;
      RECT 7.295000 1.190000 7.625000 1.520000 ;
      RECT 8.225000 1.190000 8.555000 1.520000 ;
    LAYER mcon ;
      RECT 2.010000 1.210000 2.180000 1.380000 ;
      RECT 2.890000 1.210000 3.060000 1.380000 ;
      RECT 3.750000 1.210000 3.920000 1.380000 ;
      RECT 4.590000 1.210000 4.760000 1.380000 ;
      RECT 5.505000 1.210000 5.675000 1.380000 ;
      RECT 6.445000 1.210000 6.615000 1.380000 ;
      RECT 7.375000 1.210000 7.545000 1.380000 ;
      RECT 8.305000 1.210000 8.475000 1.380000 ;
    LAYER met1 ;
      RECT 1.940000 1.180000 8.640000 1.410000 ;
  END
END sky130_fd_sc_ms__clkbuf_16

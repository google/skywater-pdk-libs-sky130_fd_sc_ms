* File: sky130_fd_sc_ms__o221a_1.pex.spice
* Created: Wed Sep  2 12:22:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O221A_1%A_83_264# 1 2 3 12 16 19 20 21 24 26 30 33
+ 35 36 40 42 46
c96 40 0 4.75931e-20 $X=1.89 $Y=2.115
c97 19 0 1.2498e-19 $X=0.7 $Y=1.95
r98 42 44 15.698 $w=4.33e-07 $l=4.25e-07 $layer=LI1_cond $X=3.987 $Y=0.525
+ $X2=3.987 $Y2=0.95
r99 36 49 40.9837 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.485
+ $X2=0.6 $Y2=1.65
r100 36 48 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.485
+ $X2=0.6 $Y2=1.32
r101 35 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=1.485
+ $X2=0.62 $Y2=1.65
r102 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.485 $X2=0.62 $Y2=1.485
r103 33 46 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.12 $Y=1.96
+ $X2=4.04 $Y2=2.045
r104 33 44 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.12 $Y=1.96
+ $X2=4.12 $Y2=0.95
r105 28 46 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.13
+ $X2=4.04 $Y2=2.045
r106 28 30 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.04 $Y=2.13
+ $X2=4.04 $Y2=2.815
r107 27 40 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.055 $Y=2.045
+ $X2=1.89 $Y2=2.04
r108 26 46 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.045
+ $X2=4.04 $Y2=2.045
r109 26 27 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=3.875 $Y=2.045
+ $X2=2.055 $Y2=2.045
r110 22 40 0.89609 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.89 $Y=2.13 $X2=1.89
+ $Y2=2.04
r111 22 24 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.89 $Y=2.13
+ $X2=1.89 $Y2=2.815
r112 20 40 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.725 $Y=2.035
+ $X2=1.89 $Y2=2.04
r113 20 21 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.725 $Y=2.035
+ $X2=0.785 $Y2=2.035
r114 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.95
+ $X2=0.785 $Y2=2.035
r115 19 38 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.7 $Y=1.95 $X2=0.7
+ $Y2=1.65
r116 16 48 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.57 $Y=0.74
+ $X2=0.57 $Y2=1.32
r117 12 49 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.65
r118 3 46 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.96 $X2=4.04 $Y2=2.125
r119 3 30 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.96 $X2=4.04 $Y2=2.815
r120 2 40 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=1.96 $X2=1.89 $Y2=2.115
r121 2 24 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=1.96 $X2=1.89 $Y2=2.815
r122 1 42 91 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=2 $X=3.725
+ $Y=0.37 $X2=3.935 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%A1 3 7 9 12
c39 12 0 9.50927e-20 $X=1.17 $Y=1.615
c40 7 0 4.75931e-20 $X=1.245 $Y=2.46
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.78
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.45
r43 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r44 7 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.245 $Y=2.46
+ $X2=1.245 $Y2=1.78
r45 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.15 $Y=0.79 $X2=1.15
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%A2 3 7 9 12
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.78
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.45
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r38 7 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.665 $Y=2.46
+ $X2=1.665 $Y2=1.78
r39 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.65 $Y=0.79 $X2=1.65
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%B2 5 7 8 9 11 12 15 17
c44 5 0 3.89885e-20 $X=2.235 $Y=2.46
r45 15 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.615
+ $X2=2.31 $Y2=1.78
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.615 $X2=2.31 $Y2=1.615
r47 12 16 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.31 $Y2=1.615
r48 9 11 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.72 $Y=1.1 $X2=2.72
+ $Y2=0.69
r49 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.645 $Y=1.175
+ $X2=2.72 $Y2=1.1
r50 7 8 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.645 $Y=1.175
+ $X2=2.475 $Y2=1.175
r51 5 17 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.235 $Y=2.46
+ $X2=2.235 $Y2=1.78
r52 1 8 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.31 $Y=1.25
+ $X2=2.475 $Y2=1.175
r53 1 15 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.31 $Y=1.25
+ $X2=2.31 $Y2=1.615
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%B1 3 7 9 13
c36 9 0 3.89885e-20 $X=3.12 $Y=1.665
r37 13 15 11.1231 $w=2.6e-07 $l=6e-08 $layer=POLY_cond $X=3.09 $Y=1.625 $X2=3.15
+ $Y2=1.625
r38 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.625 $X2=3.09 $Y2=1.625
r39 5 15 15.628 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.46 $X2=3.15
+ $Y2=1.625
r40 5 7 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.15 $Y=1.46 $X2=3.15
+ $Y2=0.69
r41 1 13 52.8346 $w=2.6e-07 $l=3.5812e-07 $layer=POLY_cond $X=2.805 $Y=1.79
+ $X2=3.09 $Y2=1.625
r42 1 3 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=2.805 $Y=1.79
+ $X2=2.805 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%C1 2 5 8 10 11 12 16 18
c37 18 0 4.4527e-20 $X=3.7 $Y=1.12
c38 16 0 1.66579e-19 $X=3.66 $Y=1.285
r39 16 18 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=3.7 $Y=1.285
+ $X2=3.7 $Y2=1.12
r40 11 12 12.8802 $w=3.38e-07 $l=3.8e-07 $layer=LI1_cond $X=3.655 $Y=1.285
+ $X2=3.655 $Y2=1.665
r41 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.66
+ $Y=1.285 $X2=3.66 $Y2=1.285
r42 8 10 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=3.815 $Y=2.46
+ $X2=3.815 $Y2=1.79
r43 5 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.65 $Y=0.69 $X2=3.65
+ $Y2=1.12
r44 2 10 45.5979 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=3.7 $Y=1.585 $X2=3.7
+ $Y2=1.79
r45 1 16 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=3.7 $Y=1.325 $X2=3.7
+ $Y2=1.285
r46 1 2 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=3.7 $Y=1.325 $X2=3.7
+ $Y2=1.585
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%X 1 2 11 13 15 16 17 23 29
r23 21 29 0.0853661 $w=4.03e-07 $l=3e-09 $layer=LI1_cond $X=0.317 $Y=0.928
+ $X2=0.317 $Y2=0.925
r24 17 31 8.55498 $w=4.03e-07 $l=1.61e-07 $layer=LI1_cond $X=0.317 $Y=0.969
+ $X2=0.317 $Y2=1.13
r25 17 21 1.16667 $w=4.03e-07 $l=4.1e-08 $layer=LI1_cond $X=0.317 $Y=0.969
+ $X2=0.317 $Y2=0.928
r26 17 29 1.16667 $w=4.03e-07 $l=4.1e-08 $layer=LI1_cond $X=0.317 $Y=0.884
+ $X2=0.317 $Y2=0.925
r27 16 17 9.36182 $w=4.03e-07 $l=3.29e-07 $layer=LI1_cond $X=0.317 $Y=0.555
+ $X2=0.317 $Y2=0.884
r28 16 23 1.13822 $w=4.03e-07 $l=4e-08 $layer=LI1_cond $X=0.317 $Y=0.555
+ $X2=0.317 $Y2=0.515
r29 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.2 $Y=1.82 $X2=0.2
+ $Y2=1.13
r30 11 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=1.82
r31 11 13 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r32 2 13 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r33 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r34 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.37 $X2=0.355 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%VPWR 1 2 11 15 17 19 29 30 33 36
r42 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 27 36 14.9939 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.285 $Y2=3.33
r47 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 26 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 20 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.06 $Y=3.33 $X2=0.87
+ $Y2=3.33
r54 20 22 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 19 36 14.9939 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.285 $Y2=3.33
r56 19 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 13 36 3.22441 $w=8.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=3.245
+ $X2=3.285 $Y2=3.33
r60 13 15 12.2456 $w=8.38e-07 $l=8.6e-07 $layer=LI1_cond $X=3.285 $Y=3.245
+ $X2=3.285 $Y2=2.385
r61 9 33 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245 $X2=0.87
+ $Y2=3.33
r62 9 11 25.1718 $w=3.78e-07 $l=8.3e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.415
r63 2 15 150 $w=1.7e-07 $l=8.30753e-07 $layer=licon1_PDIFF $count=4 $X=2.895
+ $Y=1.96 $X2=3.54 $Y2=2.385
r64 1 11 300 $w=1.7e-07 $l=6.99107e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.87 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%VGND 1 2 11 17 20 21 22 32 33 36
c44 11 0 9.50927e-20 $X=0.855 $Y=0.515
r45 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r47 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r48 27 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r49 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.855
+ $Y2=0
r51 24 26 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.68
+ $Y2=0
r52 22 33 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r53 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r54 22 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r55 20 26 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.68
+ $Y2=0
r56 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.865
+ $Y2=0
r57 19 29 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.16
+ $Y2=0
r58 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.865
+ $Y2=0
r59 15 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.865 $Y=0.085
+ $X2=1.865 $Y2=0
r60 15 17 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=1.865 $Y=0.085
+ $X2=1.865 $Y2=0.735
r61 11 13 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.855 $Y=0.515
+ $X2=0.855 $Y2=0.965
r62 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.085
+ $X2=0.855 $Y2=0
r63 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.855 $Y=0.085
+ $X2=0.855 $Y2=0.515
r64 2 17 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.47 $X2=1.865 $Y2=0.735
r65 1 13 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.37 $X2=0.855 $Y2=0.965
r66 1 11 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.37 $X2=0.855 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%A_245_94# 1 2 9 11 12 15
c36 11 0 2.11106e-19 $X=2.77 $Y=1.195
r37 13 15 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.935 $Y=1.11
+ $X2=2.935 $Y2=0.81
r38 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.77 $Y=1.195
+ $X2=2.935 $Y2=1.11
r39 11 12 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=2.77 $Y=1.195
+ $X2=1.53 $Y2=1.195
r40 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.365 $Y=1.11
+ $X2=1.53 $Y2=1.195
r41 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.365 $Y=1.11
+ $X2=1.365 $Y2=0.615
r42 2 15 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.37 $X2=2.935 $Y2=0.81
r43 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.225
+ $Y=0.47 $X2=1.365 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_1%A_456_74# 1 2 9 11 12 15
r22 13 15 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.435 $Y=0.425
+ $X2=3.435 $Y2=0.525
r23 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.27 $Y=0.34
+ $X2=3.435 $Y2=0.425
r24 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=0.34
+ $X2=2.59 $Y2=0.34
r25 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.425 $Y=0.425
+ $X2=2.59 $Y2=0.34
r26 7 9 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.425 $Y=0.425 $X2=2.425
+ $Y2=0.515
r27 2 15 91 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=2 $X=3.225
+ $Y=0.37 $X2=3.435 $Y2=0.525
r28 1 9 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=2.28
+ $Y=0.37 $X2=2.505 $Y2=0.515
.ends


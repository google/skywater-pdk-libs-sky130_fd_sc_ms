* File: sky130_fd_sc_ms__a31o_2.spice
* Created: Fri Aug 28 17:06:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a31o_2.pex.spice"
.subckt sky130_fd_sc_ms__a31o_2  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_97_296#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_97_296#_M1008_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.23495 AS=0.1036 PD=1.375 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1001 A_371_74# N_A3_M1001_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.23495 PD=0.98 PS=1.375 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1006 A_449_74# N_A2_M1006_g A_371_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75001.9
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1011 N_A_97_296#_M1011_d N_A1_M1011_g A_449_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1554 PD=1.16 PS=1.16 NRD=9.72 NRS=25.128 M=1 R=4.93333
+ SA=75002.5 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_97_296#_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75003
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1002_d N_A_97_296#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1003 N_X_M1002_d N_A_97_296#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.306943 PD=1.39 PS=1.7434 NRD=0 NRS=14.6568 M=1 R=6.22222
+ SA=90000.6 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1004 N_A_365_368#_M1004_d N_A3_M1004_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.274057 PD=1.27 PS=1.5566 NRD=0 NRS=33.1551 M=1 R=5.55556
+ SA=90001.3 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_365_368#_M1004_d VPB PSHORT L=0.18 W=1
+ AD=0.23 AS=0.135 PD=1.46 PS=1.27 NRD=19.7 NRS=0 M=1 R=5.55556 SA=90001.8
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1009 N_A_365_368#_M1009_d N_A1_M1009_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.23 PD=1.32 PS=1.46 NRD=0 NRS=15.7403 M=1 R=5.55556 SA=90002.4
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_97_296#_M1010_d N_B1_M1010_g N_A_365_368#_M1009_d VPB PSHORT L=0.18
+ W=1 AD=0.29 AS=0.16 PD=2.58 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__a31o_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__maj3_1.spice
* Created: Wed Sep  2 12:11:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__maj3_1.pex.spice"
.subckt sky130_fd_sc_ms__maj3_1  VNB VPB B C A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_84_74#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.148965 AS=0.2081 PD=1.21725 PS=2.05 NRD=14.592 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1011 A_223_120# N_A_M1011_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.128835 PD=0.88 PS=1.05275 NRD=12.18 NRS=4.68 M=1 R=4.26667 SA=75000.8
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_84_74#_M1004_d N_B_M1004_g A_223_120# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1222 AS=0.0768 PD=1.08 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.1
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 A_403_136# N_B_M1013_g N_A_84_74#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1222 PD=0.88 PS=1.08 NRD=12.18 NRS=15.468 M=1 R=4.26667
+ SA=75001.5 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g A_403_136# VNB NLOWVT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=13.116 NRS=12.18 M=1 R=4.26667 SA=75001.9
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 A_595_136# N_A_M1005_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64 AD=0.0864
+ AS=0.1344 PD=0.91 PS=1.06 NRD=15 NRS=13.116 M=1 R=4.26667 SA=75002.4
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_84_74#_M1008_d N_C_M1008_g A_595_136# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1733 AS=0.0864 PD=1.85 PS=0.91 NRD=0 NRS=15 M=1 R=4.26667 SA=75002.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_84_74#_M1001_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.187547 AS=0.3136 PD=1.52679 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1006 A_229_384# N_A_M1006_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.167453 PD=1.24 PS=1.36321 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1010 N_A_84_74#_M1010_d N_B_M1010_g A_229_384# VPB PSHORT L=0.18 W=1 AD=0.15
+ AS=0.12 PD=1.3 PS=1.24 NRD=4.9053 NRS=12.7853 M=1 R=5.55556 SA=90001.1
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1009 A_409_384# N_B_M1009_g N_A_84_74#_M1010_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.15 PD=1.24 PS=1.3 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90001.6 SB=90001.6
+ A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_C_M1012_g A_409_384# VPB PSHORT L=0.18 W=1 AD=0.18
+ AS=0.12 PD=1.36 PS=1.24 NRD=6.8753 NRS=12.7853 M=1 R=5.55556 SA=90002
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 A_601_384# N_A_M1000_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.18 PD=1.24 PS=1.36 NRD=12.7853 NRS=8.8453 M=1 R=5.55556 SA=90002.6
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_84_74#_M1003_d N_C_M1003_g A_601_384# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90003 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__maj3_1.pxi.spice"
*
.ends
*
*

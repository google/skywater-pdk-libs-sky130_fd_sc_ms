* File: sky130_fd_sc_ms__o21ba_1.pxi.spice
* Created: Wed Sep  2 12:22:10 2020
* 
x_PM_SKY130_FD_SC_MS__O21BA_1%A1 N_A1_c_75_n N_A1_c_80_n N_A1_M1002_g
+ N_A1_M1008_g A1 A1 N_A1_c_77_n N_A1_c_78_n PM_SKY130_FD_SC_MS__O21BA_1%A1
x_PM_SKY130_FD_SC_MS__O21BA_1%A2 N_A2_M1003_g N_A2_M1009_g N_A2_c_104_n
+ N_A2_c_105_n N_A2_c_106_n A2 A2 N_A2_c_108_n PM_SKY130_FD_SC_MS__O21BA_1%A2
x_PM_SKY130_FD_SC_MS__O21BA_1%A_281_244# N_A_281_244#_M1006_s
+ N_A_281_244#_M1007_s N_A_281_244#_M1004_g N_A_281_244#_M1005_g
+ N_A_281_244#_c_145_n N_A_281_244#_c_146_n N_A_281_244#_c_147_n
+ N_A_281_244#_c_148_n N_A_281_244#_c_154_n N_A_281_244#_c_155_n
+ N_A_281_244#_c_149_n N_A_281_244#_c_150_n N_A_281_244#_c_151_n
+ PM_SKY130_FD_SC_MS__O21BA_1%A_281_244#
x_PM_SKY130_FD_SC_MS__O21BA_1%B1_N N_B1_N_M1007_g N_B1_N_M1006_g B1_N
+ N_B1_N_c_203_n N_B1_N_c_204_n PM_SKY130_FD_SC_MS__O21BA_1%B1_N
x_PM_SKY130_FD_SC_MS__O21BA_1%A_203_392# N_A_203_392#_M1005_d
+ N_A_203_392#_M1003_d N_A_203_392#_M1000_g N_A_203_392#_M1001_g
+ N_A_203_392#_c_239_n N_A_203_392#_c_240_n N_A_203_392#_c_247_n
+ N_A_203_392#_c_241_n N_A_203_392#_c_249_n N_A_203_392#_c_253_n
+ N_A_203_392#_c_242_n N_A_203_392#_c_243_n N_A_203_392#_c_244_n
+ PM_SKY130_FD_SC_MS__O21BA_1%A_203_392#
x_PM_SKY130_FD_SC_MS__O21BA_1%VPWR N_VPWR_M1002_s N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n VPWR
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_319_n N_VPWR_c_328_n
+ N_VPWR_c_329_n PM_SKY130_FD_SC_MS__O21BA_1%VPWR
x_PM_SKY130_FD_SC_MS__O21BA_1%X N_X_M1001_d N_X_M1000_d N_X_c_364_n N_X_c_365_n
+ X X X X N_X_c_366_n PM_SKY130_FD_SC_MS__O21BA_1%X
x_PM_SKY130_FD_SC_MS__O21BA_1%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1009_d
+ N_A_27_74#_c_390_n N_A_27_74#_c_394_n N_A_27_74#_c_391_n N_A_27_74#_c_392_n
+ PM_SKY130_FD_SC_MS__O21BA_1%A_27_74#
x_PM_SKY130_FD_SC_MS__O21BA_1%VGND N_VGND_M1008_d N_VGND_M1006_d N_VGND_c_417_n
+ N_VGND_c_418_n VGND N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n PM_SKY130_FD_SC_MS__O21BA_1%VGND
cc_1 VNB N_A1_c_75_n 0.0298684f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.625
cc_2 VNB A1 0.0231282f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A1_c_77_n 0.020516f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_4 VNB N_A1_c_78_n 0.0261918f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.13
cc_5 VNB N_A2_c_104_n 0.019683f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A2_c_105_n 0.022135f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A2_c_106_n 0.0016372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A2 0.00689173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_c_108_n 0.0160326f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_10 VNB N_A_281_244#_M1004_g 0.00864087f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_281_244#_M1005_g 0.0268815f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_12 VNB N_A_281_244#_c_145_n 0.0116334f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_13 VNB N_A_281_244#_c_146_n 0.00211765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_281_244#_c_147_n 0.00647567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_281_244#_c_148_n 0.0367177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_281_244#_c_149_n 0.00327435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_281_244#_c_150_n 0.00421238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_281_244#_c_151_n 0.0388575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_N_M1007_g 0.00686837f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.89
cc_20 VNB B1_N 0.00365732f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_21 VNB N_B1_N_c_203_n 0.0328137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_N_c_204_n 0.0229476f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_23 VNB N_A_203_392#_M1000_g 5.81932e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_A_203_392#_M1001_g 0.0299727f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_25 VNB N_A_203_392#_c_239_n 0.0176071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_203_392#_c_240_n 0.00623122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_203_392#_c_241_n 2.56499e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_203_392#_c_242_n 0.00393771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_203_392#_c_243_n 0.00302585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_203_392#_c_244_n 0.0349911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_319_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_364_n 0.0267037f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_X_c_365_n 0.01394f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_34 VNB N_X_c_366_n 0.0249686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_390_n 0.0193497f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_A_27_74#_c_391_n 0.00752814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_392_n 0.00252555f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_38 VNB N_VGND_c_417_n 0.00970653f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_39 VNB N_VGND_c_418_n 0.0172154f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_40 VNB N_VGND_c_419_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_41 VNB N_VGND_c_420_n 0.0543292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_421_n 0.0190372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_422_n 0.24119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_423_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_424_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A1_c_75_n 0.0264224f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.625
cc_47 VPB N_A1_c_80_n 0.0202235f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.89
cc_48 VPB A1 0.00808948f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_49 VPB N_A2_M1003_g 0.0233718f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.89
cc_50 VPB N_A2_c_106_n 0.0134208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB A2 0.00506394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_281_244#_M1004_g 0.0334424f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_53 VPB N_A_281_244#_c_146_n 0.00414068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_281_244#_c_154_n 0.00944815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_281_244#_c_155_n 0.00902131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_B1_N_M1007_g 0.0296654f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.89
cc_57 VPB N_A_203_392#_M1000_g 0.0302143f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_58 VPB N_A_203_392#_c_240_n 0.00601893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_203_392#_c_247_n 0.0169246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_203_392#_c_241_n 0.00319328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_203_392#_c_249_n 0.00331921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_320_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_63 VPB N_VPWR_c_321_n 0.0480138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_322_n 0.0215074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_323_n 0.020334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_324_n 0.0323805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_325_n 0.0320766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_326_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_319_n 0.0757841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_328_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_329_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB X 0.0136968f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.295
cc_73 VPB X 0.0415472f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_366_n 0.00750262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 N_A1_c_75_n N_A2_M1003_g 0.067779f $X=0.395 $Y=1.625 $X2=0 $Y2=0
cc_76 N_A1_c_78_n N_A2_c_104_n 0.0218539f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_77 N_A1_c_75_n N_A2_c_105_n 0.0154493f $X=0.395 $Y=1.625 $X2=0 $Y2=0
cc_78 A1 A2 0.0348017f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_77_n A2 0.00260358f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_80 A1 N_A2_c_108_n 0.00246986f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A1_c_77_n N_A2_c_108_n 0.0154493f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_82 N_A1_c_75_n N_VPWR_c_321_n 0.0013539f $X=0.395 $Y=1.625 $X2=0 $Y2=0
cc_83 N_A1_c_80_n N_VPWR_c_321_n 0.0254086f $X=0.505 $Y=1.89 $X2=0 $Y2=0
cc_84 A1 N_VPWR_c_321_n 0.0255131f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A1_c_80_n N_VPWR_c_324_n 0.00460063f $X=0.505 $Y=1.89 $X2=0 $Y2=0
cc_86 N_A1_c_80_n N_VPWR_c_319_n 0.00908371f $X=0.505 $Y=1.89 $X2=0 $Y2=0
cc_87 N_A1_c_78_n N_A_27_74#_c_390_n 0.00684796f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_88 A1 N_A_27_74#_c_394_n 0.00787831f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A1_c_78_n N_A_27_74#_c_394_n 0.00967287f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_90 A1 N_A_27_74#_c_391_n 0.0254243f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A1_c_77_n N_A_27_74#_c_391_n 0.00137692f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_92 N_A1_c_78_n N_A_27_74#_c_391_n 7.15033e-19 $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_93 N_A1_c_78_n N_A_27_74#_c_392_n 5.85113e-19 $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_94 N_A1_c_78_n N_VGND_c_417_n 0.00488987f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_95 N_A1_c_78_n N_VGND_c_419_n 0.00434272f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_96 N_A1_c_78_n N_VGND_c_422_n 0.00439339f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_97 N_A2_M1003_g N_A_281_244#_M1004_g 0.0205576f $X=0.925 $Y=2.46 $X2=0 $Y2=0
cc_98 N_A2_c_105_n N_A_281_244#_M1004_g 0.0152062f $X=1 $Y=1.635 $X2=0 $Y2=0
cc_99 N_A2_c_104_n N_A_281_244#_M1005_g 0.0109162f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_100 A2 N_A_281_244#_M1005_g 7.79834e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A2_c_108_n N_A_281_244#_M1005_g 0.00380119f $X=1 $Y=1.295 $X2=0 $Y2=0
cc_102 A2 N_A_281_244#_c_145_n 0.00560722f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A2_c_108_n N_A_281_244#_c_145_n 0.0152062f $X=1 $Y=1.295 $X2=0 $Y2=0
cc_104 A2 N_A_203_392#_c_240_n 0.0357245f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A2_c_108_n N_A_203_392#_c_240_n 2.2434e-19 $X=1 $Y=1.295 $X2=0 $Y2=0
cc_106 N_A2_M1003_g N_A_203_392#_c_249_n 0.00313467f $X=0.925 $Y=2.46 $X2=0
+ $Y2=0
cc_107 N_A2_c_106_n N_A_203_392#_c_253_n 7.87638e-19 $X=1 $Y=1.8 $X2=0 $Y2=0
cc_108 A2 N_A_203_392#_c_253_n 0.0219906f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A2_M1003_g N_VPWR_c_321_n 0.00349819f $X=0.925 $Y=2.46 $X2=0 $Y2=0
cc_110 N_A2_M1003_g N_VPWR_c_322_n 5.73176e-19 $X=0.925 $Y=2.46 $X2=0 $Y2=0
cc_111 N_A2_M1003_g N_VPWR_c_324_n 0.00553757f $X=0.925 $Y=2.46 $X2=0 $Y2=0
cc_112 N_A2_M1003_g N_VPWR_c_319_n 0.0109071f $X=0.925 $Y=2.46 $X2=0 $Y2=0
cc_113 N_A2_c_104_n N_A_27_74#_c_390_n 5.85113e-19 $X=1 $Y=1.13 $X2=0 $Y2=0
cc_114 N_A2_c_104_n N_A_27_74#_c_394_n 0.00974567f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_115 A2 N_A_27_74#_c_394_n 0.0347531f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A2_c_108_n N_A_27_74#_c_394_n 9.46749e-19 $X=1 $Y=1.295 $X2=0 $Y2=0
cc_117 N_A2_c_104_n N_A_27_74#_c_392_n 0.00669591f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_118 N_A2_c_104_n N_VGND_c_417_n 0.00488987f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_119 N_A2_c_104_n N_VGND_c_420_n 0.00434272f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_120 N_A2_c_104_n N_VGND_c_422_n 0.00435917f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_121 N_A_281_244#_c_146_n N_B1_N_M1007_g 0.00835568f $X=2.14 $Y=1.82 $X2=0
+ $Y2=0
cc_122 N_A_281_244#_c_155_n N_B1_N_M1007_g 0.00661147f $X=2.52 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_281_244#_c_148_n B1_N 0.00131019f $X=2.14 $Y=1.385 $X2=0 $Y2=0
cc_124 N_A_281_244#_c_155_n B1_N 0.00974338f $X=2.52 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_281_244#_c_149_n B1_N 0.0235839f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_126 N_A_281_244#_c_150_n B1_N 0.0143996f $X=2.555 $Y=0.845 $X2=0 $Y2=0
cc_127 N_A_281_244#_c_147_n N_B1_N_c_203_n 0.00114872f $X=2.14 $Y=1.385 $X2=0
+ $Y2=0
cc_128 N_A_281_244#_c_148_n N_B1_N_c_203_n 0.0212168f $X=2.14 $Y=1.385 $X2=0
+ $Y2=0
cc_129 N_A_281_244#_c_155_n N_B1_N_c_203_n 9.86294e-19 $X=2.52 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_281_244#_c_150_n N_B1_N_c_203_n 0.00105115f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_131 N_A_281_244#_c_149_n N_B1_N_c_204_n 0.00438837f $X=2.14 $Y=1.22 $X2=0
+ $Y2=0
cc_132 N_A_281_244#_c_150_n N_B1_N_c_204_n 0.00422447f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_133 N_A_281_244#_M1005_g N_A_203_392#_c_239_n 0.00745905f $X=1.51 $Y=0.69
+ $X2=0 $Y2=0
cc_134 N_A_281_244#_c_150_n N_A_203_392#_c_239_n 0.0264642f $X=2.555 $Y=0.845
+ $X2=0 $Y2=0
cc_135 N_A_281_244#_M1004_g N_A_203_392#_c_240_n 0.0134829f $X=1.495 $Y=2.46
+ $X2=0 $Y2=0
cc_136 N_A_281_244#_c_147_n N_A_203_392#_c_240_n 0.0414317f $X=2.14 $Y=1.385
+ $X2=0 $Y2=0
cc_137 N_A_281_244#_c_148_n N_A_203_392#_c_240_n 2.99159e-19 $X=2.14 $Y=1.385
+ $X2=0 $Y2=0
cc_138 N_A_281_244#_c_154_n N_A_203_392#_c_240_n 0.0117446f $X=2.305 $Y=1.985
+ $X2=0 $Y2=0
cc_139 N_A_281_244#_c_149_n N_A_203_392#_c_240_n 0.00863714f $X=2.14 $Y=1.22
+ $X2=0 $Y2=0
cc_140 N_A_281_244#_c_151_n N_A_203_392#_c_240_n 0.0203485f $X=1.975 $Y=1.385
+ $X2=0 $Y2=0
cc_141 N_A_281_244#_M1007_s N_A_203_392#_c_247_n 0.0107941f $X=2.305 $Y=1.84
+ $X2=0 $Y2=0
cc_142 N_A_281_244#_c_154_n N_A_203_392#_c_247_n 0.0277408f $X=2.305 $Y=1.985
+ $X2=0 $Y2=0
cc_143 N_A_281_244#_c_155_n N_A_203_392#_c_247_n 0.0248385f $X=2.52 $Y=1.985
+ $X2=0 $Y2=0
cc_144 N_A_281_244#_c_155_n N_A_203_392#_c_241_n 0.0143474f $X=2.52 $Y=1.985
+ $X2=0 $Y2=0
cc_145 N_A_281_244#_M1004_g N_A_203_392#_c_253_n 0.0325821f $X=1.495 $Y=2.46
+ $X2=0 $Y2=0
cc_146 N_A_281_244#_c_154_n N_A_203_392#_c_253_n 0.0152281f $X=2.305 $Y=1.985
+ $X2=0 $Y2=0
cc_147 N_A_281_244#_c_151_n N_A_203_392#_c_253_n 4.1398e-19 $X=1.975 $Y=1.385
+ $X2=0 $Y2=0
cc_148 N_A_281_244#_c_149_n N_A_203_392#_c_242_n 0.00146638f $X=2.14 $Y=1.22
+ $X2=0 $Y2=0
cc_149 N_A_281_244#_c_151_n N_A_203_392#_c_242_n 0.00677504f $X=1.975 $Y=1.385
+ $X2=0 $Y2=0
cc_150 N_A_281_244#_M1004_g N_VPWR_c_322_n 0.00955167f $X=1.495 $Y=2.46 $X2=0
+ $Y2=0
cc_151 N_A_281_244#_M1004_g N_VPWR_c_324_n 0.00460063f $X=1.495 $Y=2.46 $X2=0
+ $Y2=0
cc_152 N_A_281_244#_M1004_g N_VPWR_c_319_n 0.00461999f $X=1.495 $Y=2.46 $X2=0
+ $Y2=0
cc_153 N_A_281_244#_M1005_g N_A_27_74#_c_394_n 0.00205241f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_154 N_A_281_244#_M1005_g N_A_27_74#_c_392_n 0.00454372f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_155 N_A_281_244#_M1005_g N_VGND_c_420_n 0.00451267f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_156 N_A_281_244#_c_150_n N_VGND_c_420_n 0.00927306f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_157 N_A_281_244#_M1005_g N_VGND_c_422_n 0.00881535f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_158 N_A_281_244#_c_150_n N_VGND_c_422_n 0.0165534f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_159 N_B1_N_M1007_g N_A_203_392#_M1000_g 0.0239852f $X=2.75 $Y=2.26 $X2=0
+ $Y2=0
cc_160 B1_N N_A_203_392#_M1001_g 7.87159e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B1_N_c_204_n N_A_203_392#_M1001_g 0.0181853f $X=2.68 $Y=1.22 $X2=0
+ $Y2=0
cc_162 N_B1_N_M1007_g N_A_203_392#_c_247_n 0.020286f $X=2.75 $Y=2.26 $X2=0 $Y2=0
cc_163 N_B1_N_M1007_g N_A_203_392#_c_241_n 0.00989557f $X=2.75 $Y=2.26 $X2=0
+ $Y2=0
cc_164 N_B1_N_M1007_g N_A_203_392#_c_243_n 0.00222581f $X=2.75 $Y=2.26 $X2=0
+ $Y2=0
cc_165 B1_N N_A_203_392#_c_243_n 0.0156452f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B1_N_c_203_n N_A_203_392#_c_243_n 0.00140768f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_167 N_B1_N_M1007_g N_A_203_392#_c_244_n 0.00494446f $X=2.75 $Y=2.26 $X2=0
+ $Y2=0
cc_168 B1_N N_A_203_392#_c_244_n 2.75885e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B1_N_c_203_n N_A_203_392#_c_244_n 0.0122189f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_170 N_B1_N_M1007_g N_VPWR_c_323_n 0.00385696f $X=2.75 $Y=2.26 $X2=0 $Y2=0
cc_171 N_B1_N_M1007_g N_VPWR_c_325_n 0.00482866f $X=2.75 $Y=2.26 $X2=0 $Y2=0
cc_172 N_B1_N_M1007_g N_VPWR_c_319_n 0.00555093f $X=2.75 $Y=2.26 $X2=0 $Y2=0
cc_173 N_B1_N_c_204_n N_X_c_364_n 6.61818e-19 $X=2.68 $Y=1.22 $X2=0 $Y2=0
cc_174 N_B1_N_M1007_g X 9.03352e-19 $X=2.75 $Y=2.26 $X2=0 $Y2=0
cc_175 N_B1_N_c_204_n N_VGND_c_418_n 0.00650911f $X=2.68 $Y=1.22 $X2=0 $Y2=0
cc_176 N_B1_N_c_204_n N_VGND_c_420_n 0.00434489f $X=2.68 $Y=1.22 $X2=0 $Y2=0
cc_177 N_B1_N_c_204_n N_VGND_c_422_n 0.00487769f $X=2.68 $Y=1.22 $X2=0 $Y2=0
cc_178 N_A_203_392#_c_240_n N_VPWR_M1004_d 5.31322e-19 $X=1.7 $Y=1.97 $X2=0
+ $Y2=0
cc_179 N_A_203_392#_c_247_n N_VPWR_M1004_d 0.0045773f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_180 N_A_203_392#_c_253_n N_VPWR_M1004_d 0.0122394f $X=1.785 $Y=2.23 $X2=0
+ $Y2=0
cc_181 N_A_203_392#_c_247_n N_VPWR_M1007_d 0.0106453f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_182 N_A_203_392#_c_241_n N_VPWR_M1007_d 0.00914173f $X=3.14 $Y=2.32 $X2=0
+ $Y2=0
cc_183 N_A_203_392#_c_249_n N_VPWR_c_321_n 0.0066941f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_184 N_A_203_392#_c_249_n N_VPWR_c_322_n 0.0127976f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_185 N_A_203_392#_c_253_n N_VPWR_c_322_n 0.0224354f $X=1.785 $Y=2.23 $X2=0
+ $Y2=0
cc_186 N_A_203_392#_M1000_g N_VPWR_c_323_n 0.00534567f $X=3.335 $Y=2.4 $X2=0
+ $Y2=0
cc_187 N_A_203_392#_c_247_n N_VPWR_c_323_n 0.024198f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_188 N_A_203_392#_c_249_n N_VPWR_c_324_n 0.0142934f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_189 N_A_203_392#_M1000_g N_VPWR_c_326_n 0.005209f $X=3.335 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_203_392#_M1000_g N_VPWR_c_319_n 0.00990469f $X=3.335 $Y=2.4 $X2=0
+ $Y2=0
cc_191 N_A_203_392#_c_247_n N_VPWR_c_319_n 0.0354692f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_192 N_A_203_392#_c_249_n N_VPWR_c_319_n 0.0119825f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_193 N_A_203_392#_c_253_n N_VPWR_c_319_n 0.00657271f $X=1.785 $Y=2.23 $X2=0
+ $Y2=0
cc_194 N_A_203_392#_M1001_g N_X_c_364_n 0.00806387f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_203_392#_M1001_g N_X_c_365_n 0.00386394f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_203_392#_c_243_n N_X_c_365_n 0.00175157f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_197 N_A_203_392#_c_244_n N_X_c_365_n 4.73526e-19 $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_198 N_A_203_392#_M1000_g X 0.00320667f $X=3.335 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_203_392#_c_241_n X 0.0196895f $X=3.14 $Y=2.32 $X2=0 $Y2=0
cc_200 N_A_203_392#_c_243_n X 0.00151667f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_201 N_A_203_392#_M1000_g X 0.0145882f $X=3.335 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_203_392#_M1001_g N_X_c_366_n 0.00477624f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_203_392#_c_241_n N_X_c_366_n 0.00535845f $X=3.14 $Y=2.32 $X2=0 $Y2=0
cc_204 N_A_203_392#_c_243_n N_X_c_366_n 0.0249376f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_205 N_A_203_392#_c_244_n N_X_c_366_n 0.0102032f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_206 N_A_203_392#_c_239_n N_A_27_74#_c_392_n 0.0172628f $X=1.78 $Y=0.515 $X2=0
+ $Y2=0
cc_207 N_A_203_392#_M1001_g N_VGND_c_418_n 0.00703428f $X=3.34 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_203_392#_c_243_n N_VGND_c_418_n 0.00834888f $X=3.25 $Y=1.485 $X2=0
+ $Y2=0
cc_209 N_A_203_392#_c_244_n N_VGND_c_418_n 0.00283306f $X=3.25 $Y=1.485 $X2=0
+ $Y2=0
cc_210 N_A_203_392#_c_239_n N_VGND_c_420_n 0.0146357f $X=1.78 $Y=0.515 $X2=0
+ $Y2=0
cc_211 N_A_203_392#_M1001_g N_VGND_c_421_n 0.00434272f $X=3.34 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_203_392#_M1001_g N_VGND_c_422_n 0.00828734f $X=3.34 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_203_392#_c_239_n N_VGND_c_422_n 0.0121141f $X=1.78 $Y=0.515 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_323_n X 0.0129586f $X=3.06 $Y=2.78 $X2=0 $Y2=0
cc_215 N_VPWR_c_326_n X 0.0158876f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_319_n X 0.0130823f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_217 N_X_c_364_n N_VGND_c_418_n 0.0259022f $X=3.555 $Y=0.515 $X2=0 $Y2=0
cc_218 N_X_c_364_n N_VGND_c_421_n 0.0161257f $X=3.555 $Y=0.515 $X2=0 $Y2=0
cc_219 N_X_c_364_n N_VGND_c_422_n 0.013291f $X=3.555 $Y=0.515 $X2=0 $Y2=0
cc_220 N_A_27_74#_c_394_n N_VGND_M1008_d 0.0125077f $X=1.115 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_221 N_A_27_74#_c_390_n N_VGND_c_417_n 0.0109215f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_222 N_A_27_74#_c_394_n N_VGND_c_417_n 0.0243105f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_223 N_A_27_74#_c_392_n N_VGND_c_417_n 0.0109215f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_390_n N_VGND_c_419_n 0.0144497f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_392_n N_VGND_c_420_n 0.0144232f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_226 N_A_27_74#_c_390_n N_VGND_c_422_n 0.0119539f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_227 N_A_27_74#_c_394_n N_VGND_c_422_n 0.0116461f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_228 N_A_27_74#_c_392_n N_VGND_c_422_n 0.0119105f $X=1.28 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__or2_1.spice
* Created: Wed Sep  2 12:27:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or2_1.pex.spice"
.subckt sky130_fd_sc_ms__or2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_A_63_368#_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.130625 AS=0.2695 PD=1.025 PS=2.08 NRD=34.908 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_63_368#_M1003_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.130625 PD=0.997674 PS=1.025 NRD=17.448 NRS=7.632 M=1
+ R=3.66667 SA=75001 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1000 N_X_M1000_d N_A_63_368#_M1000_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_155_368# N_B_M1001_g N_A_63_368#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1008 AS=0.2352 PD=1.08 PS=2.24 NRD=15.2281 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_155_368# VPB PSHORT L=0.18 W=0.84 AD=0.2742
+ AS=0.1008 PD=1.48286 PS=1.08 NRD=63.6507 NRS=15.2281 M=1 R=4.66667 SA=90000.6
+ SB=90001 A=0.1512 P=2.04 MULT=1
MM1004 N_X_M1004_d N_A_63_368#_M1004_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3656 PD=2.8 PS=1.97714 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__or2_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a21bo_2.pxi.spice
* Created: Fri Aug 28 16:58:00 2020
* 
x_PM_SKY130_FD_SC_MS__A21BO_2%B1_N N_B1_N_M1001_g N_B1_N_c_74_n N_B1_N_M1010_g
+ B1_N N_B1_N_c_75_n N_B1_N_c_76_n PM_SKY130_FD_SC_MS__A21BO_2%B1_N
x_PM_SKY130_FD_SC_MS__A21BO_2%A_187_244# N_A_187_244#_M1003_d
+ N_A_187_244#_M1006_s N_A_187_244#_M1002_g N_A_187_244#_c_104_n
+ N_A_187_244#_M1000_g N_A_187_244#_M1004_g N_A_187_244#_c_106_n
+ N_A_187_244#_M1005_g N_A_187_244#_c_119_p N_A_187_244#_c_107_n
+ N_A_187_244#_c_108_n N_A_187_244#_c_109_n N_A_187_244#_c_110_n
+ N_A_187_244#_c_114_n N_A_187_244#_c_123_p
+ PM_SKY130_FD_SC_MS__A21BO_2%A_187_244#
x_PM_SKY130_FD_SC_MS__A21BO_2%A_32_368# N_A_32_368#_M1010_s N_A_32_368#_M1001_s
+ N_A_32_368#_M1003_g N_A_32_368#_c_207_n N_A_32_368#_M1006_g
+ N_A_32_368#_c_201_n N_A_32_368#_c_202_n N_A_32_368#_c_203_n
+ N_A_32_368#_c_210_n N_A_32_368#_c_217_n N_A_32_368#_c_211_n
+ N_A_32_368#_c_204_n N_A_32_368#_c_246_n N_A_32_368#_c_205_n
+ N_A_32_368#_c_255_n N_A_32_368#_c_206_n N_A_32_368#_c_266_p
+ PM_SKY130_FD_SC_MS__A21BO_2%A_32_368#
x_PM_SKY130_FD_SC_MS__A21BO_2%A1 N_A1_M1011_g N_A1_M1007_g A1 N_A1_c_300_n
+ N_A1_c_301_n PM_SKY130_FD_SC_MS__A21BO_2%A1
x_PM_SKY130_FD_SC_MS__A21BO_2%A2 N_A2_M1009_g N_A2_M1008_g A2 N_A2_c_340_n
+ PM_SKY130_FD_SC_MS__A21BO_2%A2
x_PM_SKY130_FD_SC_MS__A21BO_2%VPWR N_VPWR_M1001_d N_VPWR_M1004_s N_VPWR_M1007_d
+ N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n VPWR N_VPWR_c_368_n
+ N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_364_n N_VPWR_c_373_n
+ N_VPWR_c_374_n N_VPWR_c_375_n PM_SKY130_FD_SC_MS__A21BO_2%VPWR
x_PM_SKY130_FD_SC_MS__A21BO_2%X N_X_M1000_s N_X_M1002_d N_X_c_422_n N_X_c_423_n
+ N_X_c_425_n X PM_SKY130_FD_SC_MS__A21BO_2%X
x_PM_SKY130_FD_SC_MS__A21BO_2%A_507_392# N_A_507_392#_M1006_d
+ N_A_507_392#_M1008_d N_A_507_392#_c_462_n N_A_507_392#_c_457_n
+ N_A_507_392#_c_458_n N_A_507_392#_c_459_n
+ PM_SKY130_FD_SC_MS__A21BO_2%A_507_392#
x_PM_SKY130_FD_SC_MS__A21BO_2%VGND N_VGND_M1010_d N_VGND_M1005_d N_VGND_M1009_d
+ N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n
+ N_VGND_c_487_n VGND N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n
+ N_VGND_c_491_n PM_SKY130_FD_SC_MS__A21BO_2%VGND
cc_1 VNB N_B1_N_M1001_g 0.00958212f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.26
cc_2 VNB N_B1_N_c_74_n 0.0228559f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.22
cc_3 VNB N_B1_N_c_75_n 0.0225328f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_4 VNB N_B1_N_c_76_n 0.0534441f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.385
cc_5 VNB N_A_187_244#_M1002_g 0.0142239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_187_244#_c_104_n 0.0176121f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_7 VNB N_A_187_244#_M1004_g 0.00653034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_187_244#_c_106_n 0.019167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_187_244#_c_107_n 0.00881618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_187_244#_c_108_n 0.00390742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_187_244#_c_109_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_187_244#_c_110_n 0.0469464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_32_368#_M1003_g 0.0221011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_32_368#_c_201_n 0.0465265f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_15 VNB N_A_32_368#_c_202_n 0.00860503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_32_368#_c_203_n 0.00372942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_32_368#_c_204_n 0.00426191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_32_368#_c_205_n 0.00620465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_32_368#_c_206_n 0.0225067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_M1011_g 0.0204236f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.26
cc_21 VNB N_A1_M1007_g 0.00318739f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.835
cc_22 VNB N_A1_c_300_n 0.02979f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_23 VNB N_A1_c_301_n 0.0159715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_M1009_g 0.0408671f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.26
cc_25 VNB A2 0.00472574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_340_n 0.0348817f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.385
cc_27 VNB N_VPWR_c_364_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_422_n 0.00239017f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.835
cc_29 VNB N_X_c_423_n 0.00285947f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_VGND_c_482_n 0.0157102f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_31 VNB N_VGND_c_483_n 0.0124379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_484_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_485_n 0.037498f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.365
cc_34 VNB N_VGND_c_486_n 0.0259864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_487_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_488_n 0.0189193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_489_n 0.0312656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_490_n 0.01106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_491_n 0.243653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_B1_N_M1001_g 0.0320826f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.26
cc_41 VPB N_A_187_244#_M1002_g 0.0237612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_187_244#_M1004_g 0.0247803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_187_244#_c_108_n 6.19153e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_187_244#_c_114_n 0.0178285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_32_368#_c_207_n 0.00617707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_32_368#_M1006_g 0.0233023f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.385
cc_47 VPB N_A_32_368#_c_203_n 0.00372942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_32_368#_c_210_n 0.0187054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_32_368#_c_211_n 0.0224256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_32_368#_c_204_n 0.00325106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_32_368#_c_205_n 0.0177629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A1_M1007_g 0.0281888f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.835
cc_53 VPB N_A1_c_301_n 0.00540584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A2_M1008_g 0.0318997f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.835
cc_55 VPB A2 0.00276779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A2_c_340_n 0.0233136f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.385
cc_57 VPB N_VPWR_c_365_n 0.0164504f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_58 VPB N_VPWR_c_366_n 0.011178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_367_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.365
cc_60 VPB N_VPWR_c_368_n 0.0208665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_369_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_370_n 0.0303553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_371_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_364_n 0.0838259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_373_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_374_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_375_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_423_n 0.00162883f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_69 VPB N_X_c_425_n 0.00254834f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_70 VPB N_A_507_392#_c_457_n 0.0148093f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_71 VPB N_A_507_392#_c_458_n 0.0300702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_507_392#_c_459_n 0.00178465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 N_B1_N_M1001_g N_A_187_244#_M1002_g 0.0345778f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_74 N_B1_N_c_74_n N_A_187_244#_c_104_n 0.0180021f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_75 N_B1_N_c_76_n N_A_187_244#_c_110_n 0.0205347f $X=0.65 $Y=1.385 $X2=0 $Y2=0
cc_76 N_B1_N_M1001_g N_A_32_368#_c_210_n 0.00742872f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_77 N_B1_N_c_75_n N_A_32_368#_c_210_n 0.0196109f $X=0.345 $Y=1.385 $X2=0 $Y2=0
cc_78 N_B1_N_c_76_n N_A_32_368#_c_210_n 0.00528718f $X=0.65 $Y=1.385 $X2=0 $Y2=0
cc_79 N_B1_N_M1001_g N_A_32_368#_c_217_n 0.017322f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_80 N_B1_N_c_76_n N_A_32_368#_c_217_n 0.00135613f $X=0.65 $Y=1.385 $X2=0 $Y2=0
cc_81 N_B1_N_M1001_g N_A_32_368#_c_211_n 0.0081913f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_82 N_B1_N_M1001_g N_A_32_368#_c_204_n 0.00997485f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_83 N_B1_N_c_74_n N_A_32_368#_c_204_n 0.00946285f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_84 N_B1_N_c_75_n N_A_32_368#_c_204_n 0.0268756f $X=0.345 $Y=1.385 $X2=0 $Y2=0
cc_85 N_B1_N_c_76_n N_A_32_368#_c_204_n 0.00861295f $X=0.65 $Y=1.385 $X2=0 $Y2=0
cc_86 N_B1_N_c_74_n N_A_32_368#_c_206_n 0.018243f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_87 N_B1_N_c_75_n N_A_32_368#_c_206_n 0.0204716f $X=0.345 $Y=1.385 $X2=0 $Y2=0
cc_88 N_B1_N_c_76_n N_A_32_368#_c_206_n 0.00331213f $X=0.65 $Y=1.385 $X2=0 $Y2=0
cc_89 N_B1_N_M1001_g N_VPWR_c_365_n 0.00387296f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_90 N_B1_N_M1001_g N_VPWR_c_368_n 0.0046462f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_91 N_B1_N_M1001_g N_VPWR_c_364_n 0.00555093f $X=0.51 $Y=2.26 $X2=0 $Y2=0
cc_92 N_B1_N_c_74_n N_X_c_422_n 0.00117035f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_93 N_B1_N_c_74_n N_X_c_423_n 4.56618e-19 $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_94 N_B1_N_c_76_n N_X_c_423_n 2.83559e-19 $X=0.65 $Y=1.385 $X2=0 $Y2=0
cc_95 N_B1_N_c_74_n N_VGND_c_482_n 0.00400491f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_96 N_B1_N_c_74_n N_VGND_c_486_n 0.00432822f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_97 N_B1_N_c_74_n N_VGND_c_491_n 0.00487769f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_98 N_A_187_244#_c_106_n N_A_32_368#_M1003_g 0.0084396f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_99 N_A_187_244#_c_119_p N_A_32_368#_M1003_g 0.00596357f $X=2.385 $Y=1.005
+ $X2=0 $Y2=0
cc_100 N_A_187_244#_c_107_n N_A_32_368#_M1003_g 0.0010596f $X=1.735 $Y=1.005
+ $X2=0 $Y2=0
cc_101 N_A_187_244#_c_108_n N_A_32_368#_M1003_g 0.00527003f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_102 N_A_187_244#_c_109_n N_A_32_368#_M1003_g 0.0122808f $X=2.645 $Y=0.515
+ $X2=0 $Y2=0
cc_103 N_A_187_244#_c_123_p N_A_32_368#_M1003_g 0.0068369f $X=2.597 $Y=1.005
+ $X2=0 $Y2=0
cc_104 N_A_187_244#_c_108_n N_A_32_368#_c_207_n 0.00152841f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_105 N_A_187_244#_c_114_n N_A_32_368#_c_207_n 0.00305606f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_106 N_A_187_244#_c_114_n N_A_32_368#_M1006_g 0.032028f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_107 N_A_187_244#_M1004_g N_A_32_368#_c_201_n 0.00167994f $X=1.475 $Y=2.4
+ $X2=0 $Y2=0
cc_108 N_A_187_244#_c_119_p N_A_32_368#_c_201_n 0.00602892f $X=2.385 $Y=1.005
+ $X2=0 $Y2=0
cc_109 N_A_187_244#_c_107_n N_A_32_368#_c_201_n 0.00180262f $X=1.735 $Y=1.005
+ $X2=0 $Y2=0
cc_110 N_A_187_244#_c_110_n N_A_32_368#_c_201_n 0.018977f $X=1.525 $Y=1.385
+ $X2=0 $Y2=0
cc_111 N_A_187_244#_c_114_n N_A_32_368#_c_201_n 0.00530616f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_112 N_A_187_244#_c_108_n N_A_32_368#_c_202_n 0.00903297f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_113 N_A_187_244#_c_108_n N_A_32_368#_c_203_n 0.00353279f $X=2.47 $Y=1.76
+ $X2=0 $Y2=0
cc_114 N_A_187_244#_M1002_g N_A_32_368#_c_211_n 7.22282e-19 $X=1.025 $Y=2.4
+ $X2=0 $Y2=0
cc_115 N_A_187_244#_c_104_n N_A_32_368#_c_204_n 5.80921e-19 $X=1.185 $Y=1.22
+ $X2=0 $Y2=0
cc_116 N_A_187_244#_c_110_n N_A_32_368#_c_204_n 0.0100161f $X=1.525 $Y=1.385
+ $X2=0 $Y2=0
cc_117 N_A_187_244#_M1002_g N_A_32_368#_c_246_n 0.0191438f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_118 N_A_187_244#_M1004_g N_A_32_368#_c_246_n 0.0221395f $X=1.475 $Y=2.4 $X2=0
+ $Y2=0
cc_119 N_A_187_244#_c_114_n N_A_32_368#_c_246_n 0.0113609f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_120 N_A_187_244#_M1004_g N_A_32_368#_c_205_n 0.00838506f $X=1.475 $Y=2.4
+ $X2=0 $Y2=0
cc_121 N_A_187_244#_c_119_p N_A_32_368#_c_205_n 0.0286626f $X=2.385 $Y=1.005
+ $X2=0 $Y2=0
cc_122 N_A_187_244#_c_107_n N_A_32_368#_c_205_n 0.0350515f $X=1.735 $Y=1.005
+ $X2=0 $Y2=0
cc_123 N_A_187_244#_c_108_n N_A_32_368#_c_205_n 0.0314791f $X=2.47 $Y=1.76 $X2=0
+ $Y2=0
cc_124 N_A_187_244#_c_110_n N_A_32_368#_c_205_n 9.88986e-19 $X=1.525 $Y=1.385
+ $X2=0 $Y2=0
cc_125 N_A_187_244#_c_114_n N_A_32_368#_c_205_n 0.0183437f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_126 N_A_187_244#_c_114_n N_A_32_368#_c_255_n 0.0174708f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_127 N_A_187_244#_c_104_n N_A_32_368#_c_206_n 0.00105802f $X=1.185 $Y=1.22
+ $X2=0 $Y2=0
cc_128 N_A_187_244#_c_108_n N_A1_M1011_g 0.00286552f $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_129 N_A_187_244#_c_109_n N_A1_M1011_g 0.0111096f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_130 N_A_187_244#_c_123_p N_A1_M1011_g 0.00346711f $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_131 N_A_187_244#_c_108_n N_A1_M1007_g 4.44452e-19 $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_132 N_A_187_244#_c_114_n N_A1_M1007_g 0.00403551f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_133 N_A_187_244#_c_108_n N_A1_c_300_n 0.00177514f $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_134 N_A_187_244#_c_123_p N_A1_c_300_n 7.83088e-19 $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_135 N_A_187_244#_c_108_n N_A1_c_301_n 0.0395719f $X=2.47 $Y=1.76 $X2=0 $Y2=0
cc_136 N_A_187_244#_c_114_n N_A1_c_301_n 0.00172161f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_137 N_A_187_244#_c_123_p N_A1_c_301_n 0.00451909f $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_138 N_A_187_244#_c_109_n N_A2_M1009_g 0.00172432f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_139 N_A_187_244#_c_123_p N_A2_M1009_g 5.12803e-19 $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_140 N_A_187_244#_M1002_g N_VPWR_c_365_n 0.0137777f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_141 N_A_187_244#_M1004_g N_VPWR_c_365_n 0.00149196f $X=1.475 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_187_244#_M1002_g N_VPWR_c_366_n 0.00149196f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_143 N_A_187_244#_M1004_g N_VPWR_c_366_n 0.0137777f $X=1.475 $Y=2.4 $X2=0
+ $Y2=0
cc_144 N_A_187_244#_c_114_n N_VPWR_c_366_n 0.0310049f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_145 N_A_187_244#_M1002_g N_VPWR_c_369_n 0.00460063f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_146 N_A_187_244#_M1004_g N_VPWR_c_369_n 0.00460063f $X=1.475 $Y=2.4 $X2=0
+ $Y2=0
cc_147 N_A_187_244#_c_114_n N_VPWR_c_370_n 0.0157979f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_148 N_A_187_244#_M1002_g N_VPWR_c_364_n 0.00908554f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_149 N_A_187_244#_M1004_g N_VPWR_c_364_n 0.00908554f $X=1.475 $Y=2.4 $X2=0
+ $Y2=0
cc_150 N_A_187_244#_c_114_n N_VPWR_c_364_n 0.0129376f $X=2.22 $Y=2.225 $X2=0
+ $Y2=0
cc_151 N_A_187_244#_c_104_n N_X_c_422_n 0.0201735f $X=1.185 $Y=1.22 $X2=0 $Y2=0
cc_152 N_A_187_244#_c_106_n N_X_c_422_n 0.0101064f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_153 N_A_187_244#_c_107_n N_X_c_422_n 0.0177631f $X=1.735 $Y=1.005 $X2=0 $Y2=0
cc_154 N_A_187_244#_c_110_n N_X_c_422_n 0.00101837f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_155 N_A_187_244#_M1002_g N_X_c_423_n 0.00953176f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_187_244#_c_104_n N_X_c_423_n 0.00468919f $X=1.185 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A_187_244#_M1004_g N_X_c_423_n 0.00419426f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_187_244#_c_106_n N_X_c_423_n 5.48773e-19 $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A_187_244#_c_107_n N_X_c_423_n 0.0312442f $X=1.735 $Y=1.005 $X2=0 $Y2=0
cc_160 N_A_187_244#_c_110_n N_X_c_423_n 0.00950173f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_161 N_A_187_244#_M1002_g N_X_c_425_n 0.00570912f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_187_244#_M1004_g N_X_c_425_n 0.00419833f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_187_244#_c_107_n N_X_c_425_n 0.00290413f $X=1.735 $Y=1.005 $X2=0
+ $Y2=0
cc_164 N_A_187_244#_c_110_n N_X_c_425_n 0.00578305f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_165 N_A_187_244#_c_114_n N_A_507_392#_c_459_n 0.0277129f $X=2.22 $Y=2.225
+ $X2=0 $Y2=0
cc_166 N_A_187_244#_c_119_p N_VGND_M1005_d 0.0154162f $X=2.385 $Y=1.005 $X2=0
+ $Y2=0
cc_167 N_A_187_244#_c_104_n N_VGND_c_482_n 0.00487752f $X=1.185 $Y=1.22 $X2=0
+ $Y2=0
cc_168 N_A_187_244#_c_110_n N_VGND_c_482_n 0.00290042f $X=1.525 $Y=1.385 $X2=0
+ $Y2=0
cc_169 N_A_187_244#_c_106_n N_VGND_c_483_n 0.00422881f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_170 N_A_187_244#_c_119_p N_VGND_c_483_n 0.0448286f $X=2.385 $Y=1.005 $X2=0
+ $Y2=0
cc_171 N_A_187_244#_c_109_n N_VGND_c_483_n 0.0158686f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_172 N_A_187_244#_c_109_n N_VGND_c_485_n 0.0157759f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_173 N_A_187_244#_c_123_p N_VGND_c_485_n 0.00499344f $X=2.597 $Y=1.005 $X2=0
+ $Y2=0
cc_174 N_A_187_244#_c_104_n N_VGND_c_488_n 0.00421809f $X=1.185 $Y=1.22 $X2=0
+ $Y2=0
cc_175 N_A_187_244#_c_106_n N_VGND_c_488_n 0.00433139f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_176 N_A_187_244#_c_109_n N_VGND_c_489_n 0.0144922f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_177 N_A_187_244#_c_104_n N_VGND_c_491_n 0.00443777f $X=1.185 $Y=1.22 $X2=0
+ $Y2=0
cc_178 N_A_187_244#_c_106_n N_VGND_c_491_n 0.00819075f $X=1.615 $Y=1.22 $X2=0
+ $Y2=0
cc_179 N_A_187_244#_c_109_n N_VGND_c_491_n 0.0118826f $X=2.645 $Y=0.515 $X2=0
+ $Y2=0
cc_180 N_A_32_368#_M1003_g N_A1_M1011_g 0.0130291f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_32_368#_c_207_n N_A1_M1007_g 0.027922f $X=2.445 $Y=1.82 $X2=0 $Y2=0
cc_182 N_A_32_368#_c_203_n N_A1_M1007_g 0.00571367f $X=2.445 $Y=1.73 $X2=0 $Y2=0
cc_183 N_A_32_368#_c_202_n N_A1_c_300_n 0.0206661f $X=2.43 $Y=1.425 $X2=0 $Y2=0
cc_184 N_A_32_368#_c_202_n N_A1_c_301_n 3.61775e-19 $X=2.43 $Y=1.425 $X2=0 $Y2=0
cc_185 N_A_32_368#_c_203_n N_A1_c_301_n 4.76375e-19 $X=2.445 $Y=1.73 $X2=0 $Y2=0
cc_186 N_A_32_368#_c_217_n N_VPWR_M1001_d 6.29515e-19 $X=0.68 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_32_368#_c_204_n N_VPWR_M1001_d 0.00873042f $X=0.765 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_32_368#_c_246_n N_VPWR_M1001_d 0.00131722f $X=1.605 $Y=2.325
+ $X2=-0.19 $Y2=-0.245
cc_189 N_A_32_368#_c_266_p N_VPWR_M1001_d 0.00185913f $X=0.765 $Y=2.325
+ $X2=-0.19 $Y2=-0.245
cc_190 N_A_32_368#_c_246_n N_VPWR_M1004_s 0.00467309f $X=1.605 $Y=2.325 $X2=0
+ $Y2=0
cc_191 N_A_32_368#_c_205_n N_VPWR_M1004_s 0.00113495f $X=1.707 $Y=1.89 $X2=0
+ $Y2=0
cc_192 N_A_32_368#_c_255_n N_VPWR_M1004_s 0.00686721f $X=1.707 $Y=2.24 $X2=0
+ $Y2=0
cc_193 N_A_32_368#_c_217_n N_VPWR_c_365_n 0.00183477f $X=0.68 $Y=2.325 $X2=0
+ $Y2=0
cc_194 N_A_32_368#_c_211_n N_VPWR_c_365_n 0.00497738f $X=0.45 $Y=2.325 $X2=0
+ $Y2=0
cc_195 N_A_32_368#_c_246_n N_VPWR_c_365_n 0.00440852f $X=1.605 $Y=2.325 $X2=0
+ $Y2=0
cc_196 N_A_32_368#_c_266_p N_VPWR_c_365_n 0.0152373f $X=0.765 $Y=2.325 $X2=0
+ $Y2=0
cc_197 N_A_32_368#_M1006_g N_VPWR_c_366_n 0.00368778f $X=2.445 $Y=2.46 $X2=0
+ $Y2=0
cc_198 N_A_32_368#_c_246_n N_VPWR_c_366_n 0.0191357f $X=1.605 $Y=2.325 $X2=0
+ $Y2=0
cc_199 N_A_32_368#_M1006_g N_VPWR_c_367_n 7.10319e-19 $X=2.445 $Y=2.46 $X2=0
+ $Y2=0
cc_200 N_A_32_368#_c_211_n N_VPWR_c_368_n 0.006683f $X=0.45 $Y=2.325 $X2=0 $Y2=0
cc_201 N_A_32_368#_M1006_g N_VPWR_c_370_n 0.0048691f $X=2.445 $Y=2.46 $X2=0
+ $Y2=0
cc_202 N_A_32_368#_M1006_g N_VPWR_c_364_n 0.00878547f $X=2.445 $Y=2.46 $X2=0
+ $Y2=0
cc_203 N_A_32_368#_c_211_n N_VPWR_c_364_n 0.010015f $X=0.45 $Y=2.325 $X2=0 $Y2=0
cc_204 N_A_32_368#_c_246_n N_X_M1002_d 0.00761462f $X=1.605 $Y=2.325 $X2=0 $Y2=0
cc_205 N_A_32_368#_c_204_n N_X_c_422_n 0.00229049f $X=0.765 $Y=2.24 $X2=0 $Y2=0
cc_206 N_A_32_368#_c_206_n N_X_c_422_n 0.0187392f $X=0.435 $Y=0.775 $X2=0 $Y2=0
cc_207 N_A_32_368#_c_204_n N_X_c_423_n 0.0562054f $X=0.765 $Y=2.24 $X2=0 $Y2=0
cc_208 N_A_32_368#_c_205_n N_X_c_423_n 0.00438884f $X=1.707 $Y=1.89 $X2=0 $Y2=0
cc_209 N_A_32_368#_c_204_n N_X_c_425_n 0.0186884f $X=0.765 $Y=2.24 $X2=0 $Y2=0
cc_210 N_A_32_368#_c_246_n N_X_c_425_n 0.020291f $X=1.605 $Y=2.325 $X2=0 $Y2=0
cc_211 N_A_32_368#_c_205_n N_X_c_425_n 0.00319331f $X=1.707 $Y=1.89 $X2=0 $Y2=0
cc_212 N_A_32_368#_M1006_g N_A_507_392#_c_459_n 8.26109e-19 $X=2.445 $Y=2.46
+ $X2=0 $Y2=0
cc_213 N_A_32_368#_c_204_n N_VGND_M1010_d 8.56368e-19 $X=0.765 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_32_368#_c_206_n N_VGND_M1010_d 0.00257106f $X=0.435 $Y=0.775
+ $X2=-0.19 $Y2=-0.245
cc_215 N_A_32_368#_c_206_n N_VGND_c_482_n 0.0124903f $X=0.435 $Y=0.775 $X2=0
+ $Y2=0
cc_216 N_A_32_368#_M1003_g N_VGND_c_483_n 0.0042292f $X=2.43 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_32_368#_c_206_n N_VGND_c_486_n 0.00797936f $X=0.435 $Y=0.775 $X2=0
+ $Y2=0
cc_218 N_A_32_368#_M1003_g N_VGND_c_489_n 0.00434272f $X=2.43 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_32_368#_M1003_g N_VGND_c_491_n 0.00822841f $X=2.43 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_32_368#_c_206_n N_VGND_c_491_n 0.0179874f $X=0.435 $Y=0.775 $X2=0
+ $Y2=0
cc_221 N_A1_M1011_g N_A2_M1009_g 0.0375784f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_c_300_n N_A2_M1009_g 0.019932f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_223 N_A1_c_301_n N_A2_M1009_g 0.00865654f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_224 N_A1_c_301_n A2 0.0270452f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_225 N_A1_M1007_g N_A2_c_340_n 0.0514121f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_226 N_A1_M1007_g N_VPWR_c_367_n 0.0117786f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_227 N_A1_M1007_g N_VPWR_c_370_n 0.00460063f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_228 N_A1_M1007_g N_VPWR_c_364_n 0.00908665f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_229 N_A1_M1007_g N_A_507_392#_c_462_n 0.0152168f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_230 N_A1_c_301_n N_A_507_392#_c_462_n 0.0202388f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_231 N_A1_M1007_g N_A_507_392#_c_457_n 7.15258e-19 $X=2.895 $Y=2.46 $X2=0
+ $Y2=0
cc_232 N_A1_M1007_g N_A_507_392#_c_458_n 7.4508e-19 $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_233 N_A1_M1007_g N_A_507_392#_c_459_n 8.34606e-19 $X=2.895 $Y=2.46 $X2=0
+ $Y2=0
cc_234 N_A1_c_300_n N_A_507_392#_c_459_n 4.71617e-19 $X=2.88 $Y=1.425 $X2=0
+ $Y2=0
cc_235 N_A1_c_301_n N_A_507_392#_c_459_n 0.0014591f $X=2.88 $Y=1.425 $X2=0 $Y2=0
cc_236 N_A1_M1011_g N_VGND_c_485_n 0.00277908f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1011_g N_VGND_c_489_n 0.00434272f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_M1011_g N_VGND_c_491_n 0.00821825f $X=2.86 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A2_M1008_g N_VPWR_c_367_n 0.0035371f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_240 N_A2_M1008_g N_VPWR_c_371_n 0.005209f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_241 N_A2_M1008_g N_VPWR_c_364_n 0.00986083f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_242 N_A2_M1008_g N_A_507_392#_c_462_n 0.0174429f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_243 N_A2_M1008_g N_A_507_392#_c_457_n 0.00394102f $X=3.345 $Y=2.46 $X2=0
+ $Y2=0
cc_244 A2 N_A_507_392#_c_457_n 0.0276657f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A2_c_340_n N_A_507_392#_c_457_n 0.00236651f $X=3.57 $Y=1.615 $X2=0
+ $Y2=0
cc_246 N_A2_M1008_g N_A_507_392#_c_458_n 0.0105176f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_247 N_A2_M1009_g N_VGND_c_485_n 0.0203366f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_248 A2 N_VGND_c_485_n 0.0126785f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A2_c_340_n N_VGND_c_485_n 0.00193914f $X=3.57 $Y=1.615 $X2=0 $Y2=0
cc_250 N_A2_M1009_g N_VGND_c_489_n 0.00383152f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1009_g N_VGND_c_491_n 0.00757998f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_252 N_VPWR_M1007_d N_A_507_392#_c_462_n 0.00384175f $X=2.985 $Y=1.96 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_367_n N_A_507_392#_c_462_n 0.014901f $X=3.12 $Y=2.71 $X2=0 $Y2=0
cc_254 N_VPWR_c_367_n N_A_507_392#_c_458_n 0.0184665f $X=3.12 $Y=2.71 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_371_n N_A_507_392#_c_458_n 0.014549f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_364_n N_A_507_392#_c_458_n 0.0119743f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_367_n N_A_507_392#_c_459_n 0.017687f $X=3.12 $Y=2.71 $X2=0 $Y2=0
cc_258 N_VPWR_c_370_n N_A_507_392#_c_459_n 0.00749631f $X=2.955 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_364_n N_A_507_392#_c_459_n 0.0062048f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_260 N_X_c_422_n N_VGND_M1010_d 0.00215131f $X=1.105 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_261 N_X_c_423_n N_VGND_M1010_d 6.05713e-19 $X=1.105 $Y=1.82 $X2=-0.19
+ $Y2=-0.245
cc_262 N_X_c_422_n N_VGND_c_482_n 0.0157951f $X=1.105 $Y=1.04 $X2=0 $Y2=0
cc_263 N_X_c_422_n N_VGND_c_483_n 0.0160262f $X=1.105 $Y=1.04 $X2=0 $Y2=0
cc_264 N_X_c_422_n N_VGND_c_488_n 0.0147221f $X=1.105 $Y=1.04 $X2=0 $Y2=0
cc_265 N_X_c_422_n N_VGND_c_491_n 0.0180091f $X=1.105 $Y=1.04 $X2=0 $Y2=0

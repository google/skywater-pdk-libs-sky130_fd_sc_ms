* NGSPICE file created from sky130_fd_sc_ms__ha_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__ha_2 A B VGND VNB VPB VPWR COUT SUM
M1000 COUT a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.01665e+12p ps=1.023e+07u
M1001 a_278_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.083e+11p pd=4.09e+06u as=0p ps=0u
M1002 SUM a_394_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.9664e+12p ps=1.448e+07u
M1003 VPWR a_394_388# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 SUM a_394_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=0p ps=0u
M1005 a_310_388# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1006 COUT a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1007 VGND B a_278_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_27_74# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1010 a_394_388# B a_310_388# VPB pshort w=1e+06u l=180000u
+  ad=9.6e+11p pd=3.92e+06u as=0p ps=0u
M1011 VPWR a_27_74# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_394_388# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_74# a_394_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1015 VPWR A a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_114_74# B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_278_74# a_27_74# a_394_388# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.01625e+11p ps=2.05e+06u
.ends


* File: sky130_fd_sc_ms__o211a_4.spice
* Created: Fri Aug 28 17:53:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o211a_4.pex.spice"
.subckt sky130_fd_sc_ms__o211a_4  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_91_48#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_91_48#_M1013_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1013_d N_A_91_48#_M1016_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_91_48#_M1017_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_510_125#_M1014_d N_B1_M1014_g N_A_597_125#_M1014_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1817 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1015 N_A_597_125#_M1014_s N_C1_M1015_g N_A_91_48#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1020 N_A_597_125#_M1020_d N_C1_M1020_g N_A_91_48#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_510_125#_M1019_d N_B1_M1019_g N_A_597_125#_M1020_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1152 AS=0.112 PD=1 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_A1_M1012_g N_A_510_125#_M1019_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0992 AS=0.1152 PD=0.95 PS=1 NRD=0.936 NRS=14.988 M=1 R=4.26667 SA=75002.1
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 N_A_510_125#_M1011_d N_A2_M1011_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1072 AS=0.0992 PD=0.975 PS=0.95 NRD=10.308 NRS=4.68 M=1 R=4.26667
+ SA=75002.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1021 N_A_510_125#_M1011_d N_A2_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1072 AS=0.112 PD=0.975 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1021_s N_A1_M1022_g N_A_510_125#_M1022_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75003.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_X_M1004_d N_A_91_48#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90004.8 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1004_d N_A_91_48#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1008_d N_A_91_48#_M1008_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.2
+ SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1008_d N_A_91_48#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.301943 PD=1.39 PS=1.88571 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.7 SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1009_s N_B1_M1010_g N_A_91_48#_M1010_s VPB PSHORT L=0.18 W=0.84
+ AD=0.226457 AS=0.1134 PD=1.41429 PS=1.11 NRD=48.659 NRS=0 M=1 R=4.66667
+ SA=90002.4 SB=90003.7 A=0.1512 P=2.04 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_A_91_48#_M1010_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1617 AS=0.1134 PD=1.225 PS=1.11 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90002.8 SB=90003.2 A=0.1512 P=2.04 MULT=1
MM1007 N_VPWR_M1000_d N_C1_M1007_g N_A_91_48#_M1007_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1617 AS=0.1134 PD=1.225 PS=1.11 NRD=14.0658 NRS=0 M=1 R=4.66667
+ SA=90003.4 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1023 N_VPWR_M1023_d N_B1_M1023_g N_A_91_48#_M1007_s VPB PSHORT L=0.18 W=0.84
+ AD=0.179413 AS=0.1134 PD=1.28283 PS=1.11 NRD=19.3454 NRS=0 M=1 R=4.66667
+ SA=90003.9 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1023_d N_A1_M1005_g N_A_971_391#_M1005_s VPB PSHORT L=0.18 W=1
+ AD=0.213587 AS=0.135 PD=1.52717 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90003.8 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1001 N_A_971_391#_M1005_s N_A2_M1001_g N_A_91_48#_M1001_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90004.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1003 N_A_971_391#_M1003_d N_A2_M1003_g N_A_91_48#_M1001_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90004.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_971_391#_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.33 AS=0.135 PD=2.66 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90005.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ms__o211a_4.pxi.spice"
*
.ends
*
*

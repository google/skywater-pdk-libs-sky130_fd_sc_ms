* File: sky130_fd_sc_ms__sdfrtp_4.spice
* Created: Wed Sep  2 12:30:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfrtp_4.pex.spice"
.subckt sky130_fd_sc_ms__sdfrtp_4  VNB VPB SCE D SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1042 N_VGND_M1042_d N_SCE_M1042_g N_A_27_74#_M1042_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 noxref_25 N_A_27_74#_M1007_g N_noxref_24_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.07665 AS=0.1197 PD=0.785 PS=1.41 NRD=36.42 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 N_A_415_81#_M1008_d N_D_M1008_g noxref_25 VNB NLOWVT L=0.15 W=0.42
+ AD=0.1155 AS=0.07665 PD=0.97 PS=0.785 NRD=77.136 NRS=36.42 M=1 R=2.8
+ SA=75000.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1025 noxref_26 N_SCE_M1025_g N_A_415_81#_M1008_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=0.97 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_noxref_24_M1005_d N_SCD_M1005_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0693 AS=0.0441 PD=0.75 PS=0.63 NRD=8.568 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_RESET_B_M1013_g N_noxref_24_M1005_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0693 PD=1.41 PS=0.75 NRD=5.712 NRS=5.712 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_CLK_M1038_g N_A_834_93#_M1038_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.16425 AS=0.27955 PD=1.27 PS=2.44 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75000.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1041 N_A_1037_387#_M1041_d N_A_834_93#_M1041_g N_VGND_M1038_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1924 AS=0.16425 PD=2 PS=1.27 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_1233_138#_M1027_d N_A_834_93#_M1027_g N_A_415_81#_M1027_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1017 A_1319_138# N_A_1037_387#_M1017_g N_A_1233_138#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1000 A_1397_138# N_A_1367_112#_M1000_g A_1319_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_RESET_B_M1034_g A_1397_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20551 AS=0.0504 PD=1.19845 PS=0.66 NRD=124.08 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1028 N_A_1367_112#_M1028_d N_A_1233_138#_M1028_g N_VGND_M1034_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.124942 AS=0.36209 PD=1.14217 PS=2.11155 NRD=0 NRS=70.428
+ M=1 R=4.93333 SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1006 N_A_1745_74#_M1006_d N_A_1037_387#_M1006_g N_A_1367_112#_M1028_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.261434 AS=0.108058 PD=1.85962 PS=0.987826
+ NRD=101.244 NRS=0 M=1 R=4.26667 SA=75001.9 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1036 A_1955_74# N_A_834_93#_M1036_g N_A_1745_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.171566 PD=0.66 PS=1.22038 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75002.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_2003_48#_M1032_g A_1955_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=15.708 NRS=18.564 M=1 R=2.8 SA=75002.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1045 A_2141_74# N_RESET_B_M1045_g N_VGND_M1032_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75003.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_2003_48#_M1030_d N_A_1745_74#_M1030_g A_2141_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1512 AS=0.0441 PD=1.56 PS=0.63 NRD=9.996 NRS=14.28 M=1 R=2.8
+ SA=75003.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_1745_74#_M1011_g N_A_2339_74#_M1011_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1011_d N_A_2339_74#_M1009_g N_Q_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_2339_74#_M1020_g N_Q_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3293 AS=0.1036 PD=1.63 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1020_d N_A_2339_74#_M1033_g N_Q_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3293 AS=0.1036 PD=1.63 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1037 N_VGND_M1037_d N_A_2339_74#_M1037_g N_Q_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_SCE_M1004_g N_A_27_74#_M1004_s VPB PSHORT L=0.18 W=0.64
+ AD=0.3008 AS=0.1792 PD=1.58 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90003.3 A=0.1152 P=1.64 MULT=1
MM1039 A_343_464# N_SCE_M1039_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.3008 PD=0.88 PS=1.58 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90001.3
+ SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1021 N_A_415_81#_M1021_d N_D_M1021_g A_343_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.7
+ SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1024 A_517_464# N_A_27_74#_M1024_g N_A_415_81#_M1021_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1216 AS=0.0864 PD=1.02 PS=0.91 NRD=41.5473 NRS=0 M=1 R=3.55556
+ SA=90002.2 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1043 N_VPWR_M1043_d N_SCD_M1043_g A_517_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1248 AS=0.1216 PD=1.03 PS=1.02 NRD=0 NRS=41.5473 M=1 R=3.55556 SA=90002.7
+ SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1035 N_A_415_81#_M1035_d N_RESET_B_M1035_g N_VPWR_M1043_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1824 AS=0.1248 PD=1.85 PS=1.03 NRD=0 NRS=33.8446 M=1 R=3.55556
+ SA=90003.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1026 N_VPWR_M1026_d N_CLK_M1026_g N_A_834_93#_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1040 N_A_1037_387#_M1040_d N_A_834_93#_M1040_g N_VPWR_M1026_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1016 N_A_1233_138#_M1016_d N_A_1037_387#_M1016_g N_A_415_81#_M1016_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1012 A_1345_463# N_A_834_93#_M1012_g N_A_1233_138#_M1016_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_1367_112#_M1002_g A_1345_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.133025 AS=0.0441 PD=1.115 PS=0.63 NRD=122.751 NRS=23.443 M=1 R=2.33333
+ SA=90001.1 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1003 N_A_1233_138#_M1003_d N_RESET_B_M1003_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.133025 PD=1.4 PS=1.115 NRD=0 NRS=122.751 M=1 R=2.33333
+ SA=90001.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1018 N_A_1367_112#_M1018_d N_A_1233_138#_M1018_g N_VPWR_M1018_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1022 N_A_1745_74#_M1022_d N_A_834_93#_M1022_g N_A_1367_112#_M1018_d VPB PSHORT
+ L=0.18 W=1 AD=0.286602 AS=0.135 PD=2.47183 PS=1.27 NRD=33.4703 NRS=0 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1014 A_1985_508# N_A_1037_387#_M1014_g N_A_1745_74#_M1022_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.120373 PD=0.66 PS=1.03817 NRD=30.4759 NRS=39.8531 M=1
+ R=2.33333 SA=90000.8 SB=90002.8 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_2003_48#_M1010_g A_1985_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.10605 AS=0.0504 PD=0.925 PS=0.66 NRD=68.0044 NRS=30.4759 M=1 R=2.33333
+ SA=90001.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1031 N_A_2003_48#_M1031_d N_RESET_B_M1031_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.42 AD=0.07455 AS=0.10605 PD=0.775 PS=0.925 NRD=0 NRS=37.5088 M=1 R=2.33333
+ SA=90001.9 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1044 N_VPWR_M1044_d N_A_1745_74#_M1044_g N_A_2003_48#_M1031_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1134 AS=0.07455 PD=1.00333 PS=0.775 NRD=53.9386 NRS=37.5088
+ M=1 R=2.33333 SA=90002.5 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1001 N_VPWR_M1044_d N_A_1745_74#_M1001_g N_A_2339_74#_M1001_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.2268 AS=0.1134 PD=2.00667 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.8 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1046 N_VPWR_M1046_d N_A_1745_74#_M1046_g N_A_2339_74#_M1001_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1614 AS=0.1134 PD=1.26429 PS=1.11 NRD=18.7544 NRS=0 M=1
+ R=4.66667 SA=90001.2 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1015 N_Q_M1015_d N_A_2339_74#_M1015_g N_VPWR_M1046_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2152 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.4
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1019 N_Q_M1015_d N_A_2339_74#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.8
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1023 N_Q_M1023_d N_A_2339_74#_M1023_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1029 N_Q_M1023_d N_A_2339_74#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX47_noxref VNB VPB NWDIODE A=28.5069 P=34.48
c_159 VNB 0 1.59743e-19 $X=0 $Y=0
c_2400 A_1397_138# 0 1.57165e-19 $X=6.985 $Y=0.69
*
.include "sky130_fd_sc_ms__sdfrtp_4.pxi.spice"
*
.ends
*
*

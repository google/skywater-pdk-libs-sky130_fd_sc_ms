* File: sky130_fd_sc_ms__o22a_4.pex.spice
* Created: Fri Aug 28 17:58:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O22A_4%A2 3 7 9 11 14 16 22 23
c53 23 0 1.5038e-19 $X=1.425 $Y=1.587
c54 3 0 9.05627e-20 $X=0.955 $Y=2.46
r55 23 24 4.30357 $w=3.36e-07 $l=3e-08 $layer=POLY_cond $X=1.425 $Y=1.587
+ $X2=1.455 $Y2=1.587
r56 21 23 10.7589 $w=3.36e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.587
+ $X2=1.425 $Y2=1.587
r57 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.615 $X2=1.35 $Y2=1.615
r58 16 22 0.892596 $w=6.68e-07 $l=5e-08 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.615
r59 12 24 17.3521 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.455 $Y=1.78
+ $X2=1.455 $Y2=1.587
r60 12 14 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.455 $Y=1.78
+ $X2=1.455 $Y2=2.46
r61 9 23 21.6522 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.425 $Y=1.395
+ $X2=1.425 $Y2=1.587
r62 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=1.395
+ $X2=1.425 $Y2=1
r63 5 21 50.9256 $w=3.36e-07 $l=3.55e-07 $layer=POLY_cond $X=0.995 $Y=1.587
+ $X2=1.35 $Y2=1.587
r64 5 18 5.7381 $w=3.36e-07 $l=4e-08 $layer=POLY_cond $X=0.995 $Y=1.587
+ $X2=0.955 $Y2=1.587
r65 5 7 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.995 $Y=1.45
+ $X2=0.995 $Y2=1
r66 1 18 17.3521 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.955 $Y=1.78
+ $X2=0.955 $Y2=1.587
r67 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.955 $Y=1.78
+ $X2=0.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%A1 3 6 8 9 10 13 18 19 22
r66 22 25 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.615
+ $X2=2.01 $Y2=1.78
r67 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.615
+ $X2=2.01 $Y2=1.45
r68 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.01
+ $Y=1.615 $X2=2.01 $Y2=1.615
r69 19 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=2.01 $Y2=1.615
r70 18 24 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.965 $Y=1 $X2=1.965
+ $Y2=1.45
r71 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.965 $Y=0.31
+ $X2=1.965 $Y2=1
r72 13 25 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.955 $Y=2.46
+ $X2=1.955 $Y2=1.78
r73 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.89 $Y=0.235
+ $X2=1.965 $Y2=0.31
r74 9 10 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=1.89 $Y=0.235
+ $X2=0.57 $Y2=0.235
r75 6 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.395
+ $X2=0.495 $Y2=1
r76 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.31
+ $X2=0.57 $Y2=0.235
r77 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=0.31
+ $X2=0.495 $Y2=1
r78 1 6 70.5366 $w=1.64e-07 $l=2.44949e-07 $layer=POLY_cond $X=0.505 $Y=1.635
+ $X2=0.495 $Y2=1.395
r79 1 3 320.685 $w=1.8e-07 $l=8.25e-07 $layer=POLY_cond $X=0.505 $Y=1.635
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%B2 3 7 9 11 14 16 17 24 25
c55 24 0 1.52901e-19 $X=3.34 $Y=1.615
c56 3 0 1.28833e-19 $X=2.925 $Y=1
r57 25 26 3.50291 $w=3.44e-07 $l=2.5e-08 $layer=POLY_cond $X=3.43 $Y=1.587
+ $X2=3.455 $Y2=1.587
r58 23 25 12.6105 $w=3.44e-07 $l=9e-08 $layer=POLY_cond $X=3.34 $Y=1.587
+ $X2=3.43 $Y2=1.587
r59 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.34
+ $Y=1.615 $X2=3.34 $Y2=1.615
r60 21 23 53.9448 $w=3.44e-07 $l=3.85e-07 $layer=POLY_cond $X=2.955 $Y=1.587
+ $X2=3.34 $Y2=1.587
r61 17 24 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.12 $Y=1.615
+ $X2=3.34 $Y2=1.615
r62 16 17 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=3.12 $Y2=1.615
r63 12 26 17.902 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.455 $Y=1.78
+ $X2=3.455 $Y2=1.587
r64 12 14 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.455 $Y=1.78
+ $X2=3.455 $Y2=2.46
r65 9 25 22.2144 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.43 $Y=1.395
+ $X2=3.43 $Y2=1.587
r66 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.43 $Y=1.395
+ $X2=3.43 $Y2=1
r67 5 21 17.902 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.955 $Y=1.78
+ $X2=2.955 $Y2=1.587
r68 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.955 $Y=1.78
+ $X2=2.955 $Y2=2.46
r69 1 21 4.20349 $w=3.44e-07 $l=3e-08 $layer=POLY_cond $X=2.925 $Y=1.587
+ $X2=2.955 $Y2=1.587
r70 1 3 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.925 $Y=1.45
+ $X2=2.925 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%B1 4 5 7 9 14 17 21 22 24
c74 22 0 1.28833e-19 $X=2.16 $Y=0.555
c75 17 0 1.52901e-19 $X=3.955 $Y=2.46
r76 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=0.405
+ $X2=2.445 $Y2=0.57
r77 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.445
+ $Y=0.405 $X2=2.445 $Y2=0.405
r78 24 27 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.445 $Y=0.235
+ $X2=2.445 $Y2=0.405
r79 22 28 9.79437 $w=3.55e-07 $l=2.85e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=2.445 $Y2=0.462
r80 20 21 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.915 $Y=1.395
+ $X2=3.915 $Y2=1.545
r81 17 21 355.669 $w=1.8e-07 $l=9.15e-07 $layer=POLY_cond $X=3.955 $Y=2.46
+ $X2=3.955 $Y2=1.545
r82 14 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.86 $Y=1 $X2=3.86
+ $Y2=1.395
r83 11 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.86 $Y=0.31
+ $X2=3.86 $Y2=1
r84 10 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=0.235
+ $X2=2.445 $Y2=0.235
r85 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.785 $Y=0.235
+ $X2=3.86 $Y2=0.31
r86 9 10 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=3.785 $Y=0.235
+ $X2=2.61 $Y2=0.235
r87 5 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.505 $Y=1.485
+ $X2=2.505 $Y2=1.395
r88 5 7 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=2.505 $Y=1.485
+ $X2=2.505 $Y2=2.46
r89 4 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.49 $Y=1 $X2=2.49
+ $Y2=1.395
r90 4 29 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.49 $Y=1 $X2=2.49
+ $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%A_209_392# 1 2 3 4 15 19 23 27 31 35 39 43 47
+ 55 58 59 61 62 64 67 71 73 76 77 79 89
c175 71 0 9.05627e-20 $X=1.23 $Y=2.115
c176 62 0 1.20589e-19 $X=3.845 $Y=1.595
c177 15 0 2.50841e-19 $X=4.505 $Y=2.4
r178 89 90 8.1319 $w=3.26e-07 $l=5.5e-08 $layer=POLY_cond $X=6.165 $Y=1.515
+ $X2=6.22 $Y2=1.515
r179 88 89 55.4448 $w=3.26e-07 $l=3.75e-07 $layer=POLY_cond $X=5.79 $Y=1.515
+ $X2=6.165 $Y2=1.515
r180 87 88 11.089 $w=3.26e-07 $l=7.5e-08 $layer=POLY_cond $X=5.715 $Y=1.515
+ $X2=5.79 $Y2=1.515
r181 84 85 54.7055 $w=3.26e-07 $l=3.7e-07 $layer=POLY_cond $X=4.99 $Y=1.515
+ $X2=5.36 $Y2=1.515
r182 83 84 8.87117 $w=3.26e-07 $l=6e-08 $layer=POLY_cond $X=4.93 $Y=1.515
+ $X2=4.99 $Y2=1.515
r183 80 83 51.7485 $w=3.26e-07 $l=3.5e-07 $layer=POLY_cond $X=4.58 $Y=1.515
+ $X2=4.93 $Y2=1.515
r184 80 81 11.089 $w=3.26e-07 $l=7.5e-08 $layer=POLY_cond $X=4.58 $Y=1.515
+ $X2=4.505 $Y2=1.515
r185 79 80 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.58
+ $Y=1.515 $X2=4.58 $Y2=1.515
r186 75 77 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0.79
+ $X2=3.81 $Y2=0.79
r187 75 76 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0.79
+ $X2=3.48 $Y2=0.79
r188 68 87 17.0031 $w=3.26e-07 $l=1.15e-07 $layer=POLY_cond $X=5.6 $Y=1.515
+ $X2=5.715 $Y2=1.515
r189 68 85 35.4847 $w=3.26e-07 $l=2.4e-07 $layer=POLY_cond $X=5.6 $Y=1.515
+ $X2=5.36 $Y2=1.515
r190 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.6
+ $Y=1.515 $X2=5.6 $Y2=1.515
r191 65 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=1.515
+ $X2=4.5 $Y2=1.515
r192 65 67 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=4.585 $Y=1.515
+ $X2=5.6 $Y2=1.515
r193 64 79 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=1.35 $X2=4.5
+ $Y2=1.515
r194 63 64 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.5 $Y=0.92 $X2=4.5
+ $Y2=1.35
r195 61 79 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.415 $Y=1.595
+ $X2=4.5 $Y2=1.515
r196 61 62 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.415 $Y=1.595
+ $X2=3.845 $Y2=1.595
r197 59 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.415 $Y=0.835
+ $X2=4.5 $Y2=0.92
r198 59 77 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.415 $Y=0.835
+ $X2=3.81 $Y2=0.835
r199 57 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.76 $Y=1.68
+ $X2=3.845 $Y2=1.595
r200 57 58 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.76 $Y=1.68
+ $X2=3.76 $Y2=1.95
r201 56 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=2.035
+ $X2=3.23 $Y2=2.035
r202 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.675 $Y=2.035
+ $X2=3.76 $Y2=1.95
r203 55 56 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.675 $Y=2.035
+ $X2=3.395 $Y2=2.035
r204 51 76 47.4444 $w=1.78e-07 $l=7.7e-07 $layer=LI1_cond $X=2.71 $Y=0.83
+ $X2=3.48 $Y2=0.83
r205 48 71 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.035
+ $X2=1.23 $Y2=2.035
r206 47 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.23 $Y2=2.035
r207 47 48 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=1.395 $Y2=2.035
r208 41 90 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.22 $Y=1.35
+ $X2=6.22 $Y2=1.515
r209 41 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.22 $Y=1.35
+ $X2=6.22 $Y2=0.74
r210 37 89 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.68
+ $X2=6.165 $Y2=1.515
r211 37 39 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.165 $Y=1.68
+ $X2=6.165 $Y2=2.4
r212 33 88 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.79 $Y=1.35
+ $X2=5.79 $Y2=1.515
r213 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.79 $Y=1.35
+ $X2=5.79 $Y2=0.74
r214 29 87 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.68
+ $X2=5.715 $Y2=1.515
r215 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.715 $Y=1.68
+ $X2=5.715 $Y2=2.4
r216 25 85 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.36 $Y=1.35
+ $X2=5.36 $Y2=1.515
r217 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.36 $Y=1.35
+ $X2=5.36 $Y2=0.74
r218 21 84 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.99 $Y=1.68
+ $X2=4.99 $Y2=1.515
r219 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.99 $Y=1.68
+ $X2=4.99 $Y2=2.4
r220 17 83 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.93 $Y=1.35
+ $X2=4.93 $Y2=1.515
r221 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.93 $Y=1.35
+ $X2=4.93 $Y2=0.74
r222 13 81 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.68
+ $X2=4.505 $Y2=1.515
r223 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.505 $Y=1.68
+ $X2=4.505 $Y2=2.4
r224 4 73 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=3.045
+ $Y=1.96 $X2=3.23 $Y2=2.115
r225 3 71 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.96 $X2=1.23 $Y2=2.115
r226 2 75 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.68 $X2=3.645 $Y2=0.83
r227 1 51 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.68 $X2=2.71 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%VPWR 1 2 3 4 5 16 18 24 28 34 36 38 43 44 46
+ 47 48 50 68 76 80
r82 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r83 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 71 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r86 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r87 68 79 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r88 68 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33 $X2=6
+ $Y2=3.33
r89 67 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r90 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r92 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 61 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 60 63 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r97 58 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r102 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 51 73 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r105 51 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r107 50 56 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 48 64 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 48 61 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 46 66 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.365 $Y2=3.33
r112 45 70 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.53 $Y=3.33 $X2=6
+ $Y2=3.33
r113 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.365 $Y2=3.33
r114 43 63 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.1 $Y=3.33 $X2=4.08
+ $Y2=3.33
r115 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=3.33
+ $X2=4.265 $Y2=3.33
r116 42 66 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.265 $Y2=3.33
r118 38 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.44 $Y=1.985
+ $X2=6.44 $Y2=2.815
r119 36 79 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r120 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.815
r121 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=3.33
r122 32 34 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=2.355
r123 28 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.265 $Y=2.015
+ $X2=4.265 $Y2=2.415
r124 26 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.265 $Y=3.245
+ $X2=4.265 $Y2=3.33
r125 26 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.265 $Y=3.245
+ $X2=4.265 $Y2=2.415
r126 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r127 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.455
r128 18 21 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=2.815
r129 16 73 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r130 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r131 5 41 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.84 $X2=6.44 $Y2=2.815
r132 5 38 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.84 $X2=6.44 $Y2=1.985
r133 4 34 300 $w=1.7e-07 $l=6.41872e-07 $layer=licon1_PDIFF $count=2 $X=5.08
+ $Y=1.84 $X2=5.365 $Y2=2.355
r134 3 31 300 $w=1.7e-07 $l=5.54189e-07 $layer=licon1_PDIFF $count=2 $X=4.045
+ $Y=1.96 $X2=4.265 $Y2=2.415
r135 3 28 600 $w=1.7e-07 $l=2.45967e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.96 $X2=4.265 $Y2=2.015
r136 2 24 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.96 $X2=2.23 $Y2=2.455
r137 1 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r138 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%A_119_392# 1 2 9 13 14 17
c26 9 0 1.5038e-19 $X=0.73 $Y=2.115
r27 15 17 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.73 $Y=2.905
+ $X2=1.73 $Y2=2.455
r28 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=1.73 $Y2=2.905
r29 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=0.895 $Y2=2.99
r30 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.73 $Y=2.115 $X2=0.73
+ $Y2=2.815
r31 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r32 7 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.73 $Y=2.905 $X2=0.73
+ $Y2=2.815
r33 2 17 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.96 $X2=1.73 $Y2=2.455
r34 1 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.815
r35 1 9 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%A_519_392# 1 2 9 11 12 15
c24 15 0 1.58786e-19 $X=3.73 $Y=2.455
c25 11 0 9.20547e-20 $X=3.565 $Y=2.99
r26 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.73 $Y=2.905
+ $X2=3.73 $Y2=2.455
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.565 $Y=2.99
+ $X2=3.73 $Y2=2.905
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.565 $Y=2.99
+ $X2=2.895 $Y2=2.99
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.73 $Y=2.905
+ $X2=2.895 $Y2=2.99
r30 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.73 $Y=2.905 $X2=2.73
+ $Y2=2.455
r31 2 15 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=3.545
+ $Y=1.96 $X2=3.73 $Y2=2.455
r32 1 9 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.96 $X2=2.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%X 1 2 3 4 13 15 17 21 23 24 27 31 33 34 38 42
r72 41 42 18.7898 $w=2.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=1.295
+ $X2=6.48 $Y2=1.295
r73 39 41 13.8636 $w=1.76e-07 $l=2e-07 $layer=LI1_cond $X=6.012 $Y=1.095
+ $X2=6.012 $Y2=1.295
r74 34 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.02 $Y=1.85
+ $X2=5.94 $Y2=1.935
r75 33 41 7.97159 $w=1.76e-07 $l=1.18933e-07 $layer=LI1_cond $X=6.02 $Y=1.41
+ $X2=6.012 $Y2=1.295
r76 33 34 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.02 $Y=1.41
+ $X2=6.02 $Y2=1.85
r77 29 39 5.6459 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.012 $Y=1.01
+ $X2=6.012 $Y2=1.095
r78 29 31 29.6757 $w=1.83e-07 $l=4.95e-07 $layer=LI1_cond $X=6.012 $Y=1.01
+ $X2=6.012 $Y2=0.515
r79 25 38 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.02 $X2=5.94
+ $Y2=1.935
r80 25 27 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=5.94 $Y=2.02
+ $X2=5.94 $Y2=2.815
r81 23 39 0.927112 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=5.92 $Y=1.095
+ $X2=6.012 $Y2=1.095
r82 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.92 $Y=1.095
+ $X2=5.23 $Y2=1.095
r83 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.105 $Y=1.01
+ $X2=5.23 $Y2=1.095
r84 19 21 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.105 $Y=1.01
+ $X2=5.105 $Y2=0.515
r85 18 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=1.935
+ $X2=4.765 $Y2=1.935
r86 17 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=1.935
+ $X2=5.94 $Y2=1.935
r87 17 18 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.775 $Y=1.935
+ $X2=4.93 $Y2=1.935
r88 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=2.02
+ $X2=4.765 $Y2=1.935
r89 13 15 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=4.765 $Y=2.02
+ $X2=4.765 $Y2=2.815
r90 4 38 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.94 $Y2=2.015
r91 4 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.94 $Y2=2.815
r92 3 36 400 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_PDIFF $count=1 $X=4.595
+ $Y=1.84 $X2=4.765 $Y2=2.015
r93 3 15 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=4.595
+ $Y=1.84 $X2=4.765 $Y2=2.815
r94 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.37 $X2=6.005 $Y2=0.515
r95 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.005
+ $Y=0.37 $X2=5.145 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%A_27_136# 1 2 3 4 5 18 20 21 24 32 35 36 38
+ 39
r62 38 39 8.29777 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=1.215
+ $X2=3.91 $Y2=1.215
r63 34 36 8.11354 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.06
+ $X2=2.375 $Y2=1.06
r64 34 35 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.06
+ $X2=2.045 $Y2=1.06
r65 31 39 42.9043 $w=1.88e-07 $l=7.35e-07 $layer=LI1_cond $X=3.175 $Y=1.185
+ $X2=3.91 $Y2=1.185
r66 31 36 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=3.175 $Y=1.185
+ $X2=2.375 $Y2=1.185
r67 27 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.195
+ $X2=1.25 $Y2=1.195
r68 27 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.375 $Y=1.195
+ $X2=2.045 $Y2=1.195
r69 22 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.11
+ $X2=1.25 $Y2=1.195
r70 22 24 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.25 $Y=1.11
+ $X2=1.25 $Y2=0.97
r71 20 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.195
+ $X2=1.25 $Y2=1.195
r72 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.195
+ $X2=0.445 $Y2=1.195
r73 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.445 $Y2=1.195
r74 16 18 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.28 $Y2=0.825
r75 5 38 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.68 $X2=4.075 $Y2=1.175
r76 4 31 182 $w=1.7e-07 $l=5.75891e-07 $layer=licon1_NDIFF $count=1 $X=3 $Y=0.68
+ $X2=3.175 $Y2=1.175
r77 3 34 182 $w=1.7e-07 $l=4.57165e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.68 $X2=2.21 $Y2=1.06
r78 2 24 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.68 $X2=1.21 $Y2=0.97
r79 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 56 61 67 70 73 76 80
r86 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r87 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r88 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r89 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r92 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r93 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r94 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=5.575
+ $Y2=0
r95 62 64 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=6
+ $Y2=0
r96 61 79 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.497
+ $Y2=0
r97 61 64 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6
+ $Y2=0
r98 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r99 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r100 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.635
+ $Y2=0
r102 57 59 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r103 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.575
+ $Y2=0
r104 56 59 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.04
+ $Y2=0
r105 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r106 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r107 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r108 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r109 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r110 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r111 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.16 $Y2=0
r112 48 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.635
+ $Y2=0
r113 48 54 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.08
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r115 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r118 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r119 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r120 43 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r121 41 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r124 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r125 36 55 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r126 36 52 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.16
+ $Y2=0
r127 32 79 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.497 $Y2=0
r128 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.515
r129 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0
r130 28 30 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0.625
r131 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=0.085
+ $X2=4.635 $Y2=0
r132 24 26 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.635 $Y=0.085
+ $X2=4.635 $Y2=0.415
r133 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r134 20 22 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.84
r135 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r136 16 18 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.84
r137 5 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.295
+ $Y=0.37 $X2=6.44 $Y2=0.515
r138 4 30 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.37 $X2=5.575 $Y2=0.625
r139 3 26 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.27 $X2=4.635 $Y2=0.415
r140 2 22 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.68 $X2=1.71 $Y2=0.84
r141 1 18 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.78 $Y2=0.84
.ends


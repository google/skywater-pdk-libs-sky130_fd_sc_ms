* File: sky130_fd_sc_ms__nor2_1.spice
* Created: Wed Sep  2 12:15:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor2_1.pex.spice"
.subckt sky130_fd_sc_ms__nor2_1  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_Y_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 A_119_368# N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g A_119_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.1344 PD=2.8 PS=1.36 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90000.6 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3852 P=7.36
c_96 A_119_368# 0 1.80995e-20 $X=0.595 $Y=1.84
*
.include "sky130_fd_sc_ms__nor2_1.pxi.spice"
*
.ends
*
*

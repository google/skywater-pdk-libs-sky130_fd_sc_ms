* File: sky130_fd_sc_ms__edfxtp_1.pxi.spice
* Created: Fri Aug 28 17:32:51 2020
* 
x_PM_SKY130_FD_SC_MS__EDFXTP_1%D N_D_M1008_g N_D_M1009_g D D N_D_c_262_n
+ N_D_c_263_n N_D_c_264_n N_D_c_268_n PM_SKY130_FD_SC_MS__EDFXTP_1%D
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_159_446# N_A_159_446#_M1010_s
+ N_A_159_446#_M1032_s N_A_159_446#_M1015_g N_A_159_446#_c_316_n
+ N_A_159_446#_M1021_g N_A_159_446#_c_317_n N_A_159_446#_c_318_n
+ N_A_159_446#_c_305_n N_A_159_446#_c_306_n N_A_159_446#_c_307_n
+ N_A_159_446#_c_335_n N_A_159_446#_c_308_n N_A_159_446#_c_309_n
+ N_A_159_446#_c_310_n N_A_159_446#_c_322_n N_A_159_446#_c_311_n
+ N_A_159_446#_c_312_n N_A_159_446#_c_313_n N_A_159_446#_c_314_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_159_446#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%DE N_DE_M1006_g N_DE_c_429_n N_DE_c_430_n
+ N_DE_c_431_n N_DE_c_432_n N_DE_M1010_g N_DE_c_438_n N_DE_M1032_g N_DE_c_439_n
+ N_DE_c_440_n N_DE_c_441_n N_DE_M1016_g N_DE_c_433_n DE N_DE_c_435_n
+ N_DE_c_436_n PM_SKY130_FD_SC_MS__EDFXTP_1%DE
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_533_61# N_A_533_61#_M1003_d N_A_533_61#_M1014_d
+ N_A_533_61#_M1022_g N_A_533_61#_M1027_g N_A_533_61#_c_517_n
+ N_A_533_61#_M1002_g N_A_533_61#_c_518_n N_A_533_61#_c_519_n
+ N_A_533_61#_M1000_g N_A_533_61#_c_531_n N_A_533_61#_c_532_n
+ N_A_533_61#_c_533_n N_A_533_61#_c_534_n N_A_533_61#_c_520_n
+ N_A_533_61#_c_535_n N_A_533_61#_c_521_n N_A_533_61#_c_522_n
+ N_A_533_61#_c_523_n N_A_533_61#_c_524_n N_A_533_61#_c_525_n
+ N_A_533_61#_c_526_n N_A_533_61#_c_527_n N_A_533_61#_c_528_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_533_61#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%CLK N_CLK_M1011_g N_CLK_c_713_n N_CLK_M1025_g CLK
+ N_CLK_c_716_n N_CLK_c_717_n PM_SKY130_FD_SC_MS__EDFXTP_1%CLK
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_958_74# N_A_958_74#_M1033_d N_A_958_74#_M1005_d
+ N_A_958_74#_M1013_g N_A_958_74#_c_753_n N_A_958_74#_M1028_g
+ N_A_958_74#_M1029_g N_A_958_74#_M1026_g N_A_958_74#_c_755_n
+ N_A_958_74#_c_756_n N_A_958_74#_c_757_n N_A_958_74#_c_778_n
+ N_A_958_74#_c_758_n N_A_958_74#_c_759_n N_A_958_74#_c_760_n
+ N_A_958_74#_c_761_n N_A_958_74#_c_847_p N_A_958_74#_c_762_n
+ N_A_958_74#_c_763_n N_A_958_74#_c_764_n N_A_958_74#_c_765_n
+ N_A_958_74#_c_766_n N_A_958_74#_c_767_n N_A_958_74#_c_768_n
+ N_A_958_74#_c_780_n N_A_958_74#_c_781_n N_A_958_74#_c_769_n
+ N_A_958_74#_c_770_n N_A_958_74#_c_771_n N_A_958_74#_c_772_n
+ N_A_958_74#_c_773_n N_A_958_74#_c_774_n N_A_958_74#_c_775_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_958_74#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_763_74# N_A_763_74#_M1011_d N_A_763_74#_M1025_d
+ N_A_763_74#_M1033_g N_A_763_74#_c_971_n N_A_763_74#_c_985_n
+ N_A_763_74#_M1005_g N_A_763_74#_M1024_g N_A_763_74#_c_973_n
+ N_A_763_74#_c_974_n N_A_763_74#_M1017_g N_A_763_74#_M1030_g
+ N_A_763_74#_M1007_g N_A_763_74#_c_976_n N_A_763_74#_c_977_n
+ N_A_763_74#_c_978_n N_A_763_74#_c_979_n N_A_763_74#_c_980_n
+ N_A_763_74#_c_993_n N_A_763_74#_c_994_n N_A_763_74#_c_981_n
+ N_A_763_74#_c_995_n N_A_763_74#_c_996_n N_A_763_74#_c_982_n
+ N_A_763_74#_c_983_n N_A_763_74#_c_999_n N_A_763_74#_c_1000_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_763_74#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_1409_64# N_A_1409_64#_M1004_d
+ N_A_1409_64#_M1023_d N_A_1409_64#_M1001_g N_A_1409_64#_M1020_g
+ N_A_1409_64#_M1018_g N_A_1409_64#_M1012_g N_A_1409_64#_c_1158_n
+ N_A_1409_64#_c_1159_n N_A_1409_64#_c_1160_n N_A_1409_64#_c_1161_n
+ N_A_1409_64#_c_1167_n N_A_1409_64#_c_1162_n N_A_1409_64#_c_1163_n
+ N_A_1409_64#_c_1177_n N_A_1409_64#_c_1178_n N_A_1409_64#_c_1164_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_1409_64#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_1156_90# N_A_1156_90#_M1024_d
+ N_A_1156_90#_M1013_d N_A_1156_90#_M1004_g N_A_1156_90#_M1023_g
+ N_A_1156_90#_c_1257_n N_A_1156_90#_c_1285_n N_A_1156_90#_c_1262_n
+ N_A_1156_90#_c_1263_n N_A_1156_90#_c_1264_n N_A_1156_90#_c_1258_n
+ N_A_1156_90#_c_1259_n N_A_1156_90#_c_1260_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_1156_90#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_1895_74# N_A_1895_74#_M1029_d
+ N_A_1895_74#_M1030_d N_A_1895_74#_M1003_g N_A_1895_74#_M1014_g
+ N_A_1895_74#_c_1355_n N_A_1895_74#_c_1356_n N_A_1895_74#_M1019_g
+ N_A_1895_74#_M1031_g N_A_1895_74#_c_1358_n N_A_1895_74#_c_1359_n
+ N_A_1895_74#_c_1360_n N_A_1895_74#_c_1422_n N_A_1895_74#_c_1367_n
+ N_A_1895_74#_c_1368_n N_A_1895_74#_c_1369_n N_A_1895_74#_c_1361_n
+ N_A_1895_74#_c_1362_n N_A_1895_74#_c_1363_n N_A_1895_74#_c_1364_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%A_1895_74#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%A_27_508# N_A_27_508#_M1009_s N_A_27_508#_M1022_d
+ N_A_27_508#_M1024_s N_A_27_508#_M1008_s N_A_27_508#_M1027_d
+ N_A_27_508#_M1013_s N_A_27_508#_c_1481_n N_A_27_508#_c_1488_n
+ N_A_27_508#_c_1489_n N_A_27_508#_c_1490_n N_A_27_508#_c_1491_n
+ N_A_27_508#_c_1492_n N_A_27_508#_c_1493_n N_A_27_508#_c_1494_n
+ N_A_27_508#_c_1495_n N_A_27_508#_c_1482_n N_A_27_508#_c_1497_n
+ N_A_27_508#_c_1498_n N_A_27_508#_c_1483_n N_A_27_508#_c_1484_n
+ N_A_27_508#_c_1499_n N_A_27_508#_c_1564_n N_A_27_508#_c_1500_n
+ N_A_27_508#_c_1485_n N_A_27_508#_c_1501_n N_A_27_508#_c_1486_n
+ N_A_27_508#_c_1502_n PM_SKY130_FD_SC_MS__EDFXTP_1%A_27_508#
x_PM_SKY130_FD_SC_MS__EDFXTP_1%VPWR N_VPWR_M1015_d N_VPWR_M1032_d N_VPWR_M1025_s
+ N_VPWR_M1005_s N_VPWR_M1020_d N_VPWR_M1018_s N_VPWR_M1000_d N_VPWR_M1031_d
+ N_VPWR_c_1654_n N_VPWR_c_1655_n N_VPWR_c_1656_n N_VPWR_c_1657_n
+ N_VPWR_c_1658_n N_VPWR_c_1659_n N_VPWR_c_1660_n N_VPWR_c_1661_n
+ N_VPWR_c_1662_n N_VPWR_c_1663_n N_VPWR_c_1664_n N_VPWR_c_1665_n
+ N_VPWR_c_1666_n N_VPWR_c_1667_n N_VPWR_c_1668_n N_VPWR_c_1669_n
+ N_VPWR_c_1670_n VPWR N_VPWR_c_1671_n N_VPWR_c_1672_n N_VPWR_c_1673_n
+ N_VPWR_c_1674_n N_VPWR_c_1675_n N_VPWR_c_1676_n N_VPWR_c_1677_n
+ N_VPWR_c_1653_n PM_SKY130_FD_SC_MS__EDFXTP_1%VPWR
x_PM_SKY130_FD_SC_MS__EDFXTP_1%Q N_Q_M1019_s N_Q_M1031_s N_Q_c_1791_n
+ N_Q_c_1792_n Q Q Q Q N_Q_c_1794_n Q PM_SKY130_FD_SC_MS__EDFXTP_1%Q
x_PM_SKY130_FD_SC_MS__EDFXTP_1%VGND N_VGND_M1006_d N_VGND_M1010_d N_VGND_M1011_s
+ N_VGND_M1033_s N_VGND_M1001_d N_VGND_M1012_s N_VGND_M1002_d N_VGND_M1019_d
+ N_VGND_c_1819_n N_VGND_c_1820_n N_VGND_c_1821_n N_VGND_c_1822_n
+ N_VGND_c_1823_n N_VGND_c_1824_n N_VGND_c_1825_n N_VGND_c_1826_n
+ N_VGND_c_1827_n N_VGND_c_1828_n N_VGND_c_1829_n N_VGND_c_1830_n
+ N_VGND_c_1831_n N_VGND_c_1832_n VGND N_VGND_c_1833_n N_VGND_c_1834_n
+ N_VGND_c_1835_n N_VGND_c_1836_n N_VGND_c_1837_n N_VGND_c_1838_n
+ N_VGND_c_1839_n N_VGND_c_1840_n N_VGND_c_1841_n N_VGND_c_1842_n
+ PM_SKY130_FD_SC_MS__EDFXTP_1%VGND
cc_1 VNB N_D_M1009_g 0.025709f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.58
cc_2 VNB N_D_c_262_n 0.0171113f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_3 VNB N_D_c_263_n 0.0117045f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_4 VNB N_D_c_264_n 0.0399559f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_5 VNB N_A_159_446#_M1021_g 0.0386628f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_6 VNB N_A_159_446#_c_305_n 0.00331491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_159_446#_c_306_n 0.0273265f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.665
cc_8 VNB N_A_159_446#_c_307_n 0.00951957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_159_446#_c_308_n 0.00319209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_159_446#_c_309_n 3.2668e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_159_446#_c_310_n 0.00674726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_159_446#_c_311_n 0.0029594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_159_446#_c_312_n 6.37728e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_159_446#_c_313_n 0.0037051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_159_446#_c_314_n 0.0279463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_DE_M1006_g 0.0227548f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_17 VNB N_DE_c_429_n 0.0256476f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.98
cc_18 VNB N_DE_c_430_n 0.0101882f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.58
cc_19 VNB N_DE_c_431_n 0.0115035f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.98
cc_20 VNB N_DE_c_432_n 0.0166758f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_DE_c_433_n 0.0236907f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_22 VNB DE 0.00159289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_DE_c_435_n 0.0148266f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.825
cc_24 VNB N_DE_c_436_n 0.0176647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_533_61#_M1022_g 0.0228356f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_26 VNB N_A_533_61#_c_517_n 0.0182482f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_27 VNB N_A_533_61#_c_518_n 0.0406862f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_28 VNB N_A_533_61#_c_519_n 0.00732576f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_29 VNB N_A_533_61#_c_520_n 0.0108941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_533_61#_c_521_n 0.028351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_533_61#_c_522_n 0.00306562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_533_61#_c_523_n 0.00462585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_533_61#_c_524_n 0.0036769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_533_61#_c_525_n 0.0603477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_533_61#_c_526_n 0.010322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_533_61#_c_527_n 0.0325649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_533_61#_c_528_n 0.010666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_CLK_c_713_n 0.0235908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_CLK_M1025_g 0.00191101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB CLK 0.00749125f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.98
cc_41 VNB N_CLK_c_716_n 0.0403775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_CLK_c_717_n 0.0204272f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_43 VNB N_A_958_74#_c_753_n 0.0184494f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_44 VNB N_A_958_74#_M1026_g 0.00355316f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_45 VNB N_A_958_74#_c_755_n 0.00945287f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.145
cc_46 VNB N_A_958_74#_c_756_n 0.0195832f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_47 VNB N_A_958_74#_c_757_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_958_74#_c_758_n 0.0134814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_958_74#_c_759_n 0.0210336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_958_74#_c_760_n 0.00189334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_958_74#_c_761_n 0.012232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_958_74#_c_762_n 0.0177357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_958_74#_c_763_n 0.00257567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_958_74#_c_764_n 0.011221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_958_74#_c_765_n 0.0049927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_958_74#_c_766_n 0.00315025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_958_74#_c_767_n 0.0115318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_958_74#_c_768_n 0.00145761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_958_74#_c_769_n 0.0357913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_958_74#_c_770_n 0.00837626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_958_74#_c_771_n 0.00984652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_958_74#_c_772_n 0.0355682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_958_74#_c_773_n 0.00360052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_958_74#_c_774_n 0.0305607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_958_74#_c_775_n 0.0188906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_763_74#_M1033_g 0.039916f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_67 VNB N_A_763_74#_c_971_n 0.0163226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_763_74#_M1024_g 0.060147f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_69 VNB N_A_763_74#_c_973_n 0.0447281f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_70 VNB N_A_763_74#_c_974_n 0.0127566f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.145
cc_71 VNB N_A_763_74#_M1007_g 0.0523977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_763_74#_c_976_n 0.00710918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_763_74#_c_977_n 0.00706889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_763_74#_c_978_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_763_74#_c_979_n 0.0118574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_763_74#_c_980_n 0.0182436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_763_74#_c_981_n 0.00148024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_763_74#_c_982_n 0.00381083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_763_74#_c_983_n 0.0178679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1409_64#_M1001_g 0.0291657f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_81 VNB N_A_1409_64#_M1020_g 0.00834433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1409_64#_M1018_g 0.00468362f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_83 VNB N_A_1409_64#_M1012_g 0.0269585f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_84 VNB N_A_1409_64#_c_1158_n 0.0548296f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.145
cc_85 VNB N_A_1409_64#_c_1159_n 0.0136506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1409_64#_c_1160_n 0.00646005f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_87 VNB N_A_1409_64#_c_1161_n 0.00782438f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.825
cc_88 VNB N_A_1409_64#_c_1162_n 0.00102187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1409_64#_c_1163_n 0.0127351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1409_64#_c_1164_n 0.0452693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1156_90#_M1004_g 0.0366237f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_92 VNB N_A_1156_90#_c_1257_n 0.02004f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_93 VNB N_A_1156_90#_c_1258_n 3.83683e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1156_90#_c_1259_n 0.0135877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1156_90#_c_1260_n 0.00354447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1895_74#_M1003_g 0.0293184f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_97 VNB N_A_1895_74#_M1014_g 0.0216858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1895_74#_c_1355_n 0.0559245f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_99 VNB N_A_1895_74#_c_1356_n 0.0215641f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_100 VNB N_A_1895_74#_M1031_g 0.0295f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_101 VNB N_A_1895_74#_c_1358_n 0.015548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1895_74#_c_1359_n 0.00329363f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.665
cc_103 VNB N_A_1895_74#_c_1360_n 0.0109396f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.825
cc_104 VNB N_A_1895_74#_c_1361_n 0.00243682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1895_74#_c_1362_n 0.00510635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1895_74#_c_1363_n 0.0384052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1895_74#_c_1364_n 0.0106154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_27_508#_c_1481_n 0.0404044f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_109 VNB N_A_27_508#_c_1482_n 0.00984382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_27_508#_c_1483_n 0.00828722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_27_508#_c_1484_n 0.0125822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_27_508#_c_1485_n 0.0297869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_27_508#_c_1486_n 0.013391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VPWR_c_1653_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_Q_c_1791_n 0.00764267f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_116 VNB N_Q_c_1792_n 0.0018251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB Q 0.00236984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_Q_c_1794_n 0.00432377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1819_n 0.00867737f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.665
cc_120 VNB N_VGND_c_1820_n 0.0111489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1821_n 0.00989189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1822_n 0.018697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1823_n 0.00789365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1824_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1825_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1826_n 0.0546602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1827_n 0.0319647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1828_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1829_n 0.0614466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1830_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1831_n 0.0298174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1832_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1833_n 0.0309056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1834_n 0.0189154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1835_n 0.020445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1836_n 0.0328797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1837_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1838_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1839_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1840_n 0.0444719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1841_n 0.0314426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1842_n 0.729984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VPB N_D_M1008_g 0.0510438f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_144 VPB N_D_c_263_n 0.00411548f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_145 VPB N_D_c_264_n 0.0118292f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_146 VPB N_D_c_268_n 0.0160786f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_147 VPB N_A_159_446#_M1015_g 0.0240866f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_148 VPB N_A_159_446#_c_316_n 0.0144439f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_149 VPB N_A_159_446#_c_317_n 0.0201231f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_150 VPB N_A_159_446#_c_318_n 0.0159417f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_151 VPB N_A_159_446#_c_306_n 0.0119695f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_152 VPB N_A_159_446#_c_308_n 0.00744243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_159_446#_c_309_n 0.00580517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_159_446#_c_322_n 0.00731159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_159_446#_c_311_n 0.00185815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_159_446#_c_313_n 0.00251827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_159_446#_c_314_n 0.00894816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_DE_c_431_n 0.0177427f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.98
cc_159 VPB N_DE_c_438_n 0.0192314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_DE_c_439_n 0.0328522f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_161 VPB N_DE_c_440_n 0.0270321f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_162 VPB N_DE_c_441_n 0.0173698f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_163 VPB N_A_533_61#_M1027_g 0.0494915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_533_61#_M1000_g 0.0224592f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_165 VPB N_A_533_61#_c_531_n 0.00967562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_533_61#_c_532_n 0.031501f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.825
cc_167 VPB N_A_533_61#_c_533_n 0.00836297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_533_61#_c_534_n 0.0100587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_533_61#_c_535_n 0.00354939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_533_61#_c_521_n 0.0654153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_533_61#_c_522_n 0.00294976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_533_61#_c_523_n 0.00262327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_533_61#_c_524_n 2.54227e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_533_61#_c_525_n 0.01285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_533_61#_c_526_n 0.00287546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_533_61#_c_527_n 0.0205345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_CLK_M1025_g 0.0291232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_958_74#_M1013_g 0.031737f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_179 VPB N_A_958_74#_M1026_g 0.0586496f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_180 VPB N_A_958_74#_c_778_n 0.00227852f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_181 VPB N_A_958_74#_c_758_n 0.00158825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_958_74#_c_780_n 0.00860942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_958_74#_c_781_n 0.0477078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_763_74#_c_971_n 0.010671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_763_74#_c_985_n 0.024314f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_186 VPB N_A_763_74#_c_973_n 0.0246448f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_187 VPB N_A_763_74#_c_974_n 0.00987168f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.145
cc_188 VPB N_A_763_74#_M1017_g 0.0256211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_763_74#_M1030_g 0.0293264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_763_74#_c_978_n 0.00340096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_763_74#_c_979_n 0.0050397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_763_74#_c_980_n 0.00533717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_763_74#_c_993_n 0.0140888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_763_74#_c_994_n 0.00339591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_763_74#_c_995_n 0.00876936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_763_74#_c_996_n 0.0331617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_763_74#_c_982_n 0.00165135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_763_74#_c_983_n 0.0159061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_763_74#_c_999_n 0.0376682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_763_74#_c_1000_n 0.0165753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1409_64#_M1020_g 0.064814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1409_64#_M1018_g 0.0420119f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_203 VPB N_A_1409_64#_c_1167_n 0.00519453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1409_64#_c_1162_n 0.0100339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_1156_90#_M1023_g 0.0246147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1156_90#_c_1262_n 0.00333807f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.145
cc_207 VPB N_A_1156_90#_c_1263_n 0.00684953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1156_90#_c_1264_n 0.00900679f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.825
cc_209 VPB N_A_1156_90#_c_1258_n 0.00167199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1156_90#_c_1259_n 0.0203348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1156_90#_c_1260_n 0.0121922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1895_74#_M1014_g 0.0575485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1895_74#_M1031_g 0.0338686f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_214 VPB N_A_1895_74#_c_1367_n 0.00725775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1895_74#_c_1368_n 0.0104845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1895_74#_c_1369_n 0.00679115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1895_74#_c_1361_n 0.00116664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_27_508#_c_1481_n 0.0244832f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_219 VPB N_A_27_508#_c_1488_n 0.0281836f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.145
cc_220 VPB N_A_27_508#_c_1489_n 0.0279518f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.295
cc_221 VPB N_A_27_508#_c_1490_n 0.0120405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_27_508#_c_1491_n 0.0168821f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.825
cc_223 VPB N_A_27_508#_c_1492_n 0.00348146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_27_508#_c_1493_n 0.00145547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_27_508#_c_1494_n 0.0212414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_27_508#_c_1495_n 0.00113173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_27_508#_c_1482_n 0.00831197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_27_508#_c_1497_n 0.0290649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_27_508#_c_1498_n 0.00161349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_27_508#_c_1499_n 0.00891819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_27_508#_c_1500_n 0.00660873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_27_508#_c_1501_n 0.0124532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_27_508#_c_1502_n 0.0153432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1654_n 0.00746943f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_235 VPB N_VPWR_c_1655_n 0.0241365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1656_n 0.0238553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1657_n 0.0243513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1658_n 0.0100759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1659_n 0.0124616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1660_n 0.011136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1661_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1662_n 0.0649725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1663_n 0.0293385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1664_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1665_n 0.0298174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1666_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1667_n 0.0314345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1668_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1669_n 0.0215854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1670_n 0.00612665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1671_n 0.0323948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1672_n 0.0590477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1673_n 0.0583199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1674_n 0.033781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1675_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1676_n 0.00613589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1677_n 0.0103609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1653_n 0.188771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB Q 0.0149243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 N_D_M1008_g N_A_159_446#_c_317_n 0.0525811f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_261 N_D_M1008_g N_A_159_446#_c_318_n 0.00843883f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_262 N_D_c_268_n N_A_159_446#_c_318_n 0.0137702f $X=0.52 $Y=1.99 $X2=0 $Y2=0
cc_263 N_D_M1009_g N_A_159_446#_c_305_n 2.08437e-19 $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_264 N_D_c_262_n N_A_159_446#_c_305_n 0.00142126f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_265 N_D_c_263_n N_A_159_446#_c_305_n 0.0513743f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_266 N_D_c_264_n N_A_159_446#_c_305_n 2.79757e-19 $X=0.52 $Y=1.825 $X2=0 $Y2=0
cc_267 N_D_c_263_n N_A_159_446#_c_306_n 0.00320031f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_268 N_D_c_264_n N_A_159_446#_c_306_n 0.0137702f $X=0.52 $Y=1.825 $X2=0 $Y2=0
cc_269 N_D_M1009_g N_A_159_446#_c_335_n 8.2231e-19 $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_270 N_D_c_263_n N_A_159_446#_c_309_n 0.0312709f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_271 N_D_c_264_n N_A_159_446#_c_309_n 3.92359e-19 $X=0.52 $Y=1.825 $X2=0 $Y2=0
cc_272 N_D_M1009_g N_DE_M1006_g 0.0377085f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_273 N_D_c_262_n N_DE_c_430_n 0.00787042f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_274 N_D_c_263_n N_DE_c_430_n 8.91711e-19 $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_275 N_D_M1008_g N_A_27_508#_c_1481_n 0.00675092f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_276 N_D_M1009_g N_A_27_508#_c_1481_n 0.0053259f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_277 N_D_c_262_n N_A_27_508#_c_1481_n 0.0245541f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_278 N_D_c_263_n N_A_27_508#_c_1481_n 0.0766518f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_279 N_D_M1008_g N_A_27_508#_c_1488_n 0.0165077f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_280 N_D_M1008_g N_A_27_508#_c_1489_n 0.01291f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_281 N_D_c_263_n N_A_27_508#_c_1489_n 0.0270499f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_282 N_D_c_268_n N_A_27_508#_c_1489_n 6.79407e-19 $X=0.52 $Y=1.99 $X2=0 $Y2=0
cc_283 N_D_M1009_g N_A_27_508#_c_1485_n 0.0103351f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_284 N_D_c_262_n N_A_27_508#_c_1485_n 0.00386592f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_285 N_D_c_263_n N_A_27_508#_c_1485_n 0.00885856f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_286 N_D_M1008_g N_A_27_508#_c_1501_n 0.00518121f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_287 N_D_c_263_n N_A_27_508#_c_1501_n 6.96185e-19 $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_288 N_D_c_268_n N_A_27_508#_c_1501_n 0.00236763f $X=0.52 $Y=1.99 $X2=0 $Y2=0
cc_289 N_D_M1008_g N_VPWR_c_1654_n 0.00180811f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_290 N_D_M1008_g N_VPWR_c_1663_n 0.005209f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_291 N_D_M1008_g N_VPWR_c_1653_n 0.00986576f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_292 N_D_M1009_g N_VGND_c_1819_n 0.00124923f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_293 N_D_M1009_g N_VGND_c_1833_n 0.00432935f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_294 N_D_M1009_g N_VGND_c_1842_n 0.00821075f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_295 N_A_159_446#_c_305_n N_DE_M1006_g 3.25298e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_296 N_A_159_446#_c_335_n N_DE_M1006_g 0.0092911f $X=1.305 $Y=0.855 $X2=0
+ $Y2=0
cc_297 N_A_159_446#_c_310_n N_DE_M1006_g 0.00290865f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_298 N_A_159_446#_c_305_n N_DE_c_429_n 0.0164959f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_299 N_A_159_446#_c_307_n N_DE_c_429_n 0.0078387f $X=1.57 $Y=0.855 $X2=0 $Y2=0
cc_300 N_A_159_446#_c_308_n N_DE_c_429_n 0.00330448f $X=1.705 $Y=1.695 $X2=0
+ $Y2=0
cc_301 N_A_159_446#_c_305_n N_DE_c_430_n 0.00292959f $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_302 N_A_159_446#_c_306_n N_DE_c_430_n 0.0182201f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_303 N_A_159_446#_c_305_n N_DE_c_431_n 9.98266e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_304 N_A_159_446#_c_306_n N_DE_c_431_n 0.0094379f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_305 N_A_159_446#_c_308_n N_DE_c_431_n 0.00510837f $X=1.705 $Y=1.695 $X2=0
+ $Y2=0
cc_306 N_A_159_446#_c_309_n N_DE_c_431_n 9.01876e-19 $X=1.305 $Y=1.695 $X2=0
+ $Y2=0
cc_307 N_A_159_446#_c_322_n N_DE_c_431_n 0.00622022f $X=1.79 $Y=2.495 $X2=0
+ $Y2=0
cc_308 N_A_159_446#_c_312_n N_DE_c_431_n 0.00563344f $X=1.79 $Y=1.695 $X2=0
+ $Y2=0
cc_309 N_A_159_446#_c_313_n N_DE_c_431_n 0.00145247f $X=2.22 $Y=1.55 $X2=0 $Y2=0
cc_310 N_A_159_446#_c_314_n N_DE_c_431_n 0.0154054f $X=2.38 $Y=1.55 $X2=0 $Y2=0
cc_311 N_A_159_446#_M1021_g N_DE_c_432_n 0.0199563f $X=2.38 $Y=0.645 $X2=0 $Y2=0
cc_312 N_A_159_446#_c_305_n N_DE_c_432_n 2.20134e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_313 N_A_159_446#_c_307_n N_DE_c_432_n 0.00377761f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_314 N_A_159_446#_c_310_n N_DE_c_432_n 7.31217e-19 $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_315 N_A_159_446#_c_322_n N_DE_c_438_n 0.0050064f $X=1.79 $Y=2.495 $X2=0 $Y2=0
cc_316 N_A_159_446#_c_316_n N_DE_c_440_n 0.00250929f $X=1.05 $Y=2.23 $X2=0 $Y2=0
cc_317 N_A_159_446#_c_318_n N_DE_c_440_n 0.0094379f $X=1.14 $Y=2.01 $X2=0 $Y2=0
cc_318 N_A_159_446#_c_322_n N_DE_c_440_n 0.0116006f $X=1.79 $Y=2.495 $X2=0 $Y2=0
cc_319 N_A_159_446#_c_311_n N_DE_c_440_n 0.00670782f $X=2.055 $Y=1.695 $X2=0
+ $Y2=0
cc_320 N_A_159_446#_c_313_n N_DE_c_440_n 0.00113269f $X=2.22 $Y=1.55 $X2=0 $Y2=0
cc_321 N_A_159_446#_c_314_n N_DE_c_440_n 0.022076f $X=2.38 $Y=1.55 $X2=0 $Y2=0
cc_322 N_A_159_446#_c_307_n N_DE_c_433_n 0.00681326f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_323 N_A_159_446#_c_311_n N_DE_c_433_n 0.00434828f $X=2.055 $Y=1.695 $X2=0
+ $Y2=0
cc_324 N_A_159_446#_c_312_n N_DE_c_433_n 0.00101655f $X=1.79 $Y=1.695 $X2=0
+ $Y2=0
cc_325 N_A_159_446#_M1021_g DE 0.00150886f $X=2.38 $Y=0.645 $X2=0 $Y2=0
cc_326 N_A_159_446#_c_305_n DE 0.0218472f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_327 N_A_159_446#_c_306_n DE 3.48291e-19 $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_328 N_A_159_446#_c_307_n DE 0.0247809f $X=1.57 $Y=0.855 $X2=0 $Y2=0
cc_329 N_A_159_446#_c_308_n DE 0.014091f $X=1.705 $Y=1.695 $X2=0 $Y2=0
cc_330 N_A_159_446#_c_312_n DE 0.0112841f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_331 N_A_159_446#_c_313_n DE 0.00348554f $X=2.22 $Y=1.55 $X2=0 $Y2=0
cc_332 N_A_159_446#_M1021_g N_DE_c_435_n 0.00817197f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_333 N_A_159_446#_c_305_n N_DE_c_435_n 0.00546415f $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_334 N_A_159_446#_c_305_n N_DE_c_436_n 3.48291e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_335 N_A_159_446#_c_306_n N_DE_c_436_n 0.00609406f $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_336 N_A_159_446#_c_308_n N_DE_c_436_n 0.00104323f $X=1.705 $Y=1.695 $X2=0
+ $Y2=0
cc_337 N_A_159_446#_c_314_n N_DE_c_436_n 0.0034012f $X=2.38 $Y=1.55 $X2=0 $Y2=0
cc_338 N_A_159_446#_M1021_g N_A_533_61#_M1022_g 0.0421816f $X=2.38 $Y=0.645
+ $X2=0 $Y2=0
cc_339 N_A_159_446#_c_313_n N_A_533_61#_c_522_n 0.00774583f $X=2.22 $Y=1.55
+ $X2=0 $Y2=0
cc_340 N_A_159_446#_c_314_n N_A_533_61#_c_522_n 0.00333561f $X=2.38 $Y=1.55
+ $X2=0 $Y2=0
cc_341 N_A_159_446#_c_313_n N_A_533_61#_c_525_n 2.95947e-19 $X=2.22 $Y=1.55
+ $X2=0 $Y2=0
cc_342 N_A_159_446#_c_314_n N_A_533_61#_c_525_n 0.0421816f $X=2.38 $Y=1.55 $X2=0
+ $Y2=0
cc_343 N_A_159_446#_M1021_g N_A_533_61#_c_526_n 0.0107379f $X=2.38 $Y=0.645
+ $X2=0 $Y2=0
cc_344 N_A_159_446#_c_313_n N_A_533_61#_c_526_n 0.0285435f $X=2.22 $Y=1.55 $X2=0
+ $Y2=0
cc_345 N_A_159_446#_c_317_n N_A_27_508#_c_1488_n 0.00208077f $X=1.05 $Y=2.305
+ $X2=0 $Y2=0
cc_346 N_A_159_446#_c_316_n N_A_27_508#_c_1489_n 0.00448415f $X=1.05 $Y=2.23
+ $X2=0 $Y2=0
cc_347 N_A_159_446#_c_317_n N_A_27_508#_c_1489_n 0.0179837f $X=1.05 $Y=2.305
+ $X2=0 $Y2=0
cc_348 N_A_159_446#_c_318_n N_A_27_508#_c_1489_n 0.00125351f $X=1.14 $Y=2.01
+ $X2=0 $Y2=0
cc_349 N_A_159_446#_c_308_n N_A_27_508#_c_1489_n 0.0103913f $X=1.705 $Y=1.695
+ $X2=0 $Y2=0
cc_350 N_A_159_446#_c_309_n N_A_27_508#_c_1489_n 0.0258112f $X=1.305 $Y=1.695
+ $X2=0 $Y2=0
cc_351 N_A_159_446#_c_322_n N_A_27_508#_c_1489_n 0.0141315f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_352 N_A_159_446#_M1015_g N_A_27_508#_c_1490_n 0.00451709f $X=0.885 $Y=2.75
+ $X2=0 $Y2=0
cc_353 N_A_159_446#_c_317_n N_A_27_508#_c_1490_n 0.00102928f $X=1.05 $Y=2.305
+ $X2=0 $Y2=0
cc_354 N_A_159_446#_c_322_n N_A_27_508#_c_1490_n 0.0284388f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_355 N_A_159_446#_c_322_n N_A_27_508#_c_1491_n 0.0127728f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_356 N_A_159_446#_M1015_g N_A_27_508#_c_1492_n 7.1147e-19 $X=0.885 $Y=2.75
+ $X2=0 $Y2=0
cc_357 N_A_159_446#_c_322_n N_A_27_508#_c_1493_n 0.0230284f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_358 N_A_159_446#_c_313_n N_A_27_508#_c_1494_n 0.013613f $X=2.22 $Y=1.55 $X2=0
+ $Y2=0
cc_359 N_A_159_446#_c_314_n N_A_27_508#_c_1494_n 0.00183975f $X=2.38 $Y=1.55
+ $X2=0 $Y2=0
cc_360 N_A_159_446#_c_322_n N_A_27_508#_c_1495_n 0.013005f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_361 N_A_159_446#_c_311_n N_A_27_508#_c_1495_n 8.44449e-19 $X=2.055 $Y=1.695
+ $X2=0 $Y2=0
cc_362 N_A_159_446#_c_313_n N_A_27_508#_c_1495_n 0.0143089f $X=2.22 $Y=1.55
+ $X2=0 $Y2=0
cc_363 N_A_159_446#_c_314_n N_A_27_508#_c_1495_n 5.27783e-19 $X=2.38 $Y=1.55
+ $X2=0 $Y2=0
cc_364 N_A_159_446#_c_335_n N_A_27_508#_c_1485_n 0.00145863f $X=1.305 $Y=0.855
+ $X2=0 $Y2=0
cc_365 N_A_159_446#_M1021_g N_A_27_508#_c_1486_n 0.00124492f $X=2.38 $Y=0.645
+ $X2=0 $Y2=0
cc_366 N_A_159_446#_M1015_g N_VPWR_c_1654_n 0.0146016f $X=0.885 $Y=2.75 $X2=0
+ $Y2=0
cc_367 N_A_159_446#_c_317_n N_VPWR_c_1654_n 0.00423427f $X=1.05 $Y=2.305 $X2=0
+ $Y2=0
cc_368 N_A_159_446#_M1015_g N_VPWR_c_1663_n 0.00460063f $X=0.885 $Y=2.75 $X2=0
+ $Y2=0
cc_369 N_A_159_446#_M1015_g N_VPWR_c_1653_n 0.00908061f $X=0.885 $Y=2.75 $X2=0
+ $Y2=0
cc_370 N_A_159_446#_c_335_n N_VGND_M1006_d 0.00220205f $X=1.305 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_371 N_A_159_446#_c_307_n N_VGND_c_1819_n 0.00351808f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_372 N_A_159_446#_c_335_n N_VGND_c_1819_n 0.0196647f $X=1.305 $Y=0.855 $X2=0
+ $Y2=0
cc_373 N_A_159_446#_c_310_n N_VGND_c_1819_n 0.0125975f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_374 N_A_159_446#_M1021_g N_VGND_c_1820_n 0.012473f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_375 N_A_159_446#_c_307_n N_VGND_c_1820_n 0.00463069f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_376 N_A_159_446#_c_310_n N_VGND_c_1820_n 0.0134516f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_377 N_A_159_446#_c_313_n N_VGND_c_1820_n 0.0101419f $X=2.22 $Y=1.55 $X2=0
+ $Y2=0
cc_378 N_A_159_446#_c_314_n N_VGND_c_1820_n 0.00165606f $X=2.38 $Y=1.55 $X2=0
+ $Y2=0
cc_379 N_A_159_446#_M1021_g N_VGND_c_1827_n 0.00441186f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_380 N_A_159_446#_c_310_n N_VGND_c_1834_n 0.00860429f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_381 N_A_159_446#_M1021_g N_VGND_c_1842_n 0.0044119f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_382 N_A_159_446#_c_307_n N_VGND_c_1842_n 0.00826433f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_383 N_A_159_446#_c_335_n N_VGND_c_1842_n 0.00271168f $X=1.305 $Y=0.855 $X2=0
+ $Y2=0
cc_384 N_A_159_446#_c_310_n N_VGND_c_1842_n 0.00870705f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_385 N_DE_c_439_n N_A_533_61#_M1027_g 0.0475288f $X=2.605 $Y=2.03 $X2=0 $Y2=0
cc_386 N_DE_c_439_n N_A_533_61#_c_525_n 0.00665363f $X=2.605 $Y=2.03 $X2=0 $Y2=0
cc_387 N_DE_c_439_n N_A_533_61#_c_526_n 0.00107062f $X=2.605 $Y=2.03 $X2=0 $Y2=0
cc_388 N_DE_c_438_n N_A_27_508#_c_1490_n 0.00358222f $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_389 N_DE_c_438_n N_A_27_508#_c_1491_n 0.0107712f $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_390 N_DE_c_438_n N_A_27_508#_c_1493_n 0.0215711f $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_391 N_DE_c_441_n N_A_27_508#_c_1493_n 0.00359987f $X=2.695 $Y=2.105 $X2=0
+ $Y2=0
cc_392 N_DE_c_439_n N_A_27_508#_c_1494_n 0.0172172f $X=2.605 $Y=2.03 $X2=0 $Y2=0
cc_393 N_DE_c_441_n N_A_27_508#_c_1494_n 0.00738909f $X=2.695 $Y=2.105 $X2=0
+ $Y2=0
cc_394 N_DE_c_438_n N_A_27_508#_c_1495_n 4.47919e-19 $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_395 N_DE_c_439_n N_A_27_508#_c_1495_n 0.0022419f $X=2.605 $Y=2.03 $X2=0 $Y2=0
cc_396 N_DE_c_440_n N_A_27_508#_c_1495_n 0.00325956f $X=2.105 $Y=2.03 $X2=0
+ $Y2=0
cc_397 N_DE_M1006_g N_A_27_508#_c_1485_n 0.00168095f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_398 N_DE_c_441_n N_A_27_508#_c_1502_n 0.00186935f $X=2.695 $Y=2.105 $X2=0
+ $Y2=0
cc_399 N_DE_c_438_n N_VPWR_c_1655_n 0.0025598f $X=2.015 $Y=2.105 $X2=0 $Y2=0
cc_400 N_DE_c_439_n N_VPWR_c_1655_n 9.92786e-19 $X=2.605 $Y=2.03 $X2=0 $Y2=0
cc_401 N_DE_c_441_n N_VPWR_c_1655_n 0.0103847f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_402 N_DE_c_438_n N_VPWR_c_1665_n 8.4712e-19 $X=2.015 $Y=2.105 $X2=0 $Y2=0
cc_403 N_DE_c_441_n N_VPWR_c_1667_n 0.00363301f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_404 N_DE_c_441_n N_VPWR_c_1653_n 0.00444302f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_405 N_DE_M1006_g N_VGND_c_1819_n 0.00953711f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_406 N_DE_c_429_n N_VGND_c_1819_n 9.9363e-19 $X=1.515 $Y=1.025 $X2=0 $Y2=0
cc_407 N_DE_c_432_n N_VGND_c_1819_n 0.00208085f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_408 N_DE_c_432_n N_VGND_c_1820_n 0.0111681f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_409 N_DE_M1006_g N_VGND_c_1833_n 0.00383152f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_410 N_DE_c_432_n N_VGND_c_1834_n 0.00441186f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_411 N_DE_M1006_g N_VGND_c_1842_n 0.00615424f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_412 N_DE_c_432_n N_VGND_c_1842_n 0.0044119f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_413 N_A_533_61#_c_521_n CLK 0.0167f $X=11.615 $Y=1.665 $X2=0 $Y2=0
cc_414 N_A_533_61#_c_525_n CLK 4.84099e-19 $X=2.83 $Y=1.21 $X2=0 $Y2=0
cc_415 N_A_533_61#_c_521_n N_CLK_c_716_n 0.00417411f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_416 N_A_533_61#_c_525_n N_CLK_c_716_n 0.0150512f $X=2.83 $Y=1.21 $X2=0 $Y2=0
cc_417 N_A_533_61#_c_525_n N_CLK_c_717_n 0.00337304f $X=2.83 $Y=1.21 $X2=0 $Y2=0
cc_418 N_A_533_61#_M1000_g N_A_958_74#_M1026_g 0.0373927f $X=10.785 $Y=2.72
+ $X2=0 $Y2=0
cc_419 N_A_533_61#_c_531_n N_A_958_74#_M1026_g 8.23648e-19 $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_420 N_A_533_61#_c_532_n N_A_958_74#_M1026_g 0.0204492f $X=10.83 $Y=2.185
+ $X2=0 $Y2=0
cc_421 N_A_533_61#_c_521_n N_A_958_74#_M1026_g 0.00564714f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_422 N_A_533_61#_c_527_n N_A_958_74#_M1026_g 0.0146467f $X=10.83 $Y=2.02 $X2=0
+ $Y2=0
cc_423 N_A_533_61#_c_521_n N_A_958_74#_c_755_n 0.00789556f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_424 N_A_533_61#_c_521_n N_A_958_74#_c_778_n 0.0140524f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_425 N_A_533_61#_c_521_n N_A_958_74#_c_758_n 0.0221532f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_426 N_A_533_61#_c_521_n N_A_958_74#_c_761_n 0.00423047f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_427 N_A_533_61#_c_521_n N_A_958_74#_c_765_n 0.00730168f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_428 N_A_533_61#_c_521_n N_A_958_74#_c_766_n 7.61262e-19 $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_429 N_A_533_61#_c_519_n N_A_958_74#_c_767_n 0.00130497f $X=10.375 $Y=0.94
+ $X2=0 $Y2=0
cc_430 N_A_533_61#_c_521_n N_A_958_74#_c_767_n 0.015916f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_431 N_A_533_61#_c_521_n N_A_958_74#_c_780_n 0.00761408f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_432 N_A_533_61#_c_521_n N_A_958_74#_c_769_n 0.00190225f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_433 N_A_533_61#_c_521_n N_A_958_74#_c_770_n 0.0098216f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_434 N_A_533_61#_c_521_n N_A_958_74#_c_771_n 0.01903f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_435 N_A_533_61#_c_521_n N_A_958_74#_c_772_n 0.00174952f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_436 N_A_533_61#_c_519_n N_A_958_74#_c_773_n 0.0019999f $X=10.375 $Y=0.94
+ $X2=0 $Y2=0
cc_437 N_A_533_61#_c_521_n N_A_958_74#_c_773_n 0.00931256f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_438 N_A_533_61#_c_527_n N_A_958_74#_c_773_n 7.22432e-19 $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_439 N_A_533_61#_c_519_n N_A_958_74#_c_774_n 0.017152f $X=10.375 $Y=0.94 $X2=0
+ $Y2=0
cc_440 N_A_533_61#_c_527_n N_A_958_74#_c_774_n 0.0205371f $X=10.83 $Y=2.02 $X2=0
+ $Y2=0
cc_441 N_A_533_61#_c_521_n N_A_763_74#_c_971_n 0.00466003f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_442 N_A_533_61#_c_521_n N_A_763_74#_c_985_n 0.00240649f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_443 N_A_533_61#_c_521_n N_A_763_74#_c_973_n 0.0172604f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_444 N_A_533_61#_c_521_n N_A_763_74#_c_974_n 0.00661656f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_445 N_A_533_61#_c_517_n N_A_763_74#_M1007_g 0.0406264f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_446 N_A_533_61#_c_521_n N_A_763_74#_c_978_n 0.0193665f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_447 N_A_533_61#_c_521_n N_A_763_74#_c_979_n 0.0523905f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_448 N_A_533_61#_c_521_n N_A_763_74#_c_994_n 0.00977116f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_449 N_A_533_61#_c_521_n N_A_763_74#_c_981_n 0.00551289f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_450 N_A_533_61#_c_521_n N_A_763_74#_c_995_n 0.00239393f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_451 N_A_533_61#_c_521_n N_A_763_74#_c_982_n 0.0217703f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_452 N_A_533_61#_c_521_n N_A_763_74#_c_983_n 0.00819353f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_453 N_A_533_61#_c_521_n N_A_1409_64#_M1020_g 0.00192057f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_454 N_A_533_61#_c_521_n N_A_1409_64#_M1018_g 0.0118048f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_455 N_A_533_61#_c_521_n N_A_1409_64#_c_1158_n 0.00379165f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_456 N_A_533_61#_c_521_n N_A_1409_64#_c_1159_n 7.57862e-19 $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_457 N_A_533_61#_c_521_n N_A_1409_64#_c_1160_n 0.0112543f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_458 N_A_533_61#_c_521_n N_A_1409_64#_c_1167_n 0.00666783f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_459 N_A_533_61#_c_521_n N_A_1409_64#_c_1162_n 0.0170068f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_460 N_A_533_61#_c_521_n N_A_1409_64#_c_1163_n 0.0135625f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_461 N_A_533_61#_c_521_n N_A_1409_64#_c_1177_n 0.0170777f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_462 N_A_533_61#_c_521_n N_A_1409_64#_c_1178_n 0.00784482f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_463 N_A_533_61#_c_521_n N_A_1409_64#_c_1164_n 0.0066297f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_464 N_A_533_61#_c_521_n N_A_1156_90#_c_1257_n 0.010891f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_465 N_A_533_61#_c_521_n N_A_1156_90#_c_1262_n 0.0151876f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_466 N_A_533_61#_c_521_n N_A_1156_90#_c_1264_n 0.00152612f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_467 N_A_533_61#_c_521_n N_A_1156_90#_c_1258_n 0.0186899f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_468 N_A_533_61#_c_521_n N_A_1156_90#_c_1259_n 0.00508221f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_469 N_A_533_61#_c_521_n N_A_1156_90#_c_1260_n 0.0554077f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_470 N_A_533_61#_c_518_n N_A_1895_74#_M1003_g 0.0054796f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_471 N_A_533_61#_c_520_n N_A_1895_74#_M1003_g 0.00230527f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_472 N_A_533_61#_c_528_n N_A_1895_74#_M1003_g 0.00646527f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_473 N_A_533_61#_M1000_g N_A_1895_74#_M1014_g 0.0124769f $X=10.785 $Y=2.72
+ $X2=0 $Y2=0
cc_474 N_A_533_61#_c_531_n N_A_1895_74#_M1014_g 0.0163634f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_475 N_A_533_61#_c_532_n N_A_1895_74#_M1014_g 0.00958672f $X=10.83 $Y=2.185
+ $X2=0 $Y2=0
cc_476 N_A_533_61#_c_533_n N_A_1895_74#_M1014_g 0.0102317f $X=11.72 $Y=2.435
+ $X2=0 $Y2=0
cc_477 N_A_533_61#_c_535_n N_A_1895_74#_M1014_g 0.00521104f $X=11.72 $Y=2.207
+ $X2=0 $Y2=0
cc_478 N_A_533_61#_c_521_n N_A_1895_74#_M1014_g 0.010206f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_479 N_A_533_61#_c_523_n N_A_1895_74#_M1014_g 0.00239059f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_480 N_A_533_61#_c_524_n N_A_1895_74#_M1014_g 0.0209862f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_481 N_A_533_61#_c_527_n N_A_1895_74#_M1014_g 0.0187228f $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_482 N_A_533_61#_c_528_n N_A_1895_74#_M1014_g 0.00816022f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_483 N_A_533_61#_c_520_n N_A_1895_74#_c_1355_n 0.00332519f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_484 N_A_533_61#_c_523_n N_A_1895_74#_c_1355_n 4.89582e-19 $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_485 N_A_533_61#_c_524_n N_A_1895_74#_c_1355_n 0.0012174f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_486 N_A_533_61#_c_528_n N_A_1895_74#_c_1355_n 0.0149104f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_487 N_A_533_61#_c_520_n N_A_1895_74#_c_1356_n 0.00180935f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_488 N_A_533_61#_c_533_n N_A_1895_74#_M1031_g 0.00104557f $X=11.72 $Y=2.435
+ $X2=0 $Y2=0
cc_489 N_A_533_61#_c_535_n N_A_1895_74#_M1031_g 4.79912e-19 $X=11.72 $Y=2.207
+ $X2=0 $Y2=0
cc_490 N_A_533_61#_c_524_n N_A_1895_74#_M1031_g 0.00135259f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_491 N_A_533_61#_c_517_n N_A_1895_74#_c_1360_n 0.00454092f $X=10.3 $Y=0.865
+ $X2=0 $Y2=0
cc_492 N_A_533_61#_c_518_n N_A_1895_74#_c_1360_n 0.0155364f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_493 N_A_533_61#_c_519_n N_A_1895_74#_c_1360_n 0.00422433f $X=10.375 $Y=0.94
+ $X2=0 $Y2=0
cc_494 N_A_533_61#_c_521_n N_A_1895_74#_c_1360_n 0.00541203f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_495 N_A_533_61#_c_531_n N_A_1895_74#_c_1367_n 0.00884557f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_496 N_A_533_61#_c_531_n N_A_1895_74#_c_1368_n 0.0202046f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_497 N_A_533_61#_c_532_n N_A_1895_74#_c_1368_n 0.00422279f $X=10.83 $Y=2.185
+ $X2=0 $Y2=0
cc_498 N_A_533_61#_c_521_n N_A_1895_74#_c_1368_n 0.0147772f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_499 N_A_533_61#_c_527_n N_A_1895_74#_c_1368_n 0.00941512f $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_500 N_A_533_61#_c_532_n N_A_1895_74#_c_1369_n 4.73647e-19 $X=10.83 $Y=2.185
+ $X2=0 $Y2=0
cc_501 N_A_533_61#_c_521_n N_A_1895_74#_c_1369_n 0.0124112f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_502 N_A_533_61#_c_527_n N_A_1895_74#_c_1369_n 5.07165e-19 $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_503 N_A_533_61#_c_521_n N_A_1895_74#_c_1361_n 0.0215477f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_504 N_A_533_61#_c_527_n N_A_1895_74#_c_1361_n 0.0132717f $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_505 N_A_533_61#_c_518_n N_A_1895_74#_c_1362_n 3.34269e-19 $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_506 N_A_533_61#_c_532_n N_A_1895_74#_c_1362_n 7.13955e-19 $X=10.83 $Y=2.185
+ $X2=0 $Y2=0
cc_507 N_A_533_61#_c_520_n N_A_1895_74#_c_1362_n 0.00103395f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_508 N_A_533_61#_c_521_n N_A_1895_74#_c_1362_n 0.0230881f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_509 N_A_533_61#_c_527_n N_A_1895_74#_c_1362_n 0.00376914f $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_510 N_A_533_61#_c_528_n N_A_1895_74#_c_1362_n 0.0256537f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_511 N_A_533_61#_c_518_n N_A_1895_74#_c_1363_n 0.0213762f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_512 N_A_533_61#_c_520_n N_A_1895_74#_c_1363_n 0.00396895f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_513 N_A_533_61#_c_521_n N_A_1895_74#_c_1363_n 0.00552909f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_514 N_A_533_61#_c_528_n N_A_1895_74#_c_1363_n 0.00465196f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_515 N_A_533_61#_c_518_n N_A_1895_74#_c_1364_n 0.00859599f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_516 N_A_533_61#_c_527_n N_A_1895_74#_c_1364_n 0.00762021f $X=10.83 $Y=2.02
+ $X2=0 $Y2=0
cc_517 N_A_533_61#_M1027_g N_A_27_508#_c_1494_n 0.00924014f $X=3.085 $Y=2.39
+ $X2=0 $Y2=0
cc_518 N_A_533_61#_c_521_n N_A_27_508#_c_1494_n 0.00761887f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_519 N_A_533_61#_c_522_n N_A_27_508#_c_1494_n 0.00466191f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_520 N_A_533_61#_c_525_n N_A_27_508#_c_1494_n 0.00316757f $X=2.83 $Y=1.21
+ $X2=0 $Y2=0
cc_521 N_A_533_61#_c_526_n N_A_27_508#_c_1494_n 0.0267574f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_522 N_A_533_61#_M1022_g N_A_27_508#_c_1482_n 0.00513151f $X=2.74 $Y=0.645
+ $X2=0 $Y2=0
cc_523 N_A_533_61#_M1027_g N_A_27_508#_c_1482_n 0.0122012f $X=3.085 $Y=2.39
+ $X2=0 $Y2=0
cc_524 N_A_533_61#_c_521_n N_A_27_508#_c_1482_n 0.0266392f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_533_61#_c_522_n N_A_27_508#_c_1482_n 4.40756e-19 $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_526 N_A_533_61#_c_525_n N_A_27_508#_c_1482_n 0.0205144f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_527 N_A_533_61#_c_526_n N_A_27_508#_c_1482_n 0.0519058f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_528 N_A_533_61#_c_521_n N_A_27_508#_c_1497_n 0.0250517f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_533_61#_c_521_n N_A_27_508#_c_1498_n 0.0133932f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_533_61#_c_521_n N_A_27_508#_c_1483_n 0.0194929f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_533_61#_c_521_n N_A_27_508#_c_1484_n 0.0020928f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_533_61#_c_521_n N_A_27_508#_c_1564_n 0.00301115f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_533_61#_M1022_g N_A_27_508#_c_1486_n 0.00946606f $X=2.74 $Y=0.645
+ $X2=0 $Y2=0
cc_534 N_A_533_61#_c_525_n N_A_27_508#_c_1486_n 0.0090921f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_535 N_A_533_61#_c_526_n N_A_27_508#_c_1486_n 0.0118563f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_536 N_A_533_61#_M1027_g N_A_27_508#_c_1502_n 0.0179192f $X=3.085 $Y=2.39
+ $X2=0 $Y2=0
cc_537 N_A_533_61#_c_521_n N_A_27_508#_c_1502_n 0.00808113f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_533_61#_c_531_n N_VPWR_M1000_d 0.00232385f $X=11.555 $Y=2.207 $X2=0
+ $Y2=0
cc_539 N_A_533_61#_M1027_g N_VPWR_c_1655_n 0.00141573f $X=3.085 $Y=2.39 $X2=0
+ $Y2=0
cc_540 N_A_533_61#_M1027_g N_VPWR_c_1656_n 0.00215112f $X=3.085 $Y=2.39 $X2=0
+ $Y2=0
cc_541 N_A_533_61#_M1000_g N_VPWR_c_1660_n 0.0210499f $X=10.785 $Y=2.72 $X2=0
+ $Y2=0
cc_542 N_A_533_61#_c_531_n N_VPWR_c_1660_n 0.0337659f $X=11.555 $Y=2.207 $X2=0
+ $Y2=0
cc_543 N_A_533_61#_c_532_n N_VPWR_c_1660_n 0.00299573f $X=10.83 $Y=2.185 $X2=0
+ $Y2=0
cc_544 N_A_533_61#_c_533_n N_VPWR_c_1660_n 0.0167985f $X=11.72 $Y=2.435 $X2=0
+ $Y2=0
cc_545 N_A_533_61#_M1027_g N_VPWR_c_1667_n 0.00398295f $X=3.085 $Y=2.39 $X2=0
+ $Y2=0
cc_546 N_A_533_61#_M1000_g N_VPWR_c_1673_n 0.00554681f $X=10.785 $Y=2.72 $X2=0
+ $Y2=0
cc_547 N_A_533_61#_c_533_n N_VPWR_c_1674_n 0.0129767f $X=11.72 $Y=2.435 $X2=0
+ $Y2=0
cc_548 N_A_533_61#_M1027_g N_VPWR_c_1653_n 0.00529631f $X=3.085 $Y=2.39 $X2=0
+ $Y2=0
cc_549 N_A_533_61#_M1000_g N_VPWR_c_1653_n 0.00539832f $X=10.785 $Y=2.72 $X2=0
+ $Y2=0
cc_550 N_A_533_61#_c_533_n N_VPWR_c_1653_n 0.0118673f $X=11.72 $Y=2.435 $X2=0
+ $Y2=0
cc_551 N_A_533_61#_c_520_n N_Q_c_1791_n 0.0319039f $X=11.62 $Y=0.57 $X2=0 $Y2=0
cc_552 N_A_533_61#_c_528_n N_Q_c_1792_n 0.0319039f $X=11.765 $Y=1.55 $X2=0 $Y2=0
cc_553 N_A_533_61#_c_533_n Q 0.0484729f $X=11.72 $Y=2.435 $X2=0 $Y2=0
cc_554 N_A_533_61#_c_534_n Q 0.0188962f $X=11.765 $Y=2.095 $X2=0 $Y2=0
cc_555 N_A_533_61#_c_535_n Q 0.018397f $X=11.72 $Y=2.207 $X2=0 $Y2=0
cc_556 N_A_533_61#_c_523_n Q 0.00740378f $X=11.76 $Y=1.665 $X2=0 $Y2=0
cc_557 N_A_533_61#_c_524_n Q 0.0188962f $X=11.76 $Y=1.665 $X2=0 $Y2=0
cc_558 N_A_533_61#_c_528_n N_Q_c_1794_n 0.0252426f $X=11.765 $Y=1.55 $X2=0 $Y2=0
cc_559 N_A_533_61#_M1022_g N_VGND_c_1820_n 0.00180764f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_560 N_A_533_61#_M1022_g N_VGND_c_1821_n 0.00309386f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_561 N_A_533_61#_c_521_n N_VGND_c_1821_n 6.4869e-19 $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_562 N_A_533_61#_c_521_n N_VGND_c_1822_n 0.00166402f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_563 N_A_533_61#_c_520_n N_VGND_c_1826_n 4.75821e-19 $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_564 N_A_533_61#_M1022_g N_VGND_c_1827_n 0.00506571f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_565 N_A_533_61#_c_520_n N_VGND_c_1836_n 0.0165341f $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_566 N_A_533_61#_c_517_n N_VGND_c_1840_n 0.00383152f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_567 N_A_533_61#_c_517_n N_VGND_c_1841_n 0.011715f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_568 N_A_533_61#_c_518_n N_VGND_c_1841_n 0.00459991f $X=10.815 $Y=0.94 $X2=0
+ $Y2=0
cc_569 N_A_533_61#_c_520_n N_VGND_c_1841_n 0.00290096f $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_570 N_A_533_61#_M1022_g N_VGND_c_1842_n 0.00525227f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_571 N_A_533_61#_c_517_n N_VGND_c_1842_n 0.00380989f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_572 N_A_533_61#_c_520_n N_VGND_c_1842_n 0.013075f $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_573 N_CLK_c_713_n N_A_763_74#_M1033_g 0.00202801f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_574 N_CLK_c_717_n N_A_763_74#_c_976_n 0.0064177f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_575 N_CLK_c_713_n N_A_763_74#_c_977_n 0.00730881f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_576 CLK N_A_763_74#_c_977_n 0.0214612f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_577 N_CLK_c_717_n N_A_763_74#_c_977_n 0.00934401f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_578 N_CLK_c_713_n N_A_763_74#_c_978_n 0.00287369f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_579 N_CLK_M1025_g N_A_763_74#_c_978_n 0.0188895f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_580 CLK N_A_763_74#_c_978_n 0.00638598f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_581 N_CLK_c_713_n N_A_763_74#_c_979_n 0.00277002f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_582 N_CLK_M1025_g N_A_763_74#_c_979_n 0.00528842f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_583 N_CLK_c_713_n N_A_763_74#_c_980_n 0.00624738f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_584 N_CLK_c_713_n N_A_763_74#_c_981_n 0.00326043f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_585 N_CLK_c_717_n N_A_763_74#_c_981_n 0.00239841f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_586 N_CLK_M1025_g N_A_763_74#_c_999_n 0.00624738f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_587 CLK N_A_27_508#_c_1482_n 0.0268019f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_588 N_CLK_c_716_n N_A_27_508#_c_1482_n 0.00214569f $X=3.615 $Y=1.385 $X2=0
+ $Y2=0
cc_589 N_CLK_c_717_n N_A_27_508#_c_1482_n 0.00316008f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_590 N_CLK_M1025_g N_A_27_508#_c_1497_n 0.0173042f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_591 N_CLK_M1025_g N_A_27_508#_c_1502_n 0.00859351f $X=4.06 $Y=2.32 $X2=0
+ $Y2=0
cc_592 CLK N_A_27_508#_c_1502_n 3.50421e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_593 N_CLK_M1025_g N_VPWR_c_1656_n 0.0195245f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_594 N_CLK_M1025_g N_VPWR_c_1671_n 0.00519349f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_595 N_CLK_M1025_g N_VPWR_c_1653_n 0.00524044f $X=4.06 $Y=2.32 $X2=0 $Y2=0
cc_596 CLK N_VGND_c_1821_n 0.0134779f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_597 N_CLK_c_716_n N_VGND_c_1821_n 0.0011191f $X=3.615 $Y=1.385 $X2=0 $Y2=0
cc_598 N_CLK_c_717_n N_VGND_c_1821_n 0.00467989f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_599 N_CLK_c_717_n N_VGND_c_1822_n 0.00380993f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_600 N_CLK_c_717_n N_VGND_c_1835_n 0.00434272f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_601 N_CLK_c_717_n N_VGND_c_1842_n 0.00830282f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_602 N_A_958_74#_c_755_n N_A_763_74#_M1033_g 0.00978502f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_603 N_A_958_74#_c_757_n N_A_763_74#_M1033_g 0.00474255f $X=5.095 $Y=0.34
+ $X2=0 $Y2=0
cc_604 N_A_958_74#_c_755_n N_A_763_74#_c_971_n 0.00640673f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_605 N_A_958_74#_c_778_n N_A_763_74#_c_985_n 0.00485767f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_606 N_A_958_74#_c_758_n N_A_763_74#_c_985_n 0.00170003f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_607 N_A_958_74#_c_780_n N_A_763_74#_c_985_n 0.00119344f $X=5.91 $Y=2.06 $X2=0
+ $Y2=0
cc_608 N_A_958_74#_c_781_n N_A_763_74#_c_985_n 0.00523175f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_609 N_A_958_74#_c_755_n N_A_763_74#_M1024_g 0.00475197f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_610 N_A_958_74#_c_756_n N_A_763_74#_M1024_g 0.0146867f $X=5.825 $Y=0.34 $X2=0
+ $Y2=0
cc_611 N_A_958_74#_c_758_n N_A_763_74#_M1024_g 0.0248347f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_612 N_A_958_74#_c_758_n N_A_763_74#_c_973_n 0.0126149f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_613 N_A_958_74#_c_780_n N_A_763_74#_c_973_n 0.00108974f $X=5.91 $Y=2.06 $X2=0
+ $Y2=0
cc_614 N_A_958_74#_c_781_n N_A_763_74#_c_973_n 0.024355f $X=6.085 $Y=2.135 $X2=0
+ $Y2=0
cc_615 N_A_958_74#_c_769_n N_A_763_74#_c_973_n 0.0158136f $X=6.67 $Y=1.145 $X2=0
+ $Y2=0
cc_616 N_A_958_74#_c_770_n N_A_763_74#_c_973_n 0.00140016f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_617 N_A_958_74#_c_778_n N_A_763_74#_c_974_n 0.00801127f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_618 N_A_958_74#_M1013_g N_A_763_74#_M1017_g 0.0174003f $X=6.385 $Y=2.75 $X2=0
+ $Y2=0
cc_619 N_A_958_74#_M1026_g N_A_763_74#_M1030_g 0.0215631f $X=10.365 $Y=2.72
+ $X2=0 $Y2=0
cc_620 N_A_958_74#_c_767_n N_A_763_74#_M1007_g 0.011158f $X=10.275 $Y=1.29 $X2=0
+ $Y2=0
cc_621 N_A_958_74#_c_771_n N_A_763_74#_M1007_g 5.09316e-19 $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_622 N_A_958_74#_c_772_n N_A_763_74#_M1007_g 0.0102681f $X=9.36 $Y=1.385 $X2=0
+ $Y2=0
cc_623 N_A_958_74#_c_773_n N_A_763_74#_M1007_g 8.46596e-19 $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_624 N_A_958_74#_c_774_n N_A_763_74#_M1007_g 0.00953531f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_625 N_A_958_74#_c_775_n N_A_763_74#_M1007_g 0.0190284f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_626 N_A_958_74#_c_755_n N_A_763_74#_c_979_n 0.00591734f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_627 N_A_958_74#_c_755_n N_A_763_74#_c_980_n 0.00264098f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_628 N_A_958_74#_M1026_g N_A_763_74#_c_994_n 4.27252e-19 $X=10.365 $Y=2.72
+ $X2=0 $Y2=0
cc_629 N_A_958_74#_c_781_n N_A_763_74#_c_996_n 0.0111993f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_630 N_A_958_74#_c_767_n N_A_763_74#_c_982_n 0.0283969f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_631 N_A_958_74#_c_773_n N_A_763_74#_c_982_n 0.00253545f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_632 N_A_958_74#_c_774_n N_A_763_74#_c_982_n 0.00164371f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_633 N_A_958_74#_c_767_n N_A_763_74#_c_983_n 0.00481612f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_634 N_A_958_74#_c_771_n N_A_763_74#_c_983_n 4.65488e-19 $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_635 N_A_958_74#_c_772_n N_A_763_74#_c_983_n 0.00547187f $X=9.36 $Y=1.385
+ $X2=0 $Y2=0
cc_636 N_A_958_74#_c_773_n N_A_763_74#_c_983_n 5.91559e-19 $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_637 N_A_958_74#_c_774_n N_A_763_74#_c_983_n 0.0217713f $X=10.44 $Y=1.42 $X2=0
+ $Y2=0
cc_638 N_A_958_74#_c_758_n N_A_763_74#_c_1000_n 2.32223e-19 $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_639 N_A_958_74#_c_781_n N_A_763_74#_c_1000_n 0.0037154f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_640 N_A_958_74#_c_753_n N_A_1409_64#_M1001_g 0.0218463f $X=6.67 $Y=0.98 $X2=0
+ $Y2=0
cc_641 N_A_958_74#_c_759_n N_A_1409_64#_M1001_g 9.04159e-19 $X=6.79 $Y=0.34
+ $X2=0 $Y2=0
cc_642 N_A_958_74#_c_760_n N_A_1409_64#_M1001_g 0.00456962f $X=6.875 $Y=0.935
+ $X2=0 $Y2=0
cc_643 N_A_958_74#_c_761_n N_A_1409_64#_M1001_g 0.0155025f $X=7.59 $Y=1.02 $X2=0
+ $Y2=0
cc_644 N_A_958_74#_c_847_p N_A_1409_64#_M1001_g 0.00183812f $X=7.675 $Y=0.935
+ $X2=0 $Y2=0
cc_645 N_A_958_74#_c_763_n N_A_1409_64#_M1001_g 2.95155e-19 $X=7.76 $Y=0.34
+ $X2=0 $Y2=0
cc_646 N_A_958_74#_c_769_n N_A_1409_64#_M1001_g 0.0205478f $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_647 N_A_958_74#_c_770_n N_A_1409_64#_M1001_g 0.00490258f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_648 N_A_958_74#_c_762_n N_A_1409_64#_M1012_g 6.63977e-19 $X=8.27 $Y=0.34
+ $X2=0 $Y2=0
cc_649 N_A_958_74#_c_764_n N_A_1409_64#_M1012_g 0.00510095f $X=8.355 $Y=0.935
+ $X2=0 $Y2=0
cc_650 N_A_958_74#_c_765_n N_A_1409_64#_M1012_g 0.0165155f $X=9.11 $Y=1.02 $X2=0
+ $Y2=0
cc_651 N_A_958_74#_c_771_n N_A_1409_64#_M1012_g 0.00621114f $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_652 N_A_958_74#_c_772_n N_A_1409_64#_M1012_g 0.0213033f $X=9.36 $Y=1.385
+ $X2=0 $Y2=0
cc_653 N_A_958_74#_c_775_n N_A_1409_64#_M1012_g 0.0321202f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_654 N_A_958_74#_c_765_n N_A_1409_64#_c_1158_n 0.00882684f $X=9.11 $Y=1.02
+ $X2=0 $Y2=0
cc_655 N_A_958_74#_c_766_n N_A_1409_64#_c_1158_n 0.00134551f $X=8.44 $Y=1.02
+ $X2=0 $Y2=0
cc_656 N_A_958_74#_c_761_n N_A_1409_64#_c_1160_n 0.0135045f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_657 N_A_958_74#_c_761_n N_A_1409_64#_c_1161_n 0.00769005f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_658 N_A_958_74#_c_762_n N_A_1409_64#_c_1161_n 0.012971f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_659 N_A_958_74#_c_764_n N_A_1409_64#_c_1161_n 0.0251105f $X=8.355 $Y=0.935
+ $X2=0 $Y2=0
cc_660 N_A_958_74#_c_766_n N_A_1409_64#_c_1161_n 0.0141515f $X=8.44 $Y=1.02
+ $X2=0 $Y2=0
cc_661 N_A_958_74#_c_766_n N_A_1409_64#_c_1163_n 0.0145877f $X=8.44 $Y=1.02
+ $X2=0 $Y2=0
cc_662 N_A_958_74#_c_765_n N_A_1409_64#_c_1177_n 0.0334569f $X=9.11 $Y=1.02
+ $X2=0 $Y2=0
cc_663 N_A_958_74#_c_771_n N_A_1409_64#_c_1177_n 0.0236381f $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_664 N_A_958_74#_c_772_n N_A_1409_64#_c_1177_n 2.66003e-19 $X=9.36 $Y=1.385
+ $X2=0 $Y2=0
cc_665 N_A_958_74#_c_761_n N_A_1409_64#_c_1178_n 0.0319684f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_666 N_A_958_74#_c_770_n N_A_1409_64#_c_1178_n 0.0028512f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_667 N_A_958_74#_c_761_n N_A_1409_64#_c_1164_n 0.00726198f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_668 N_A_958_74#_c_758_n N_A_1156_90#_M1024_d 0.00768863f $X=5.91 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_669 N_A_958_74#_c_761_n N_A_1156_90#_M1004_g 0.00553873f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_670 N_A_958_74#_c_847_p N_A_1156_90#_M1004_g 0.0131174f $X=7.675 $Y=0.935
+ $X2=0 $Y2=0
cc_671 N_A_958_74#_c_762_n N_A_1156_90#_M1004_g 0.0103073f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_958_74#_c_763_n N_A_1156_90#_M1004_g 0.00210537f $X=7.76 $Y=0.34
+ $X2=0 $Y2=0
cc_673 N_A_958_74#_c_764_n N_A_1156_90#_M1004_g 0.00339873f $X=8.355 $Y=0.935
+ $X2=0 $Y2=0
cc_674 N_A_958_74#_c_753_n N_A_1156_90#_c_1257_n 0.00363252f $X=6.67 $Y=0.98
+ $X2=0 $Y2=0
cc_675 N_A_958_74#_c_758_n N_A_1156_90#_c_1257_n 0.06434f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_676 N_A_958_74#_c_760_n N_A_1156_90#_c_1257_n 0.00426874f $X=6.875 $Y=0.935
+ $X2=0 $Y2=0
cc_677 N_A_958_74#_c_769_n N_A_1156_90#_c_1257_n 0.00231928f $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_678 N_A_958_74#_c_770_n N_A_1156_90#_c_1257_n 0.0294985f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_679 N_A_958_74#_c_753_n N_A_1156_90#_c_1285_n 0.00607399f $X=6.67 $Y=0.98
+ $X2=0 $Y2=0
cc_680 N_A_958_74#_c_758_n N_A_1156_90#_c_1285_n 0.0133947f $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_681 N_A_958_74#_c_759_n N_A_1156_90#_c_1285_n 0.0310197f $X=6.79 $Y=0.34
+ $X2=0 $Y2=0
cc_682 N_A_958_74#_c_769_n N_A_1156_90#_c_1285_n 4.46549e-19 $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_683 N_A_958_74#_c_770_n N_A_1156_90#_c_1285_n 0.00682255f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_684 N_A_958_74#_c_758_n N_A_1156_90#_c_1262_n 0.0122725f $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_685 N_A_958_74#_c_780_n N_A_1156_90#_c_1262_n 0.00555219f $X=5.91 $Y=2.06
+ $X2=0 $Y2=0
cc_686 N_A_958_74#_c_781_n N_A_1156_90#_c_1262_n 0.0035112f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_687 N_A_958_74#_c_769_n N_A_1156_90#_c_1262_n 0.00149648f $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_688 N_A_958_74#_c_770_n N_A_1156_90#_c_1262_n 0.0145923f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_689 N_A_958_74#_M1013_g N_A_1156_90#_c_1263_n 0.00773467f $X=6.385 $Y=2.75
+ $X2=0 $Y2=0
cc_690 N_A_958_74#_M1013_g N_A_1156_90#_c_1264_n 0.0107935f $X=6.385 $Y=2.75
+ $X2=0 $Y2=0
cc_691 N_A_958_74#_c_758_n N_A_1156_90#_c_1264_n 7.8612e-19 $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_692 N_A_958_74#_c_780_n N_A_1156_90#_c_1264_n 0.0319585f $X=5.91 $Y=2.06
+ $X2=0 $Y2=0
cc_693 N_A_958_74#_c_781_n N_A_1156_90#_c_1264_n 0.00585766f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_694 N_A_958_74#_c_761_n N_A_1156_90#_c_1260_n 0.00326485f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_695 N_A_958_74#_c_775_n N_A_1895_74#_c_1359_n 0.00968523f $X=9.36 $Y=1.22
+ $X2=0 $Y2=0
cc_696 N_A_958_74#_c_767_n N_A_1895_74#_c_1360_n 0.0306291f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_697 N_A_958_74#_c_773_n N_A_1895_74#_c_1360_n 0.021501f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_698 N_A_958_74#_c_774_n N_A_1895_74#_c_1360_n 3.74086e-19 $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_699 N_A_958_74#_c_767_n N_A_1895_74#_c_1422_n 0.020247f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_700 N_A_958_74#_c_771_n N_A_1895_74#_c_1422_n 6.75349e-19 $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_701 N_A_958_74#_c_775_n N_A_1895_74#_c_1422_n 0.00314181f $X=9.36 $Y=1.22
+ $X2=0 $Y2=0
cc_702 N_A_958_74#_M1026_g N_A_1895_74#_c_1367_n 0.0111547f $X=10.365 $Y=2.72
+ $X2=0 $Y2=0
cc_703 N_A_958_74#_M1026_g N_A_1895_74#_c_1368_n 0.00596987f $X=10.365 $Y=2.72
+ $X2=0 $Y2=0
cc_704 N_A_958_74#_c_773_n N_A_1895_74#_c_1368_n 0.0116227f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_705 N_A_958_74#_c_774_n N_A_1895_74#_c_1368_n 0.00105037f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_706 N_A_958_74#_M1026_g N_A_1895_74#_c_1369_n 0.0176305f $X=10.365 $Y=2.72
+ $X2=0 $Y2=0
cc_707 N_A_958_74#_c_767_n N_A_1895_74#_c_1369_n 0.00357633f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_708 N_A_958_74#_c_773_n N_A_1895_74#_c_1369_n 0.00771291f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_709 N_A_958_74#_M1026_g N_A_1895_74#_c_1361_n 0.00231398f $X=10.365 $Y=2.72
+ $X2=0 $Y2=0
cc_710 N_A_958_74#_c_773_n N_A_1895_74#_c_1361_n 0.0187515f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_711 N_A_958_74#_c_774_n N_A_1895_74#_c_1361_n 0.00131611f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_712 N_A_958_74#_c_773_n N_A_1895_74#_c_1364_n 0.0111691f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_713 N_A_958_74#_c_774_n N_A_1895_74#_c_1364_n 4.90605e-19 $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_714 N_A_958_74#_c_778_n N_A_27_508#_c_1498_n 0.0138332f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_715 N_A_958_74#_c_758_n N_A_27_508#_c_1498_n 0.0041226f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_716 N_A_958_74#_c_778_n N_A_27_508#_c_1483_n 0.011918f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_717 N_A_958_74#_c_758_n N_A_27_508#_c_1483_n 0.0123714f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_718 N_A_958_74#_c_755_n N_A_27_508#_c_1484_n 0.0360689f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_719 N_A_958_74#_c_756_n N_A_27_508#_c_1484_n 0.0229863f $X=5.825 $Y=0.34
+ $X2=0 $Y2=0
cc_720 N_A_958_74#_c_758_n N_A_27_508#_c_1484_n 0.0561201f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_721 N_A_958_74#_M1005_d N_A_27_508#_c_1499_n 0.00568043f $X=5.5 $Y=1.84 $X2=0
+ $Y2=0
cc_722 N_A_958_74#_M1013_g N_A_27_508#_c_1499_n 7.77652e-19 $X=6.385 $Y=2.75
+ $X2=0 $Y2=0
cc_723 N_A_958_74#_c_778_n N_A_27_508#_c_1499_n 0.00923409f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_724 N_A_958_74#_c_780_n N_A_27_508#_c_1499_n 0.0284908f $X=5.91 $Y=2.06 $X2=0
+ $Y2=0
cc_725 N_A_958_74#_c_781_n N_A_27_508#_c_1499_n 0.00233063f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_726 N_A_958_74#_M1005_d N_A_27_508#_c_1564_n 0.0058186f $X=5.5 $Y=1.84 $X2=0
+ $Y2=0
cc_727 N_A_958_74#_M1013_g N_A_27_508#_c_1564_n 0.00501053f $X=6.385 $Y=2.75
+ $X2=0 $Y2=0
cc_728 N_A_958_74#_c_778_n N_A_27_508#_c_1564_n 0.00637529f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_729 N_A_958_74#_M1013_g N_A_27_508#_c_1500_n 7.6107e-19 $X=6.385 $Y=2.75
+ $X2=0 $Y2=0
cc_730 N_A_958_74#_M1026_g N_VPWR_c_1660_n 0.00167758f $X=10.365 $Y=2.72 $X2=0
+ $Y2=0
cc_731 N_A_958_74#_M1013_g N_VPWR_c_1672_n 0.0048691f $X=6.385 $Y=2.75 $X2=0
+ $Y2=0
cc_732 N_A_958_74#_M1026_g N_VPWR_c_1673_n 0.00667211f $X=10.365 $Y=2.72 $X2=0
+ $Y2=0
cc_733 N_A_958_74#_M1013_g N_VPWR_c_1653_n 0.00878547f $X=6.385 $Y=2.75 $X2=0
+ $Y2=0
cc_734 N_A_958_74#_M1026_g N_VPWR_c_1653_n 0.00643509f $X=10.365 $Y=2.72 $X2=0
+ $Y2=0
cc_735 N_A_958_74#_c_761_n N_VGND_M1001_d 0.00494641f $X=7.59 $Y=1.02 $X2=0
+ $Y2=0
cc_736 N_A_958_74#_c_847_p N_VGND_M1001_d 0.00544252f $X=7.675 $Y=0.935 $X2=0
+ $Y2=0
cc_737 N_A_958_74#_c_765_n N_VGND_M1012_s 0.0068916f $X=9.11 $Y=1.02 $X2=0 $Y2=0
cc_738 N_A_958_74#_c_755_n N_VGND_c_1822_n 0.0259603f $X=4.93 $Y=0.515 $X2=0
+ $Y2=0
cc_739 N_A_958_74#_c_757_n N_VGND_c_1822_n 0.0112234f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_740 N_A_958_74#_c_759_n N_VGND_c_1823_n 0.0122752f $X=6.79 $Y=0.34 $X2=0
+ $Y2=0
cc_741 N_A_958_74#_c_760_n N_VGND_c_1823_n 0.0208855f $X=6.875 $Y=0.935 $X2=0
+ $Y2=0
cc_742 N_A_958_74#_c_761_n N_VGND_c_1823_n 0.0177503f $X=7.59 $Y=1.02 $X2=0
+ $Y2=0
cc_743 N_A_958_74#_c_847_p N_VGND_c_1823_n 0.025461f $X=7.675 $Y=0.935 $X2=0
+ $Y2=0
cc_744 N_A_958_74#_c_763_n N_VGND_c_1823_n 0.014745f $X=7.76 $Y=0.34 $X2=0 $Y2=0
cc_745 N_A_958_74#_c_762_n N_VGND_c_1824_n 0.0146661f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_746 N_A_958_74#_c_764_n N_VGND_c_1824_n 0.0258447f $X=8.355 $Y=0.935 $X2=0
+ $Y2=0
cc_747 N_A_958_74#_c_765_n N_VGND_c_1824_n 0.0154151f $X=9.11 $Y=1.02 $X2=0
+ $Y2=0
cc_748 N_A_958_74#_c_775_n N_VGND_c_1824_n 0.00180636f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_749 N_A_958_74#_c_753_n N_VGND_c_1829_n 8.05596e-19 $X=6.67 $Y=0.98 $X2=0
+ $Y2=0
cc_750 N_A_958_74#_c_756_n N_VGND_c_1829_n 0.0469671f $X=5.825 $Y=0.34 $X2=0
+ $Y2=0
cc_751 N_A_958_74#_c_757_n N_VGND_c_1829_n 0.0235688f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_752 N_A_958_74#_c_759_n N_VGND_c_1829_n 0.063341f $X=6.79 $Y=0.34 $X2=0 $Y2=0
cc_753 N_A_958_74#_c_768_n N_VGND_c_1829_n 0.0121867f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_754 N_A_958_74#_c_762_n N_VGND_c_1831_n 0.0449818f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_755 N_A_958_74#_c_763_n N_VGND_c_1831_n 0.0121867f $X=7.76 $Y=0.34 $X2=0
+ $Y2=0
cc_756 N_A_958_74#_c_775_n N_VGND_c_1840_n 0.00434272f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_757 N_A_958_74#_c_756_n N_VGND_c_1842_n 0.0274384f $X=5.825 $Y=0.34 $X2=0
+ $Y2=0
cc_758 N_A_958_74#_c_757_n N_VGND_c_1842_n 0.0127152f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_759 N_A_958_74#_c_759_n N_VGND_c_1842_n 0.0364914f $X=6.79 $Y=0.34 $X2=0
+ $Y2=0
cc_760 N_A_958_74#_c_762_n N_VGND_c_1842_n 0.025776f $X=8.27 $Y=0.34 $X2=0 $Y2=0
cc_761 N_A_958_74#_c_763_n N_VGND_c_1842_n 0.00660921f $X=7.76 $Y=0.34 $X2=0
+ $Y2=0
cc_762 N_A_958_74#_c_768_n N_VGND_c_1842_n 0.00660921f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_763 N_A_958_74#_c_775_n N_VGND_c_1842_n 0.00822691f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_764 N_A_958_74#_c_760_n A_1349_90# 0.00579581f $X=6.875 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_765 N_A_958_74#_c_765_n A_1797_74# 0.00378025f $X=9.11 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_766 N_A_958_74#_c_771_n A_1797_74# 0.00761182f $X=9.285 $Y=1.29 $X2=-0.19
+ $Y2=-0.245
cc_767 N_A_763_74#_c_993_n N_A_1409_64#_M1023_d 0.00768578f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_768 N_A_763_74#_c_973_n N_A_1409_64#_M1020_g 0.0125636f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_769 N_A_763_74#_M1017_g N_A_1409_64#_M1020_g 0.0274184f $X=6.835 $Y=2.75
+ $X2=0 $Y2=0
cc_770 N_A_763_74#_c_993_n N_A_1409_64#_M1020_g 0.0164131f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_771 N_A_763_74#_c_995_n N_A_1409_64#_M1020_g 0.00981771f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_772 N_A_763_74#_c_996_n N_A_1409_64#_M1020_g 0.0196743f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_773 N_A_763_74#_c_993_n N_A_1409_64#_M1018_g 0.0230891f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_774 N_A_763_74#_c_994_n N_A_1409_64#_M1018_g 0.0145515f $X=9.715 $Y=2.41
+ $X2=0 $Y2=0
cc_775 N_A_763_74#_c_982_n N_A_1409_64#_c_1159_n 0.00294553f $X=9.9 $Y=1.635
+ $X2=0 $Y2=0
cc_776 N_A_763_74#_c_993_n N_A_1409_64#_c_1167_n 0.0335536f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_777 N_A_763_74#_c_993_n N_A_1156_90#_M1023_g 0.018103f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_778 N_A_763_74#_c_973_n N_A_1156_90#_c_1257_n 0.00673678f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_779 N_A_763_74#_c_973_n N_A_1156_90#_c_1262_n 0.0119426f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_780 N_A_763_74#_M1017_g N_A_1156_90#_c_1263_n 0.0106519f $X=6.835 $Y=2.75
+ $X2=0 $Y2=0
cc_781 N_A_763_74#_c_995_n N_A_1156_90#_c_1263_n 0.00452884f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_782 N_A_763_74#_c_996_n N_A_1156_90#_c_1263_n 0.00270314f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_783 N_A_763_74#_c_973_n N_A_1156_90#_c_1264_n 0.00102203f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_784 N_A_763_74#_M1017_g N_A_1156_90#_c_1264_n 0.00147536f $X=6.835 $Y=2.75
+ $X2=0 $Y2=0
cc_785 N_A_763_74#_c_995_n N_A_1156_90#_c_1264_n 0.0341444f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_786 N_A_763_74#_c_1000_n N_A_1156_90#_c_1264_n 0.00950617f $X=6.862 $Y=2
+ $X2=0 $Y2=0
cc_787 N_A_763_74#_c_993_n N_A_1156_90#_c_1258_n 0.00552924f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_788 N_A_763_74#_c_993_n N_A_1156_90#_c_1259_n 0.00161236f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_789 N_A_763_74#_c_973_n N_A_1156_90#_c_1260_n 0.0052678f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_790 N_A_763_74#_c_993_n N_A_1156_90#_c_1260_n 0.0165064f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_791 N_A_763_74#_c_995_n N_A_1156_90#_c_1260_n 0.0220457f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_792 N_A_763_74#_c_996_n N_A_1156_90#_c_1260_n 0.00138798f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_793 N_A_763_74#_c_1000_n N_A_1156_90#_c_1260_n 0.00772026f $X=6.862 $Y=2
+ $X2=0 $Y2=0
cc_794 N_A_763_74#_M1007_g N_A_1895_74#_c_1359_n 0.00369459f $X=9.91 $Y=0.58
+ $X2=0 $Y2=0
cc_795 N_A_763_74#_M1007_g N_A_1895_74#_c_1360_n 0.0121459f $X=9.91 $Y=0.58
+ $X2=0 $Y2=0
cc_796 N_A_763_74#_M1030_g N_A_1895_74#_c_1367_n 0.00106024f $X=9.83 $Y=2.46
+ $X2=0 $Y2=0
cc_797 N_A_763_74#_M1030_g N_A_1895_74#_c_1369_n 0.00138628f $X=9.83 $Y=2.46
+ $X2=0 $Y2=0
cc_798 N_A_763_74#_c_994_n N_A_1895_74#_c_1369_n 0.0141024f $X=9.715 $Y=2.41
+ $X2=0 $Y2=0
cc_799 N_A_763_74#_c_982_n N_A_1895_74#_c_1369_n 0.0056188f $X=9.9 $Y=1.635
+ $X2=0 $Y2=0
cc_800 N_A_763_74#_c_983_n N_A_1895_74#_c_1369_n 0.00290424f $X=9.9 $Y=1.635
+ $X2=0 $Y2=0
cc_801 N_A_763_74#_M1025_d N_A_27_508#_c_1497_n 0.00698137f $X=4.15 $Y=1.76
+ $X2=0 $Y2=0
cc_802 N_A_763_74#_c_971_n N_A_27_508#_c_1497_n 0.00248816f $X=5.32 $Y=1.655
+ $X2=0 $Y2=0
cc_803 N_A_763_74#_c_978_n N_A_27_508#_c_1497_n 0.0111569f $X=4.12 $Y=1.805
+ $X2=0 $Y2=0
cc_804 N_A_763_74#_c_979_n N_A_27_508#_c_1497_n 0.056864f $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_805 N_A_763_74#_c_999_n N_A_27_508#_c_1497_n 0.00862812f $X=4.735 $Y=1.655
+ $X2=0 $Y2=0
cc_806 N_A_763_74#_c_971_n N_A_27_508#_c_1498_n 0.00590951f $X=5.32 $Y=1.655
+ $X2=0 $Y2=0
cc_807 N_A_763_74#_c_985_n N_A_27_508#_c_1498_n 0.00702545f $X=5.41 $Y=1.73
+ $X2=0 $Y2=0
cc_808 N_A_763_74#_c_979_n N_A_27_508#_c_1498_n 0.0292713f $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_809 N_A_763_74#_c_999_n N_A_27_508#_c_1498_n 0.00148825f $X=4.735 $Y=1.655
+ $X2=0 $Y2=0
cc_810 N_A_763_74#_c_971_n N_A_27_508#_c_1483_n 0.00546736f $X=5.32 $Y=1.655
+ $X2=0 $Y2=0
cc_811 N_A_763_74#_M1024_g N_A_27_508#_c_1483_n 0.00334012f $X=5.705 $Y=0.66
+ $X2=0 $Y2=0
cc_812 N_A_763_74#_c_974_n N_A_27_508#_c_1483_n 0.011932f $X=5.78 $Y=1.655 $X2=0
+ $Y2=0
cc_813 N_A_763_74#_c_979_n N_A_27_508#_c_1483_n 0.0104131f $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_814 N_A_763_74#_c_980_n N_A_27_508#_c_1483_n 7.30496e-19 $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_815 N_A_763_74#_M1033_g N_A_27_508#_c_1484_n 0.00970544f $X=4.715 $Y=0.74
+ $X2=0 $Y2=0
cc_816 N_A_763_74#_M1024_g N_A_27_508#_c_1484_n 0.0222528f $X=5.705 $Y=0.66
+ $X2=0 $Y2=0
cc_817 N_A_763_74#_c_974_n N_A_27_508#_c_1484_n 0.00196875f $X=5.78 $Y=1.655
+ $X2=0 $Y2=0
cc_818 N_A_763_74#_c_979_n N_A_27_508#_c_1484_n 3.79465e-19 $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_819 N_A_763_74#_c_985_n N_A_27_508#_c_1564_n 0.0320751f $X=5.41 $Y=1.73 $X2=0
+ $Y2=0
cc_820 N_A_763_74#_c_985_n N_A_27_508#_c_1500_n 0.00752696f $X=5.41 $Y=1.73
+ $X2=0 $Y2=0
cc_821 N_A_763_74#_c_993_n N_VPWR_M1020_d 0.00639897f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_822 N_A_763_74#_c_993_n N_VPWR_M1018_s 0.0117572f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_823 N_A_763_74#_c_985_n N_VPWR_c_1657_n 0.00536186f $X=5.41 $Y=1.73 $X2=0
+ $Y2=0
cc_824 N_A_763_74#_M1017_g N_VPWR_c_1658_n 0.0012037f $X=6.835 $Y=2.75 $X2=0
+ $Y2=0
cc_825 N_A_763_74#_c_993_n N_VPWR_c_1658_n 0.0211156f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_826 N_A_763_74#_c_993_n N_VPWR_c_1659_n 0.0212012f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_827 N_A_763_74#_c_993_n N_VPWR_c_1669_n 0.00977184f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_828 N_A_763_74#_c_985_n N_VPWR_c_1672_n 0.00499824f $X=5.41 $Y=1.73 $X2=0
+ $Y2=0
cc_829 N_A_763_74#_M1017_g N_VPWR_c_1672_n 0.005209f $X=6.835 $Y=2.75 $X2=0
+ $Y2=0
cc_830 N_A_763_74#_c_993_n N_VPWR_c_1672_n 0.00350068f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_831 N_A_763_74#_c_995_n N_VPWR_c_1672_n 0.00227549f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_832 N_A_763_74#_M1030_g N_VPWR_c_1673_n 0.00504357f $X=9.83 $Y=2.46 $X2=0
+ $Y2=0
cc_833 N_A_763_74#_c_993_n N_VPWR_c_1673_n 0.0124331f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_834 N_A_763_74#_c_985_n N_VPWR_c_1653_n 0.00547071f $X=5.41 $Y=1.73 $X2=0
+ $Y2=0
cc_835 N_A_763_74#_M1017_g N_VPWR_c_1653_n 0.00984084f $X=6.835 $Y=2.75 $X2=0
+ $Y2=0
cc_836 N_A_763_74#_M1030_g N_VPWR_c_1653_n 0.00913029f $X=9.83 $Y=2.46 $X2=0
+ $Y2=0
cc_837 N_A_763_74#_c_993_n N_VPWR_c_1653_n 0.0536685f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_838 N_A_763_74#_c_995_n N_VPWR_c_1653_n 0.00470026f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_839 N_A_763_74#_c_993_n A_1385_508# 0.00151223f $X=9.63 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_840 N_A_763_74#_c_995_n A_1385_508# 0.00292236f $X=6.875 $Y=2.165 $X2=-0.19
+ $Y2=-0.245
cc_841 N_A_763_74#_c_993_n A_1797_392# 0.0386712f $X=9.63 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_842 N_A_763_74#_c_994_n A_1797_392# 0.0078024f $X=9.715 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_843 N_A_763_74#_c_976_n N_VGND_c_1821_n 0.024306f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_844 N_A_763_74#_M1033_g N_VGND_c_1822_n 0.00473533f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_845 N_A_763_74#_c_976_n N_VGND_c_1822_n 0.0534949f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_846 N_A_763_74#_c_979_n N_VGND_c_1822_n 0.0122043f $X=4.735 $Y=1.635 $X2=0
+ $Y2=0
cc_847 N_A_763_74#_c_980_n N_VGND_c_1822_n 3.36125e-19 $X=4.735 $Y=1.635 $X2=0
+ $Y2=0
cc_848 N_A_763_74#_M1033_g N_VGND_c_1829_n 0.00430908f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_849 N_A_763_74#_M1024_g N_VGND_c_1829_n 8.05596e-19 $X=5.705 $Y=0.66 $X2=0
+ $Y2=0
cc_850 N_A_763_74#_c_976_n N_VGND_c_1835_n 0.0145488f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_851 N_A_763_74#_M1007_g N_VGND_c_1840_n 0.00461464f $X=9.91 $Y=0.58 $X2=0
+ $Y2=0
cc_852 N_A_763_74#_M1007_g N_VGND_c_1841_n 0.00147769f $X=9.91 $Y=0.58 $X2=0
+ $Y2=0
cc_853 N_A_763_74#_M1033_g N_VGND_c_1842_n 0.0082568f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_854 N_A_763_74#_M1007_g N_VGND_c_1842_n 0.00463846f $X=9.91 $Y=0.58 $X2=0
+ $Y2=0
cc_855 N_A_763_74#_c_976_n N_VGND_c_1842_n 0.0119924f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_856 N_A_1409_64#_M1001_g N_A_1156_90#_M1004_g 0.0132329f $X=7.12 $Y=0.66
+ $X2=0 $Y2=0
cc_857 N_A_1409_64#_c_1158_n N_A_1156_90#_M1004_g 0.00723897f $X=8.805 $Y=1.44
+ $X2=0 $Y2=0
cc_858 N_A_1409_64#_c_1160_n N_A_1156_90#_M1004_g 0.0143234f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_859 N_A_1409_64#_c_1161_n N_A_1156_90#_M1004_g 0.00891563f $X=8.015 $Y=0.85
+ $X2=0 $Y2=0
cc_860 N_A_1409_64#_c_1163_n N_A_1156_90#_M1004_g 5.12204e-19 $X=8.44 $Y=1.44
+ $X2=0 $Y2=0
cc_861 N_A_1409_64#_c_1164_n N_A_1156_90#_M1004_g 0.0169447f $X=7.34 $Y=1.365
+ $X2=0 $Y2=0
cc_862 N_A_1409_64#_M1020_g N_A_1156_90#_M1023_g 0.0335606f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_863 N_A_1409_64#_c_1167_n N_A_1156_90#_M1023_g 0.00446827f $X=8.27 $Y=2.155
+ $X2=0 $Y2=0
cc_864 N_A_1409_64#_c_1162_n N_A_1156_90#_M1023_g 0.00554531f $X=8.355 $Y=2.07
+ $X2=0 $Y2=0
cc_865 N_A_1409_64#_M1020_g N_A_1156_90#_c_1263_n 0.00153499f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_866 N_A_1409_64#_M1020_g N_A_1156_90#_c_1258_n 3.28132e-19 $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_867 N_A_1409_64#_c_1160_n N_A_1156_90#_c_1258_n 0.0139504f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_868 N_A_1409_64#_c_1167_n N_A_1156_90#_c_1258_n 0.00284462f $X=8.27 $Y=2.155
+ $X2=0 $Y2=0
cc_869 N_A_1409_64#_c_1162_n N_A_1156_90#_c_1258_n 0.0113679f $X=8.355 $Y=2.07
+ $X2=0 $Y2=0
cc_870 N_A_1409_64#_c_1163_n N_A_1156_90#_c_1258_n 0.00702578f $X=8.44 $Y=1.44
+ $X2=0 $Y2=0
cc_871 N_A_1409_64#_M1020_g N_A_1156_90#_c_1259_n 0.0165867f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_872 N_A_1409_64#_c_1158_n N_A_1156_90#_c_1259_n 0.0037983f $X=8.805 $Y=1.44
+ $X2=0 $Y2=0
cc_873 N_A_1409_64#_c_1160_n N_A_1156_90#_c_1259_n 0.00220559f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_874 N_A_1409_64#_c_1162_n N_A_1156_90#_c_1259_n 0.0028377f $X=8.355 $Y=2.07
+ $X2=0 $Y2=0
cc_875 N_A_1409_64#_c_1163_n N_A_1156_90#_c_1259_n 0.00328914f $X=8.44 $Y=1.44
+ $X2=0 $Y2=0
cc_876 N_A_1409_64#_M1020_g N_A_1156_90#_c_1260_n 0.0137102f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_877 N_A_1409_64#_c_1160_n N_A_1156_90#_c_1260_n 0.0143302f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_878 N_A_1409_64#_c_1178_n N_A_1156_90#_c_1260_n 0.0201775f $X=7.46 $Y=1.367
+ $X2=0 $Y2=0
cc_879 N_A_1409_64#_c_1164_n N_A_1156_90#_c_1260_n 0.00655078f $X=7.34 $Y=1.365
+ $X2=0 $Y2=0
cc_880 N_A_1409_64#_M1012_g N_A_1895_74#_c_1359_n 0.00159894f $X=8.91 $Y=0.74
+ $X2=0 $Y2=0
cc_881 N_A_1409_64#_M1012_g N_A_1895_74#_c_1422_n 5.21752e-19 $X=8.91 $Y=0.74
+ $X2=0 $Y2=0
cc_882 N_A_1409_64#_M1020_g N_VPWR_c_1658_n 0.00967292f $X=7.34 $Y=2.75 $X2=0
+ $Y2=0
cc_883 N_A_1409_64#_M1018_g N_VPWR_c_1659_n 0.0185022f $X=8.895 $Y=2.46 $X2=0
+ $Y2=0
cc_884 N_A_1409_64#_M1020_g N_VPWR_c_1672_n 0.00360022f $X=7.34 $Y=2.75 $X2=0
+ $Y2=0
cc_885 N_A_1409_64#_M1018_g N_VPWR_c_1673_n 0.00337485f $X=8.895 $Y=2.46 $X2=0
+ $Y2=0
cc_886 N_A_1409_64#_M1020_g N_VPWR_c_1653_n 0.00467883f $X=7.34 $Y=2.75 $X2=0
+ $Y2=0
cc_887 N_A_1409_64#_M1018_g N_VPWR_c_1653_n 0.00443342f $X=8.895 $Y=2.46 $X2=0
+ $Y2=0
cc_888 N_A_1409_64#_M1001_g N_VGND_c_1823_n 0.00752223f $X=7.12 $Y=0.66 $X2=0
+ $Y2=0
cc_889 N_A_1409_64#_M1012_g N_VGND_c_1824_n 0.0133979f $X=8.91 $Y=0.74 $X2=0
+ $Y2=0
cc_890 N_A_1409_64#_M1001_g N_VGND_c_1829_n 0.00432588f $X=7.12 $Y=0.66 $X2=0
+ $Y2=0
cc_891 N_A_1409_64#_M1012_g N_VGND_c_1840_n 0.00383152f $X=8.91 $Y=0.74 $X2=0
+ $Y2=0
cc_892 N_A_1409_64#_M1001_g N_VGND_c_1842_n 0.00437282f $X=7.12 $Y=0.66 $X2=0
+ $Y2=0
cc_893 N_A_1409_64#_M1012_g N_VGND_c_1842_n 0.00758168f $X=8.91 $Y=0.74 $X2=0
+ $Y2=0
cc_894 N_A_1156_90#_c_1263_n N_A_27_508#_c_1499_n 0.0073808f $X=6.61 $Y=2.75
+ $X2=0 $Y2=0
cc_895 N_A_1156_90#_c_1263_n N_A_27_508#_c_1500_n 0.0117853f $X=6.61 $Y=2.75
+ $X2=0 $Y2=0
cc_896 N_A_1156_90#_M1023_g N_VPWR_c_1658_n 0.00430567f $X=7.885 $Y=2.445 $X2=0
+ $Y2=0
cc_897 N_A_1156_90#_c_1263_n N_VPWR_c_1658_n 0.00580551f $X=6.61 $Y=2.75 $X2=0
+ $Y2=0
cc_898 N_A_1156_90#_M1023_g N_VPWR_c_1659_n 0.0063586f $X=7.885 $Y=2.445 $X2=0
+ $Y2=0
cc_899 N_A_1156_90#_M1023_g N_VPWR_c_1669_n 0.00481391f $X=7.885 $Y=2.445 $X2=0
+ $Y2=0
cc_900 N_A_1156_90#_c_1263_n N_VPWR_c_1672_n 0.0154817f $X=6.61 $Y=2.75 $X2=0
+ $Y2=0
cc_901 N_A_1156_90#_M1023_g N_VPWR_c_1653_n 0.00619157f $X=7.885 $Y=2.445 $X2=0
+ $Y2=0
cc_902 N_A_1156_90#_c_1263_n N_VPWR_c_1653_n 0.0127081f $X=6.61 $Y=2.75 $X2=0
+ $Y2=0
cc_903 N_A_1156_90#_M1004_g N_VGND_c_1823_n 0.00129371f $X=7.8 $Y=0.77 $X2=0
+ $Y2=0
cc_904 N_A_1156_90#_M1004_g N_VGND_c_1831_n 8.23937e-19 $X=7.8 $Y=0.77 $X2=0
+ $Y2=0
cc_905 N_A_1895_74#_M1014_g N_VPWR_c_1660_n 0.00729563f $X=11.495 $Y=2.61 $X2=0
+ $Y2=0
cc_906 N_A_1895_74#_c_1367_n N_VPWR_c_1660_n 0.00760545f $X=10.055 $Y=2.105
+ $X2=0 $Y2=0
cc_907 N_A_1895_74#_M1031_g N_VPWR_c_1662_n 0.00649215f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_908 N_A_1895_74#_c_1367_n N_VPWR_c_1673_n 0.0120294f $X=10.055 $Y=2.105 $X2=0
+ $Y2=0
cc_909 N_A_1895_74#_M1014_g N_VPWR_c_1674_n 0.00636575f $X=11.495 $Y=2.61 $X2=0
+ $Y2=0
cc_910 N_A_1895_74#_M1031_g N_VPWR_c_1674_n 0.005209f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_911 N_A_1895_74#_M1014_g N_VPWR_c_1653_n 0.00643509f $X=11.495 $Y=2.61 $X2=0
+ $Y2=0
cc_912 N_A_1895_74#_M1031_g N_VPWR_c_1653_n 0.00991105f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_913 N_A_1895_74#_c_1367_n N_VPWR_c_1653_n 0.00926813f $X=10.055 $Y=2.105
+ $X2=0 $Y2=0
cc_914 N_A_1895_74#_c_1356_n N_Q_c_1791_n 0.00837961f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_915 N_A_1895_74#_c_1355_n N_Q_c_1792_n 0.00274954f $X=12.32 $Y=1.26 $X2=0
+ $Y2=0
cc_916 N_A_1895_74#_c_1356_n N_Q_c_1792_n 0.00214314f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_917 N_A_1895_74#_M1014_g Q 0.00265655f $X=11.495 $Y=2.61 $X2=0 $Y2=0
cc_918 N_A_1895_74#_M1031_g Q 0.0354022f $X=12.465 $Y=2.4 $X2=0 $Y2=0
cc_919 N_A_1895_74#_c_1355_n N_Q_c_1794_n 0.0167995f $X=12.32 $Y=1.26 $X2=0
+ $Y2=0
cc_920 N_A_1895_74#_c_1356_n N_Q_c_1794_n 0.00326896f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_921 N_A_1895_74#_M1031_g N_Q_c_1794_n 0.00920291f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_922 N_A_1895_74#_c_1358_n N_Q_c_1794_n 0.00652656f $X=12.437 $Y=1.26 $X2=0
+ $Y2=0
cc_923 N_A_1895_74#_c_1359_n N_VGND_c_1824_n 0.0109084f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_924 N_A_1895_74#_c_1356_n N_VGND_c_1826_n 0.0196825f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_925 N_A_1895_74#_c_1358_n N_VGND_c_1826_n 0.00213924f $X=12.437 $Y=1.26 $X2=0
+ $Y2=0
cc_926 N_A_1895_74#_M1003_g N_VGND_c_1836_n 0.00461464f $X=11.405 $Y=0.58 $X2=0
+ $Y2=0
cc_927 N_A_1895_74#_c_1356_n N_VGND_c_1836_n 0.00434272f $X=12.395 $Y=1.185
+ $X2=0 $Y2=0
cc_928 N_A_1895_74#_c_1359_n N_VGND_c_1840_n 0.0145243f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_929 N_A_1895_74#_M1003_g N_VGND_c_1841_n 0.00540028f $X=11.405 $Y=0.58 $X2=0
+ $Y2=0
cc_930 N_A_1895_74#_c_1359_n N_VGND_c_1841_n 0.00520222f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_931 N_A_1895_74#_c_1360_n N_VGND_c_1841_n 0.0313981f $X=10.775 $Y=0.92 $X2=0
+ $Y2=0
cc_932 N_A_1895_74#_c_1362_n N_VGND_c_1841_n 0.0175339f $X=11.34 $Y=1.17 $X2=0
+ $Y2=0
cc_933 N_A_1895_74#_c_1363_n N_VGND_c_1841_n 0.00268565f $X=11.34 $Y=1.17 $X2=0
+ $Y2=0
cc_934 N_A_1895_74#_c_1364_n N_VGND_c_1841_n 0.0151641f $X=10.86 $Y=1.085 $X2=0
+ $Y2=0
cc_935 N_A_1895_74#_M1003_g N_VGND_c_1842_n 0.00917524f $X=11.405 $Y=0.58 $X2=0
+ $Y2=0
cc_936 N_A_1895_74#_c_1356_n N_VGND_c_1842_n 0.00828933f $X=12.395 $Y=1.185
+ $X2=0 $Y2=0
cc_937 N_A_1895_74#_c_1359_n N_VGND_c_1842_n 0.0119829f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_938 N_A_1895_74#_c_1360_n N_VGND_c_1842_n 0.0191617f $X=10.775 $Y=0.92 $X2=0
+ $Y2=0
cc_939 N_A_1895_74#_c_1364_n N_VGND_c_1842_n 6.25089e-19 $X=10.86 $Y=1.085 $X2=0
+ $Y2=0
cc_940 N_A_27_508#_c_1493_n N_VPWR_M1032_d 0.00650381f $X=2.13 $Y=2.905 $X2=0
+ $Y2=0
cc_941 N_A_27_508#_c_1497_n N_VPWR_M1025_s 0.0070834f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_942 N_A_27_508#_c_1497_n N_VPWR_M1005_s 0.00194622f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_943 N_A_27_508#_c_1498_n N_VPWR_M1005_s 0.0110601f $X=5.215 $Y=2.31 $X2=0
+ $Y2=0
cc_944 N_A_27_508#_c_1564_n N_VPWR_M1005_s 0.00153606f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_945 N_A_27_508#_c_1488_n N_VPWR_c_1654_n 0.0138414f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_946 N_A_27_508#_c_1489_n N_VPWR_c_1654_n 0.0201388f $X=1.365 $Y=2.265 $X2=0
+ $Y2=0
cc_947 N_A_27_508#_c_1490_n N_VPWR_c_1654_n 0.0292992f $X=1.45 $Y=2.905 $X2=0
+ $Y2=0
cc_948 N_A_27_508#_c_1492_n N_VPWR_c_1654_n 0.0146661f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_949 N_A_27_508#_c_1491_n N_VPWR_c_1655_n 0.0147456f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_950 N_A_27_508#_c_1493_n N_VPWR_c_1655_n 0.0465116f $X=2.13 $Y=2.905 $X2=0
+ $Y2=0
cc_951 N_A_27_508#_c_1494_n N_VPWR_c_1655_n 0.0174776f $X=3.1 $Y=2.035 $X2=0
+ $Y2=0
cc_952 N_A_27_508#_c_1502_n N_VPWR_c_1655_n 0.0111167f $X=3.31 $Y=2.39 $X2=0
+ $Y2=0
cc_953 N_A_27_508#_c_1497_n N_VPWR_c_1656_n 0.0214974f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_954 N_A_27_508#_c_1497_n N_VPWR_c_1657_n 0.00876485f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_955 N_A_27_508#_c_1564_n N_VPWR_c_1657_n 0.0116705f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_956 N_A_27_508#_c_1488_n N_VPWR_c_1663_n 0.0154414f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_957 N_A_27_508#_c_1491_n N_VPWR_c_1665_n 0.0449818f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_958 N_A_27_508#_c_1492_n N_VPWR_c_1665_n 0.0121867f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_959 N_A_27_508#_c_1502_n N_VPWR_c_1667_n 0.0062845f $X=3.31 $Y=2.39 $X2=0
+ $Y2=0
cc_960 N_A_27_508#_c_1499_n N_VPWR_c_1672_n 0.00681477f $X=5.995 $Y=2.605 $X2=0
+ $Y2=0
cc_961 N_A_27_508#_c_1564_n N_VPWR_c_1672_n 0.00254381f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_962 N_A_27_508#_c_1500_n N_VPWR_c_1672_n 0.0107588f $X=6.16 $Y=2.75 $X2=0
+ $Y2=0
cc_963 N_A_27_508#_c_1488_n N_VPWR_c_1653_n 0.0127129f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_964 N_A_27_508#_c_1491_n N_VPWR_c_1653_n 0.025776f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_965 N_A_27_508#_c_1492_n N_VPWR_c_1653_n 0.00660921f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_966 N_A_27_508#_c_1497_n N_VPWR_c_1653_n 0.0425703f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_967 N_A_27_508#_c_1499_n N_VPWR_c_1653_n 0.0109468f $X=5.995 $Y=2.605 $X2=0
+ $Y2=0
cc_968 N_A_27_508#_c_1564_n N_VPWR_c_1653_n 0.0103201f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_969 N_A_27_508#_c_1500_n N_VPWR_c_1653_n 0.00904147f $X=6.16 $Y=2.75 $X2=0
+ $Y2=0
cc_970 N_A_27_508#_c_1502_n N_VPWR_c_1653_n 0.0105777f $X=3.31 $Y=2.39 $X2=0
+ $Y2=0
cc_971 N_A_27_508#_c_1485_n N_VGND_c_1819_n 0.00841519f $X=0.365 $Y=0.575 $X2=0
+ $Y2=0
cc_972 N_A_27_508#_c_1486_n N_VGND_c_1820_n 0.01581f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_973 N_A_27_508#_c_1482_n N_VGND_c_1821_n 0.00998528f $X=3.185 $Y=1.95 $X2=0
+ $Y2=0
cc_974 N_A_27_508#_c_1486_n N_VGND_c_1821_n 0.0369819f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_975 N_A_27_508#_c_1486_n N_VGND_c_1827_n 0.0163765f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_976 N_A_27_508#_c_1485_n N_VGND_c_1833_n 0.0199786f $X=0.365 $Y=0.575 $X2=0
+ $Y2=0
cc_977 N_A_27_508#_c_1485_n N_VGND_c_1842_n 0.0162038f $X=0.365 $Y=0.575 $X2=0
+ $Y2=0
cc_978 N_A_27_508#_c_1486_n N_VGND_c_1842_n 0.0167347f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_979 N_VPWR_c_1662_n Q 0.0395687f $X=12.69 $Y=1.985 $X2=0 $Y2=0
cc_980 N_VPWR_c_1674_n Q 0.014549f $X=12.605 $Y=3.33 $X2=0 $Y2=0
cc_981 N_VPWR_c_1653_n Q 0.0119743f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_982 N_Q_c_1791_n N_VGND_c_1826_n 0.0308109f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_983 N_Q_c_1791_n N_VGND_c_1836_n 0.0145639f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_984 N_Q_c_1791_n N_VGND_c_1842_n 0.0119984f $X=12.18 $Y=0.515 $X2=0 $Y2=0

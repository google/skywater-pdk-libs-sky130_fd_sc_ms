* NGSPICE file created from sky130_fd_sc_ms__fa_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_315_75# B a_237_75# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_69_260# CIN a_315_75# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1002 a_936_75# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.65875e+12p ps=1.244e+07u
M1003 a_321_389# B a_220_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6175e+11p pd=3.07e+06u as=3.43375e+11p ps=2.86e+06u
M1004 a_69_260# CIN a_321_389# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 VPWR CIN a_512_347# VPB pshort w=1e+06u l=180000u
+  ad=2.0852e+12p pd=1.495e+07u as=6.3e+11p ps=5.26e+06u
M1006 a_512_347# a_465_249# a_69_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 COUT a_465_249# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1008 VGND CIN a_501_75# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.096e+11p ps=3.84e+06u
M1009 a_1110_347# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.35e+11p pd=5.47e+06u as=0p ps=0u
M1010 a_501_75# a_465_249# a_69_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_237_75# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_512_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_465_249# B a_919_347# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=3.25e+11p ps=2.65e+06u
M1014 VGND B a_501_75# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1100_75# B VGND VNB nlowvt w=640000u l=150000u
+  ad=8.888e+11p pd=5.27e+06u as=0p ps=0u
M1016 a_501_75# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_465_249# B a_936_75# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1018 COUT a_465_249# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1019 a_919_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1110_347# CIN a_465_249# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_69_260# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1022 VPWR A a_1110_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A a_1100_75# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1100_75# CIN a_465_249# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B a_512_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_69_260# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1027 a_220_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ms__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__nand3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.430000 2.295000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265000 1.430000 1.595000 1.550000 ;
        RECT 1.265000 1.550000 1.795000 1.680000 ;
        RECT 1.425000 1.680000 1.795000 1.950000 ;
        RECT 1.425000 1.950000 2.825000 2.120000 ;
        RECT 2.655000 1.320000 3.065000 1.650000 ;
        RECT 2.655000 1.650000 2.825000 1.950000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.735000 1.550000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.120000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.820000 1.095000 2.290000 ;
        RECT 0.565000 2.290000 2.795000 2.460000 ;
        RECT 0.565000 2.460000 0.895000 2.980000 ;
        RECT 0.925000 1.090000 2.275000 1.260000 ;
        RECT 0.925000 1.260000 1.095000 1.820000 ;
        RECT 1.515000 2.460000 1.845000 2.980000 ;
        RECT 1.945000 0.935000 2.275000 1.090000 ;
        RECT 2.525000 2.460000 2.795000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.100000  0.350000 0.350000 0.750000 ;
      RECT 0.100000  0.750000 3.260000 0.765000 ;
      RECT 0.100000  0.765000 1.370000 0.920000 ;
      RECT 0.100000  0.920000 0.430000 1.010000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.530000  0.085000 0.860000 0.580000 ;
      RECT 1.040000  0.330000 1.210000 0.595000 ;
      RECT 1.040000  0.595000 3.260000 0.750000 ;
      RECT 1.065000  2.630000 1.315000 3.245000 ;
      RECT 1.455000  0.255000 2.765000 0.425000 ;
      RECT 2.015000  2.630000 2.345000 3.245000 ;
      RECT 2.930000  0.765000 3.260000 1.150000 ;
      RECT 2.945000  0.405000 3.260000 0.595000 ;
      RECT 2.995000  1.820000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ms__nand3_2
END LIBRARY

* File: sky130_fd_sc_ms__nand3b_2.pxi.spice
* Created: Fri Aug 28 17:44:01 2020
* 
x_PM_SKY130_FD_SC_MS__NAND3B_2%A_N N_A_N_M1002_g N_A_N_M1000_g A_N N_A_N_c_72_n
+ N_A_N_c_73_n PM_SKY130_FD_SC_MS__NAND3B_2%A_N
x_PM_SKY130_FD_SC_MS__NAND3B_2%C N_C_c_103_n N_C_M1001_g N_C_M1003_g N_C_c_104_n
+ N_C_M1008_g N_C_M1013_g C C N_C_c_106_n PM_SKY130_FD_SC_MS__NAND3B_2%C
x_PM_SKY130_FD_SC_MS__NAND3B_2%A_27_94# N_A_27_94#_M1002_s N_A_27_94#_M1000_s
+ N_A_27_94#_M1004_g N_A_27_94#_c_163_n N_A_27_94#_M1006_g N_A_27_94#_M1005_g
+ N_A_27_94#_M1007_g N_A_27_94#_c_165_n N_A_27_94#_c_174_n N_A_27_94#_c_166_n
+ N_A_27_94#_c_167_n N_A_27_94#_c_168_n N_A_27_94#_c_169_n N_A_27_94#_c_176_n
+ N_A_27_94#_c_205_n N_A_27_94#_c_170_n N_A_27_94#_c_171_n
+ PM_SKY130_FD_SC_MS__NAND3B_2%A_27_94#
x_PM_SKY130_FD_SC_MS__NAND3B_2%B N_B_c_277_n N_B_M1009_g N_B_c_273_n N_B_M1010_g
+ N_B_c_274_n N_B_M1012_g N_B_c_275_n N_B_M1011_g B B B
+ PM_SKY130_FD_SC_MS__NAND3B_2%B
x_PM_SKY130_FD_SC_MS__NAND3B_2%VPWR N_VPWR_M1000_d N_VPWR_M1013_d N_VPWR_M1005_s
+ N_VPWR_M1012_s N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n
+ N_VPWR_c_325_n N_VPWR_c_326_n VPWR N_VPWR_c_327_n N_VPWR_c_315_n
+ PM_SKY130_FD_SC_MS__NAND3B_2%VPWR
x_PM_SKY130_FD_SC_MS__NAND3B_2%Y N_Y_M1006_d N_Y_M1003_s N_Y_M1004_d N_Y_M1009_d
+ N_Y_c_382_n N_Y_c_377_n N_Y_c_388_n N_Y_c_378_n N_Y_c_397_n N_Y_c_398_n
+ N_Y_c_413_n N_Y_c_379_n N_Y_c_401_n Y PM_SKY130_FD_SC_MS__NAND3B_2%Y
x_PM_SKY130_FD_SC_MS__NAND3B_2%VGND N_VGND_M1002_d N_VGND_M1008_s N_VGND_c_441_n
+ N_VGND_c_442_n VGND N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n PM_SKY130_FD_SC_MS__NAND3B_2%VGND
x_PM_SKY130_FD_SC_MS__NAND3B_2%A_206_74# N_A_206_74#_M1001_d N_A_206_74#_M1010_d
+ N_A_206_74#_c_490_n N_A_206_74#_c_487_n N_A_206_74#_c_488_n
+ N_A_206_74#_c_489_n N_A_206_74#_c_507_n N_A_206_74#_c_503_n
+ PM_SKY130_FD_SC_MS__NAND3B_2%A_206_74#
x_PM_SKY130_FD_SC_MS__NAND3B_2%A_403_54# N_A_403_54#_M1006_s N_A_403_54#_M1007_s
+ N_A_403_54#_M1011_s N_A_403_54#_c_529_n N_A_403_54#_c_530_n
+ PM_SKY130_FD_SC_MS__NAND3B_2%A_403_54#
cc_1 VNB N_A_N_M1002_g 0.0391626f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.79
cc_2 VNB N_A_N_c_72_n 0.00895418f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_3 VNB N_A_N_c_73_n 0.0306784f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.615
cc_4 VNB N_C_c_103_n 0.0152719f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.45
cc_5 VNB N_C_c_104_n 0.0171557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB C 0.00358799f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_7 VNB N_C_c_106_n 0.0794805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_94#_c_163_n 0.0182994f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_9 VNB N_A_27_94#_M1007_g 0.0185822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_94#_c_165_n 0.0266041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_94#_c_166_n 0.0022042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_94#_c_167_n 0.0104221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_94#_c_168_n 0.00531239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_94#_c_169_n 0.0110158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_94#_c_170_n 0.00729475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_94#_c_171_n 0.0492504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_273_n 0.0165885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_274_n 0.0403075f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.46
cc_19 VNB N_B_c_275_n 0.0205306f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_20 VNB B 0.0223755f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_21 VNB N_VPWR_c_315_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.00108338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_441_n 0.0093225f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_VGND_c_442_n 0.0108515f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_25 VNB N_VGND_c_443_n 0.0174171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_444_n 0.0166891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_445_n 0.0644788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_446_n 0.261576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_447_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_448_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_206_74#_c_487_n 0.00214855f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A_206_74#_c_488_n 0.00617097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_206_74#_c_489_n 0.00550897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_403_54#_c_529_n 0.0324263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_403_54#_c_530_n 0.0265018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_N_M1000_g 0.0314483f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_37 VPB N_A_N_c_72_n 0.00811757f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_38 VPB N_A_N_c_73_n 0.0241559f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.615
cc_39 VPB N_C_M1003_g 0.0219397f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_40 VPB N_C_M1013_g 0.021907f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_41 VPB C 0.00618035f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_42 VPB N_C_c_106_n 0.0058192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_27_94#_M1004_g 0.0215268f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_44 VPB N_A_27_94#_M1005_g 0.0220969f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_45 VPB N_A_27_94#_c_174_n 0.0353343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_94#_c_168_n 0.00158431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_94#_c_176_n 0.00910826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_94#_c_170_n 0.001031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_94#_c_171_n 0.0127164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B_c_277_n 0.0185999f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.45
cc_51 VPB N_B_c_274_n 0.0125841f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_52 VPB N_B_M1012_g 0.0260532f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_53 VPB B 0.0148353f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_54 VPB N_VPWR_c_316_n 0.00885173f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.78
cc_55 VPB N_VPWR_c_317_n 0.00578998f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_56 VPB N_VPWR_c_318_n 0.00914506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_319_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_320_n 0.0487491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_321_n 0.0259932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_322_n 0.00468662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_323_n 0.0202526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_324_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_325_n 0.0186844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_326_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_327_n 0.0212417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_315_n 0.0752481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_Y_c_377_n 0.00270215f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.78
cc_68 VPB N_Y_c_378_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_Y_c_379_n 0.00276474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB Y 0.00320025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 N_A_N_M1002_g N_C_c_103_n 0.021804f $X=0.48 $Y=0.79 $X2=-0.19 $Y2=-0.245
cc_72 N_A_N_M1000_g N_C_M1003_g 0.0129542f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_73 N_A_N_c_73_n C 5.01606e-19 $X=0.48 $Y=1.615 $X2=0 $Y2=0
cc_74 N_A_N_M1002_g N_C_c_106_n 0.00438823f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_75 N_A_N_c_73_n N_C_c_106_n 0.0129542f $X=0.48 $Y=1.615 $X2=0 $Y2=0
cc_76 N_A_N_M1002_g N_A_27_94#_c_165_n 4.43891e-19 $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_77 N_A_N_M1000_g N_A_27_94#_c_174_n 0.0124794f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_78 N_A_N_M1002_g N_A_27_94#_c_166_n 0.0157512f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_79 N_A_N_c_72_n N_A_27_94#_c_166_n 0.0132391f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_80 N_A_N_c_73_n N_A_27_94#_c_166_n 0.0064453f $X=0.48 $Y=1.615 $X2=0 $Y2=0
cc_81 N_A_N_c_72_n N_A_27_94#_c_167_n 0.0178519f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_82 N_A_N_c_73_n N_A_27_94#_c_167_n 0.00299816f $X=0.48 $Y=1.615 $X2=0 $Y2=0
cc_83 N_A_N_M1002_g N_A_27_94#_c_168_n 0.00598746f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_84 N_A_N_M1000_g N_A_27_94#_c_168_n 0.0088582f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_85 N_A_N_c_72_n N_A_27_94#_c_168_n 0.0247013f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_86 N_A_N_c_73_n N_A_27_94#_c_168_n 0.00547512f $X=0.48 $Y=1.615 $X2=0 $Y2=0
cc_87 N_A_N_M1000_g N_A_27_94#_c_176_n 0.0158473f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_88 N_A_N_c_72_n N_A_27_94#_c_176_n 0.0184134f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_89 N_A_N_c_73_n N_A_27_94#_c_176_n 0.00798369f $X=0.48 $Y=1.615 $X2=0 $Y2=0
cc_90 N_A_N_M1000_g N_VPWR_c_316_n 0.00308476f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_91 N_A_N_M1000_g N_VPWR_c_321_n 0.005209f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_92 N_A_N_M1000_g N_VPWR_c_315_n 0.00987008f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_93 N_A_N_M1000_g N_Y_c_377_n 6.22261e-19 $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_94 N_A_N_M1002_g N_VGND_c_441_n 0.0125975f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_95 N_A_N_M1002_g N_VGND_c_443_n 0.00421418f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_96 N_A_N_M1002_g N_VGND_c_446_n 0.00432128f $X=0.48 $Y=0.79 $X2=0 $Y2=0
cc_97 N_C_M1013_g N_A_27_94#_M1004_g 0.0262605f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_98 C N_A_27_94#_M1004_g 0.00235175f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_99 N_C_c_106_n N_A_27_94#_c_163_n 0.00235466f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_100 N_C_M1003_g N_A_27_94#_c_174_n 6.32856e-19 $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_101 N_C_M1003_g N_A_27_94#_c_168_n 0.0034271f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_102 C N_A_27_94#_c_168_n 0.0267651f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_103 N_C_c_106_n N_A_27_94#_c_168_n 0.0076931f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_104 N_C_c_103_n N_A_27_94#_c_169_n 0.00771139f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_105 N_C_c_104_n N_A_27_94#_c_169_n 0.00671798f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_106 C N_A_27_94#_c_169_n 0.051126f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_107 N_C_c_106_n N_A_27_94#_c_169_n 0.0310057f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_108 N_C_M1003_g N_A_27_94#_c_176_n 0.00149833f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_109 N_C_c_103_n N_A_27_94#_c_205_n 0.00184514f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_110 N_C_c_106_n N_A_27_94#_c_205_n 0.00108279f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_111 C N_A_27_94#_c_170_n 0.0168746f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_112 N_C_c_106_n N_A_27_94#_c_170_n 0.0030545f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_113 C N_A_27_94#_c_171_n 0.00104708f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_C_c_106_n N_A_27_94#_c_171_n 0.0183764f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_115 N_C_M1003_g N_VPWR_c_316_n 0.00312369f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_116 N_C_M1013_g N_VPWR_c_317_n 0.00342668f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_117 N_C_M1003_g N_VPWR_c_323_n 0.005209f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_118 N_C_M1013_g N_VPWR_c_323_n 0.005209f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_119 N_C_M1003_g N_VPWR_c_315_n 0.00982981f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_120 N_C_M1013_g N_VPWR_c_315_n 0.00982602f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_121 N_C_M1003_g N_Y_c_382_n 0.00308089f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_122 N_C_M1013_g N_Y_c_382_n 8.84614e-19 $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_123 C N_Y_c_382_n 0.0270344f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_124 N_C_c_106_n N_Y_c_382_n 8.24477e-19 $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_125 N_C_M1003_g N_Y_c_377_n 0.0120585f $X=1.2 $Y=2.4 $X2=0 $Y2=0
cc_126 N_C_M1013_g N_Y_c_377_n 0.0117745f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_127 N_C_M1013_g N_Y_c_388_n 0.0131783f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_128 C N_Y_c_388_n 0.011149f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_C_c_103_n N_VGND_c_441_n 0.00556327f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_130 N_C_c_103_n N_VGND_c_442_n 3.69172e-19 $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_131 N_C_c_104_n N_VGND_c_442_n 0.00769205f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_132 N_C_c_103_n N_VGND_c_444_n 0.00433834f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_133 N_C_c_104_n N_VGND_c_444_n 0.00281141f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_134 N_C_c_103_n N_VGND_c_446_n 0.00825089f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_135 N_C_c_104_n N_VGND_c_446_n 0.00365066f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_136 N_C_c_103_n N_A_206_74#_c_490_n 0.00221999f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_137 N_C_c_106_n N_A_206_74#_c_490_n 6.05025e-19 $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_138 N_C_c_103_n N_A_206_74#_c_487_n 0.00498672f $X=0.955 $Y=1.185 $X2=0 $Y2=0
cc_139 N_C_c_104_n N_A_206_74#_c_487_n 2.93125e-19 $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_140 N_C_c_104_n N_A_206_74#_c_488_n 0.0118272f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_141 N_C_c_106_n N_A_206_74#_c_488_n 0.00166748f $X=1.615 $Y=1.515 $X2=0 $Y2=0
cc_142 N_C_c_104_n N_A_206_74#_c_489_n 0.00212344f $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_143 N_C_c_104_n N_A_403_54#_c_529_n 4.19228e-19 $X=1.385 $Y=1.185 $X2=0 $Y2=0
cc_144 N_A_27_94#_M1007_g N_B_c_273_n 0.0272472f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_145 N_A_27_94#_M1005_g N_B_c_274_n 0.0255282f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_27_94#_M1007_g N_B_c_274_n 0.0122044f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_147 N_A_27_94#_M1005_g B 4.0143e-19 $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_27_94#_M1007_g B 0.00344966f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_149 N_A_27_94#_c_168_n N_VPWR_M1000_d 0.00140859f $X=0.805 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_27_94#_c_176_n N_VPWR_M1000_d 0.00263856f $X=0.805 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_27_94#_c_174_n N_VPWR_c_316_n 0.0238827f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_152 N_A_27_94#_c_176_n N_VPWR_c_316_n 0.00386873f $X=0.805 $Y=2.035 $X2=0
+ $Y2=0
cc_153 N_A_27_94#_M1004_g N_VPWR_c_317_n 0.0130546f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_27_94#_M1005_g N_VPWR_c_317_n 5.60811e-19 $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_27_94#_M1005_g N_VPWR_c_318_n 0.00670269f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_27_94#_c_174_n N_VPWR_c_321_n 0.014549f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_157 N_A_27_94#_M1004_g N_VPWR_c_325_n 0.00460063f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_27_94#_M1005_g N_VPWR_c_325_n 0.005209f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_27_94#_M1004_g N_VPWR_c_315_n 0.00908554f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_27_94#_M1005_g N_VPWR_c_315_n 0.00984153f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_27_94#_c_174_n N_VPWR_c_315_n 0.0119743f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_162 N_A_27_94#_c_176_n N_Y_c_382_n 0.00794526f $X=0.805 $Y=2.035 $X2=0 $Y2=0
cc_163 N_A_27_94#_M1004_g N_Y_c_377_n 8.00171e-19 $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_27_94#_c_174_n N_Y_c_377_n 0.00435609f $X=0.47 $Y=2.815 $X2=0 $Y2=0
cc_165 N_A_27_94#_M1004_g N_Y_c_388_n 0.0151885f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_27_94#_c_170_n N_Y_c_388_n 0.0141353f $X=2.19 $Y=1.175 $X2=0 $Y2=0
cc_167 N_A_27_94#_c_171_n N_Y_c_388_n 3.54977e-19 $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A_27_94#_M1005_g N_Y_c_378_n 0.0127744f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_27_94#_c_171_n N_Y_c_397_n 0.00466734f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A_27_94#_M1005_g N_Y_c_398_n 0.0130547f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_27_94#_c_171_n N_Y_c_398_n 0.00358503f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A_27_94#_M1005_g N_Y_c_379_n 8.96373e-19 $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A_27_94#_c_163_n N_Y_c_401_n 0.00600238f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_174 N_A_27_94#_M1007_g N_Y_c_401_n 0.00207245f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_175 N_A_27_94#_c_170_n N_Y_c_401_n 0.0051356f $X=2.19 $Y=1.175 $X2=0 $Y2=0
cc_176 N_A_27_94#_M1004_g Y 0.00332508f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_27_94#_c_163_n Y 0.00157436f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_178 N_A_27_94#_M1005_g Y 0.00807389f $X=2.645 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_27_94#_M1007_g Y 0.00539959f $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_180 N_A_27_94#_c_170_n Y 0.0319153f $X=2.19 $Y=1.175 $X2=0 $Y2=0
cc_181 N_A_27_94#_c_171_n Y 0.016958f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A_27_94#_c_166_n N_VGND_M1002_d 0.00116505f $X=0.72 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_27_94#_c_205_n N_VGND_M1002_d 0.00112241f $X=0.805 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_27_94#_c_169_n N_VGND_M1008_s 0.00205663f $X=2.025 $Y=1.175 $X2=0
+ $Y2=0
cc_185 N_A_27_94#_c_165_n N_VGND_c_441_n 0.0168919f $X=0.265 $Y=0.615 $X2=0
+ $Y2=0
cc_186 N_A_27_94#_c_166_n N_VGND_c_441_n 0.0100896f $X=0.72 $Y=1.175 $X2=0 $Y2=0
cc_187 N_A_27_94#_c_205_n N_VGND_c_441_n 0.00855018f $X=0.805 $Y=1.175 $X2=0
+ $Y2=0
cc_188 N_A_27_94#_c_163_n N_VGND_c_442_n 0.00241358f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_189 N_A_27_94#_c_165_n N_VGND_c_443_n 0.00787252f $X=0.265 $Y=0.615 $X2=0
+ $Y2=0
cc_190 N_A_27_94#_c_163_n N_VGND_c_445_n 7.84925e-19 $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_191 N_A_27_94#_M1007_g N_VGND_c_445_n 7.84925e-19 $X=2.85 $Y=0.87 $X2=0 $Y2=0
cc_192 N_A_27_94#_c_165_n N_VGND_c_446_n 0.0085887f $X=0.265 $Y=0.615 $X2=0
+ $Y2=0
cc_193 N_A_27_94#_c_169_n N_A_206_74#_M1001_d 0.00176461f $X=2.025 $Y=1.175
+ $X2=-0.19 $Y2=-0.245
cc_194 N_A_27_94#_c_169_n N_A_206_74#_c_490_n 0.0151918f $X=2.025 $Y=1.175 $X2=0
+ $Y2=0
cc_195 N_A_27_94#_c_169_n N_A_206_74#_c_488_n 0.0479995f $X=2.025 $Y=1.175 $X2=0
+ $Y2=0
cc_196 N_A_27_94#_c_163_n N_A_206_74#_c_489_n 0.00301228f $X=2.42 $Y=1.35 $X2=0
+ $Y2=0
cc_197 N_A_27_94#_c_170_n N_A_206_74#_c_489_n 0.00682868f $X=2.19 $Y=1.175 $X2=0
+ $Y2=0
cc_198 N_A_27_94#_c_171_n N_A_206_74#_c_489_n 3.24197e-19 $X=2.645 $Y=1.515
+ $X2=0 $Y2=0
cc_199 N_A_27_94#_c_163_n N_A_206_74#_c_503_n 0.0159728f $X=2.42 $Y=1.35 $X2=0
+ $Y2=0
cc_200 N_A_27_94#_M1007_g N_A_206_74#_c_503_n 0.0149272f $X=2.85 $Y=0.87 $X2=0
+ $Y2=0
cc_201 N_A_27_94#_c_170_n N_A_206_74#_c_503_n 0.00950299f $X=2.19 $Y=1.175 $X2=0
+ $Y2=0
cc_202 N_A_27_94#_c_171_n N_A_206_74#_c_503_n 0.001279f $X=2.645 $Y=1.515 $X2=0
+ $Y2=0
cc_203 N_A_27_94#_c_170_n N_A_403_54#_M1006_s 0.0033664f $X=2.19 $Y=1.175
+ $X2=-0.19 $Y2=-0.245
cc_204 N_A_27_94#_c_163_n N_A_403_54#_c_529_n 0.0103526f $X=2.42 $Y=1.35 $X2=0
+ $Y2=0
cc_205 N_A_27_94#_M1007_g N_A_403_54#_c_529_n 0.00963483f $X=2.85 $Y=0.87 $X2=0
+ $Y2=0
cc_206 N_B_c_277_n N_VPWR_c_318_n 0.0103551f $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_207 N_B_c_277_n N_VPWR_c_320_n 7.87307e-19 $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_208 N_B_M1012_g N_VPWR_c_320_n 0.0177701f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_209 B N_VPWR_c_320_n 0.0254127f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_210 N_B_c_277_n N_VPWR_c_327_n 0.005209f $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_211 N_B_M1012_g N_VPWR_c_327_n 0.00460063f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_212 N_B_c_277_n N_VPWR_c_315_n 0.0098563f $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_213 N_B_M1012_g N_VPWR_c_315_n 0.00909135f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B_c_277_n N_Y_c_378_n 8.77012e-19 $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_215 N_B_c_277_n N_Y_c_397_n 0.0138786f $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_216 B N_Y_c_397_n 0.0255673f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_217 N_B_c_277_n N_Y_c_413_n 8.84614e-19 $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_218 N_B_c_274_n N_Y_c_413_n 9.18264e-19 $X=3.815 $Y=1.68 $X2=0 $Y2=0
cc_219 B N_Y_c_413_n 0.0251484f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B_c_277_n N_Y_c_379_n 0.0135087f $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_221 N_B_M1012_g N_Y_c_379_n 2.01597e-19 $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B_c_273_n N_Y_c_401_n 8.93946e-19 $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_223 N_B_c_277_n Y 0.00316694f $X=3.305 $Y=1.77 $X2=0 $Y2=0
cc_224 N_B_c_274_n Y 4.9668e-19 $X=3.815 $Y=1.68 $X2=0 $Y2=0
cc_225 B Y 0.0313541f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_226 N_B_c_273_n N_VGND_c_445_n 7.84925e-19 $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_227 N_B_c_275_n N_VGND_c_445_n 7.84925e-19 $X=3.84 $Y=1.35 $X2=0 $Y2=0
cc_228 N_B_c_273_n N_A_206_74#_c_507_n 0.0187719f $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_229 N_B_c_274_n N_A_206_74#_c_507_n 0.00484393f $X=3.815 $Y=1.68 $X2=0 $Y2=0
cc_230 N_B_c_275_n N_A_206_74#_c_507_n 0.00611925f $X=3.84 $Y=1.35 $X2=0 $Y2=0
cc_231 B N_A_206_74#_c_507_n 0.0574195f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B_c_273_n N_A_403_54#_c_529_n 0.00963483f $X=3.41 $Y=1.35 $X2=0 $Y2=0
cc_233 N_B_c_275_n N_A_403_54#_c_529_n 0.0140521f $X=3.84 $Y=1.35 $X2=0 $Y2=0
cc_234 B N_A_403_54#_c_530_n 0.020209f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_VPWR_c_316_n N_Y_c_377_n 0.0253838f $X=0.95 $Y=2.455 $X2=0 $Y2=0
cc_236 N_VPWR_c_317_n N_Y_c_377_n 0.0271924f $X=1.97 $Y=2.41 $X2=0 $Y2=0
cc_237 N_VPWR_c_323_n N_Y_c_377_n 0.0164702f $X=1.805 $Y=3.33 $X2=0 $Y2=0
cc_238 N_VPWR_c_315_n N_Y_c_377_n 0.0134964f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_M1013_d N_Y_c_388_n 0.00941308f $X=1.785 $Y=1.84 $X2=0 $Y2=0
cc_240 N_VPWR_c_317_n N_Y_c_388_n 0.0189268f $X=1.97 $Y=2.41 $X2=0 $Y2=0
cc_241 N_VPWR_c_317_n N_Y_c_378_n 0.0234083f $X=1.97 $Y=2.41 $X2=0 $Y2=0
cc_242 N_VPWR_c_318_n N_Y_c_378_n 0.0220532f $X=2.955 $Y=2.41 $X2=0 $Y2=0
cc_243 N_VPWR_c_325_n N_Y_c_378_n 0.0109793f $X=2.79 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_315_n N_Y_c_378_n 0.00901959f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_M1005_s N_Y_c_397_n 0.0122207f $X=2.735 $Y=1.84 $X2=0 $Y2=0
cc_246 N_VPWR_c_318_n N_Y_c_398_n 0.0265313f $X=2.955 $Y=2.41 $X2=0 $Y2=0
cc_247 N_VPWR_c_318_n N_Y_c_379_n 0.0404966f $X=2.955 $Y=2.41 $X2=0 $Y2=0
cc_248 N_VPWR_c_320_n N_Y_c_379_n 0.0315827f $X=4.04 $Y=2.035 $X2=0 $Y2=0
cc_249 N_VPWR_c_327_n N_Y_c_379_n 0.014549f $X=3.875 $Y=3.33 $X2=0 $Y2=0
cc_250 N_VPWR_c_315_n N_Y_c_379_n 0.0119743f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_M1005_s Y 0.00168479f $X=2.735 $Y=1.84 $X2=0 $Y2=0
cc_252 N_Y_M1006_d N_A_206_74#_c_503_n 0.00337414f $X=2.495 $Y=0.5 $X2=0 $Y2=0
cc_253 N_Y_c_401_n N_A_206_74#_c_503_n 0.0168934f $X=2.635 $Y=1.095 $X2=0 $Y2=0
cc_254 N_VGND_c_441_n N_A_206_74#_c_490_n 0.01223f $X=0.695 $Y=0.725 $X2=0 $Y2=0
cc_255 N_VGND_c_441_n N_A_206_74#_c_487_n 0.0296545f $X=0.695 $Y=0.725 $X2=0
+ $Y2=0
cc_256 N_VGND_c_442_n N_A_206_74#_c_487_n 0.0104546f $X=1.6 $Y=0.495 $X2=0 $Y2=0
cc_257 N_VGND_c_444_n N_A_206_74#_c_487_n 0.0118323f $X=1.435 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_446_n N_A_206_74#_c_487_n 0.00911095f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_M1008_s N_A_206_74#_c_488_n 0.00433153f $X=1.46 $Y=0.37 $X2=0
+ $Y2=0
cc_260 N_VGND_c_442_n N_A_206_74#_c_488_n 0.0212697f $X=1.6 $Y=0.495 $X2=0 $Y2=0
cc_261 N_VGND_c_444_n N_A_206_74#_c_488_n 0.00197156f $X=1.435 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_445_n N_A_206_74#_c_488_n 0.0024506f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_446_n N_A_206_74#_c_488_n 0.00976958f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_264 N_VGND_c_445_n N_A_206_74#_c_489_n 6.97459e-19 $X=4.08 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_446_n N_A_206_74#_c_489_n 0.00468475f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_442_n N_A_403_54#_c_529_n 0.0128051f $X=1.6 $Y=0.495 $X2=0 $Y2=0
cc_267 N_VGND_c_445_n N_A_403_54#_c_529_n 0.0990761f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_446_n N_A_403_54#_c_529_n 0.0808667f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_269 N_A_206_74#_c_489_n N_A_403_54#_M1006_s 0.00147525f $X=2.105 $Y=0.795
+ $X2=-0.19 $Y2=-0.245
cc_270 N_A_206_74#_c_503_n N_A_403_54#_M1006_s 0.00484861f $X=2.97 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_271 N_A_206_74#_c_507_n N_A_403_54#_M1007_s 0.00950662f $X=3.625 $Y=0.755
+ $X2=0 $Y2=0
cc_272 N_A_206_74#_c_489_n N_A_403_54#_c_529_n 0.11551f $X=2.105 $Y=0.795 $X2=0
+ $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__nor4_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nor4_1 A B C D VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.7975e+11p ps=6.9e+06u
M1001 a_147_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=3.136e+11p ps=2.8e+06u
M1002 a_345_368# C a_231_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=4.368e+11p ps=3.02e+06u
M1003 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_231_368# B a_147_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y D a_345_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1007 VGND D Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a311o_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__a311o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.450000 2.835000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.450000 2.295000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.260000 1.795000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.260000 3.715000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.440000 4.215000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.550000 0.995000 2.060000 ;
        RECT 0.730000 0.350000 1.060000 0.750000 ;
        RECT 0.730000 0.750000 0.995000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.105000  1.350000 0.435000 2.230000 ;
      RECT 0.105000  2.230000 1.335000 2.400000 ;
      RECT 0.215000  2.570000 0.545000 3.245000 ;
      RECT 0.300000  0.085000 0.550000 1.130000 ;
      RECT 1.115000  2.570000 1.445000 3.245000 ;
      RECT 1.165000  0.920000 4.040000 1.090000 ;
      RECT 1.165000  1.090000 1.335000 1.950000 ;
      RECT 1.165000  1.950000 4.035000 2.120000 ;
      RECT 1.165000  2.120000 1.335000 2.230000 ;
      RECT 1.230000  0.085000 1.630000 0.750000 ;
      RECT 1.635000  2.290000 3.165000 2.570000 ;
      RECT 1.635000  2.570000 1.965000 2.980000 ;
      RECT 2.135000  2.740000 2.665000 3.245000 ;
      RECT 2.630000  0.350000 3.000000 0.920000 ;
      RECT 2.835000  2.570000 3.165000 2.980000 ;
      RECT 3.170000  0.085000 3.540000 0.750000 ;
      RECT 3.705000  2.120000 4.035000 2.980000 ;
      RECT 3.710000  0.350000 4.040000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__a311o_2

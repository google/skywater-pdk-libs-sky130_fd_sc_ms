* NGSPICE file created from sky130_fd_sc_ms__sdfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_353_93# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=2.8826e+12p ps=2.42e+07u
M1001 a_1906_424# a_977_243# VPWR VPB pshort w=840000u l=180000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1002 a_305_119# D a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.129e+11p ps=3.17e+06u
M1003 a_197_119# a_867_82# a_1162_497# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 VGND RESET_B a_1579_258# VNB nlowvt w=420000u l=150000u
+  ad=2.11888e+12p pd=1.742e+07u as=1.197e+11p ps=1.41e+06u
M1005 a_977_243# a_1162_497# a_1434_78# VNB nlowvt w=550000u l=150000u
+  ad=2.09e+11p pd=1.86e+06u as=5.1045e+11p ps=4.25e+06u
M1006 a_119_119# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 Q_N a_2133_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 VPWR SCD a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.552e+11p ps=3.67e+06u
M1009 a_2392_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.947e+11p pd=4.37e+06u as=0p ps=0u
M1010 VGND a_2133_410# a_2164_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1011 a_197_119# D a_215_464# VPB pshort w=640000u l=180000u
+  ad=3.84e+11p pd=3.76e+06u as=1.536e+11p ps=1.76e+06u
M1012 VPWR a_2133_410# a_2091_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 a_27_464# a_353_93# a_197_119# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1162_497# a_867_82# a_1084_497# VPB pshort w=420000u l=180000u
+  ad=2.107e+11p pd=1.99e+06u as=8.82e+10p ps=1.26e+06u
M1015 a_1954_119# a_867_82# a_1906_424# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=0p ps=0u
M1016 VPWR a_2133_410# a_3078_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1017 a_197_119# a_662_82# a_1162_497# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND CLK_N a_662_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1019 a_867_82# a_662_82# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.219e+11p pd=2.35e+06u as=0p ps=0u
M1020 a_1162_497# a_662_82# a_1151_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 a_353_93# SCE VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1022 Q a_3078_384# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1023 a_2512_392# a_1579_258# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1024 VGND a_2133_410# a_3078_384# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1025 a_1151_119# a_977_243# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND SET_B a_1434_78# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1954_119# a_662_82# a_1876_119# VNB nlowvt w=550000u l=150000u
+  ad=4.807e+11p pd=2.9e+06u as=1.32e+11p ps=1.58e+06u
M1028 VPWR SET_B a_2133_410# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1029 VPWR CLK_N a_662_82# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1030 a_2091_508# a_662_82# a_1954_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1084_497# a_977_243# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2392_74# a_1954_119# a_2133_410# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.812e+11p ps=2.24e+06u
M1033 a_867_82# a_662_82# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1034 a_197_119# SCE a_119_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_353_93# a_305_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_215_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1531_424# a_1162_497# a_977_243# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=6.09e+11p ps=4.81e+06u
M1038 Q a_3078_384# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1039 a_2133_410# a_1579_258# a_2392_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_2164_119# a_867_82# a_1954_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_1579_258# a_1531_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1876_119# a_977_243# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Q_N a_2133_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1044 a_977_243# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1434_78# a_1579_258# a_977_243# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2133_410# a_1954_119# a_2512_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR RESET_B a_1579_258# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.529e+11p ps=3.68e+06u
.ends


* NGSPICE file created from sky130_fd_sc_ms__sdfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1370_290# a_1223_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=3.2444e+12p ps=2.643e+07u
M1001 VPWR a_2607_392# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1002 a_2000_74# a_852_119# a_1790_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.33e+11p ps=3.08e+06u
M1003 VGND RESET_B a_223_79# VNB nlowvt w=420000u l=150000u
+  ad=2.20072e+12p pd=1.854e+07u as=2.751e+11p ps=2.99e+06u
M1004 a_1790_74# a_852_119# a_1370_290# VPB pshort w=1e+06u l=180000u
+  ad=3.816e+11p pd=3.22e+06u as=0p ps=0u
M1005 Q_N a_1790_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 a_388_79# D a_310_464# VPB pshort w=640000u l=180000u
+  ad=6.96975e+11p pd=5.83e+06u as=1.536e+11p ps=1.76e+06u
M1007 a_1370_290# a_1223_119# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1008 VPWR a_1790_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR SCE a_27_79# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 a_2607_392# a_1790_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1011 VGND RESET_B a_1401_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1012 a_310_79# a_27_79# a_223_79# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1013 a_223_79# SCD a_547_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1014 a_1223_119# a_852_119# a_388_79# VNB nlowvt w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=3.906e+11p ps=3.54e+06u
M1015 a_1323_119# a_1025_119# a_1223_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_2006_373# a_1790_74# a_2158_74# VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1017 a_1790_74# a_1025_119# a_1370_290# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_2607_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1019 VPWR CLK a_852_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1020 VPWR a_1370_290# a_1328_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 VGND CLK a_852_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.95675e+11p ps=2.05e+06u
M1022 VPWR a_2006_373# a_1958_471# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 a_2006_373# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1024 a_2158_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q_N a_1790_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1026 a_388_79# D a_310_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_541_483# a_27_79# a_388_79# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1028 VPWR a_1790_74# a_2006_373# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_2607_392# a_1790_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1030 VGND SCE a_27_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1031 a_547_79# SCE a_388_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1223_119# a_1025_119# a_388_79# VPB pshort w=420000u l=180000u
+  ad=2.247e+11p pd=2.75e+06u as=0p ps=0u
M1033 a_1025_119# a_852_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1034 a_1223_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_388_79# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1025_119# a_852_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1037 VGND a_1790_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_2607_392# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_310_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1328_457# a_852_119# a_1223_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR SCD a_541_483# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1958_471# a_1025_119# a_1790_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1401_119# a_1370_290# a_1323_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 Q a_2607_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND a_2006_373# a_2000_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


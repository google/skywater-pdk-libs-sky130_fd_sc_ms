# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o2bb2a_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o2bb2a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.420000 1.315000 1.710000 ;
        RECT 1.085000 1.710000 1.315000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.430000 1.835000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.180000 4.215000 1.510000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.510000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.455000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.425000  1.300000 0.795000 1.630000 ;
      RECT 0.615000  1.950000 0.945000 3.245000 ;
      RECT 0.625000  0.085000 1.120000 0.910000 ;
      RECT 0.625000  1.080000 1.460000 1.250000 ;
      RECT 0.625000  1.250000 0.795000 1.300000 ;
      RECT 1.150000  1.950000 2.380000 2.280000 ;
      RECT 1.290000  0.255000 2.815000 0.425000 ;
      RECT 1.290000  0.425000 1.460000 1.080000 ;
      RECT 1.630000  0.595000 1.880000 1.090000 ;
      RECT 1.630000  1.090000 2.380000 1.260000 ;
      RECT 1.655000  2.450000 2.820000 3.245000 ;
      RECT 2.050000  1.260000 2.380000 1.950000 ;
      RECT 2.485000  0.425000 2.815000 0.920000 ;
      RECT 2.645000  0.920000 2.815000 1.900000 ;
      RECT 2.645000  1.900000 3.320000 2.070000 ;
      RECT 2.990000  2.070000 3.320000 2.780000 ;
      RECT 2.995000  0.340000 3.245000 0.840000 ;
      RECT 2.995000  0.840000 4.205000 1.010000 ;
      RECT 3.415000  0.085000 3.745000 0.670000 ;
      RECT 3.870000  1.900000 4.200000 3.245000 ;
      RECT 3.955000  0.340000 4.205000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__o2bb2a_1

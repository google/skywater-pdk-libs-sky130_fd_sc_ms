* File: sky130_fd_sc_ms__nor4_1.spice
* Created: Fri Aug 28 17:49:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4_1.pex.spice"
.subckt sky130_fd_sc_ms__nor4_1  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_Y_M1000_d VNB NLOWVT L=0.15 W=0.74 AD=0.1924
+ AS=0.1036 PD=1.26 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1924 PD=1.02 PS=1.26 NRD=0 NRS=27.564 M=1 R=4.93333 SA=75001.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_D_M1007_g N_Y_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.23225 AS=0.1036 PD=2.19 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_147_368# N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90001.8
+ A=0.2016 P=2.6 MULT=1
MM1005 A_231_368# N_B_M1005_g A_147_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1002 A_345_368# N_C_M1002_g A_231_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=24.6053 M=1 R=6.22222 SA=90001.2
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_D_M1006_g A_345_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90001.8 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__nor4_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_547_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_1235_119# a_837_119# a_1339_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X2 a_225_81# a_27_74# a_312_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 Q a_2495_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VGND a_837_119# a_1037_119# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_1235_119# a_1037_119# a_1354_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_837_119# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VPWR a_1824_74# a_2495_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 a_2082_446# a_1824_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X9 VPWR a_837_119# a_1037_119# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X11 a_517_483# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X12 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_2040_508# a_2082_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X14 a_390_81# SCE a_547_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 Q a_2495_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_1339_457# a_1383_349# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X17 a_390_81# a_837_119# a_1235_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_1383_349# a_837_119# a_1824_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X19 VPWR a_2495_392# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 VGND a_2495_392# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR RESET_B a_1235_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X22 a_1824_74# a_1037_119# a_2040_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X23 a_1383_349# a_1037_119# a_1824_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_2078_74# a_2082_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_1824_74# a_837_119# a_2078_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_390_81# a_27_74# a_517_483# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X27 VPWR RESET_B a_390_81# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X28 a_837_119# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VPWR a_1235_119# a_1383_349# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X30 VGND a_1824_74# a_2495_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 a_390_81# a_1037_119# a_1235_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X32 VPWR RESET_B a_2082_446# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X33 a_1354_119# a_1383_349# a_1432_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 VGND RESET_B a_2242_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 a_1432_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 a_2242_74# a_1824_74# a_2082_446# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VGND a_1235_119# a_1383_349# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 VPWR SCE a_343_483# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X39 a_343_483# D a_390_81# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X40 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X41 a_312_81# D a_390_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

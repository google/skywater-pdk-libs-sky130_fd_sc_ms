* File: sky130_fd_sc_ms__a2bb2oi_1.spice
* Created: Wed Sep  2 11:54:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2bb2oi_1.pex.spice"
.subckt sky130_fd_sc_ms__a2bb2oi_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1000 N_A_126_112#_M1000_d N_A1_N_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.5 A=0.0825 P=1.4 MULT=1
MM1009 N_VGND_M1009_d N_A2_N_M1009_g N_A_126_112#_M1000_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.209064 AS=0.077 PD=1.31318 PS=0.83 NRD=70.932 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75002 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_126_112#_M1001_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.281286 PD=1.02 PS=1.76682 NRD=0 NRS=52.716 M=1 R=4.93333
+ SA=75001.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 A_488_74# N_B2_M1007_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g A_488_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1961
+ AS=0.1184 PD=2.01 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75002.1 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1008 A_120_392# N_A1_N_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1 AD=0.105
+ AS=0.26 PD=1.21 PS=2.52 NRD=9.8303 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90000.6
+ A=0.18 P=2.36 MULT=1
MM1002 N_A_126_112#_M1002_d N_A2_N_M1002_g A_120_392# VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_402_368#_M1004_d N_A_126_112#_M1004_g N_Y_M1004_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1006_d N_B2_M1006_g N_A_402_368#_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.168 AS=0.1512 PD=1.42 PS=1.39 NRD=1.7533 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1005 N_A_402_368#_M1005_d N_B1_M1005_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.168 PD=2.76 PS=1.42 NRD=0 NRS=1.7533 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__a2bb2oi_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3b_1 A B C_N VGND VNB VPB VPWR Y
M1000 Y a_27_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.477e+11p pd=4.17e+06u as=5.8515e+11p ps=4.58e+06u
M1001 Y a_27_112# a_347_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=4.368e+11p ps=3.02e+06u
M1002 a_347_368# B a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.688e+11p ps=2.72e+06u
M1003 a_263_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.06e+11p ps=3.02e+06u
M1004 VGND C_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.695e+11p ps=2.08e+06u
M1005 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1007 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

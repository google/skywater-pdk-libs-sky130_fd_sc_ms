* File: sky130_fd_sc_ms__and3_1.pxi.spice
* Created: Wed Sep  2 11:57:38 2020
* 
x_PM_SKY130_FD_SC_MS__AND3_1%A N_A_M1006_g N_A_c_57_n N_A_M1001_g N_A_c_59_n
+ N_A_c_60_n A N_A_c_62_n PM_SKY130_FD_SC_MS__AND3_1%A
x_PM_SKY130_FD_SC_MS__AND3_1%B N_B_M1003_g N_B_M1002_g B B N_B_c_99_n
+ N_B_c_100_n PM_SKY130_FD_SC_MS__AND3_1%B
x_PM_SKY130_FD_SC_MS__AND3_1%C N_C_M1005_g N_C_M1004_g C N_C_c_145_n
+ PM_SKY130_FD_SC_MS__AND3_1%C
x_PM_SKY130_FD_SC_MS__AND3_1%A_27_398# N_A_27_398#_M1001_s N_A_27_398#_M1006_s
+ N_A_27_398#_M1003_d N_A_27_398#_c_181_n N_A_27_398#_M1007_g
+ N_A_27_398#_M1000_g N_A_27_398#_c_182_n N_A_27_398#_c_187_n
+ N_A_27_398#_c_188_n N_A_27_398#_c_189_n N_A_27_398#_c_190_n
+ N_A_27_398#_c_191_n N_A_27_398#_c_192_n N_A_27_398#_c_193_n
+ N_A_27_398#_c_183_n N_A_27_398#_c_184_n PM_SKY130_FD_SC_MS__AND3_1%A_27_398#
x_PM_SKY130_FD_SC_MS__AND3_1%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_262_n
+ N_VPWR_c_263_n VPWR N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n
+ N_VPWR_c_261_n N_VPWR_c_268_n N_VPWR_c_269_n PM_SKY130_FD_SC_MS__AND3_1%VPWR
x_PM_SKY130_FD_SC_MS__AND3_1%X N_X_M1007_d N_X_M1000_d N_X_c_300_n N_X_c_301_n X
+ X X X N_X_c_302_n PM_SKY130_FD_SC_MS__AND3_1%X
x_PM_SKY130_FD_SC_MS__AND3_1%VGND N_VGND_M1004_d N_VGND_c_324_n N_VGND_c_325_n
+ N_VGND_c_326_n VGND N_VGND_c_327_n N_VGND_c_328_n
+ PM_SKY130_FD_SC_MS__AND3_1%VGND
cc_1 VNB N_A_M1006_g 0.00748651f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_2 VNB N_A_c_57_n 0.0397668f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.57
cc_3 VNB N_A_M1001_g 0.0144312f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_4 VNB N_A_c_59_n 0.0116103f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.545
cc_5 VNB N_A_c_60_n 0.0424882f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_6 VNB A 0.00759927f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.47
cc_7 VNB N_A_c_62_n 0.0208892f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.462
cc_8 VNB B 0.00357895f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.395
cc_9 VNB N_B_c_99_n 0.0200684f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.412
cc_10 VNB N_B_c_100_n 0.016463f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_11 VNB N_C_M1004_g 0.0258025f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.57
cc_12 VNB C 0.00338947f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_13 VNB N_C_c_145_n 0.0254582f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.545
cc_14 VNB N_A_27_398#_c_181_n 0.0220597f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_15 VNB N_A_27_398#_c_182_n 0.0376576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_398#_c_183_n 0.00166255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_398#_c_184_n 0.0337128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_261_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_X_c_300_n 0.0234698f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1
cc_20 VNB N_X_c_301_n 0.0184679f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_21 VNB N_X_c_302_n 0.023805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_324_n 0.0191361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_325_n 0.0444379f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.395
cc_24 VNB N_VGND_c_326_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.545
cc_25 VNB N_VGND_c_327_n 0.0273666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_328_n 0.202229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A_M1006_g 0.0386363f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_28 VPB N_B_M1003_g 0.0258112f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.545
cc_29 VPB B 0.00357649f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.395
cc_30 VPB N_B_c_99_n 0.0107534f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=0.412
cc_31 VPB N_C_M1005_g 0.0268368f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.545
cc_32 VPB C 0.00203124f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1
cc_33 VPB N_C_c_145_n 0.016466f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.545
cc_34 VPB N_A_27_398#_M1000_g 0.0285547f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_35 VPB N_A_27_398#_c_182_n 0.0121764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_27_398#_c_187_n 0.0309311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_27_398#_c_188_n 0.00913152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_398#_c_189_n 0.0028561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_398#_c_190_n 0.00968866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_398#_c_191_n 0.0026353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_398#_c_192_n 0.00719737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_398#_c_193_n 0.00499084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_27_398#_c_183_n 7.30623e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_27_398#_c_184_n 0.00777352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_262_n 0.0170576f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1
cc_46 VPB N_VPWR_c_263_n 0.00948708f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=0.412
cc_47 VPB N_VPWR_c_264_n 0.0197293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_265_n 0.0181128f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=0.462
cc_49 VPB N_VPWR_c_266_n 0.017913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_261_n 0.0641378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_268_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_269_n 0.0140183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB X 0.00529771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB X 0.0395491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_X_c_302_n 0.00895792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 N_A_M1006_g N_B_M1003_g 0.0234122f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_57 N_A_M1006_g B 9.39698e-19 $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_58 N_A_M1001_g B 0.00222717f $X=0.53 $Y=1 $X2=0 $Y2=0
cc_59 N_A_c_59_n B 4.14418e-19 $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_60 A B 0.00728026f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_61 N_A_c_62_n B 0.00666142f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_62 N_A_M1006_g N_B_c_99_n 0.0103774f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_63 N_A_c_59_n N_B_c_99_n 0.00587736f $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_64 N_A_c_57_n N_B_c_100_n 0.0011105f $X=0.53 $Y=0.57 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_B_c_100_n 0.0251307f $X=0.53 $Y=1 $X2=0 $Y2=0
cc_66 A N_B_c_100_n 0.00718878f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_67 N_A_c_62_n N_B_c_100_n 0.00365215f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_68 N_A_c_57_n N_C_M1004_g 7.00286e-19 $X=0.53 $Y=0.57 $X2=0 $Y2=0
cc_69 A N_C_M1004_g 0.00212205f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_70 N_A_M1006_g N_A_27_398#_c_182_n 0.0162666f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_71 N_A_M1001_g N_A_27_398#_c_182_n 0.0179899f $X=0.53 $Y=1 $X2=0 $Y2=0
cc_72 N_A_c_59_n N_A_27_398#_c_182_n 0.00669835f $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_73 N_A_c_60_n N_A_27_398#_c_182_n 0.00770329f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_74 N_A_c_62_n N_A_27_398#_c_182_n 0.0263323f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_75 N_A_M1006_g N_A_27_398#_c_187_n 0.0139308f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_A_27_398#_c_188_n 0.0143302f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_77 N_A_c_59_n N_A_27_398#_c_188_n 3.2368e-19 $X=0.51 $Y=1.545 $X2=0 $Y2=0
cc_78 N_A_M1006_g N_A_27_398#_c_189_n 5.73514e-19 $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_A_27_398#_c_192_n 0.00357833f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_80 N_A_M1006_g N_VPWR_c_262_n 0.00454317f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_81 N_A_M1006_g N_VPWR_c_264_n 0.00560776f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_82 N_A_M1006_g N_VPWR_c_261_n 0.00606454f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_83 A A_233_136# 0.00220589f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_84 A N_VGND_c_324_n 0.0186975f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A_c_60_n N_VGND_c_325_n 0.0116176f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_86 N_A_c_62_n N_VGND_c_325_n 0.0795377f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_87 N_A_c_57_n N_VGND_c_328_n 0.0073025f $X=0.53 $Y=0.57 $X2=0 $Y2=0
cc_88 N_A_c_60_n N_VGND_c_328_n 0.00773969f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_89 N_A_c_62_n N_VGND_c_328_n 0.043082f $X=1.085 $Y=0.462 $X2=0 $Y2=0
cc_90 B N_C_M1004_g 0.0068958f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B_c_99_n N_C_M1004_g 6.80675e-19 $X=1.01 $Y=1.595 $X2=0 $Y2=0
cc_92 N_B_c_100_n N_C_M1004_g 0.0325782f $X=1.01 $Y=1.43 $X2=0 $Y2=0
cc_93 B C 0.0268673f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B_c_99_n C 2.72576e-19 $X=1.01 $Y=1.595 $X2=0 $Y2=0
cc_95 N_B_M1003_g N_C_c_145_n 0.0244455f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_96 B N_C_c_145_n 0.00244375f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_99_n N_C_c_145_n 0.0163959f $X=1.01 $Y=1.595 $X2=0 $Y2=0
cc_98 N_B_M1003_g N_A_27_398#_c_182_n 8.41888e-19 $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_99 B N_A_27_398#_c_182_n 0.0261437f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B_c_99_n N_A_27_398#_c_182_n 0.00102333f $X=1.01 $Y=1.595 $X2=0 $Y2=0
cc_101 N_B_c_100_n N_A_27_398#_c_182_n 0.00223336f $X=1.01 $Y=1.43 $X2=0 $Y2=0
cc_102 N_B_M1003_g N_A_27_398#_c_187_n 5.72628e-19 $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_103 N_B_M1003_g N_A_27_398#_c_188_n 0.0134232f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_104 B N_A_27_398#_c_188_n 0.0212186f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_99_n N_A_27_398#_c_188_n 7.9189e-19 $X=1.01 $Y=1.595 $X2=0 $Y2=0
cc_106 N_B_M1003_g N_A_27_398#_c_189_n 0.0120102f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_107 N_B_M1003_g N_A_27_398#_c_193_n 0.00134389f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_108 B N_A_27_398#_c_193_n 0.0182023f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B_c_99_n N_A_27_398#_c_193_n 2.22764e-19 $X=1.01 $Y=1.595 $X2=0 $Y2=0
cc_110 N_B_M1003_g N_VPWR_c_262_n 0.00307419f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_111 N_B_M1003_g N_VPWR_c_263_n 5.45191e-19 $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_VPWR_c_265_n 0.00560776f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_113 N_B_M1003_g N_VPWR_c_261_n 0.00606454f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_114 B A_121_136# 0.00405918f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_115 B A_233_136# 0.00359387f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_116 N_B_c_100_n N_VGND_c_325_n 4.93445e-19 $X=1.01 $Y=1.43 $X2=0 $Y2=0
cc_117 N_C_M1004_g N_A_27_398#_c_181_n 0.0219279f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_118 N_C_M1005_g N_A_27_398#_M1000_g 0.00552396f $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_119 N_C_c_145_n N_A_27_398#_M1000_g 0.0018199f $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_120 N_C_M1005_g N_A_27_398#_c_189_n 8.96491e-19 $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_121 N_C_M1005_g N_A_27_398#_c_190_n 0.0183059f $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_122 C N_A_27_398#_c_190_n 0.0243652f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_123 N_C_c_145_n N_A_27_398#_c_190_n 0.0015396f $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_124 N_C_M1005_g N_A_27_398#_c_191_n 0.0028648f $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_125 N_C_c_145_n N_A_27_398#_c_191_n 8.24616e-19 $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_126 N_C_M1004_g N_A_27_398#_c_183_n 5.59322e-19 $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_127 C N_A_27_398#_c_183_n 0.0180069f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_128 N_C_c_145_n N_A_27_398#_c_183_n 8.98411e-19 $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_129 C N_A_27_398#_c_184_n 8.96262e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_130 N_C_c_145_n N_A_27_398#_c_184_n 0.0113677f $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_131 N_C_M1005_g N_VPWR_c_263_n 0.01176f $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_132 N_C_M1005_g N_VPWR_c_265_n 0.00502805f $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_133 N_C_M1005_g N_VPWR_c_261_n 0.00525594f $X=1.505 $Y=2.41 $X2=0 $Y2=0
cc_134 N_C_M1004_g N_VGND_c_324_n 0.00515513f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_135 C N_VGND_c_324_n 0.00681967f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_C_c_145_n N_VGND_c_324_n 8.79027e-19 $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_137 N_C_M1004_g N_VGND_c_325_n 0.00428744f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_138 N_C_M1004_g N_VGND_c_328_n 0.00476395f $X=1.565 $Y=0.92 $X2=0 $Y2=0
cc_139 N_A_27_398#_c_188_n N_VPWR_M1006_d 0.00279273f $X=1.115 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_140 N_A_27_398#_c_190_n N_VPWR_M1005_d 0.0110593f $X=2.07 $Y=2.035 $X2=0
+ $Y2=0
cc_141 N_A_27_398#_c_191_n N_VPWR_M1005_d 0.00241578f $X=2.155 $Y=1.95 $X2=0
+ $Y2=0
cc_142 N_A_27_398#_c_187_n N_VPWR_c_262_n 0.021803f $X=0.28 $Y=2.135 $X2=0 $Y2=0
cc_143 N_A_27_398#_c_188_n N_VPWR_c_262_n 0.0208278f $X=1.115 $Y=2.035 $X2=0
+ $Y2=0
cc_144 N_A_27_398#_c_189_n N_VPWR_c_262_n 0.0213364f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_145 N_A_27_398#_M1000_g N_VPWR_c_263_n 0.0182374f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_27_398#_c_189_n N_VPWR_c_263_n 0.0242512f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_147 N_A_27_398#_c_190_n N_VPWR_c_263_n 0.049958f $X=2.07 $Y=2.035 $X2=0 $Y2=0
cc_148 N_A_27_398#_c_183_n N_VPWR_c_263_n 0.00123778f $X=2.235 $Y=1.515 $X2=0
+ $Y2=0
cc_149 N_A_27_398#_c_184_n N_VPWR_c_263_n 5.2873e-19 $X=2.375 $Y=1.515 $X2=0
+ $Y2=0
cc_150 N_A_27_398#_c_187_n N_VPWR_c_264_n 0.00949319f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_151 N_A_27_398#_c_189_n N_VPWR_c_265_n 0.00818063f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_152 N_A_27_398#_M1000_g N_VPWR_c_266_n 0.00475445f $X=2.375 $Y=2.4 $X2=0
+ $Y2=0
cc_153 N_A_27_398#_M1000_g N_VPWR_c_261_n 0.00942403f $X=2.375 $Y=2.4 $X2=0
+ $Y2=0
cc_154 N_A_27_398#_c_187_n N_VPWR_c_261_n 0.0110977f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_155 N_A_27_398#_c_189_n N_VPWR_c_261_n 0.00957104f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_156 N_A_27_398#_c_181_n N_X_c_300_n 0.00624223f $X=2.145 $Y=1.35 $X2=0 $Y2=0
cc_157 N_A_27_398#_c_181_n N_X_c_301_n 0.00220367f $X=2.145 $Y=1.35 $X2=0 $Y2=0
cc_158 N_A_27_398#_c_183_n N_X_c_301_n 0.0131627f $X=2.235 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A_27_398#_c_184_n N_X_c_301_n 0.00386616f $X=2.375 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A_27_398#_M1000_g X 8.99587e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_27_398#_c_181_n N_X_c_302_n 0.00426097f $X=2.145 $Y=1.35 $X2=0 $Y2=0
cc_162 N_A_27_398#_c_191_n N_X_c_302_n 0.00735838f $X=2.155 $Y=1.95 $X2=0 $Y2=0
cc_163 N_A_27_398#_c_183_n N_X_c_302_n 0.0223685f $X=2.235 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A_27_398#_c_184_n N_X_c_302_n 0.0118525f $X=2.375 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A_27_398#_c_181_n N_VGND_c_324_n 0.0089425f $X=2.145 $Y=1.35 $X2=0
+ $Y2=0
cc_166 N_A_27_398#_c_181_n N_VGND_c_327_n 0.00467453f $X=2.145 $Y=1.35 $X2=0
+ $Y2=0
cc_167 N_A_27_398#_c_181_n N_VGND_c_328_n 0.00505379f $X=2.145 $Y=1.35 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_263_n X 0.0297014f $X=2.145 $Y=2.375 $X2=0 $Y2=0
cc_169 N_VPWR_c_266_n X 0.0126277f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_170 N_VPWR_c_261_n X 0.0104521f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_171 N_X_c_300_n N_VGND_c_324_n 0.0206774f $X=2.36 $Y=0.645 $X2=0 $Y2=0
cc_172 N_X_c_300_n N_VGND_c_327_n 0.0093375f $X=2.36 $Y=0.645 $X2=0 $Y2=0
cc_173 N_X_c_300_n N_VGND_c_328_n 0.0109911f $X=2.36 $Y=0.645 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o32a_1.spice
* Created: Fri Aug 28 18:03:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o32a_1.pex.spice"
.subckt sky130_fd_sc_ms__o32a_1  VNB VPB A1 A2 A3 B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_83_264#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157545 AS=0.2109 PD=1.24406 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_251_74#_M1010_d N_A1_M1010_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.136255 PD=0.92 PS=1.07594 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.8 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_251_74#_M1010_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.0896 PD=1.06 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1008 N_A_251_74#_M1008_d N_A3_M1008_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1344 PD=0.99 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.8
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_83_264#_M1006_d N_B2_M1006_g N_A_251_74#_M1008_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1424 AS=0.112 PD=1.085 PS=0.99 NRD=14.988 NRS=13.116 M=1 R=4.26667
+ SA=75002.3 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1000 N_A_251_74#_M1000_d N_B1_M1000_g N_A_83_264#_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2144 AS=0.1424 PD=1.95 PS=1.085 NRD=0 NRS=15.936 M=1 R=4.26667
+ SA=75002.9 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_83_264#_M1003_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.274506 AS=0.3136 PD=1.69057 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1005 A_251_368# N_A1_M1005_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.245094 PD=1.24 PS=1.50943 NRD=12.7853 NRS=31.0078 M=1 R=5.55556
+ SA=90000.8 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1009 A_335_368# N_A2_M1009_g A_251_368# VPB PSHORT L=0.18 W=1 AD=0.18 AS=0.12
+ PD=1.36 PS=1.24 NRD=24.6053 NRS=12.7853 M=1 R=5.55556 SA=90001.3 SB=90001.9
+ A=0.18 P=2.36 MULT=1
MM1011 N_A_83_264#_M1011_d N_A3_M1011_g A_335_368# VPB PSHORT L=0.18 W=1 AD=0.18
+ AS=0.18 PD=1.36 PS=1.36 NRD=7.8603 NRS=24.6053 M=1 R=5.55556 SA=90001.8
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1001 A_551_368# N_B2_M1001_g N_A_83_264#_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.2075 AS=0.18 PD=1.415 PS=1.36 NRD=30.0228 NRS=7.8603 M=1 R=5.55556
+ SA=90002.3 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g A_551_368# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.2075 PD=2.56 PS=1.415 NRD=0 NRS=30.0228 M=1 R=5.55556 SA=90002.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o32a_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a22oi_2.pxi.spice
* Created: Fri Aug 28 17:03:26 2020
* 
x_PM_SKY130_FD_SC_MS__A22OI_2%A1 N_A1_M1002_g N_A1_M1000_g N_A1_M1013_g
+ N_A1_M1008_g N_A1_c_85_n N_A1_c_92_n N_A1_c_101_p N_A1_c_125_p N_A1_c_93_n A1
+ A1 N_A1_c_86_n N_A1_c_87_n N_A1_c_88_n PM_SKY130_FD_SC_MS__A22OI_2%A1
x_PM_SKY130_FD_SC_MS__A22OI_2%A2 N_A2_M1001_g N_A2_M1009_g N_A2_M1011_g
+ N_A2_M1004_g A2 N_A2_c_179_n N_A2_c_176_n PM_SKY130_FD_SC_MS__A22OI_2%A2
x_PM_SKY130_FD_SC_MS__A22OI_2%B1 N_B1_M1005_g N_B1_M1003_g N_B1_M1006_g
+ N_B1_M1015_g N_B1_c_229_n N_B1_c_230_n B1 N_B1_c_231_n N_B1_c_232_n
+ N_B1_c_233_n PM_SKY130_FD_SC_MS__A22OI_2%B1
x_PM_SKY130_FD_SC_MS__A22OI_2%B2 N_B2_M1007_g N_B2_M1010_g N_B2_M1014_g
+ N_B2_M1012_g B2 N_B2_c_310_n N_B2_c_307_n PM_SKY130_FD_SC_MS__A22OI_2%B2
x_PM_SKY130_FD_SC_MS__A22OI_2%A_66_368# N_A_66_368#_M1000_d N_A_66_368#_M1009_d
+ N_A_66_368#_M1008_d N_A_66_368#_M1010_d N_A_66_368#_M1015_s
+ N_A_66_368#_c_356_n N_A_66_368#_c_357_n N_A_66_368#_c_369_n
+ N_A_66_368#_c_373_n N_A_66_368#_c_376_n N_A_66_368#_c_358_n
+ N_A_66_368#_c_359_n N_A_66_368#_c_388_n N_A_66_368#_c_360_n
+ N_A_66_368#_c_361_n N_A_66_368#_c_362_n N_A_66_368#_c_363_n
+ N_A_66_368#_c_380_n N_A_66_368#_c_364_n PM_SKY130_FD_SC_MS__A22OI_2%A_66_368#
x_PM_SKY130_FD_SC_MS__A22OI_2%VPWR N_VPWR_M1000_s N_VPWR_M1011_s N_VPWR_c_435_n
+ N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n VPWR N_VPWR_c_439_n
+ N_VPWR_c_440_n N_VPWR_c_434_n N_VPWR_c_442_n PM_SKY130_FD_SC_MS__A22OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A22OI_2%Y N_Y_M1002_d N_Y_M1013_d N_Y_M1006_s N_Y_M1003_d
+ N_Y_M1012_s N_Y_c_488_n N_Y_c_489_n N_Y_c_490_n N_Y_c_491_n N_Y_c_492_n
+ N_Y_c_498_n N_Y_c_517_n N_Y_c_562_n N_Y_c_532_n N_Y_c_565_n N_Y_c_499_n
+ N_Y_c_493_n N_Y_c_494_n N_Y_c_501_n N_Y_c_544_n N_Y_c_495_n Y
+ PM_SKY130_FD_SC_MS__A22OI_2%Y
x_PM_SKY130_FD_SC_MS__A22OI_2%A_148_74# N_A_148_74#_M1002_s N_A_148_74#_M1004_d
+ N_A_148_74#_c_588_n N_A_148_74#_c_586_n N_A_148_74#_c_592_n
+ N_A_148_74#_c_587_n PM_SKY130_FD_SC_MS__A22OI_2%A_148_74#
x_PM_SKY130_FD_SC_MS__A22OI_2%VGND N_VGND_M1001_s N_VGND_M1007_d N_VGND_c_615_n
+ N_VGND_c_616_n VGND N_VGND_c_617_n N_VGND_c_618_n N_VGND_c_619_n
+ N_VGND_c_620_n N_VGND_c_621_n N_VGND_c_622_n PM_SKY130_FD_SC_MS__A22OI_2%VGND
x_PM_SKY130_FD_SC_MS__A22OI_2%A_558_74# N_A_558_74#_M1005_d N_A_558_74#_M1014_s
+ N_A_558_74#_c_681_n N_A_558_74#_c_677_n N_A_558_74#_c_684_n
+ N_A_558_74#_c_685_n N_A_558_74#_c_678_n PM_SKY130_FD_SC_MS__A22OI_2%A_558_74#
cc_1 VNB N_A1_M1002_g 0.0308884f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.74
cc_2 VNB N_A1_M1013_g 0.0260601f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=0.74
cc_3 VNB N_A1_c_85_n 0.00242771f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.78
cc_4 VNB N_A1_c_86_n 0.0300305f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_5 VNB N_A1_c_87_n 0.0365887f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=1.515
cc_6 VNB N_A1_c_88_n 0.0179151f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.605
cc_7 VNB N_A2_M1001_g 0.0231888f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.74
cc_8 VNB N_A2_M1004_g 0.0237266f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.4
cc_9 VNB N_A2_c_176_n 0.0365157f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_B1_M1003_g 0.00629005f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.4
cc_11 VNB N_B1_M1006_g 0.0251344f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=0.74
cc_12 VNB N_B1_M1015_g 0.00180715f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.4
cc_13 VNB N_B1_c_229_n 0.0185467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_230_n 0.0342053f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.95
cc_15 VNB N_B1_c_231_n 0.0305851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_232_n 0.0201156f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_B1_c_233_n 0.00214676f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.515
cc_18 VNB N_B2_M1007_g 0.0221741f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.74
cc_19 VNB N_B2_M1014_g 0.0221293f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=0.74
cc_20 VNB N_B2_c_307_n 0.0342126f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_VPWR_c_434_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_22 VNB N_Y_c_488_n 0.0300805f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.95
cc_23 VNB N_Y_c_489_n 0.0188679f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.035
cc_24 VNB N_Y_c_490_n 0.00962716f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.95
cc_25 VNB N_Y_c_491_n 0.0040003f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.515
cc_26 VNB N_Y_c_492_n 0.00365168f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_Y_c_493_n 0.0306385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_494_n 0.0251863f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.605
cc_29 VNB N_Y_c_495_n 0.0190306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.00397591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_148_74#_c_586_n 0.00214855f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.35
cc_32 VNB N_A_148_74#_c_587_n 0.00237992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_615_n 0.00640788f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.35
cc_34 VNB N_VGND_c_616_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=1.68
cc_35 VNB N_VGND_c_617_n 0.0338243f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.78
cc_36 VNB N_VGND_c_618_n 0.0486589f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.515
cc_37 VNB N_VGND_c_619_n 0.0327812f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_38 VNB N_VGND_c_620_n 0.284644f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.515
cc_39 VNB N_VGND_c_621_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.515
cc_40 VNB N_VGND_c_622_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=1.515
cc_41 VNB N_A_558_74#_c_677_n 0.00344625f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.35
cc_42 VNB N_A_558_74#_c_678_n 0.00214855f $X=-0.19 $Y=-0.245 $X2=2.34 $Y2=2.4
cc_43 VPB N_A1_M1000_g 0.0265123f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=2.4
cc_44 VPB N_A1_M1008_g 0.0232505f $X=-0.19 $Y=1.66 $X2=2.34 $Y2=2.4
cc_45 VPB N_A1_c_85_n 7.32556e-19 $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.78
cc_46 VPB N_A1_c_92_n 5.62538e-19 $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.95
cc_47 VPB N_A1_c_93_n 0.00245065f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.515
cc_48 VPB N_A1_c_86_n 0.00577294f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.515
cc_49 VPB N_A1_c_87_n 0.0124838f $X=-0.19 $Y=1.66 $X2=2.34 $Y2=1.515
cc_50 VPB N_A1_c_88_n 0.0147178f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.605
cc_51 VPB N_A2_M1009_g 0.02138f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=2.4
cc_52 VPB N_A2_M1011_g 0.0243516f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=0.74
cc_53 VPB N_A2_c_179_n 0.00268643f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.515
cc_54 VPB N_A2_c_176_n 0.00522055f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_55 VPB N_B1_M1003_g 0.0211631f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=2.4
cc_56 VPB N_B1_M1015_g 0.0254599f $X=-0.19 $Y=1.66 $X2=2.34 $Y2=2.4
cc_57 VPB N_B2_M1010_g 0.0210178f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=2.4
cc_58 VPB N_B2_M1012_g 0.0203474f $X=-0.19 $Y=1.66 $X2=2.34 $Y2=2.4
cc_59 VPB N_B2_c_310_n 0.0028769f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.515
cc_60 VPB N_B2_c_307_n 0.00471557f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_A_66_368#_c_356_n 0.0130665f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.95
cc_62 VPB N_A_66_368#_c_357_n 0.0218419f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.515
cc_63 VPB N_A_66_368#_c_358_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.35
cc_64 VPB N_A_66_368#_c_359_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.68
cc_65 VPB N_A_66_368#_c_360_n 0.0116218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_66_368#_c_361_n 0.0241251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_66_368#_c_362_n 0.00717518f $X=-0.19 $Y=1.66 $X2=0.672 $Y2=1.605
cc_68 VPB N_A_66_368#_c_363_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_66_368#_c_364_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_435_n 0.00554449f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=1.35
cc_71 VPB N_VPWR_c_436_n 0.0115818f $X=-0.19 $Y=1.66 $X2=2.34 $Y2=1.68
cc_72 VPB N_VPWR_c_437_n 0.0235962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_438_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.78
cc_74 VPB N_VPWR_c_439_n 0.0196495f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=1.515
cc_75 VPB N_VPWR_c_440_n 0.0629081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_434_n 0.0778901f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.515
cc_77 VPB N_VPWR_c_442_n 0.0103572f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.35
cc_78 VPB N_Y_c_492_n 5.58997e-19 $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_79 VPB N_Y_c_498_n 0.00417126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_Y_c_499_n 0.0152154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_Y_c_494_n 0.0147012f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.605
cc_82 VPB N_Y_c_501_n 0.00301358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 N_A1_M1002_g N_A2_M1001_g 0.0206959f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A1_M1000_g N_A2_M1009_g 0.0483699f $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A1_c_85_n N_A2_M1009_g 6.51776e-19 $X=0.795 $Y=1.78 $X2=0 $Y2=0
cc_86 N_A1_c_92_n N_A2_M1009_g 0.00352898f $X=0.795 $Y=1.95 $X2=0 $Y2=0
cc_87 N_A1_c_101_p N_A2_M1009_g 0.0119526f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A1_M1008_g N_A2_M1011_g 0.0223475f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A1_c_101_p N_A2_M1011_g 0.0183029f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A1_c_93_n N_A2_M1011_g 0.0054532f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A1_M1013_g N_A2_M1004_g 0.0335526f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A1_c_85_n N_A2_c_179_n 0.0297103f $X=0.795 $Y=1.78 $X2=0 $Y2=0
cc_93 N_A1_c_101_p N_A2_c_179_n 0.0257705f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A1_c_93_n N_A2_c_179_n 0.0126308f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_95 N_A1_c_86_n N_A2_c_179_n 3.48721e-19 $X=0.605 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A1_c_87_n N_A2_c_179_n 6.56057e-19 $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A1_c_85_n N_A2_c_176_n 0.00192936f $X=0.795 $Y=1.78 $X2=0 $Y2=0
cc_98 N_A1_c_101_p N_A2_c_176_n 4.89879e-19 $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A1_c_93_n N_A2_c_176_n 0.00114719f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A1_c_86_n N_A2_c_176_n 0.0184134f $X=0.605 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A1_c_87_n N_A2_c_176_n 0.0239289f $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A1_c_87_n N_B1_M1003_g 0.0244645f $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A1_c_87_n N_B1_c_231_n 0.0124139f $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A1_M1013_g N_B1_c_232_n 0.0168061f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A1_c_101_p N_A_66_368#_M1009_d 0.00352567f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A1_c_86_n N_A_66_368#_c_356_n 5.95205e-19 $X=0.605 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A1_c_88_n N_A_66_368#_c_356_n 0.0213917f $X=0.71 $Y=1.605 $X2=0 $Y2=0
cc_108 N_A1_M1000_g N_A_66_368#_c_357_n 4.69176e-19 $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A1_M1000_g N_A_66_368#_c_369_n 0.0153283f $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A1_c_101_p N_A_66_368#_c_369_n 0.0175781f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A1_c_125_p N_A_66_368#_c_369_n 0.00884832f $X=0.88 $Y=2.035 $X2=0 $Y2=0
cc_112 N_A1_c_88_n N_A_66_368#_c_369_n 0.00446394f $X=0.71 $Y=1.605 $X2=0 $Y2=0
cc_113 N_A1_M1008_g N_A_66_368#_c_373_n 0.0186353f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A1_c_101_p N_A_66_368#_c_373_n 0.0466604f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A1_c_87_n N_A_66_368#_c_373_n 9.24518e-19 $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A1_M1008_g N_A_66_368#_c_376_n 0.0106757f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A1_M1008_g N_A_66_368#_c_359_n 0.00345561f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A1_M1000_g N_A_66_368#_c_363_n 5.87944e-19 $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A1_c_101_p N_A_66_368#_c_363_n 0.0171986f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A1_M1008_g N_A_66_368#_c_380_n 0.00966041f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A1_c_92_n N_VPWR_M1000_s 0.00125604f $X=0.795 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A1_c_101_p N_VPWR_M1000_s 0.00497879f $X=1.88 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A1_c_125_p N_VPWR_M1000_s 5.77118e-19 $X=0.88 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A1_c_101_p N_VPWR_M1011_s 0.0140357f $X=1.88 $Y=2.035 $X2=0 $Y2=0
cc_125 N_A1_c_93_n N_VPWR_M1011_s 0.00294627f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A1_M1000_g N_VPWR_c_435_n 0.0111267f $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A1_M1008_g N_VPWR_c_436_n 0.00475889f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A1_M1000_g N_VPWR_c_437_n 0.00460063f $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A1_M1008_g N_VPWR_c_440_n 0.00517089f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A1_M1000_g N_VPWR_c_434_n 0.00912769f $X=0.68 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A1_M1008_g N_VPWR_c_434_n 0.00979287f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A1_M1002_g N_Y_c_488_n 0.00159319f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A1_M1002_g N_Y_c_489_n 0.0151989f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A1_M1013_g N_Y_c_489_n 0.00858988f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A1_c_85_n N_Y_c_489_n 0.01399f $X=0.795 $Y=1.78 $X2=0 $Y2=0
cc_136 N_A1_c_93_n N_Y_c_489_n 0.0123843f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A1_c_86_n N_Y_c_489_n 0.00222096f $X=0.605 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A1_c_87_n N_Y_c_489_n 0.00174068f $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_c_88_n N_Y_c_489_n 0.0126866f $X=0.71 $Y=1.605 $X2=0 $Y2=0
cc_140 N_A1_c_86_n N_Y_c_490_n 0.00243921f $X=0.605 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A1_c_88_n N_Y_c_490_n 0.0218126f $X=0.71 $Y=1.605 $X2=0 $Y2=0
cc_142 N_A1_M1013_g N_Y_c_491_n 0.00348259f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1013_g N_Y_c_492_n 0.00179761f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_M1008_g N_Y_c_492_n 7.45474e-19 $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A1_c_93_n N_Y_c_492_n 0.0208052f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A1_c_87_n N_Y_c_492_n 0.0113174f $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A1_M1008_g N_Y_c_517_n 0.00500553f $X=2.34 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A1_c_93_n N_Y_c_517_n 0.011908f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A1_M1013_g Y 0.0166605f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A1_c_93_n Y 0.0144482f $X=2.045 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A1_c_87_n Y 0.01163f $X=2.34 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A1_M1002_g N_A_148_74#_c_588_n 0.00219352f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1002_g N_A_148_74#_c_586_n 0.00576372f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_M1013_g N_A_148_74#_c_587_n 0.00605667f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_M1002_g N_VGND_c_615_n 5.4581e-19 $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A1_M1002_g N_VGND_c_617_n 0.00433834f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_M1013_g N_VGND_c_618_n 0.00433139f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A1_M1002_g N_VGND_c_620_n 0.00825175f $X=0.665 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A1_M1013_g N_VGND_c_620_n 0.00641761f $X=2.025 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1009_g N_A_66_368#_c_369_n 0.0126573f $X=1.13 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A2_M1011_g N_A_66_368#_c_373_n 0.0139537f $X=1.58 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A2_M1009_g N_A_66_368#_c_363_n 0.00955292f $X=1.13 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A2_M1011_g N_A_66_368#_c_363_n 0.0135294f $X=1.58 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A2_M1009_g N_VPWR_c_435_n 0.002979f $X=1.13 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A2_M1011_g N_VPWR_c_436_n 0.00692139f $X=1.58 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A2_M1009_g N_VPWR_c_439_n 0.005209f $X=1.13 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A2_M1011_g N_VPWR_c_439_n 0.005209f $X=1.58 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A2_M1009_g N_VPWR_c_434_n 0.00982376f $X=1.13 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A2_M1011_g N_VPWR_c_434_n 0.00983964f $X=1.58 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A2_M1001_g N_Y_c_489_n 0.0117193f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1004_g N_Y_c_489_n 0.0154194f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_c_179_n N_Y_c_489_n 0.027474f $X=1.215 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A2_c_176_n N_Y_c_489_n 0.00471133f $X=1.595 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A2_M1004_g Y 0.00106882f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A2_M1001_g N_A_148_74#_c_586_n 2.93125e-19 $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A2_M1001_g N_A_148_74#_c_592_n 0.0101634f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A2_M1004_g N_A_148_74#_c_592_n 0.00916065f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_M1001_g N_A_148_74#_c_587_n 6.14282e-19 $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A2_M1004_g N_A_148_74#_c_587_n 0.00813518f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_VGND_c_615_n 0.00662966f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A2_M1004_g N_VGND_c_615_n 0.00435463f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A2_M1001_g N_VGND_c_617_n 0.00281141f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A2_M1004_g N_VGND_c_618_n 0.00330305f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A2_M1001_g N_VGND_c_620_n 0.00365164f $X=1.095 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A2_M1004_g N_VGND_c_620_n 0.00427788f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B1_c_229_n N_B2_M1007_g 0.00681238f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_187 N_B1_c_231_n N_B2_M1007_g 0.0213999f $X=2.805 $Y=1.385 $X2=0 $Y2=0
cc_188 N_B1_c_232_n N_B2_M1007_g 0.0174342f $X=2.805 $Y=1.22 $X2=0 $Y2=0
cc_189 N_B1_c_233_n N_B2_M1007_g 0.00668713f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_190 N_B1_M1006_g N_B2_M1014_g 0.0197692f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B1_c_229_n N_B2_M1014_g 0.0123163f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_192 N_B1_c_233_n N_B2_M1014_g 2.93543e-19 $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_193 N_B1_M1003_g N_B2_c_310_n 5.35648e-19 $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_194 N_B1_M1015_g N_B2_c_310_n 8.18683e-19 $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_195 N_B1_c_229_n N_B2_c_310_n 0.0407683f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_196 N_B1_c_233_n N_B2_c_310_n 0.00929155f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_197 N_B1_M1003_g N_B2_c_307_n 0.0314466f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_198 N_B1_M1015_g N_B2_c_307_n 0.0311655f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_199 N_B1_c_229_n N_B2_c_307_n 0.00758898f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_200 N_B1_c_230_n N_B2_c_307_n 0.0161738f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_201 N_B1_c_233_n N_B2_c_307_n 0.00793465f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_202 N_B1_M1003_g N_A_66_368#_c_376_n 0.00661328f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_203 N_B1_M1003_g N_A_66_368#_c_358_n 0.0117719f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_204 N_B1_M1003_g N_A_66_368#_c_359_n 0.001916f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_205 N_B1_M1003_g N_A_66_368#_c_388_n 5.71427e-19 $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_206 N_B1_M1015_g N_A_66_368#_c_388_n 5.73047e-19 $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_207 N_B1_M1015_g N_A_66_368#_c_360_n 0.0145133f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_208 N_B1_M1015_g N_A_66_368#_c_361_n 0.0097355f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_209 N_B1_M1003_g N_A_66_368#_c_380_n 0.00517963f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_210 N_B1_M1003_g N_VPWR_c_440_n 0.00333896f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B1_M1015_g N_VPWR_c_440_n 0.00333896f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_212 N_B1_M1003_g N_VPWR_c_434_n 0.00423185f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_213 N_B1_M1015_g N_VPWR_c_434_n 0.004269f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B1_c_232_n N_Y_c_491_n 0.008029f $X=2.805 $Y=1.22 $X2=0 $Y2=0
cc_215 N_B1_M1003_g N_Y_c_492_n 0.0035869f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_216 N_B1_M1003_g N_Y_c_498_n 0.0154467f $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_217 N_B1_c_231_n N_Y_c_498_n 0.0036114f $X=2.805 $Y=1.385 $X2=0 $Y2=0
cc_218 N_B1_c_233_n N_Y_c_498_n 0.0155945f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_219 N_B1_c_233_n N_Y_c_532_n 0.00322024f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_220 N_B1_M1015_g N_Y_c_499_n 0.017015f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B1_c_229_n N_Y_c_499_n 0.0127181f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_222 N_B1_c_230_n N_Y_c_499_n 5.11344e-19 $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_223 N_B1_M1006_g N_Y_c_493_n 0.00205177f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_224 N_B1_M1006_g N_Y_c_494_n 0.00300603f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B1_M1015_g N_Y_c_494_n 0.00991194f $X=4.17 $Y=2.4 $X2=0 $Y2=0
cc_226 N_B1_c_229_n N_Y_c_494_n 0.0317617f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_227 N_B1_c_230_n N_Y_c_494_n 0.00232633f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_228 N_B1_M1003_g N_Y_c_501_n 2.61968e-19 $X=2.79 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B1_c_231_n N_Y_c_501_n 9.08531e-19 $X=2.805 $Y=1.385 $X2=0 $Y2=0
cc_230 N_B1_c_233_n N_Y_c_501_n 0.0177732f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_231 N_B1_c_229_n N_Y_c_544_n 0.00696332f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_232 N_B1_c_229_n N_Y_c_495_n 0.0130294f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_233 N_B1_c_230_n N_Y_c_495_n 9.80105e-19 $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_234 N_B1_c_231_n Y 0.008029f $X=2.805 $Y=1.385 $X2=0 $Y2=0
cc_235 N_B1_c_233_n Y 0.0371385f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_236 N_B1_c_229_n N_VGND_M1007_d 0.00176891f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_237 N_B1_M1006_g N_VGND_c_616_n 5.4581e-19 $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_c_232_n N_VGND_c_616_n 4.80547e-19 $X=2.805 $Y=1.22 $X2=0 $Y2=0
cc_239 N_B1_c_232_n N_VGND_c_618_n 0.00461464f $X=2.805 $Y=1.22 $X2=0 $Y2=0
cc_240 N_B1_M1006_g N_VGND_c_619_n 0.00433834f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B1_M1006_g N_VGND_c_620_n 0.00825215f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B1_c_232_n N_VGND_c_620_n 0.0091238f $X=2.805 $Y=1.22 $X2=0 $Y2=0
cc_243 N_B1_c_233_n N_A_558_74#_M1005_d 0.0030251f $X=3.235 $Y=1.32 $X2=-0.19
+ $Y2=-0.245
cc_244 N_B1_c_229_n N_A_558_74#_M1014_s 0.00180465f $X=3.905 $Y=1.175 $X2=0
+ $Y2=0
cc_245 N_B1_c_231_n N_A_558_74#_c_681_n 7.34751e-19 $X=2.805 $Y=1.385 $X2=0
+ $Y2=0
cc_246 N_B1_c_233_n N_A_558_74#_c_681_n 0.0238114f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_247 N_B1_c_232_n N_A_558_74#_c_677_n 0.00294932f $X=2.805 $Y=1.22 $X2=0 $Y2=0
cc_248 N_B1_c_233_n N_A_558_74#_c_684_n 0.0329906f $X=3.235 $Y=1.32 $X2=0 $Y2=0
cc_249 N_B1_M1006_g N_A_558_74#_c_685_n 0.00219251f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B1_c_229_n N_A_558_74#_c_685_n 0.0163105f $X=3.905 $Y=1.175 $X2=0 $Y2=0
cc_251 N_B1_M1006_g N_A_558_74#_c_678_n 0.00576372f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B2_M1010_g N_A_66_368#_c_358_n 0.0117719f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_253 N_B2_M1010_g N_A_66_368#_c_388_n 0.0095266f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_254 N_B2_M1012_g N_A_66_368#_c_388_n 0.00939395f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_255 N_B2_M1012_g N_A_66_368#_c_360_n 0.0115958f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B2_M1012_g N_A_66_368#_c_361_n 5.73047e-19 $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B2_M1010_g N_A_66_368#_c_380_n 6.21136e-19 $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B2_M1010_g N_A_66_368#_c_364_n 0.00194226f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_259 N_B2_M1012_g N_A_66_368#_c_364_n 0.00194226f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B2_M1010_g N_VPWR_c_440_n 0.00333896f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B2_M1012_g N_VPWR_c_440_n 0.00333896f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B2_M1010_g N_VPWR_c_434_n 0.00423074f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_263 N_B2_M1012_g N_VPWR_c_434_n 0.00422796f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_264 N_B2_M1010_g N_Y_c_532_n 0.0185166f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_265 N_B2_M1012_g N_Y_c_532_n 0.0164173f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_266 N_B2_c_310_n N_Y_c_532_n 0.0226485f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_267 N_B2_c_307_n N_Y_c_532_n 4.88468e-19 $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_268 N_B2_M1010_g N_Y_c_501_n 0.00204508f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_269 N_B2_c_310_n N_Y_c_501_n 0.00343856f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_270 N_B2_M1007_g N_VGND_c_616_n 0.0067459f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_271 N_B2_M1014_g N_VGND_c_616_n 0.00662193f $X=3.685 $Y=0.74 $X2=0 $Y2=0
cc_272 N_B2_M1007_g N_VGND_c_618_n 0.00281141f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_273 N_B2_M1014_g N_VGND_c_619_n 0.00281141f $X=3.685 $Y=0.74 $X2=0 $Y2=0
cc_274 N_B2_M1007_g N_VGND_c_620_n 0.00366095f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_275 N_B2_M1014_g N_VGND_c_620_n 0.00365164f $X=3.685 $Y=0.74 $X2=0 $Y2=0
cc_276 N_B2_M1007_g N_A_558_74#_c_677_n 3.54606e-19 $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_277 N_B2_M1007_g N_A_558_74#_c_684_n 0.00983086f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_278 N_B2_M1014_g N_A_558_74#_c_684_n 0.00983086f $X=3.685 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B2_M1014_g N_A_558_74#_c_678_n 2.93125e-19 $X=3.685 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_66_368#_c_369_n N_VPWR_M1000_s 0.00330866f $X=1.19 $Y=2.375 $X2=-0.19
+ $Y2=1.66
cc_281 N_A_66_368#_c_373_n N_VPWR_M1011_s 0.0116704f $X=2.4 $Y=2.375 $X2=0 $Y2=0
cc_282 N_A_66_368#_c_357_n N_VPWR_c_435_n 0.0117266f $X=0.455 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_66_368#_c_369_n N_VPWR_c_435_n 0.0148589f $X=1.19 $Y=2.375 $X2=0
+ $Y2=0
cc_284 N_A_66_368#_c_363_n N_VPWR_c_435_n 0.0122069f $X=1.355 $Y=2.375 $X2=0
+ $Y2=0
cc_285 N_A_66_368#_c_373_n N_VPWR_c_436_n 0.0379131f $X=2.4 $Y=2.375 $X2=0 $Y2=0
cc_286 N_A_66_368#_c_359_n N_VPWR_c_436_n 0.0122917f $X=2.73 $Y=2.99 $X2=0 $Y2=0
cc_287 N_A_66_368#_c_363_n N_VPWR_c_436_n 0.0139844f $X=1.355 $Y=2.375 $X2=0
+ $Y2=0
cc_288 N_A_66_368#_c_357_n N_VPWR_c_437_n 0.011066f $X=0.455 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_66_368#_c_363_n N_VPWR_c_439_n 0.0144776f $X=1.355 $Y=2.375 $X2=0
+ $Y2=0
cc_290 N_A_66_368#_c_358_n N_VPWR_c_440_n 0.0377252f $X=3.33 $Y=2.99 $X2=0 $Y2=0
cc_291 N_A_66_368#_c_359_n N_VPWR_c_440_n 0.0234458f $X=2.73 $Y=2.99 $X2=0 $Y2=0
cc_292 N_A_66_368#_c_360_n N_VPWR_c_440_n 0.0593439f $X=4.23 $Y=2.99 $X2=0 $Y2=0
cc_293 N_A_66_368#_c_364_n N_VPWR_c_440_n 0.0234458f $X=3.495 $Y=2.99 $X2=0
+ $Y2=0
cc_294 N_A_66_368#_c_357_n N_VPWR_c_434_n 0.00915947f $X=0.455 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_66_368#_c_358_n N_VPWR_c_434_n 0.0211866f $X=3.33 $Y=2.99 $X2=0 $Y2=0
cc_296 N_A_66_368#_c_359_n N_VPWR_c_434_n 0.0125551f $X=2.73 $Y=2.99 $X2=0 $Y2=0
cc_297 N_A_66_368#_c_360_n N_VPWR_c_434_n 0.032751f $X=4.23 $Y=2.99 $X2=0 $Y2=0
cc_298 N_A_66_368#_c_363_n N_VPWR_c_434_n 0.0118404f $X=1.355 $Y=2.375 $X2=0
+ $Y2=0
cc_299 N_A_66_368#_c_364_n N_VPWR_c_434_n 0.0125551f $X=3.495 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_66_368#_c_358_n N_Y_M1003_d 0.00197722f $X=3.33 $Y=2.99 $X2=0 $Y2=0
cc_301 N_A_66_368#_c_360_n N_Y_M1012_s 0.00165831f $X=4.23 $Y=2.99 $X2=0 $Y2=0
cc_302 N_A_66_368#_M1008_d N_Y_c_498_n 9.77978e-19 $X=2.43 $Y=1.84 $X2=0 $Y2=0
cc_303 N_A_66_368#_c_380_n N_Y_c_498_n 0.00969683f $X=2.565 $Y=2.15 $X2=0 $Y2=0
cc_304 N_A_66_368#_M1008_d N_Y_c_517_n 6.97173e-19 $X=2.43 $Y=1.84 $X2=0 $Y2=0
cc_305 N_A_66_368#_c_373_n N_Y_c_517_n 7.41494e-19 $X=2.4 $Y=2.375 $X2=0 $Y2=0
cc_306 N_A_66_368#_c_380_n N_Y_c_517_n 0.00809274f $X=2.565 $Y=2.15 $X2=0 $Y2=0
cc_307 N_A_66_368#_c_358_n N_Y_c_562_n 0.014157f $X=3.33 $Y=2.99 $X2=0 $Y2=0
cc_308 N_A_66_368#_M1010_d N_Y_c_532_n 0.00314031f $X=3.36 $Y=1.84 $X2=0 $Y2=0
cc_309 N_A_66_368#_c_388_n N_Y_c_532_n 0.0170259f $X=3.495 $Y=2.385 $X2=0 $Y2=0
cc_310 N_A_66_368#_c_360_n N_Y_c_565_n 0.0118736f $X=4.23 $Y=2.99 $X2=0 $Y2=0
cc_311 N_A_66_368#_M1015_s N_Y_c_499_n 0.00923595f $X=4.26 $Y=1.84 $X2=0 $Y2=0
cc_312 N_A_66_368#_c_361_n N_Y_c_499_n 0.0220676f $X=4.395 $Y=2.385 $X2=0 $Y2=0
cc_313 N_Y_c_489_n N_A_148_74#_M1002_s 0.00176461f $X=2.04 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_314 N_Y_c_489_n N_A_148_74#_M1004_d 0.00226577f $X=2.04 $Y=1.175 $X2=0 $Y2=0
cc_315 N_Y_c_489_n N_A_148_74#_c_588_n 0.0151918f $X=2.04 $Y=1.175 $X2=0 $Y2=0
cc_316 N_Y_c_488_n N_A_148_74#_c_586_n 0.014433f $X=0.45 $Y=0.515 $X2=0 $Y2=0
cc_317 N_Y_c_489_n N_A_148_74#_c_592_n 0.0357133f $X=2.04 $Y=1.175 $X2=0 $Y2=0
cc_318 N_Y_c_489_n N_A_148_74#_c_587_n 0.0126057f $X=2.04 $Y=1.175 $X2=0 $Y2=0
cc_319 N_Y_c_491_n N_A_148_74#_c_587_n 0.011762f $X=2.345 $Y=0.515 $X2=0 $Y2=0
cc_320 Y N_A_148_74#_c_587_n 0.00754706f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_321 N_Y_c_489_n N_VGND_M1001_s 0.00251484f $X=2.04 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_322 N_Y_c_488_n N_VGND_c_617_n 0.011066f $X=0.45 $Y=0.515 $X2=0 $Y2=0
cc_323 N_Y_c_491_n N_VGND_c_618_n 0.0179822f $X=2.345 $Y=0.515 $X2=0 $Y2=0
cc_324 N_Y_c_493_n N_VGND_c_619_n 0.0206595f $X=4.33 $Y=0.515 $X2=0 $Y2=0
cc_325 N_Y_c_488_n N_VGND_c_620_n 0.00915947f $X=0.45 $Y=0.515 $X2=0 $Y2=0
cc_326 N_Y_c_491_n N_VGND_c_620_n 0.0148841f $X=2.345 $Y=0.515 $X2=0 $Y2=0
cc_327 N_Y_c_493_n N_VGND_c_620_n 0.0171001f $X=4.33 $Y=0.515 $X2=0 $Y2=0
cc_328 Y N_VGND_c_620_n 0.00357548f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_329 N_Y_c_491_n N_A_558_74#_c_677_n 0.0118811f $X=2.345 $Y=0.515 $X2=0 $Y2=0
cc_330 N_Y_c_493_n N_A_558_74#_c_678_n 0.0145046f $X=4.33 $Y=0.515 $X2=0 $Y2=0
cc_331 N_A_148_74#_c_592_n N_VGND_M1001_s 0.00472947f $X=1.645 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_332 N_A_148_74#_c_586_n N_VGND_c_615_n 0.0104546f $X=0.88 $Y=0.495 $X2=0
+ $Y2=0
cc_333 N_A_148_74#_c_592_n N_VGND_c_615_n 0.0203034f $X=1.645 $Y=0.835 $X2=0
+ $Y2=0
cc_334 N_A_148_74#_c_587_n N_VGND_c_615_n 0.00947296f $X=1.81 $Y=0.535 $X2=0
+ $Y2=0
cc_335 N_A_148_74#_c_586_n N_VGND_c_617_n 0.0118323f $X=0.88 $Y=0.495 $X2=0
+ $Y2=0
cc_336 N_A_148_74#_c_592_n N_VGND_c_617_n 0.00197156f $X=1.645 $Y=0.835 $X2=0
+ $Y2=0
cc_337 N_A_148_74#_c_592_n N_VGND_c_618_n 0.00189877f $X=1.645 $Y=0.835 $X2=0
+ $Y2=0
cc_338 N_A_148_74#_c_587_n N_VGND_c_618_n 0.0140714f $X=1.81 $Y=0.535 $X2=0
+ $Y2=0
cc_339 N_A_148_74#_c_586_n N_VGND_c_620_n 0.00911095f $X=0.88 $Y=0.495 $X2=0
+ $Y2=0
cc_340 N_A_148_74#_c_592_n N_VGND_c_620_n 0.00914714f $X=1.645 $Y=0.835 $X2=0
+ $Y2=0
cc_341 N_A_148_74#_c_587_n N_VGND_c_620_n 0.0117516f $X=1.81 $Y=0.535 $X2=0
+ $Y2=0
cc_342 N_VGND_c_616_n N_A_558_74#_c_677_n 0.01098f $X=3.47 $Y=0.495 $X2=0 $Y2=0
cc_343 N_VGND_c_618_n N_A_558_74#_c_677_n 0.0143052f $X=3.305 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_620_n N_A_558_74#_c_677_n 0.0110855f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_M1007_d N_A_558_74#_c_684_n 0.0033542f $X=3.33 $Y=0.37 $X2=0 $Y2=0
cc_346 N_VGND_c_616_n N_A_558_74#_c_684_n 0.0165203f $X=3.47 $Y=0.495 $X2=0
+ $Y2=0
cc_347 N_VGND_c_618_n N_A_558_74#_c_684_n 0.00189877f $X=3.305 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_619_n N_A_558_74#_c_684_n 0.00197156f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_620_n N_A_558_74#_c_684_n 0.00912085f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_616_n N_A_558_74#_c_678_n 0.0104546f $X=3.47 $Y=0.495 $X2=0
+ $Y2=0
cc_351 N_VGND_c_619_n N_A_558_74#_c_678_n 0.0118323f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_620_n N_A_558_74#_c_678_n 0.00911095f $X=4.56 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__nor3b_4.pex.spice
* Created: Fri Aug 28 17:48:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR3B_4%B 3 7 11 15 19 23 27 31 33 34 35 36 55
c83 15 0 9.05221e-20 $X=0.995 $Y=0.74
r84 54 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.98 $Y=1.515
+ $X2=1.995 $Y2=1.515
r85 52 54 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.65 $Y=1.515
+ $X2=1.98 $Y2=1.515
r86 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r87 50 52 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.565 $Y=1.515
+ $X2=1.65 $Y2=1.515
r88 49 50 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.455 $Y=1.515
+ $X2=1.565 $Y2=1.515
r89 48 49 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=1.005 $Y=1.515
+ $X2=1.455 $Y2=1.515
r90 47 48 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.515
+ $X2=1.005 $Y2=1.515
r91 45 47 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=0.63 $Y=1.515
+ $X2=0.995 $Y2=1.515
r92 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.515 $X2=0.63 $Y2=1.515
r93 43 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.555 $Y=1.515
+ $X2=0.63 $Y2=1.515
r94 41 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.54 $Y=1.515
+ $X2=0.555 $Y2=1.515
r95 36 53 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.65
+ $Y2=1.565
r96 35 53 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.65 $Y2=1.565
r97 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r98 34 46 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.63
+ $Y2=1.565
r99 33 46 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.63 $Y2=1.565
r100 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=1.515
r101 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.995 $Y=1.35
+ $X2=1.995 $Y2=0.74
r102 25 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.68
+ $X2=1.98 $Y2=1.515
r103 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.98 $Y=1.68
+ $X2=1.98 $Y2=2.4
r104 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=1.35
+ $X2=1.565 $Y2=1.515
r105 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.565 $Y=1.35
+ $X2=1.565 $Y2=0.74
r106 17 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.515
r107 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r108 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r109 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r110 9 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=1.515
r111 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=2.4
r112 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.68
+ $X2=0.555 $Y2=1.515
r113 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.555 $Y=1.68
+ $X2=0.555 $Y2=2.4
r114 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.35
+ $X2=0.54 $Y2=1.515
r115 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.54 $Y=1.35 $X2=0.54
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%A_468_264# 1 2 9 13 17 21 25 29 33 37 39 47
+ 53 55 57 58 63 65 76
c151 76 0 2.5976e-19 $X=3.855 $Y=1.485
c152 65 0 1.69815e-19 $X=7.4 $Y=0.5
c153 9 0 7.99092e-20 $X=2.43 $Y=2.4
r154 75 76 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.78 $Y=1.485
+ $X2=3.855 $Y2=1.485
r155 72 73 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.33 $Y=1.485
+ $X2=3.425 $Y2=1.485
r156 71 72 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=2.925 $Y=1.485
+ $X2=3.33 $Y2=1.485
r157 70 71 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.88 $Y=1.485
+ $X2=2.925 $Y2=1.485
r158 66 68 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.43 $Y=1.485
+ $X2=2.495 $Y2=1.485
r159 57 65 8.35471 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=7.48 $Y=1.01
+ $X2=7.48 $Y2=0.68
r160 57 58 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.48 $Y=1.01
+ $X2=7.48 $Y2=1.72
r161 56 63 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.055 $Y=1.805
+ $X2=6.92 $Y2=1.805
r162 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.395 $Y=1.805
+ $X2=7.48 $Y2=1.72
r163 55 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.395 $Y=1.805
+ $X2=7.055 $Y2=1.805
r164 51 63 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=1.89
+ $X2=6.92 $Y2=1.805
r165 51 53 4.05489 $w=2.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.92 $Y=1.89
+ $X2=6.92 $Y2=1.985
r166 48 61 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.195 $Y=1.805
+ $X2=4.042 $Y2=1.805
r167 47 63 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.785 $Y=1.805
+ $X2=6.92 $Y2=1.805
r168 47 48 168.973 $w=1.68e-07 $l=2.59e-06 $layer=LI1_cond $X=6.785 $Y=1.805
+ $X2=4.195 $Y2=1.805
r169 46 75 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.765 $Y=1.485
+ $X2=3.78 $Y2=1.485
r170 46 73 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.765 $Y=1.485
+ $X2=3.425 $Y2=1.485
r171 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.765
+ $Y=1.485 $X2=3.765 $Y2=1.485
r172 42 70 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.745 $Y=1.485
+ $X2=2.88 $Y2=1.485
r173 42 68 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.745 $Y=1.485
+ $X2=2.495 $Y2=1.485
r174 41 45 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=2.745 $Y=1.485
+ $X2=3.765 $Y2=1.485
r175 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.745
+ $Y=1.485 $X2=2.745 $Y2=1.485
r176 39 61 12.0912 $w=3.03e-07 $l=3.2e-07 $layer=LI1_cond $X=4.042 $Y=1.485
+ $X2=4.042 $Y2=1.805
r177 39 45 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.89 $Y=1.485
+ $X2=3.765 $Y2=1.485
r178 35 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.32
+ $X2=3.855 $Y2=1.485
r179 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.855 $Y=1.32
+ $X2=3.855 $Y2=0.74
r180 31 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.65
+ $X2=3.78 $Y2=1.485
r181 31 33 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.78 $Y=1.65
+ $X2=3.78 $Y2=2.4
r182 27 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.32
+ $X2=3.425 $Y2=1.485
r183 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.425 $Y=1.32
+ $X2=3.425 $Y2=0.74
r184 23 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.65
+ $X2=3.33 $Y2=1.485
r185 23 25 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.33 $Y=1.65
+ $X2=3.33 $Y2=2.4
r186 19 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.32
+ $X2=2.925 $Y2=1.485
r187 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.925 $Y=1.32
+ $X2=2.925 $Y2=0.74
r188 15 70 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.65
+ $X2=2.88 $Y2=1.485
r189 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.88 $Y=1.65
+ $X2=2.88 $Y2=2.4
r190 11 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.32
+ $X2=2.495 $Y2=1.485
r191 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.495 $Y=1.32
+ $X2=2.495 $Y2=0.74
r192 7 66 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.65
+ $X2=2.43 $Y2=1.485
r193 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.43 $Y=1.65 $X2=2.43
+ $Y2=2.4
r194 2 53 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.815
+ $Y=1.84 $X2=6.95 $Y2=1.985
r195 1 65 45.5 $w=1.7e-07 $l=8.32466e-07 $layer=licon1_NDIFF $count=4 $X=6.63
+ $Y=0.37 $X2=7.4 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%A 1 3 6 8 10 13 15 17 20 22 24 27 37 47 50
c92 50 0 1.78853e-19 $X=6.365 $Y=1.365
c93 47 0 1.83401e-19 $X=6.055 $Y=1.385
c94 22 0 1.69815e-19 $X=6.055 $Y=1.22
r95 44 45 20.3344 $w=3.2e-07 $l=1.35e-07 $layer=POLY_cond $X=5.555 $Y=1.385
+ $X2=5.69 $Y2=1.385
r96 43 44 47.4469 $w=3.2e-07 $l=3.15e-07 $layer=POLY_cond $X=5.24 $Y=1.385
+ $X2=5.555 $Y2=1.385
r97 42 43 57.9906 $w=3.2e-07 $l=3.85e-07 $layer=POLY_cond $X=4.855 $Y=1.385
+ $X2=5.24 $Y2=1.385
r98 41 42 9.79062 $w=3.2e-07 $l=6.5e-08 $layer=POLY_cond $X=4.79 $Y=1.385
+ $X2=4.855 $Y2=1.385
r99 37 50 3.7435 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.48 $Y=1.365
+ $X2=6.365 $Y2=1.365
r100 36 47 13.5562 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=5.965 $Y=1.385
+ $X2=6.055 $Y2=1.385
r101 36 45 41.4219 $w=3.2e-07 $l=2.75e-07 $layer=POLY_cond $X=5.965 $Y=1.385
+ $X2=5.69 $Y2=1.385
r102 35 50 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.965 $Y=1.385
+ $X2=6.365 $Y2=1.385
r103 35 36 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.965
+ $Y=1.385 $X2=5.965 $Y2=1.385
r104 32 41 27.8656 $w=3.2e-07 $l=1.85e-07 $layer=POLY_cond $X=4.605 $Y=1.385
+ $X2=4.79 $Y2=1.385
r105 32 39 27.1125 $w=3.2e-07 $l=1.8e-07 $layer=POLY_cond $X=4.605 $Y=1.385
+ $X2=4.425 $Y2=1.385
r106 31 35 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=4.605 $Y=1.385
+ $X2=5.965 $Y2=1.385
r107 31 32 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.385 $X2=4.605 $Y2=1.385
r108 25 47 12.8031 $w=3.2e-07 $l=2.03101e-07 $layer=POLY_cond $X=6.14 $Y=1.55
+ $X2=6.055 $Y2=1.385
r109 25 27 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.14 $Y=1.55
+ $X2=6.14 $Y2=2.4
r110 22 47 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.055 $Y=1.22
+ $X2=6.055 $Y2=1.385
r111 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.055 $Y=1.22
+ $X2=6.055 $Y2=0.74
r112 18 45 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.69 $Y=1.55
+ $X2=5.69 $Y2=1.385
r113 18 20 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.69 $Y=1.55
+ $X2=5.69 $Y2=2.4
r114 15 44 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.555 $Y=1.22
+ $X2=5.555 $Y2=1.385
r115 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.555 $Y=1.22
+ $X2=5.555 $Y2=0.74
r116 11 43 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.55
+ $X2=5.24 $Y2=1.385
r117 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.24 $Y=1.55
+ $X2=5.24 $Y2=2.4
r118 8 42 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=1.385
r119 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=0.74
r120 4 41 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.55
+ $X2=4.79 $Y2=1.385
r121 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.79 $Y=1.55 $X2=4.79
+ $Y2=2.4
r122 1 39 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.22
+ $X2=4.425 $Y2=1.385
r123 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.425 $Y=1.22
+ $X2=4.425 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%C_N 1 3 4 6 7 9 10 15
c38 10 0 1.83401e-19 $X=6.96 $Y=1.295
r39 15 17 26.3594 $w=4.48e-07 $l=2.45e-07 $layer=POLY_cond $X=6.93 $Y=1.49
+ $X2=7.175 $Y2=1.49
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.385 $X2=6.93 $Y2=1.385
r41 13 15 22.0558 $w=4.48e-07 $l=2.05e-07 $layer=POLY_cond $X=6.725 $Y=1.49
+ $X2=6.93 $Y2=1.49
r42 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.93 $Y=1.295 $X2=6.93
+ $Y2=1.385
r43 7 17 24.1837 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=7.175 $Y=1.76
+ $X2=7.175 $Y2=1.49
r44 7 9 133.889 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=7.175 $Y=1.76 $X2=7.175
+ $Y2=2.26
r45 4 13 24.1837 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=6.725 $Y=1.76
+ $X2=6.725 $Y2=1.49
r46 4 6 133.889 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=6.725 $Y=1.76 $X2=6.725
+ $Y2=2.26
r47 1 13 18.2902 $w=4.48e-07 $l=3.44674e-07 $layer=POLY_cond $X=6.555 $Y=1.22
+ $X2=6.725 $Y2=1.49
r48 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.555 $Y=1.22 $X2=6.555
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%A_27_368# 1 2 3 4 5 18 22 23 26 28 32 34 35
+ 43 44 45
c63 28 0 7.99092e-20 $X=2.04 $Y=2.99
c64 3 0 7.54847e-20 $X=2.07 $Y=1.84
r65 45 48 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.005 $Y=2.665
+ $X2=4.005 $Y2=2.745
r66 42 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=2.745
+ $X2=3.27 $Y2=2.745
r67 42 43 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=2.745
+ $X2=2.94 $Y2=2.745
r68 38 39 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.205 $Y=2.745
+ $X2=2.205 $Y2=2.99
r69 35 38 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.205 $Y=2.665
+ $X2=2.205 $Y2=2.745
r70 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=2.665
+ $X2=4.005 $Y2=2.665
r71 32 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.84 $Y=2.665
+ $X2=3.27 $Y2=2.665
r72 31 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=2.665
+ $X2=2.205 $Y2=2.665
r73 31 43 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.37 $Y=2.665
+ $X2=2.94 $Y2=2.665
r74 29 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.99
+ $X2=1.23 $Y2=2.99
r75 28 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=2.99
+ $X2=2.205 $Y2=2.99
r76 28 29 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.04 $Y=2.99
+ $X2=1.315 $Y2=2.99
r77 24 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.99
r78 24 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.455
r79 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.23 $Y2=2.99
r80 22 23 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.445 $Y2=2.99
r81 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r82 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r83 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r84 5 48 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.84 $X2=4.005 $Y2=2.745
r85 4 42 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.84 $X2=3.105 $Y2=2.745
r86 3 38 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=2.07
+ $Y=1.84 $X2=2.205 $Y2=2.745
r87 2 26 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.455
r88 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r89 1 18 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%A_129_368# 1 2 3 4 15 17 21 23 25 27 30 33
+ 37
c66 17 0 8.09075e-20 $X=4.795 $Y=2.325
r67 33 35 10.8284 $w=3.38e-07 $l=3e-07 $layer=LI1_cond $X=1.697 $Y=2.325
+ $X2=1.697 $Y2=2.625
r68 32 33 10.4675 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=1.697 $Y=2.035
+ $X2=1.697 $Y2=2.325
r69 25 42 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=2.23
+ $X2=5.945 $Y2=2.145
r70 25 27 10.8842 $w=2.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.945 $Y=2.23
+ $X2=5.945 $Y2=2.485
r71 24 37 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=5.1 $Y=2.145
+ $X2=4.947 $Y2=2.145
r72 23 42 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.81 $Y=2.145
+ $X2=5.945 $Y2=2.145
r73 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.81 $Y=2.145
+ $X2=5.1 $Y2=2.145
r74 21 40 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.015 $Y=2.485
+ $X2=5.015 $Y2=2.41
r75 18 33 4.76605 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.87 $Y=2.325
+ $X2=1.697 $Y2=2.325
r76 17 40 5.45178 $w=3.03e-07 $l=8.5e-08 $layer=LI1_cond $X=4.947 $Y=2.325
+ $X2=4.947 $Y2=2.41
r77 17 37 6.8013 $w=3.03e-07 $l=1.8e-07 $layer=LI1_cond $X=4.947 $Y=2.325
+ $X2=4.947 $Y2=2.145
r78 17 18 190.829 $w=1.68e-07 $l=2.925e-06 $layer=LI1_cond $X=4.795 $Y=2.325
+ $X2=1.87 $Y2=2.325
r79 16 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r80 15 32 4.76605 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.525 $Y=2.035
+ $X2=1.697 $Y2=2.035
r81 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.525 $Y=2.035
+ $X2=0.945 $Y2=2.035
r82 4 42 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=1.84 $X2=5.915 $Y2=2.145
r83 4 27 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=5.78
+ $Y=1.84 $X2=5.915 $Y2=2.485
r84 3 37 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.84 $X2=5.015 $Y2=2.145
r85 3 21 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=4.88
+ $Y=1.84 $X2=5.015 $Y2=2.485
r86 2 35 600 $w=1.7e-07 $l=8.5443e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.69 $Y2=2.625
r87 2 32 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.69 $Y2=2.035
r88 1 30 300 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=2 $X=0.645
+ $Y=1.84 $X2=0.78 $Y2=2.075
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%Y 1 2 3 4 5 6 7 8 27 30 33 35 37 41 45 47 51
+ 53 57 59 63 66 69 71 72 73 74
c137 69 0 9.05221e-20 $X=2.275 $Y=1.08
c138 41 0 7.54847e-20 $X=3.555 $Y=1.985
r139 70 74 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.82
+ $X2=2.16 $Y2=1.665
r140 68 74 24.3015 $w=2.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.16 $Y=1.18
+ $X2=2.16 $Y2=1.665
r141 68 69 6.65862 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.08
+ $X2=2.275 $Y2=1.08
r142 61 63 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.77 $Y=0.88
+ $X2=5.77 $Y2=0.515
r143 60 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0.965
+ $X2=4.64 $Y2=0.965
r144 59 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.605 $Y=0.965
+ $X2=5.77 $Y2=0.88
r145 59 60 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.605 $Y=0.965
+ $X2=4.805 $Y2=0.965
r146 55 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.88
+ $X2=4.64 $Y2=0.965
r147 55 57 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.64 $Y=0.88
+ $X2=4.64 $Y2=0.515
r148 54 72 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.805 $Y=0.965
+ $X2=3.64 $Y2=1.015
r149 53 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0.965
+ $X2=4.64 $Y2=0.965
r150 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.475 $Y=0.965
+ $X2=3.805 $Y2=0.965
r151 49 72 0.89609 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.64 $Y2=1.015
r152 49 51 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.64 $Y2=0.515
r153 48 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=1.065
+ $X2=2.71 $Y2=1.065
r154 47 72 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.475 $Y=1.065
+ $X2=3.64 $Y2=1.015
r155 47 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.475 $Y=1.065
+ $X2=2.795 $Y2=1.065
r156 43 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.98
+ $X2=2.71 $Y2=1.065
r157 43 45 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.71 $Y=0.98
+ $X2=2.71 $Y2=0.515
r158 39 41 41.4879 $w=2.48e-07 $l=9e-07 $layer=LI1_cond $X=2.655 $Y=1.945
+ $X2=3.555 $Y2=1.945
r159 37 70 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=2.275 $Y=1.945
+ $X2=2.16 $Y2=1.82
r160 37 39 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=2.275 $Y=1.945
+ $X2=2.655 $Y2=1.945
r161 35 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.065
+ $X2=2.71 $Y2=1.065
r162 35 69 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.625 $Y=1.065
+ $X2=2.275 $Y2=1.065
r163 31 68 21.0727 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=1.08
+ $X2=2.16 $Y2=1.08
r164 31 66 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=1.08
+ $X2=1.615 $Y2=1.08
r165 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.78 $Y=0.98
+ $X2=1.78 $Y2=0.515
r166 30 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.945 $Y=1.095
+ $X2=1.615 $Y2=1.095
r167 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r168 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.515
r169 8 41 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.555 $Y2=1.985
r170 7 39 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.84 $X2=2.655 $Y2=1.985
r171 6 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.63
+ $Y=0.37 $X2=5.77 $Y2=0.515
r172 5 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.5
+ $Y=0.37 $X2=4.64 $Y2=0.515
r173 4 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.37 $X2=3.64 $Y2=0.515
r174 3 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.515
r175 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.64
+ $Y=0.37 $X2=1.78 $Y2=0.515
r176 1 27 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%VPWR 1 2 3 4 15 19 23 27 29 31 33 41 46 51
+ 57 60 63 67
r94 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 55 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r99 55 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r100 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r101 52 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.415 $Y2=3.33
r102 52 54 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 51 66 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.235 $Y=3.33
+ $X2=7.457 $Y2=3.33
r104 51 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=3.33
+ $X2=6.96 $Y2=3.33
r105 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r106 50 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r107 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r108 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=3.33
+ $X2=5.465 $Y2=3.33
r109 47 49 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.63 $Y=3.33 $X2=6
+ $Y2=3.33
r110 46 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6.415 $Y2=3.33
r111 46 49 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=3.33 $X2=6
+ $Y2=3.33
r112 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r115 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.565 $Y2=3.33
r116 42 44 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 41 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.465 $Y2=3.33
r118 41 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 40 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r121 35 39 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r122 35 36 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r123 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.565 $Y2=3.33
r124 33 39 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33 $X2=4.08
+ $Y2=3.33
r125 31 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 31 36 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=0.24 $Y2=3.33
r127 27 66 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.457 $Y2=3.33
r128 27 29 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=2.16
r129 23 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.415 $Y=2.145
+ $X2=6.415 $Y2=2.825
r130 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=3.33
r131 21 26 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.415 $Y=3.245
+ $X2=6.415 $Y2=2.825
r132 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=3.33
r133 17 19 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=2.485
r134 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=3.33
r135 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=2.745
r136 4 29 300 $w=1.7e-07 $l=3.81576e-07 $layer=licon1_PDIFF $count=2 $X=7.265
+ $Y=1.84 $X2=7.4 $Y2=2.16
r137 3 26 600 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=1.84 $X2=6.415 $Y2=2.825
r138 3 23 300 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=2 $X=6.23
+ $Y=1.84 $X2=6.415 $Y2=2.145
r139 2 19 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=5.33
+ $Y=1.84 $X2=5.465 $Y2=2.485
r140 1 15 600 $w=1.7e-07 $l=9.74808e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.84 $X2=4.565 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_4%VGND 1 2 3 4 5 6 7 22 24 28 30 34 38 42 44
+ 48 52 55 56 57 59 64 69 82 83 89 92 95 98 101
r109 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r110 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r111 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r112 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r113 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r114 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r115 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r116 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r117 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r119 79 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r120 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r121 77 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r122 77 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r123 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r124 74 101 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.435 $Y=0
+ $X2=5.205 $Y2=0
r125 74 76 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.435 $Y=0 $X2=6
+ $Y2=0
r126 73 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r127 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r128 70 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r129 70 72 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r130 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r131 69 72 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.6
+ $Y2=0
r132 68 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r133 68 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r134 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r135 65 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r136 65 67 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.64 $Y2=0
r137 64 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r138 64 67 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r139 63 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r140 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r141 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r142 60 86 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r143 60 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r144 59 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r145 59 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r146 57 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r147 57 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r148 55 76 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=6
+ $Y2=0
r149 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=6.27
+ $Y2=0
r150 54 79 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.48
+ $Y2=0
r151 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.27
+ $Y2=0
r152 50 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0
r153 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0.515
r154 46 101 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=0.085
+ $X2=5.205 $Y2=0
r155 46 48 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=5.205 $Y=0.085
+ $X2=5.205 $Y2=0.515
r156 45 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r157 44 101 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=5.205 $Y2=0
r158 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=4.305 $Y2=0
r159 40 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r160 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.53
r161 36 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r162 36 38 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.645
r163 32 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r164 32 34 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.645
r165 31 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r166 30 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r167 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.445 $Y2=0
r168 26 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r169 26 28 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.675
r170 22 86 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r171 22 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r172 7 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.13
+ $Y=0.37 $X2=6.27 $Y2=0.515
r173 6 48 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.37 $X2=5.205 $Y2=0.515
r174 5 42 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.14 $Y2=0.53
r175 4 38 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.14 $Y2=0.645
r176 3 34 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.28 $Y2=0.645
r177 2 28 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.675
r178 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__a221o_4.pex.spice
* Created: Wed Sep  2 11:52:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A221O_4%A1 4 5 7 9 10 14 15 17 19 22 27 28 33
c67 14 0 1.82203e-19 $X=1.125 $Y=0.995
c68 5 0 1.22861e-20 $X=0.71 $Y=1.48
r69 33 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.6 $Y=0.4 $X2=1.6
+ $Y2=0.49
r70 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6 $Y=0.4
+ $X2=1.6 $Y2=0.4
r71 27 38 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.68 $Y=0.41
+ $X2=1.68 $Y2=0.565
r72 27 34 2.97405 $w=3.08e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=0.41 $X2=1.6
+ $Y2=0.41
r73 27 28 21.0727 $w=1.68e-07 $l=3.23e-07 $layer=LI1_cond $X=1.68 $Y=0.602
+ $X2=1.68 $Y2=0.925
r74 27 38 2.4139 $w=1.68e-07 $l=3.7e-08 $layer=LI1_cond $X=1.68 $Y=0.602
+ $X2=1.68 $Y2=0.565
r75 20 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.2 $Y=0.49
+ $X2=1.125 $Y2=0.49
r76 19 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=0.49
+ $X2=1.6 $Y2=0.49
r77 19 20 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=1.435 $Y=0.49 $X2=1.2
+ $Y2=0.49
r78 15 23 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.28 $Y=1.465
+ $X2=1.125 $Y2=1.465
r79 15 17 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=1.28 $Y=1.54
+ $X2=1.28 $Y2=2.38
r80 12 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.125 $Y=1.39
+ $X2=1.125 $Y2=1.465
r81 12 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.125 $Y=1.39
+ $X2=1.125 $Y2=0.995
r82 11 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.125 $Y=0.565
+ $X2=1.125 $Y2=0.49
r83 11 14 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.125 $Y=0.565
+ $X2=1.125 $Y2=0.995
r84 9 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.05 $Y=0.49
+ $X2=1.125 $Y2=0.49
r85 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.05 $Y=0.49 $X2=0.77
+ $Y2=0.49
r86 5 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.71 $Y=1.48 $X2=0.71
+ $Y2=1.39
r87 5 7 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=0.71 $Y=1.48 $X2=0.71
+ $Y2=2.38
r88 4 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.695 $Y=0.995
+ $X2=0.695 $Y2=1.39
r89 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.695 $Y=0.565
+ $X2=0.77 $Y2=0.49
r90 1 4 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.695 $Y=0.565
+ $X2=0.695 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%A2 3 8 11 13 15 20 22 25
c64 13 0 1.08291e-19 $X=2.89 $Y=1.33
r65 25 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.44 $Y=0.34
+ $X2=2.44 $Y2=0.505
r66 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=0.34 $X2=2.44 $Y2=0.34
r67 22 26 6.90263 $w=3.8e-07 $l=2.7037e-07 $layer=LI1_cond $X=2.64 $Y=0.555
+ $X2=2.515 $Y2=0.34
r68 13 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.89 $Y=1.33
+ $X2=2.89 $Y2=1.405
r69 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.89 $Y=1.33
+ $X2=2.89 $Y2=0.935
r70 9 20 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.625 $Y=1.405
+ $X2=2.89 $Y2=1.405
r71 9 18 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.405
+ $X2=2.46 $Y2=1.405
r72 9 11 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=2.625 $Y=1.48 $X2=2.625
+ $Y2=2.38
r73 8 28 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.46 $Y=0.935
+ $X2=2.46 $Y2=0.505
r74 6 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.46 $Y=1.33 $X2=2.46
+ $Y2=1.405
r75 6 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.46 $Y=1.33 $X2=2.46
+ $Y2=0.935
r76 1 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.175 $Y=1.405
+ $X2=2.46 $Y2=1.405
r77 1 3 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=2.175 $Y=1.48 $X2=2.175
+ $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%A_154_135# 1 2 3 4 13 15 16 18 21 23 25 28
+ 30 32 33 35 37 39 42 45 46 47 51 55 58 61 63 67 72 73 77 78
c208 58 0 1.9796e-19 $X=6.005 $Y=1.6
c209 55 0 1.2395e-19 $X=5.775 $Y=0.745
c210 47 0 1.86464e-19 $X=3.795 $Y=1.55
c211 37 0 1.44963e-19 $X=4.67 $Y=1.35
c212 33 0 1.41556e-19 $X=4.585 $Y=1.69
r213 79 80 21.8406 $w=3.2e-07 $l=1.45e-07 $layer=POLY_cond $X=3.235 $Y=1.565
+ $X2=3.38 $Y2=1.565
r214 71 83 7.53125 $w=3.2e-07 $l=5e-08 $layer=POLY_cond $X=3.76 $Y=1.565
+ $X2=3.81 $Y2=1.565
r215 70 72 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=1.55
+ $X2=3.595 $Y2=1.55
r216 70 71 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.515 $X2=3.76 $Y2=1.515
r217 65 67 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.28 $Y=1.6
+ $X2=8.28 $Y2=0.76
r218 64 78 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=1.685
+ $X2=6.085 $Y2=1.685
r219 63 65 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.115 $Y=1.685
+ $X2=8.28 $Y2=1.6
r220 63 64 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=8.115 $Y=1.685
+ $X2=6.25 $Y2=1.685
r221 59 78 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=1.77
+ $X2=6.085 $Y2=1.685
r222 59 61 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.085 $Y=1.77
+ $X2=6.085 $Y2=2.105
r223 58 78 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.005 $Y=1.6
+ $X2=6.085 $Y2=1.685
r224 57 77 3.70735 $w=2.5e-07 $l=1.92873e-07 $layer=LI1_cond $X=6.005 $Y=1.3
+ $X2=5.85 $Y2=1.215
r225 57 58 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.005 $Y=1.3
+ $X2=6.005 $Y2=1.6
r226 53 77 3.70735 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=5.775 $Y=1.13
+ $X2=5.85 $Y2=1.215
r227 53 55 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.775 $Y=1.13
+ $X2=5.775 $Y2=0.745
r228 52 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=1.215
+ $X2=4.795 $Y2=1.215
r229 51 77 2.76166 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.61 $Y=1.215
+ $X2=5.85 $Y2=1.215
r230 51 52 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.61 $Y=1.215
+ $X2=4.88 $Y2=1.215
r231 50 85 30.125 $w=3.2e-07 $l=2e-07 $layer=POLY_cond $X=4.44 $Y=1.565 $X2=4.24
+ $Y2=1.565
r232 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.44
+ $Y=1.515 $X2=4.44 $Y2=1.515
r233 47 70 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.795 $Y=1.55
+ $X2=3.76 $Y2=1.55
r234 47 49 18.5831 $w=3.98e-07 $l=6.45e-07 $layer=LI1_cond $X=3.795 $Y=1.55
+ $X2=4.44 $Y2=1.55
r235 46 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.795 $Y=1.55
+ $X2=4.795 $Y2=1.215
r236 46 49 7.77899 $w=3.98e-07 $l=2.7e-07 $layer=LI1_cond $X=4.71 $Y=1.55
+ $X2=4.44 $Y2=1.55
r237 45 72 164.406 $w=1.68e-07 $l=2.52e-06 $layer=LI1_cond $X=1.075 $Y=1.665
+ $X2=3.595 $Y2=1.665
r238 40 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.91 $Y=1.58
+ $X2=1.075 $Y2=1.665
r239 40 42 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.91 $Y=1.58
+ $X2=0.91 $Y2=1.165
r240 37 88 20.4921 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.67 $Y=1.35
+ $X2=4.67 $Y2=1.565
r241 37 39 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.67 $Y=1.35
+ $X2=4.67 $Y2=0.87
r242 33 88 12.8031 $w=3.2e-07 $l=8.5e-08 $layer=POLY_cond $X=4.585 $Y=1.565
+ $X2=4.67 $Y2=1.565
r243 33 50 21.8406 $w=3.2e-07 $l=1.45e-07 $layer=POLY_cond $X=4.585 $Y=1.565
+ $X2=4.44 $Y2=1.565
r244 33 35 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=4.585 $Y=1.69
+ $X2=4.585 $Y2=2.4
r245 30 85 20.4921 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.24 $Y=1.35
+ $X2=4.24 $Y2=1.565
r246 30 32 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.24 $Y=1.35
+ $X2=4.24 $Y2=0.87
r247 26 85 15.8156 $w=3.2e-07 $l=1.05e-07 $layer=POLY_cond $X=4.135 $Y=1.565
+ $X2=4.24 $Y2=1.565
r248 26 83 48.9531 $w=3.2e-07 $l=3.25e-07 $layer=POLY_cond $X=4.135 $Y=1.565
+ $X2=3.81 $Y2=1.565
r249 26 28 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=4.135 $Y=1.69
+ $X2=4.135 $Y2=2.4
r250 23 83 20.4921 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=3.81 $Y2=1.565
r251 23 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=3.81 $Y2=0.87
r252 19 71 11.2969 $w=3.2e-07 $l=7.5e-08 $layer=POLY_cond $X=3.685 $Y=1.565
+ $X2=3.76 $Y2=1.565
r253 19 80 45.9406 $w=3.2e-07 $l=3.05e-07 $layer=POLY_cond $X=3.685 $Y=1.565
+ $X2=3.38 $Y2=1.565
r254 19 21 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=3.685 $Y=1.69
+ $X2=3.685 $Y2=2.4
r255 16 80 20.4921 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=1.565
r256 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=0.87
r257 13 79 16.2157 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.235 $Y=1.78
+ $X2=3.235 $Y2=1.565
r258 13 15 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.235 $Y=1.78
+ $X2=3.235 $Y2=2.4
r259 4 61 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=1.96 $X2=6.085 $Y2=2.105
r260 3 67 182 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_NDIFF $count=1 $X=8.14
+ $Y=0.38 $X2=8.28 $Y2=0.76
r261 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.635
+ $Y=0.6 $X2=5.775 $Y2=0.745
r262 1 42 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=0.77
+ $Y=0.675 $X2=0.91 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%C1 3 7 11 13 14 15 17 20 21
c68 20 0 2.81466e-20 $X=5.52 $Y=1.665
c69 15 0 1.9796e-19 $X=6.31 $Y=1.715
c70 11 0 5.30963e-20 $X=5.99 $Y=0.92
r71 26 28 43.2755 $w=3.23e-07 $l=2.9e-07 $layer=POLY_cond $X=5.57 $Y=1.62
+ $X2=5.86 $Y2=1.62
r72 24 26 1.49226 $w=3.23e-07 $l=1e-08 $layer=POLY_cond $X=5.56 $Y=1.62 $X2=5.57
+ $Y2=1.62
r73 20 21 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.57 $Y=1.635 $X2=5.57
+ $Y2=2.035
r74 20 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.635 $X2=5.57 $Y2=1.635
r75 15 19 54.3311 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=6.31 $Y=1.715 $X2=6.31
+ $Y2=1.515
r76 15 17 289.589 $w=1.8e-07 $l=7.45e-07 $layer=POLY_cond $X=6.31 $Y=1.715
+ $X2=6.31 $Y2=2.46
r77 13 19 4.22461 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.22 $Y=1.515 $X2=6.31
+ $Y2=1.515
r78 13 14 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.22 $Y=1.515
+ $X2=6.065 $Y2=1.515
r79 9 14 25.1311 $w=3.23e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.99 $Y=1.44
+ $X2=6.065 $Y2=1.515
r80 9 28 19.3994 $w=3.23e-07 $l=2.3622e-07 $layer=POLY_cond $X=5.99 $Y=1.44
+ $X2=5.86 $Y2=1.62
r81 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.99 $Y=1.44 $X2=5.99
+ $Y2=0.92
r82 5 28 16.4327 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=5.86 $Y=1.8 $X2=5.86
+ $Y2=1.62
r83 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.86 $Y=1.8 $X2=5.86
+ $Y2=2.46
r84 1 24 20.7134 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.56 $Y=1.44 $X2=5.56
+ $Y2=1.62
r85 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.56 $Y=1.44 $X2=5.56
+ $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%B2 3 6 8 10 11 14 18 21 23 26 30 32 37 39 42
c93 42 0 1.2395e-19 $X=6.635 $Y=0.505
r94 35 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.635 $Y=0.34
+ $X2=6.635 $Y2=0.505
r95 35 39 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=6.635 $Y=0.34
+ $X2=6.635 $Y2=0.2
r96 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.635
+ $Y=0.34 $X2=6.635 $Y2=0.34
r97 32 37 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=6.945 $Y=0.38
+ $X2=6.945 $Y2=0.555
r98 32 34 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=6.845 $Y=0.38
+ $X2=6.635 $Y2=0.38
r99 28 30 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.475 $Y=1.405
+ $X2=7.575 $Y2=1.405
r100 23 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.575 $Y=1.33
+ $X2=7.575 $Y2=1.405
r101 22 23 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=7.575 $Y=0.275
+ $X2=7.575 $Y2=1.33
r102 21 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.475 $Y=1.625
+ $X2=7.475 $Y2=1.7
r103 20 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.475 $Y=1.48
+ $X2=7.475 $Y2=1.405
r104 20 21 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.475 $Y=1.48
+ $X2=7.475 $Y2=1.625
r105 16 26 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=7.21 $Y=1.7
+ $X2=7.475 $Y2=1.7
r106 16 24 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.21 $Y=1.7
+ $X2=7.085 $Y2=1.7
r107 16 18 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=7.21 $Y=1.775
+ $X2=7.21 $Y2=2.46
r108 12 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.085 $Y=1.625
+ $X2=7.085 $Y2=1.7
r109 12 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.085 $Y=1.625
+ $X2=7.085 $Y2=0.935
r110 10 24 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.01 $Y=1.7
+ $X2=7.085 $Y2=1.7
r111 10 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.01 $Y=1.7
+ $X2=6.85 $Y2=1.7
r112 9 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=0.2
+ $X2=6.635 $Y2=0.2
r113 8 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.5 $Y=0.2
+ $X2=7.575 $Y2=0.275
r114 8 9 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=7.5 $Y=0.2 $X2=6.8
+ $Y2=0.2
r115 4 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.76 $Y=1.775
+ $X2=6.85 $Y2=1.7
r116 4 6 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=6.76 $Y=1.775
+ $X2=6.76 $Y2=2.46
r117 3 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.655 $Y=0.935
+ $X2=6.655 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%B1 3 7 11 15 17 22 23 27 35
c51 7 0 3.65222e-20 $X=8.065 $Y=0.7
r52 28 35 0.810495 $w=5.38e-07 $l=2e-08 $layer=LI1_cond $X=9.115 $Y=1.48
+ $X2=9.095 $Y2=1.48
r53 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.115
+ $Y=1.465 $X2=9.115 $Y2=1.465
r54 23 28 5.42665 $w=5.38e-07 $l=2.45e-07 $layer=LI1_cond $X=9.36 $Y=1.48
+ $X2=9.115 $Y2=1.48
r55 22 35 5.7146 $w=4.48e-07 $l=2.15e-07 $layer=LI1_cond $X=8.88 $Y=1.525
+ $X2=9.095 $Y2=1.525
r56 20 21 8.23292 $w=3.22e-07 $l=5.5e-08 $layer=POLY_cond $X=8.44 $Y=1.51
+ $X2=8.495 $Y2=1.51
r57 17 27 72.1676 $w=4.2e-07 $l=5.45e-07 $layer=POLY_cond $X=8.57 $Y=1.51
+ $X2=9.115 $Y2=1.51
r58 17 21 11.3528 $w=4.2e-07 $l=7.5e-08 $layer=POLY_cond $X=8.57 $Y=1.51
+ $X2=8.495 $Y2=1.51
r59 13 21 20.6399 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.495 $Y=1.3
+ $X2=8.495 $Y2=1.51
r60 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.495 $Y=1.3 $X2=8.495
+ $Y2=0.7
r61 9 20 16.3606 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.44 $Y=1.72 $X2=8.44
+ $Y2=1.51
r62 9 11 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=8.44 $Y=1.72 $X2=8.44
+ $Y2=2.46
r63 5 20 56.1335 $w=3.22e-07 $l=3.75e-07 $layer=POLY_cond $X=8.065 $Y=1.51
+ $X2=8.44 $Y2=1.51
r64 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.065 $Y=1.38
+ $X2=8.065 $Y2=0.7
r65 1 5 17.2143 $w=3.22e-07 $l=2.61247e-07 $layer=POLY_cond $X=7.95 $Y=1.72
+ $X2=8.065 $Y2=1.51
r66 1 3 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=7.95 $Y=1.72 $X2=7.95
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%VPWR 1 2 3 4 5 18 22 26 30 33 34 36 37 39 40
+ 42 43 44 50 68 69 72
r89 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r90 72 75 11.0682 $w=6.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.73 $Y=2.71
+ $X2=1.73 $Y2=3.33
r91 68 69 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r92 66 69 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=9.36 $Y2=3.33
r93 65 68 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=9.36 $Y2=3.33
r94 65 66 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r98 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r99 57 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 54 75 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.73 $Y2=3.33
r102 54 56 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 50 75 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.73 $Y2=3.33
r106 50 52 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 48 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r109 44 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 44 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 42 62 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.81 $Y2=3.33
r113 41 65 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.975 $Y=3.33
+ $X2=5.04 $Y2=3.33
r114 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=3.33
+ $X2=4.81 $Y2=3.33
r115 39 59 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.91 $Y2=3.33
r117 38 62 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=3.91 $Y2=3.33
r119 36 56 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.01 $Y2=3.33
r121 35 59 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r122 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.01 $Y2=3.33
r123 33 47 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=3.33 $X2=0.24
+ $Y2=3.33
r124 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.485 $Y2=3.33
r125 32 52 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.65 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=3.33
+ $X2=0.485 $Y2=3.33
r127 28 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=3.245
+ $X2=4.81 $Y2=3.33
r128 28 30 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.81 $Y=3.245
+ $X2=4.81 $Y2=2.8
r129 24 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=3.245
+ $X2=3.91 $Y2=3.33
r130 24 26 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.91 $Y=3.245
+ $X2=3.91 $Y2=2.8
r131 20 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=3.33
r132 20 22 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=2.8
r133 16 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.485 $Y=3.245
+ $X2=0.485 $Y2=3.33
r134 16 18 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=0.485 $Y=3.245
+ $X2=0.485 $Y2=2.345
r135 5 30 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=4.675
+ $Y=1.84 $X2=4.81 $Y2=2.8
r136 4 26 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=3.775
+ $Y=1.84 $X2=3.91 $Y2=2.8
r137 3 22 600 $w=1.7e-07 $l=1.05726e-06 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.88 $X2=3.01 $Y2=2.8
r138 2 72 300 $w=1.7e-07 $l=1.06245e-06 $layer=licon1_PDIFF $count=2 $X=1.37
+ $Y=1.88 $X2=1.9 $Y2=2.71
r139 1 18 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.36
+ $Y=1.88 $X2=0.485 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%A_160_376# 1 2 3 4 15 19 21 22 23 28 30 33
+ 37
r88 33 35 5.04967 $w=3.02e-07 $l=1.25e-07 $layer=LI1_cond $X=6.985 $Y=2.445
+ $X2=6.985 $Y2=2.57
r89 24 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.15 $Y=2.025
+ $X2=6.985 $Y2=2.025
r90 23 37 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.01 $Y=2.025
+ $X2=8.195 $Y2=2.025
r91 23 24 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=8.01 $Y=2.025
+ $X2=7.15 $Y2=2.025
r92 22 33 3.2529 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=2.36
+ $X2=6.985 $Y2=2.445
r93 21 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=2.11
+ $X2=6.985 $Y2=2.025
r94 21 22 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.985 $Y=2.11
+ $X2=6.985 $Y2=2.36
r95 20 30 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=2.565 $Y=2.445
+ $X2=2.4 $Y2=2.395
r96 19 33 4.10007 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.82 $Y=2.445
+ $X2=6.985 $Y2=2.445
r97 19 20 277.599 $w=1.68e-07 $l=4.255e-06 $layer=LI1_cond $X=6.82 $Y=2.445
+ $X2=2.565 $Y2=2.445
r98 16 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=2.345
+ $X2=1.055 $Y2=2.345
r99 15 30 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=2.235 $Y=2.345
+ $X2=2.4 $Y2=2.395
r100 15 16 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=2.235 $Y=2.345
+ $X2=1.22 $Y2=2.345
r101 4 37 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=8.04
+ $Y=1.96 $X2=8.195 $Y2=2.105
r102 3 35 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=6.85
+ $Y=1.96 $X2=6.985 $Y2=2.57
r103 3 32 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.85
+ $Y=1.96 $X2=6.985 $Y2=2.105
r104 2 30 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=2.265
+ $Y=1.88 $X2=2.4 $Y2=2.345
r105 1 28 300 $w=1.7e-07 $l=5.78619e-07 $layer=licon1_PDIFF $count=2 $X=0.8
+ $Y=1.88 $X2=1.055 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%X 1 2 3 4 14 15 19 21 25 27 31 34 35 36 37
+ 40 42 46
c120 34 0 2.4855e-20 $X=2.85 $Y=2.055
c121 31 0 1.44963e-19 $X=4.455 $Y=0.645
r122 46 49 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=3.12 $Y=1.095
+ $X2=3.12 $Y2=1.295
r123 42 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r124 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.295
r125 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.295
+ $X2=0.24 $Y2=1.295
r126 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=3.12 $Y2=1.295
r127 36 37 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=0.385 $Y2=1.295
r128 33 40 31.3164 $w=2.28e-07 $l=6.25e-07 $layer=LI1_cond $X=0.24 $Y=1.92
+ $X2=0.24 $Y2=1.295
r129 29 31 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=4.415 $Y=1.01
+ $X2=4.415 $Y2=0.645
r130 28 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=1.095
+ $X2=3.595 $Y2=1.095
r131 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.29 $Y=1.095
+ $X2=4.415 $Y2=1.01
r132 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.29 $Y=1.095
+ $X2=3.76 $Y2=1.095
r133 23 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=1.01
+ $X2=3.595 $Y2=1.095
r134 23 25 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.595 $Y=1.01
+ $X2=3.595 $Y2=0.645
r135 22 46 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.235 $Y=1.095
+ $X2=3.12 $Y2=1.095
r136 21 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=1.095
+ $X2=3.595 $Y2=1.095
r137 21 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.43 $Y=1.095
+ $X2=3.235 $Y2=1.095
r138 17 19 38.4148 $w=2.68e-07 $l=9e-07 $layer=LI1_cond $X=3.46 $Y=2.055
+ $X2=4.36 $Y2=2.055
r139 15 34 13.0976 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.12 $Y=2.055
+ $X2=2.85 $Y2=2.055
r140 15 17 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.12 $Y=2.055
+ $X2=3.46 $Y2=2.055
r141 14 33 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.005
+ $X2=0.24 $Y2=1.92
r142 14 34 162.775 $w=1.68e-07 $l=2.495e-06 $layer=LI1_cond $X=0.355 $Y=2.005
+ $X2=2.85 $Y2=2.005
r143 4 19 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=4.225
+ $Y=1.84 $X2=4.36 $Y2=2.05
r144 3 17 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.84 $X2=3.46 $Y2=2.05
r145 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.315
+ $Y=0.5 $X2=4.455 $Y2=0.645
r146 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.5 $X2=3.595 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%A_1102_392# 1 2 3 4 13 17 21 23 27 33 34
r42 32 33 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=2.887
+ $X2=6.7 $Y2=2.887
r43 27 30 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.705 $Y=2.105
+ $X2=8.705 $Y2=2.815
r44 25 30 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.705 $Y=2.905
+ $X2=8.705 $Y2=2.815
r45 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=2.99
+ $X2=7.59 $Y2=2.99
r46 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.58 $Y=2.99
+ $X2=8.705 $Y2=2.905
r47 23 24 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.58 $Y=2.99
+ $X2=7.755 $Y2=2.99
r48 19 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=2.905
+ $X2=7.59 $Y2=2.99
r49 19 21 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=7.59 $Y=2.905
+ $X2=7.59 $Y2=2.38
r50 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.425 $Y=2.99
+ $X2=7.59 $Y2=2.99
r51 17 33 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.425 $Y=2.99
+ $X2=6.7 $Y2=2.99
r52 13 32 0.6761 $w=3.73e-07 $l=2.2e-08 $layer=LI1_cond $X=6.513 $Y=2.887
+ $X2=6.535 $Y2=2.887
r53 13 15 26.9825 $w=3.73e-07 $l=8.78e-07 $layer=LI1_cond $X=6.513 $Y=2.887
+ $X2=5.635 $Y2=2.887
r54 4 30 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.53
+ $Y=1.96 $X2=8.665 $Y2=2.815
r55 4 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.53
+ $Y=1.96 $X2=8.665 $Y2=2.105
r56 3 21 300 $w=1.7e-07 $l=5.46077e-07 $layer=licon1_PDIFF $count=2 $X=7.3
+ $Y=1.96 $X2=7.59 $Y2=2.38
r57 2 32 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=6.4
+ $Y=1.96 $X2=6.535 $Y2=2.8
r58 1 15 600 $w=1.7e-07 $l=9.00333e-07 $layer=licon1_PDIFF $count=1 $X=5.51
+ $Y=1.96 $X2=5.635 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%A_71_135# 1 2 3 10 15 16 17 20 24
c53 20 0 1.08291e-19 $X=2.675 $Y=1.055
c54 17 0 1.22861e-20 $X=1.425 $Y=1.325
c55 15 0 1.82203e-19 $X=1.34 $Y=1.035
r56 18 20 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=2.635 $Y=1.24
+ $X2=2.635 $Y2=1.055
r57 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.51 $Y=1.325
+ $X2=2.635 $Y2=1.24
r58 16 17 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=2.51 $Y=1.325
+ $X2=1.425 $Y2=1.325
r59 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.34 $Y=1.24
+ $X2=1.425 $Y2=1.325
r60 13 15 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.34 $Y=1.24
+ $X2=1.34 $Y2=1.035
r61 12 15 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.34 $Y=0.905
+ $X2=1.34 $Y2=1.035
r62 11 24 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=0.82
+ $X2=0.44 $Y2=0.82
r63 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.255 $Y=0.82
+ $X2=1.34 $Y2=0.905
r64 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.255 $Y=0.82
+ $X2=0.565 $Y2=0.82
r65 3 20 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.615 $X2=2.675 $Y2=1.055
r66 2 15 182 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.675 $X2=1.34 $Y2=1.035
r67 1 24 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.355
+ $Y=0.675 $X2=0.48 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%VGND 1 2 3 4 5 6 20 23 27 31 34 37 41 44 45
+ 49 52 53 55 56 60 62 71 79 87 93 94 97 100 103
c142 41 0 3.65222e-20 $X=7.3 $Y=0.925
c143 23 0 1.13409e-19 $X=3.165 $Y=0.66
r144 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r145 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r146 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r147 94 104 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=7.44 $Y2=0
r148 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r149 91 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=7.34 $Y2=0
r150 91 93 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=9.36 $Y2=0
r151 90 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r152 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r153 87 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.215 $Y=0
+ $X2=7.34 $Y2=0
r154 87 89 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.215 $Y=0
+ $X2=6.96 $Y2=0
r155 86 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r156 86 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r157 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r158 83 100 13.8654 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=5.08
+ $Y2=0
r159 83 85 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.44 $Y=0 $X2=6
+ $Y2=0
r160 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r161 79 100 13.8654 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=5.08
+ $Y2=0
r162 79 81 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=4.56
+ $Y2=0
r163 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r164 78 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r165 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r166 75 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.125
+ $Y2=0
r167 75 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.6
+ $Y2=0
r168 74 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r169 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r170 71 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.125
+ $Y2=0
r171 71 73 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.64
+ $Y2=0
r172 70 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r173 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r174 66 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=1.68 $Y2=0
r175 65 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r176 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r177 62 101 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=5.04 $Y2=0
r178 62 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r179 55 85 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6
+ $Y2=0
r180 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.215
+ $Y2=0
r181 54 89 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.3 $Y=0 $X2=6.96
+ $Y2=0
r182 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=0 $X2=6.215
+ $Y2=0
r183 52 77 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=3.6
+ $Y2=0
r184 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.94 $Y=0 $X2=4.025
+ $Y2=0
r185 51 81 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=4.56
+ $Y2=0
r186 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=0 $X2=4.025
+ $Y2=0
r187 44 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0
+ $X2=1.68 $Y2=0
r188 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.02
+ $Y2=0
r189 43 73 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.105 $Y=0
+ $X2=2.64 $Y2=0
r190 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.02
+ $Y2=0
r191 39 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.34 $Y=0.085
+ $X2=7.34 $Y2=0
r192 39 41 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=7.34 $Y=0.085
+ $X2=7.34 $Y2=0.925
r193 35 60 1.50363 $w=2.5e-07 $l=1.43e-07 $layer=LI1_cond $X=6.4 $Y=0.96 $X2=6.4
+ $Y2=0.817
r194 35 37 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=6.4 $Y=0.96
+ $X2=6.4 $Y2=1.115
r195 34 60 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=6.215 $Y=0.817
+ $X2=6.4 $Y2=0.817
r196 33 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.215 $Y=0.085
+ $X2=6.215 $Y2=0
r197 33 34 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.215 $Y=0.085
+ $X2=6.215 $Y2=0.675
r198 29 100 2.92113 $w=7.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=0.085
+ $X2=5.08 $Y2=0
r199 29 31 11.7947 $w=7.18e-07 $l=7.1e-07 $layer=LI1_cond $X=5.08 $Y=0.085
+ $X2=5.08 $Y2=0.795
r200 25 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=0.085
+ $X2=4.025 $Y2=0
r201 25 27 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.025 $Y=0.085
+ $X2=4.025 $Y2=0.66
r202 21 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=0.085
+ $X2=3.125 $Y2=0
r203 21 23 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=3.125 $Y=0.085
+ $X2=3.125 $Y2=0.66
r204 20 49 6.56455 $w=3.93e-07 $l=2.25e-07 $layer=LI1_cond $X=2.02 $Y=0.872
+ $X2=2.245 $Y2=0.872
r205 19 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r206 19 20 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.675
r207 6 41 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.615 $X2=7.3 $Y2=0.925
r208 5 34 182 $w=1.7e-07 $l=2.995e-07 $layer=licon1_NDIFF $count=1 $X=6.065
+ $Y=0.6 $X2=6.295 $Y2=0.76
r209 5 37 182 $w=1.7e-07 $l=6.77016e-07 $layer=licon1_NDIFF $count=1 $X=6.065
+ $Y=0.6 $X2=6.44 $Y2=1.115
r210 4 31 91 $w=1.7e-07 $l=7.32803e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.5 $X2=5.345 $Y2=0.795
r211 3 27 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.5 $X2=4.025 $Y2=0.66
r212 2 23 182 $w=1.7e-07 $l=2.21359e-07 $layer=licon1_NDIFF $count=1 $X=2.965
+ $Y=0.615 $X2=3.165 $Y2=0.66
r213 1 49 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.615 $X2=2.245 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_4%A_1346_123# 1 2 3 12 14 15 19 20 21 24
c51 12 0 5.30963e-20 $X=6.87 $Y=1.055
r52 22 24 4.22562 $w=2.98e-07 $l=1.1e-07 $layer=LI1_cond $X=8.775 $Y=0.425
+ $X2=8.775 $Y2=0.535
r53 20 22 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.625 $Y=0.34
+ $X2=8.775 $Y2=0.425
r54 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.625 $Y=0.34
+ $X2=7.935 $Y2=0.34
r55 17 19 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=7.81 $Y=1.26
+ $X2=7.81 $Y2=0.525
r56 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.81 $Y=0.425
+ $X2=7.935 $Y2=0.34
r57 16 19 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=7.81 $Y=0.425 $X2=7.81
+ $Y2=0.525
r58 14 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.685 $Y=1.345
+ $X2=7.81 $Y2=1.26
r59 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.685 $Y=1.345
+ $X2=7.035 $Y2=1.345
r60 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.87 $Y=1.26
+ $X2=7.035 $Y2=1.345
r61 10 12 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.87 $Y=1.26
+ $X2=6.87 $Y2=1.055
r62 3 24 91 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=2 $X=8.57
+ $Y=0.38 $X2=8.735 $Y2=0.535
r63 2 19 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=7.725
+ $Y=0.38 $X2=7.85 $Y2=0.525
r64 1 12 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=6.73
+ $Y=0.615 $X2=6.87 $Y2=1.055
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
M1000 a_815_508# a_220_419# a_672_392# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=4.915e+11p ps=3.07e+06u
M1001 Q a_863_441# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=1.31878e+12p ps=1.016e+07u
M1002 Q a_863_441# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.48785e+12p ps=1.153e+07u
M1003 VGND a_220_419# a_369_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_588_392# a_27_115# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1005 VGND D a_27_115# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 a_863_441# a_672_392# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1007 a_871_139# a_369_392# a_672_392# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.786e+11p ps=2.52e+06u
M1008 a_672_392# a_369_392# a_588_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_220_419# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 VPWR a_863_441# a_815_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_220_419# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=3.066e+11p pd=2.41e+06u as=0p ps=0u
M1012 VGND a_863_441# a_871_139# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_863_441# a_672_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1014 VPWR D a_27_115# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1015 VPWR a_220_419# a_369_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1016 a_655_79# a_27_115# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1017 a_672_392# a_220_419# a_655_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

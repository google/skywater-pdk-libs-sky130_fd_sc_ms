* File: sky130_fd_sc_ms__and4b_4.pex.spice
* Created: Fri Aug 28 17:14:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4B_4%A_N 3 7 8 11 13
r35 11 14 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.385
+ $X2=0.585 $Y2=1.55
r36 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.385
+ $X2=0.585 $Y2=1.22
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.385 $X2=0.59 $Y2=1.385
r38 8 12 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.37 $X2=0.59
+ $Y2=1.37
r39 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.535 $Y=0.79
+ $X2=0.535 $Y2=1.22
r40 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.505 $Y=2.34
+ $X2=0.505 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%A_199_294# 1 2 3 4 5 18 22 28 32 36 40 44 48
+ 50 51 60 61 62 69 70 73 75 78 80 85 92
c159 80 0 3.04181e-19 $X=6.08 $Y=2.08
c160 75 0 8.69299e-20 $X=3.515 $Y=2.085
c161 60 0 2.26005e-19 $X=2.66 $Y=1.95
r162 91 92 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.575 $Y=1.485
+ $X2=2.59 $Y2=1.485
r163 88 89 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=2.015 $Y=1.485
+ $X2=2.16 $Y2=1.485
r164 84 86 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.52 $Y=1.485
+ $X2=1.535 $Y2=1.485
r165 84 85 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.52 $Y=1.485
+ $X2=1.445 $Y2=1.485
r166 79 80 3.65747 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=2.08
+ $X2=6.08 $Y2=2.08
r167 77 79 7.40856 $w=2.78e-07 $l=1.8e-07 $layer=LI1_cond $X=5.815 $Y=2.08
+ $X2=5.995 $Y2=2.08
r168 77 78 6.95017 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=2.08
+ $X2=5.65 $Y2=2.08
r169 73 80 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.715 $Y=2.095
+ $X2=6.08 $Y2=2.095
r170 70 79 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.995 $Y=1.94
+ $X2=5.995 $Y2=2.08
r171 69 83 10.8397 $w=2.87e-07 $l=3.34201e-07 $layer=LI1_cond $X=5.995 $Y=1.3
+ $X2=6.25 $Y2=1.117
r172 69 70 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.995 $Y=1.3
+ $X2=5.995 $Y2=1.94
r173 68 78 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=4.895 $Y=2.095
+ $X2=5.65 $Y2=2.095
r174 68 75 63.6149 $w=2.48e-07 $l=1.38e-06 $layer=LI1_cond $X=4.895 $Y=2.095
+ $X2=3.515 $Y2=2.095
r175 62 64 25.8233 $w=2.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.745 $Y=2.085
+ $X2=3.35 $Y2=2.085
r176 61 75 5.8439 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.38 $Y=2.085
+ $X2=3.515 $Y2=2.085
r177 61 64 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=3.38 $Y=2.085
+ $X2=3.35 $Y2=2.085
r178 60 62 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.66 $Y=1.95
+ $X2=2.745 $Y2=2.085
r179 59 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.66 $Y=1.65 $X2=2.66
+ $Y2=1.95
r180 58 91 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.33 $Y=1.485
+ $X2=2.575 $Y2=1.485
r181 58 89 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.33 $Y=1.485
+ $X2=2.16 $Y2=1.485
r182 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.485 $X2=2.33 $Y2=1.485
r183 54 88 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.65 $Y=1.485
+ $X2=2.015 $Y2=1.485
r184 54 86 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.65 $Y=1.485
+ $X2=1.535 $Y2=1.485
r185 53 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.65 $Y=1.485
+ $X2=2.33 $Y2=1.485
r186 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.485 $X2=1.65 $Y2=1.485
r187 51 59 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.575 $Y=1.485
+ $X2=2.66 $Y2=1.65
r188 51 57 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.575 $Y=1.485
+ $X2=2.33 $Y2=1.485
r189 46 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.32
+ $X2=2.59 $Y2=1.485
r190 46 48 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.59 $Y=1.32
+ $X2=2.59 $Y2=0.74
r191 42 91 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.65
+ $X2=2.575 $Y2=1.485
r192 42 44 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.575 $Y=1.65
+ $X2=2.575 $Y2=2.4
r193 38 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.32
+ $X2=2.16 $Y2=1.485
r194 38 40 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.16 $Y=1.32
+ $X2=2.16 $Y2=0.74
r195 34 88 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.65
+ $X2=2.015 $Y2=1.485
r196 34 36 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.015 $Y=1.65
+ $X2=2.015 $Y2=2.4
r197 30 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.535 $Y=1.65
+ $X2=1.535 $Y2=1.485
r198 30 32 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=1.535 $Y=1.65
+ $X2=1.535 $Y2=2.4
r199 26 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.32
+ $X2=1.52 $Y2=1.485
r200 26 28 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.52 $Y=1.32
+ $X2=1.52 $Y2=0.74
r201 25 50 6.66866 $w=1.5e-07 $l=2.14243e-07 $layer=POLY_cond $X=1.175 $Y=1.395
+ $X2=0.995 $Y2=1.47
r202 25 85 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.175 $Y=1.395
+ $X2=1.445 $Y2=1.395
r203 20 50 18.8402 $w=1.65e-07 $l=1.91703e-07 $layer=POLY_cond $X=1.09 $Y=1.32
+ $X2=0.995 $Y2=1.47
r204 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.09 $Y=1.32
+ $X2=1.09 $Y2=0.74
r205 16 50 18.8402 $w=1.65e-07 $l=1.27279e-07 $layer=POLY_cond $X=1.085 $Y=1.56
+ $X2=0.995 $Y2=1.47
r206 16 18 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=1.085 $Y=1.56
+ $X2=1.085 $Y2=2.4
r207 5 73 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.58
+ $Y=1.96 $X2=6.715 $Y2=2.135
r208 4 77 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=5.68
+ $Y=1.96 $X2=5.815 $Y2=2.12
r209 3 68 300 $w=1.7e-07 $l=7.77592e-07 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=1.96 $X2=4.895 $Y2=2.135
r210 2 64 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.96 $X2=3.35 $Y2=2.125
r211 1 83 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=6.11
+ $Y=0.625 $X2=6.25 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%D 3 5 6 9 11 13 14 16 17 18 19 26
c59 9 0 8.69299e-20 $X=4.11 $Y=2.46
r60 26 28 19.042 $w=4.05e-07 $l=1.6e-07 $layer=POLY_cond $X=4.585 $Y=1.572
+ $X2=4.745 $Y2=1.572
r61 24 26 51.1753 $w=4.05e-07 $l=4.3e-07 $layer=POLY_cond $X=4.155 $Y=1.572
+ $X2=4.585 $Y2=1.572
r62 23 24 5.35556 $w=4.05e-07 $l=4.5e-08 $layer=POLY_cond $X=4.11 $Y=1.572
+ $X2=4.155 $Y2=1.572
r63 18 19 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.635
+ $X2=5.04 $Y2=1.635
r64 18 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.585
+ $Y=1.635 $X2=4.585 $Y2=1.635
r65 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.635
+ $X2=4.56 $Y2=1.635
r66 14 28 26.1659 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=4.745 $Y=1.345
+ $X2=4.745 $Y2=1.572
r67 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.745 $Y=1.345
+ $X2=4.745 $Y2=0.945
r68 11 24 26.1659 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=4.155 $Y=1.345
+ $X2=4.155 $Y2=1.572
r69 11 13 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.155 $Y=1.345
+ $X2=4.155 $Y2=0.945
r70 7 23 21.7585 $w=1.8e-07 $l=2.28e-07 $layer=POLY_cond $X=4.11 $Y=1.8 $X2=4.11
+ $Y2=1.572
r71 7 9 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.11 $Y=1.8 $X2=4.11
+ $Y2=2.46
r72 5 23 30.7588 $w=4.05e-07 $l=1.92819e-07 $layer=POLY_cond $X=4.02 $Y=1.725
+ $X2=4.11 $Y2=1.572
r73 5 6 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.02 $Y=1.725
+ $X2=3.665 $Y2=1.725
r74 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.575 $Y=1.8
+ $X2=3.665 $Y2=1.725
r75 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.575 $Y=1.8 $X2=3.575
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%C 3 7 8 11 13 15 17 24 25 26 28 29 32 33 34
c85 34 0 1.18606e-19 $X=3.08 $Y=1.35
c86 32 0 1.71934e-19 $X=3.08 $Y=1.515
c87 17 0 1.36857e-19 $X=5.12 $Y=2.46
c88 15 0 1.1549e-19 $X=5.12 $Y=1.825
r89 32 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.515
+ $X2=3.08 $Y2=1.68
r90 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.515
+ $X2=3.08 $Y2=1.35
r91 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.515 $X2=3.08 $Y2=1.515
r92 29 33 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.08 $Y=1.665
+ $X2=3.08 $Y2=1.515
r93 27 28 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=5.155 $Y=1.34
+ $X2=5.155 $Y2=1.49
r94 26 28 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.135 $Y=1.735
+ $X2=5.135 $Y2=1.49
r95 24 27 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.175 $Y=0.945
+ $X2=5.175 $Y2=1.34
r96 21 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.175 $Y=0.255
+ $X2=5.175 $Y2=0.945
r97 15 26 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.12 $Y=1.825 $X2=5.12
+ $Y2=1.735
r98 15 17 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.12 $Y=1.825
+ $X2=5.12 $Y2=2.46
r99 14 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.755 $Y=0.18
+ $X2=3.68 $Y2=0.18
r100 13 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.1 $Y=0.18
+ $X2=5.175 $Y2=0.255
r101 13 14 689.67 $w=1.5e-07 $l=1.345e-06 $layer=POLY_cond $X=5.1 $Y=0.18
+ $X2=3.755 $Y2=0.18
r102 9 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.68 $Y=0.255
+ $X2=3.68 $Y2=0.18
r103 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.68 $Y=0.255
+ $X2=3.68 $Y2=0.945
r104 7 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.605 $Y=0.18
+ $X2=3.68 $Y2=0.18
r105 7 8 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.605 $Y=0.18
+ $X2=3.245 $Y2=0.18
r106 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.17 $Y=0.255
+ $X2=3.245 $Y2=0.18
r107 5 34 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=3.17 $Y=0.255
+ $X2=3.17 $Y2=1.35
r108 3 35 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=3.125 $Y=2.46
+ $X2=3.125 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%A_27_368# 1 2 9 13 17 21 23 29 30 33 34 35
+ 37 38 40 41 42 50 55
c133 21 0 1.67323e-19 $X=6.49 $Y=2.46
c134 13 0 5.7483e-20 $X=6.035 $Y=0.945
r135 55 56 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.465 $Y=1.635
+ $X2=6.49 $Y2=1.635
r136 52 53 0.737003 $w=3.27e-07 $l=5e-09 $layer=POLY_cond $X=6.035 $Y=1.635
+ $X2=6.04 $Y2=1.635
r137 48 55 7.37003 $w=3.27e-07 $l=5e-08 $layer=POLY_cond $X=6.415 $Y=1.635
+ $X2=6.465 $Y2=1.635
r138 48 53 55.2752 $w=3.27e-07 $l=3.75e-07 $layer=POLY_cond $X=6.415 $Y=1.635
+ $X2=6.04 $Y2=1.635
r139 47 50 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.415 $Y=1.635
+ $X2=6.59 $Y2=1.635
r140 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.635 $X2=6.415 $Y2=1.635
r141 42 44 7.04271 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.265 $Y=2.475
+ $X2=0.265 $Y2=2.695
r142 40 41 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=1.82
r143 38 41 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.17 $Y=1.02 $X2=0.17
+ $Y2=1.82
r144 36 37 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=7.435 $Y=1.3
+ $X2=7.435 $Y2=2.39
r145 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.35 $Y=1.215
+ $X2=7.435 $Y2=1.3
r146 34 35 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.35 $Y=1.215
+ $X2=6.675 $Y2=1.215
r147 33 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.59 $Y=1.47
+ $X2=6.59 $Y2=1.635
r148 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.59 $Y=1.3
+ $X2=6.675 $Y2=1.215
r149 32 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.59 $Y=1.3
+ $X2=6.59 $Y2=1.47
r150 31 42 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.475
+ $X2=0.265 $Y2=2.475
r151 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.35 $Y=2.475
+ $X2=7.435 $Y2=2.39
r152 30 31 450.487 $w=1.68e-07 $l=6.905e-06 $layer=LI1_cond $X=7.35 $Y=2.475
+ $X2=0.445 $Y2=2.475
r153 29 42 2.72105 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.265 $Y2=2.475
r154 28 40 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=1.985
r155 28 29 12.4848 $w=3.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=2.39
r156 23 38 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.245 $Y=0.86
+ $X2=0.245 $Y2=1.02
r157 23 25 4.38438 $w=3.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.245 $Y=0.86
+ $X2=0.245 $Y2=0.745
r158 19 56 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.49 $Y=1.8
+ $X2=6.49 $Y2=1.635
r159 19 21 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.49 $Y=1.8
+ $X2=6.49 $Y2=2.46
r160 15 55 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.47
+ $X2=6.465 $Y2=1.635
r161 15 17 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.465 $Y=1.47
+ $X2=6.465 $Y2=0.945
r162 11 52 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.035 $Y=1.47
+ $X2=6.035 $Y2=1.635
r163 11 13 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.035 $Y=1.47
+ $X2=6.035 $Y2=0.945
r164 7 53 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.8
+ $X2=6.04 $Y2=1.635
r165 7 9 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.04 $Y=1.8 $X2=6.04
+ $Y2=2.46
r166 2 44 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.695
r167 2 40 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r168 1 25 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.47 $X2=0.32 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%B 1 3 8 9 10 13 18 20 27
c64 8 0 2.3468e-20 $X=5.605 $Y=0.945
r65 25 27 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=7.015 $Y=1.635
+ $X2=7.115 $Y2=1.635
r66 22 25 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.94 $Y=1.635
+ $X2=7.015 $Y2=1.635
r67 20 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.015
+ $Y=1.635 $X2=7.015 $Y2=1.635
r68 16 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.47
+ $X2=7.115 $Y2=1.635
r69 16 18 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=7.115 $Y=1.47
+ $X2=7.115 $Y2=0.945
r70 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.115 $Y=0.255
+ $X2=7.115 $Y2=0.945
r71 11 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.8
+ $X2=6.94 $Y2=1.635
r72 11 13 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.94 $Y=1.8 $X2=6.94
+ $Y2=2.46
r73 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.04 $Y=0.18
+ $X2=7.115 $Y2=0.255
r74 9 10 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=7.04 $Y=0.18
+ $X2=5.68 $Y2=0.18
r75 8 19 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.605 $Y=0.945
+ $X2=5.605 $Y2=1.395
r76 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=0.255
+ $X2=5.68 $Y2=0.18
r77 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.605 $Y=0.255
+ $X2=5.605 $Y2=0.945
r78 1 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.59 $Y=1.485 $X2=5.59
+ $Y2=1.395
r79 1 3 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=5.59 $Y=1.485
+ $X2=5.59 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%VPWR 1 2 3 4 5 6 7 26 30 32 36 40 44 48 51
+ 52 54 55 57 58 59 61 79 84 87 90 95 96
r94 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 93 95 10.5953 $w=5.93e-07 $l=5.15e-07 $layer=LI1_cond $X=7.34 $Y=2.815
+ $X2=7.34 $Y2=3.33
r96 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 82 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r101 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 79 95 8.24118 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=7 $Y=3.33 $X2=7.34
+ $Y2=3.33
r103 79 81 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=7 $Y=3.33 $X2=6.96
+ $Y2=3.33
r104 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r105 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r107 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 69 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 66 90 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=2.807 $Y2=3.33
r114 66 68 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 65 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r118 62 84 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.837 $Y2=3.33
r119 62 64 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 61 87 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.775 $Y2=3.33
r121 61 64 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 59 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 59 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 57 77 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.1 $Y=3.33 $X2=6
+ $Y2=3.33
r125 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.1 $Y=3.33
+ $X2=6.265 $Y2=3.33
r126 56 81 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.265 $Y2=3.33
r128 54 74 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.04 $Y2=3.33
r129 54 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.355 $Y2=3.33
r130 53 77 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.53 $Y=3.33 $X2=6
+ $Y2=3.33
r131 53 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.355 $Y2=3.33
r132 51 68 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=3.33
+ $X2=3.6 $Y2=3.33
r133 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.72 $Y=3.33
+ $X2=3.885 $Y2=3.33
r134 50 71 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.05 $Y=3.33 $X2=4.08
+ $Y2=3.33
r135 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=3.33
+ $X2=3.885 $Y2=3.33
r136 46 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.265 $Y=3.245
+ $X2=6.265 $Y2=3.33
r137 46 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.265 $Y=3.245
+ $X2=6.265 $Y2=2.815
r138 42 55 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.355 $Y=3.245
+ $X2=5.355 $Y2=3.33
r139 42 44 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.355 $Y=3.245
+ $X2=5.355 $Y2=2.815
r140 38 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=3.245
+ $X2=3.885 $Y2=3.33
r141 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.885 $Y=3.245
+ $X2=3.885 $Y2=2.815
r142 34 90 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.807 $Y=3.245
+ $X2=2.807 $Y2=3.33
r143 34 36 14.3638 $w=3.43e-07 $l=4.3e-07 $layer=LI1_cond $X=2.807 $Y=3.245
+ $X2=2.807 $Y2=2.815
r144 33 87 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.775 $Y2=3.33
r145 32 90 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.807 $Y2=3.33
r146 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=1.955 $Y2=3.33
r147 28 87 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r148 28 30 13.7653 $w=3.58e-07 $l=4.3e-07 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=2.815
r149 24 84 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.837 $Y=3.245
+ $X2=0.837 $Y2=3.33
r150 24 26 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=0.837 $Y=3.245
+ $X2=0.837 $Y2=2.815
r151 7 93 600 $w=1.7e-07 $l=9.71995e-07 $layer=licon1_PDIFF $count=1 $X=7.03
+ $Y=1.96 $X2=7.28 $Y2=2.815
r152 6 48 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.13
+ $Y=1.96 $X2=6.265 $Y2=2.815
r153 5 44 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.21
+ $Y=1.96 $X2=5.355 $Y2=2.815
r154 4 40 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=1.96 $X2=3.885 $Y2=2.815
r155 3 36 600 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.84 $X2=2.805 $Y2=2.815
r156 2 30 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.84 $X2=1.775 $Y2=2.815
r157 1 26 600 $w=1.7e-07 $l=1.0884e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.835 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%X 1 2 3 4 15 17 21 23 24 25 26 27 36 42 44
c62 17 0 1.18606e-19 $X=2.21 $Y=1.065
r63 34 42 1.64635 $w=3.83e-07 $l=5.5e-08 $layer=LI1_cond $X=1.277 $Y=0.98
+ $X2=1.277 $Y2=0.925
r64 27 44 4.75094 $w=2.3e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.2
+ $Y2=1.82
r65 26 44 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.82
r66 25 26 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r67 25 43 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.15
r68 24 34 3.0793 $w=3.07e-07 $l=8.5e-08 $layer=LI1_cond $X=1.277 $Y=1.065
+ $X2=1.277 $Y2=0.98
r69 24 43 3.0793 $w=3.07e-07 $l=1.17346e-07 $layer=LI1_cond $X=1.277 $Y=1.065
+ $X2=1.2 $Y2=1.15
r70 24 42 0.449004 $w=3.83e-07 $l=1.5e-08 $layer=LI1_cond $X=1.277 $Y=0.91
+ $X2=1.277 $Y2=0.925
r71 23 24 10.6264 $w=3.83e-07 $l=3.55e-07 $layer=LI1_cond $X=1.277 $Y=0.555
+ $X2=1.277 $Y2=0.91
r72 23 36 1.19734 $w=3.83e-07 $l=4e-08 $layer=LI1_cond $X=1.277 $Y=0.555
+ $X2=1.277 $Y2=0.515
r73 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.375 $Y=0.98
+ $X2=2.375 $Y2=0.515
r74 18 24 3.54158 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.47 $Y=1.065
+ $X2=1.277 $Y2=1.065
r75 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.21 $Y=1.065
+ $X2=2.375 $Y2=0.98
r76 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.21 $Y=1.065
+ $X2=1.47 $Y2=1.065
r77 13 27 2.73179 $w=4e-07 $l=1.15e-07 $layer=LI1_cond $X=1.315 $Y=2.02 $X2=1.2
+ $Y2=2.02
r78 13 15 26.6502 $w=3.98e-07 $l=9.25e-07 $layer=LI1_cond $X=1.315 $Y=2.02
+ $X2=2.24 $Y2=2.02
r79 4 15 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=2.105
+ $Y=1.84 $X2=2.24 $Y2=2.02
r80 3 27 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.84 $X2=1.31 $Y2=2.02
r81 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.235
+ $Y=0.37 $X2=2.375 $Y2=0.515
r82 1 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.165
+ $Y=0.37 $X2=1.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%VGND 1 2 3 4 15 17 21 25 29 32 33 34 36 45
+ 54 55 58 61 64
r83 64 65 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r84 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r85 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r86 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 55 65 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=4.56
+ $Y2=0
r88 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r89 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=4.45
+ $Y2=0
r90 52 54 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=4.615 $Y=0
+ $X2=7.44 $Y2=0
r91 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r92 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r93 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r94 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r95 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.45
+ $Y2=0
r96 45 50 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.08
+ $Y2=0
r97 44 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r98 44 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r99 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r100 41 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.835
+ $Y2=0
r101 41 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.64
+ $Y2=0
r102 39 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r103 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r104 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r105 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r106 34 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r107 34 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r108 32 43 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.64
+ $Y2=0
r109 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.875
+ $Y2=0
r110 31 47 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.12
+ $Y2=0
r111 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.875
+ $Y2=0
r112 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r113 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.535
r114 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r115 23 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.515
r116 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0
r117 19 21 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0.645
r118 18 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r119 17 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.835
+ $Y2=0
r120 17 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.67 $Y=0
+ $X2=0.915 $Y2=0
r121 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r122 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.595
r123 4 29 182 $w=1.7e-07 $l=2.61151e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.625 $X2=4.45 $Y2=0.535
r124 3 25 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.37 $X2=2.875 $Y2=0.515
r125 2 21 182 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.37 $X2=1.835 $Y2=0.645
r126 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.61
+ $Y=0.47 $X2=0.75 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%A_664_125# 1 2 3 12 14 15 19 20 21 24
c59 14 0 1.1549e-19 $X=5.305 $Y=1.215
r60 22 24 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.33 $Y=0.425
+ $X2=7.33 $Y2=0.78
r61 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.165 $Y=0.34
+ $X2=7.33 $Y2=0.425
r62 20 21 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=7.165 $Y=0.34
+ $X2=5.475 $Y2=0.34
r63 17 19 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.39 $Y=1.13
+ $X2=5.39 $Y2=0.77
r64 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.39 $Y=0.425
+ $X2=5.475 $Y2=0.34
r65 16 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.39 $Y=0.425
+ $X2=5.39 $Y2=0.77
r66 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.305 $Y=1.215
+ $X2=5.39 $Y2=1.13
r67 14 15 109.278 $w=1.68e-07 $l=1.675e-06 $layer=LI1_cond $X=5.305 $Y=1.215
+ $X2=3.63 $Y2=1.215
r68 10 15 22.9197 $w=8.4e-08 $l=2.03101e-07 $layer=LI1_cond $X=3.465 $Y=1.13
+ $X2=3.63 $Y2=1.215
r69 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.465 $Y=1.13
+ $X2=3.465 $Y2=0.89
r70 3 24 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=7.19
+ $Y=0.625 $X2=7.33 $Y2=0.78
r71 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.25
+ $Y=0.625 $X2=5.39 $Y2=0.77
r72 1 12 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.625 $X2=3.465 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%A_751_125# 1 2 7 12 14
r24 14 16 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.96 $Y=0.78
+ $X2=4.96 $Y2=0.875
r25 10 12 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.915 $Y=0.795
+ $X2=4.105 $Y2=0.795
r26 7 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0.875
+ $X2=4.96 $Y2=0.875
r27 7 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.795 $Y=0.875
+ $X2=4.105 $Y2=0.875
r28 2 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.625 $X2=4.96 $Y2=0.78
r29 1 10 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=3.755
+ $Y=0.625 $X2=3.915 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_4%A_1136_125# 1 2 7 9 14
c20 9 0 5.7483e-20 $X=5.78 $Y=0.68
c21 7 0 2.3468e-20 $X=6.625 $Y=0.68
r22 14 17 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.79 $Y=0.68 $X2=6.79
+ $Y2=0.77
r23 9 12 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=5.78 $Y=0.68 $X2=5.78
+ $Y2=0.78
r24 8 9 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.905 $Y=0.68 $X2=5.78
+ $Y2=0.68
r25 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=0.68
+ $X2=6.79 $Y2=0.68
r26 7 8 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.625 $Y=0.68
+ $X2=5.905 $Y2=0.68
r27 2 17 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=6.54
+ $Y=0.625 $X2=6.79 $Y2=0.77
r28 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.68
+ $Y=0.625 $X2=5.82 $Y2=0.78
.ends


* File: sky130_fd_sc_ms__fa_1.pex.spice
* Created: Fri Aug 28 17:34:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FA_1%A_69_260# 1 2 9 13 16 17 18 19 21 25 28 29 31
+ 36 41
c108 31 0 1.67865e-19 $X=1.14 $Y=1.795
c109 25 0 7.83064e-20 $X=2.245 $Y=2.59
r110 41 43 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=1.91
+ $X2=2.245 $Y2=2.035
r111 36 38 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.105 $Y=0.55
+ $X2=2.105 $Y2=0.665
r112 31 33 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.14 $Y=1.795
+ $X2=1.14 $Y2=2.035
r113 29 46 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.465
+ $X2=0.51 $Y2=1.63
r114 29 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.465
+ $X2=0.51 $Y2=1.3
r115 28 30 17.3534 $w=2.32e-07 $l=3.3e-07 $layer=LI1_cond $X=0.565 $Y=1.465
+ $X2=0.565 $Y2=1.795
r116 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.465 $X2=0.51 $Y2=1.465
r117 23 43 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=2.12
+ $X2=2.245 $Y2=2.035
r118 23 25 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.245 $Y=2.12
+ $X2=2.245 $Y2=2.59
r119 22 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.035
+ $X2=1.14 $Y2=2.035
r120 21 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=2.035
+ $X2=2.245 $Y2=2.035
r121 21 22 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.08 $Y=2.035
+ $X2=1.225 $Y2=2.035
r122 20 30 2.55969 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.705 $Y=1.795
+ $X2=0.565 $Y2=1.795
r123 19 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.795
+ $X2=1.14 $Y2=1.795
r124 19 20 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.055 $Y=1.795
+ $X2=0.705 $Y2=1.795
r125 17 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0.665
+ $X2=2.105 $Y2=0.665
r126 17 18 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.94 $Y=0.665
+ $X2=0.705 $Y2=0.665
r127 16 28 9.57122 $w=2.32e-07 $l=1.90526e-07 $layer=LI1_cond $X=0.62 $Y=1.3
+ $X2=0.565 $Y2=1.465
r128 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=0.75
+ $X2=0.705 $Y2=0.665
r129 15 16 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.62 $Y=0.75
+ $X2=0.62 $Y2=1.3
r130 13 45 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.3
r131 9 46 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=2.4
+ $X2=0.495 $Y2=1.63
r132 2 41 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.735 $X2=2.245 $Y2=1.91
r133 2 25 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.735 $X2=2.245 $Y2=2.59
r134 1 36 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.375 $X2=2.105 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%A 3 7 11 15 18 22 25 27 29 31 32 36 37 39 41 44
+ 45 48 49 51 55 58 64 67 69 71
c231 67 0 4.91364e-20 $X=4.545 $Y=1.29
c232 51 0 1.97438e-19 $X=4.545 $Y=1.012
c233 44 0 2.98399e-20 $X=5.895 $Y=1.32
c234 37 0 2.45682e-20 $X=3.465 $Y=1.29
c235 32 0 8.33772e-20 $X=3.3 $Y=1.005
c236 25 0 6.57094e-20 $X=6.055 $Y=2.235
r237 67 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.29
+ $X2=4.545 $Y2=1.455
r238 67 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.29
+ $X2=4.545 $Y2=1.125
r239 58 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.545
+ $Y=1.29 $X2=4.545 $Y2=1.29
r240 56 74 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.41
+ $X2=6.045 $Y2=1.575
r241 56 71 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=6.045 $Y=1.41
+ $X2=6.045 $Y2=1.185
r242 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.045
+ $Y=1.41 $X2=6.045 $Y2=1.41
r243 50 58 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.545 $Y=1.105
+ $X2=4.545 $Y2=1.29
r244 50 51 0.89609 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=4.545 $Y=1.105
+ $X2=4.545 $Y2=1.012
r245 48 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.385
+ $X2=1.05 $Y2=1.55
r246 48 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.385
+ $X2=1.05 $Y2=1.22
r247 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.385 $X2=1.05 $Y2=1.385
r248 45 47 18.3968 $w=2.52e-07 $l=3.8e-07 $layer=LI1_cond $X=1.05 $Y=1.005
+ $X2=1.05 $Y2=1.385
r249 44 55 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=5.895 $Y=1.447
+ $X2=6.045 $Y2=1.447
r250 43 44 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.895 $Y=1.105
+ $X2=5.895 $Y2=1.32
r251 42 51 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=4.71 $Y=1.02
+ $X2=4.545 $Y2=1.012
r252 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.81 $Y=1.02
+ $X2=5.895 $Y2=1.105
r253 41 42 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=5.81 $Y=1.02
+ $X2=4.71 $Y2=1.02
r254 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.63 $Y=1.005
+ $X2=3.465 $Y2=1.005
r255 39 51 8.61065 $w=1.7e-07 $l=1.68464e-07 $layer=LI1_cond $X=4.38 $Y=1.005
+ $X2=4.545 $Y2=1.012
r256 39 40 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.38 $Y=1.005
+ $X2=3.63 $Y2=1.005
r257 37 65 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.465 $Y=1.29
+ $X2=3.465 $Y2=1.455
r258 37 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.465 $Y=1.29
+ $X2=3.465 $Y2=1.125
r259 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.29 $X2=3.465 $Y2=1.29
r260 34 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=1.09
+ $X2=3.465 $Y2=1.005
r261 34 36 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.465 $Y=1.09
+ $X2=3.465 $Y2=1.29
r262 33 45 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=1.005
+ $X2=1.05 $Y2=1.005
r263 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=1.005
+ $X2=3.465 $Y2=1.005
r264 32 33 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=3.3 $Y=1.005
+ $X2=1.215 $Y2=1.005
r265 29 31 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=6.485 $Y=1.11
+ $X2=6.485 $Y2=0.695
r266 28 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.185
+ $X2=6.045 $Y2=1.185
r267 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.41 $Y=1.185
+ $X2=6.485 $Y2=1.11
r268 27 28 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.41 $Y=1.185
+ $X2=6.21 $Y2=1.185
r269 25 74 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.055 $Y=2.235
+ $X2=6.055 $Y2=1.575
r270 22 69 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.605 $Y=0.695
+ $X2=4.605 $Y2=1.125
r271 18 70 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=4.505 $Y=2.235
+ $X2=4.505 $Y2=1.455
r272 15 64 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.53 $Y=0.695
+ $X2=3.53 $Y2=1.125
r273 11 65 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=3.54 $Y=2.235
+ $X2=3.54 $Y2=1.455
r274 7 61 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=1.11 $Y=0.695
+ $X2=1.11 $Y2=1.22
r275 3 62 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.01 $Y=2.34
+ $X2=1.01 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%CIN 3 7 11 15 19 23 25 27 28 30 31 32 33 36 39
+ 42 45 50 51
c180 32 0 4.91364e-20 $X=4.895 $Y=1.665
c181 31 0 1.02197e-19 $X=1.825 $Y=1.665
c182 30 0 2.45682e-20 $X=3.935 $Y=1.665
c183 25 0 2.98399e-20 $X=5.155 $Y=1.425
c184 3 0 8.59909e-20 $X=1.89 $Y=0.695
r185 51 60 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=4.017 $Y=1.41
+ $X2=4.017 $Y2=1.665
r186 50 53 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.005 $Y=1.41
+ $X2=4.005 $Y2=1.575
r187 50 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.005 $Y=1.41
+ $X2=4.005 $Y2=1.245
r188 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.005
+ $Y=1.41 $X2=4.005 $Y2=1.41
r189 45 48 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.41
+ $X2=1.95 $Y2=1.575
r190 45 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.41
+ $X2=1.95 $Y2=1.245
r191 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.41 $X2=1.95 $Y2=1.41
r192 42 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r193 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r194 36 46 8.235 $w=4e-07 $l=2.7e-07 $layer=LI1_cond $X=1.68 $Y=1.52 $X2=1.95
+ $Y2=1.52
r195 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.665
r196 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r197 32 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r198 32 33 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=4.225 $Y2=1.665
r199 31 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=1.665
+ $X2=1.68 $Y2=1.665
r200 30 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r201 30 31 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=1.825 $Y2=1.665
r202 28 56 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.575
r203 28 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.245
r204 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.475
+ $Y=1.41 $X2=5.475 $Y2=1.41
r205 25 40 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.04 $Y=1.425
+ $X2=5.04 $Y2=1.665
r206 25 27 12.2927 $w=2.98e-07 $l=3.2e-07 $layer=LI1_cond $X=5.155 $Y=1.425
+ $X2=5.475 $Y2=1.425
r207 23 56 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.46 $Y=2.235
+ $X2=5.46 $Y2=1.575
r208 19 55 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.425 $Y=0.695
+ $X2=5.425 $Y2=1.245
r209 15 53 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.045 $Y=2.235
+ $X2=4.045 $Y2=1.575
r210 11 52 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.96 $Y=0.695
+ $X2=3.96 $Y2=1.245
r211 7 48 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.02 $Y=2.235
+ $X2=2.02 $Y2=1.575
r212 3 47 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.89 $Y=0.695
+ $X2=1.89 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%A_465_249# 1 2 9 13 17 19 21 22 23 24 27 28 29
+ 32 34 37 39 40 41 44 48 49 52
c187 49 0 1.99239e-19 $X=2.49 $Y=1.41
c188 48 0 1.02197e-19 $X=2.49 $Y=1.41
c189 39 0 1.09525e-19 $X=6.465 $Y=1.745
c190 13 0 1.63156e-19 $X=2.47 $Y=2.235
r191 59 61 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.235 $Y=1.065
+ $X2=6.465 $Y2=1.065
r192 52 54 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.21 $Y=0.6 $X2=5.21
+ $Y2=0.68
r193 49 66 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.41
+ $X2=2.49 $Y2=1.575
r194 49 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.41
+ $X2=2.49 $Y2=1.245
r195 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.41 $X2=2.49 $Y2=1.41
r196 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.875
+ $Y=1.385 $X2=7.875 $Y2=1.385
r197 42 44 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.875 $Y=1.15
+ $X2=7.875 $Y2=1.385
r198 41 61 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=1.065
+ $X2=6.465 $Y2=1.065
r199 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.71 $Y=1.065
+ $X2=7.875 $Y2=1.15
r200 40 41 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=7.71 $Y=1.065
+ $X2=6.55 $Y2=1.065
r201 38 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.465 $Y=1.15
+ $X2=6.465 $Y2=1.065
r202 38 39 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.465 $Y=1.15
+ $X2=6.465 $Y2=1.745
r203 37 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.98
+ $X2=6.235 $Y2=1.065
r204 36 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.235 $Y=0.765
+ $X2=6.235 $Y2=0.98
r205 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.38 $Y=1.83
+ $X2=6.465 $Y2=1.745
r206 34 35 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.38 $Y=1.83
+ $X2=5.495 $Y2=1.83
r207 33 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=0.68
+ $X2=5.21 $Y2=0.68
r208 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.15 $Y=0.68
+ $X2=6.235 $Y2=0.765
r209 32 33 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.15 $Y=0.68
+ $X2=5.375 $Y2=0.68
r210 28 35 8.77544 $w=2.85e-07 $l=3.87161e-07 $layer=LI1_cond $X=5.197 $Y=2.035
+ $X2=5.495 $Y2=1.83
r211 28 29 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=5.07 $Y=2.035 $X2=3.2
+ $Y2=2.035
r212 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=1.95
+ $X2=3.2 $Y2=2.035
r213 26 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.115 $Y=1.795
+ $X2=3.115 $Y2=1.95
r214 25 48 11.4375 $w=3.2e-07 $l=3.92301e-07 $layer=LI1_cond $X=2.75 $Y=1.71
+ $X2=2.537 $Y2=1.41
r215 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.03 $Y=1.71
+ $X2=3.115 $Y2=1.795
r216 24 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.03 $Y=1.71
+ $X2=2.75 $Y2=1.71
r217 22 45 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.055 $Y=1.385
+ $X2=7.875 $Y2=1.385
r218 22 23 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.055 $Y=1.385
+ $X2=8.145 $Y2=1.385
r219 19 23 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=8.16 $Y=1.22
+ $X2=8.145 $Y2=1.385
r220 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.16 $Y=1.22
+ $X2=8.16 $Y2=0.74
r221 15 23 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.145 $Y=1.55
+ $X2=8.145 $Y2=1.385
r222 15 17 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=8.145 $Y=1.55
+ $X2=8.145 $Y2=2.4
r223 13 66 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.47 $Y=2.235
+ $X2=2.47 $Y2=1.575
r224 9 65 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.43 $Y=0.695
+ $X2=2.43 $Y2=1.245
r225 2 28 300 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_PDIFF $count=2 $X=5.1
+ $Y=1.735 $X2=5.235 $Y2=2.035
r226 1 52 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.07
+ $Y=0.375 $X2=5.21 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%B 3 5 8 9 10 13 14 17 18 22 23 26 27 32 35 38
+ 39 40 41 42 48 49
c148 49 0 6.57094e-20 $X=7.305 $Y=1.485
c149 17 0 2.64346e-19 $X=2.955 $Y=2.235
c150 8 0 1.67865e-19 $X=1.515 $Y=2.445
c151 5 0 8.33772e-20 $X=1.515 $Y=1.805
r152 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.305
+ $Y=1.485 $X2=7.305 $Y2=1.485
r153 46 48 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.21 $Y=1.485
+ $X2=7.305 $Y2=1.485
r154 44 46 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=6.89 $Y=1.485
+ $X2=7.21 $Y2=1.485
r155 42 49 3.21335 $w=6.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.135 $Y=1.665
+ $X2=7.135 $Y2=1.485
r156 33 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.21 $Y=1.32
+ $X2=7.21 $Y2=1.485
r157 33 35 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=7.21 $Y=1.32
+ $X2=7.21 $Y2=0.695
r158 30 32 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=6.89 $Y=3.075
+ $X2=6.89 $Y2=2.31
r159 29 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.65
+ $X2=6.89 $Y2=1.485
r160 29 32 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.65
+ $X2=6.89 $Y2=2.31
r161 28 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.1 $Y=3.15 $X2=5.01
+ $Y2=3.15
r162 27 30 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.8 $Y=3.15
+ $X2=6.89 $Y2=3.075
r163 27 28 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=6.8 $Y=3.15 $X2=5.1
+ $Y2=3.15
r164 24 41 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.01 $Y=3.075
+ $X2=5.01 $Y2=3.15
r165 24 26 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=5.01 $Y=3.075
+ $X2=5.01 $Y2=2.235
r166 23 40 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.01 $Y=1.18 $X2=5.01
+ $Y2=1.09
r167 23 26 410.089 $w=1.8e-07 $l=1.055e-06 $layer=POLY_cond $X=5.01 $Y=1.18
+ $X2=5.01 $Y2=2.235
r168 22 40 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.995 $Y=0.695
+ $X2=4.995 $Y2=1.09
r169 19 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.045 $Y=3.15
+ $X2=2.955 $Y2=3.15
r170 18 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.92 $Y=3.15 $X2=5.01
+ $Y2=3.15
r171 18 19 961.436 $w=1.5e-07 $l=1.875e-06 $layer=POLY_cond $X=4.92 $Y=3.15
+ $X2=3.045 $Y2=3.15
r172 15 39 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=3.075
+ $X2=2.955 $Y2=3.15
r173 15 17 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=2.955 $Y=3.075
+ $X2=2.955 $Y2=2.235
r174 14 38 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=1.18
+ $X2=2.955 $Y2=1.09
r175 14 17 410.089 $w=1.8e-07 $l=1.055e-06 $layer=POLY_cond $X=2.955 $Y=1.18
+ $X2=2.955 $Y2=2.235
r176 13 38 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.94 $Y=0.695
+ $X2=2.94 $Y2=1.09
r177 9 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.865 $Y=3.15
+ $X2=2.955 $Y2=3.15
r178 9 10 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=2.865 $Y=3.15
+ $X2=1.605 $Y2=3.15
r179 6 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.515 $Y=3.075
+ $X2=1.605 $Y2=3.15
r180 6 8 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=1.515 $Y=3.075
+ $X2=1.515 $Y2=2.445
r181 5 37 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.515 $Y=1.805
+ $X2=1.515 $Y2=1.715
r182 5 8 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=1.515 $Y=1.805
+ $X2=1.515 $Y2=2.445
r183 3 37 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.5 $Y=0.695
+ $X2=1.5 $Y2=1.715
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%SUM 1 2 9 11 15 16 17 28
r22 21 28 2.67531 $w=2.78e-07 $l=6.5e-08 $layer=LI1_cond $X=0.225 $Y=0.99
+ $X2=0.225 $Y2=0.925
r23 17 30 7.11633 $w=2.78e-07 $l=1.3e-07 $layer=LI1_cond $X=0.225 $Y=1 $X2=0.225
+ $Y2=1.13
r24 17 21 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=0.225 $Y=1 $X2=0.225
+ $Y2=0.99
r25 17 28 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=0.225 $Y=0.915
+ $X2=0.225 $Y2=0.925
r26 16 17 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=0.225 $Y=0.515
+ $X2=0.225 $Y2=0.915
r27 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.82 $X2=0.17
+ $Y2=1.13
r28 11 13 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.22 $Y=1.985
+ $X2=0.22 $Y2=2.815
r29 9 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.955
+ $X2=0.22 $Y2=1.82
r30 9 11 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=1.955 $X2=0.22
+ $Y2=1.985
r31 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r32 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
r33 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%VPWR 1 2 3 4 5 18 24 28 32 36 41 42 43 45 50 59
+ 66 73 74 77 80 83 86
c104 4 0 1.09525e-19 $X=6.145 $Y=1.735
r105 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r107 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 74 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r111 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=7.92 $Y2=3.33
r112 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=8.4 $Y2=3.33
r113 70 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 70 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 67 83 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.472 $Y2=3.33
r117 67 69 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 66 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.92 $Y2=3.33
r119 66 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r121 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r122 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r123 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=6
+ $Y2=3.33
r124 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 59 83 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=6.12 $Y=3.33
+ $X2=6.472 $Y2=3.33
r126 59 64 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.12 $Y=3.33 $X2=6
+ $Y2=3.33
r127 58 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 55 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.245 $Y2=3.33
r130 55 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=4.08 $Y2=3.33
r131 54 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 54 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r133 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 51 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r135 51 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 50 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=3.245 $Y2=3.33
r137 50 53 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 45 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 43 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 43 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r144 41 57 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=3.33
+ $X2=4.27 $Y2=3.33
r146 40 61 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.56 $Y2=3.33
r147 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.27 $Y2=3.33
r148 36 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.92 $Y=1.985
+ $X2=7.92 $Y2=2.815
r149 34 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r150 34 39 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.815
r151 30 83 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.472 $Y=3.245
+ $X2=6.472 $Y2=3.33
r152 30 32 10.9428 $w=7.03e-07 $l=6.45e-07 $layer=LI1_cond $X=6.472 $Y=3.245
+ $X2=6.472 $Y2=2.6
r153 26 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=3.245
+ $X2=4.27 $Y2=3.33
r154 26 28 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=4.27 $Y=3.245
+ $X2=4.27 $Y2=2.47
r155 22 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=3.245
+ $X2=3.245 $Y2=3.33
r156 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.245 $Y=3.245
+ $X2=3.245 $Y2=2.795
r157 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.72 $Y=2.135
+ $X2=0.72 $Y2=2.815
r158 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r159 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.815
r160 5 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.92 $Y2=2.815
r161 5 36 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.92 $Y2=1.985
r162 4 32 300 $w=1.7e-07 $l=1.09257e-06 $layer=licon1_PDIFF $count=2 $X=6.145
+ $Y=1.735 $X2=6.66 $Y2=2.6
r163 3 28 600 $w=1.7e-07 $l=7.99656e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.735 $X2=4.27 $Y2=2.47
r164 2 24 600 $w=1.7e-07 $l=1.15568e-06 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.735 $X2=3.245 $Y2=2.795
r165 1 21 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.815
r166 1 18 300 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%A_512_347# 1 2 9 13 15 18
c34 13 0 3.49195e-19 $X=2.695 $Y=2.59
c35 9 0 1.99239e-19 $X=2.695 $Y=2.13
r36 18 21 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.765 $Y=2.375
+ $X2=3.765 $Y2=2.455
r37 16 17 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.86 $Y=2.375
+ $X2=2.735 $Y2=2.375
r38 15 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=2.375
+ $X2=3.765 $Y2=2.375
r39 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.6 $Y=2.375
+ $X2=2.86 $Y2=2.375
r40 11 17 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=2.375
r41 11 13 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=2.59
r42 7 17 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.29
+ $X2=2.735 $Y2=2.375
r43 7 9 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.735 $Y=2.29
+ $X2=2.735 $Y2=2.13
r44 2 21 600 $w=1.7e-07 $l=7.84602e-07 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=1.735 $X2=3.765 $Y2=2.455
r45 1 13 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=1.735 $X2=2.695 $Y2=2.59
r46 1 9 600 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=1.735 $X2=2.695 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%A_1110_347# 1 2 7 9 11 13 15
r28 13 20 3.10428 $w=3.2e-07 $l=1.5548e-07 $layer=LI1_cond $X=7.16 $Y=2.255
+ $X2=7.155 $Y2=2.102
r29 13 15 14.7657 $w=3.18e-07 $l=4.1e-07 $layer=LI1_cond $X=7.16 $Y=2.255
+ $X2=7.16 $Y2=2.665
r30 12 18 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.95 $Y=2.17
+ $X2=5.807 $Y2=2.17
r31 11 20 4.57783 $w=1.7e-07 $l=1.96074e-07 $layer=LI1_cond $X=6.99 $Y=2.17
+ $X2=7.155 $Y2=2.102
r32 11 12 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=6.99 $Y=2.17
+ $X2=5.95 $Y2=2.17
r33 7 18 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.807 $Y=2.255
+ $X2=5.807 $Y2=2.17
r34 7 9 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=5.807 $Y=2.255
+ $X2=5.807 $Y2=2.59
r35 2 20 600 $w=1.7e-07 $l=3.82623e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=1.81 $X2=7.155 $Y2=2.115
r36 2 15 600 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=1.81 $X2=7.155 $Y2=2.665
r37 1 18 600 $w=1.7e-07 $l=5.57696e-07 $layer=licon1_PDIFF $count=1 $X=5.55
+ $Y=1.735 $X2=5.83 $Y2=2.17
r38 1 9 600 $w=1.7e-07 $l=9.85102e-07 $layer=licon1_PDIFF $count=1 $X=5.55
+ $Y=1.735 $X2=5.83 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%COUT 1 2 7 8 9 10 11 12 13 29
r17 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=8.375 $Y=0.965
+ $X2=8.375 $Y2=0.925
r18 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=8.412 $Y=2.405
+ $X2=8.412 $Y2=2.775
r19 11 12 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=8.412 $Y=1.985
+ $X2=8.412 $Y2=2.405
r20 10 11 14.462 $w=2.53e-07 $l=3.2e-07 $layer=LI1_cond $X=8.412 $Y=1.665
+ $X2=8.412 $Y2=1.985
r21 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=8.412 $Y=1.295
+ $X2=8.412 $Y2=1.665
r22 9 45 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.412 $Y=1.295
+ $X2=8.412 $Y2=1.13
r23 8 45 5.6192 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=8.375 $Y=0.987
+ $X2=8.375 $Y2=1.13
r24 8 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=8.375 $Y=0.987
+ $X2=8.375 $Y2=0.965
r25 8 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=8.375 $Y=0.902
+ $X2=8.375 $Y2=0.925
r26 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=8.375 $Y=0.515
+ $X2=8.375 $Y2=0.902
r27 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.235
+ $Y=1.84 $X2=8.37 $Y2=2.815
r28 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.235
+ $Y=1.84 $X2=8.37 $Y2=1.985
r29 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.235
+ $Y=0.37 $X2=8.375 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%VGND 1 2 3 4 5 16 20 24 28 30 32 37 42 50 57 58
+ 69 75 78 81
r108 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r109 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r110 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r111 70 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r112 69 72 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.235 $Y=0
+ $X2=3.235 $Y2=0.325
r113 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r114 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r115 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r116 55 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=7.905
+ $Y2=0
r117 55 57 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=8.4
+ $Y2=0
r118 54 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r119 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r120 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 51 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=6.955
+ $Y2=0
r122 51 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=7.44
+ $Y2=0
r123 50 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.905
+ $Y2=0
r124 50 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.44
+ $Y2=0
r125 49 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r126 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r127 46 49 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r128 45 48 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r129 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r130 43 75 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=4.317 $Y2=0
r131 43 45 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.56
+ $Y2=0
r132 42 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=6.955
+ $Y2=0
r133 42 48 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=6.48
+ $Y2=0
r134 41 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r135 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r136 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r137 38 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r138 37 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.235
+ $Y2=0
r139 37 40 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=3.07 $Y=0 $X2=1.2
+ $Y2=0
r140 35 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r141 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r142 32 65 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=0.802 $Y=0
+ $X2=0.802 $Y2=0.325
r143 32 38 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.802 $Y=0 $X2=0.98
+ $Y2=0
r144 32 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r145 32 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r146 30 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r147 30 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r148 26 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0
r149 26 28 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0.605
r150 22 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.085
+ $X2=6.955 $Y2=0
r151 22 24 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=6.955 $Y=0.085
+ $X2=6.955 $Y2=0.305
r152 18 75 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.317 $Y=0.085
+ $X2=4.317 $Y2=0
r153 18 20 11.5831 $w=4.73e-07 $l=4.6e-07 $layer=LI1_cond $X=4.317 $Y=0.085
+ $X2=4.317 $Y2=0.545
r154 17 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.235
+ $Y2=0
r155 16 75 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=4.317
+ $Y2=0
r156 16 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.4
+ $Y2=0
r157 5 28 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=7.82
+ $Y=0.37 $X2=7.945 $Y2=0.605
r158 4 24 182 $w=1.7e-07 $l=3.88426e-07 $layer=licon1_NDIFF $count=1 $X=6.56
+ $Y=0.375 $X2=6.915 $Y2=0.305
r159 3 20 182 $w=1.7e-07 $l=3.54965e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.375 $X2=4.315 $Y2=0.545
r160 2 72 182 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.375 $X2=3.235 $Y2=0.325
r161 1 65 182 $w=1.7e-07 $l=2.51496e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.8 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%A_501_75# 1 2 7 12 14
c26 12 0 8.59909e-20 $X=2.89 $Y=0.585
r27 14 16 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.745 $Y=0.585
+ $X2=3.745 $Y2=0.665
r28 10 12 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.685 $Y=0.585
+ $X2=2.89 $Y2=0.585
r29 7 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=0.665
+ $X2=3.745 $Y2=0.665
r30 7 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.58 $Y=0.665 $X2=2.89
+ $Y2=0.665
r31 2 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.375 $X2=3.745 $Y2=0.585
r32 1 10 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.375 $X2=2.685 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__FA_1%A_1100_75# 1 2 7 12 13 14 16
r41 16 18 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.425 $Y=0.645
+ $X2=7.425 $Y2=0.725
r42 13 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=0.725
+ $X2=7.425 $Y2=0.725
r43 13 14 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.26 $Y=0.725 $X2=6.66
+ $Y2=0.725
r44 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.575 $Y=0.64
+ $X2=6.66 $Y2=0.725
r45 11 12 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.575 $Y=0.425
+ $X2=6.575 $Y2=0.64
r46 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.49 $Y=0.34
+ $X2=6.575 $Y2=0.425
r47 7 9 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.49 $Y=0.34 $X2=6.19
+ $Y2=0.34
r48 2 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=7.285
+ $Y=0.375 $X2=7.425 $Y2=0.645
r49 1 9 91 $w=1.7e-07 $l=7.07284e-07 $layer=licon1_NDIFF $count=2 $X=5.5
+ $Y=0.375 $X2=6.19 $Y2=0.34
.ends


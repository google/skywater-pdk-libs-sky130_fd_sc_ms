* File: sky130_fd_sc_ms__mux4_1.pex.spice
* Created: Wed Sep  2 12:12:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MUX4_1%A0 3 7 9 12 13
r33 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.38
+ $X2=1.155 $Y2=1.545
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.38
+ $X2=1.155 $Y2=1.215
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.38 $X2=1.155 $Y2=1.38
r36 9 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.155 $Y=1.665
+ $X2=1.155 $Y2=1.38
r37 7 14 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=1.245 $Y=0.69
+ $X2=1.245 $Y2=1.215
r38 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.2 $Y=2.205 $X2=1.2
+ $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A_27_74# 1 2 9 13 17 20 24 30 32 35 38 39 41
+ 44 45 47 51 52 55 56 58 59 61 63 64 65 67 68 69 71 73 82
c184 69 0 1.99713e-19 $X=1.695 $Y=1.2
c185 65 0 6.3344e-20 $X=1.615 $Y=0.945
c186 55 0 1.11609e-19 $X=4.665 $Y=1.445
c187 52 0 2.43471e-20 $X=4.245 $Y=1.285
c188 51 0 1.11257e-19 $X=4.245 $Y=1.285
c189 20 0 1.87958e-19 $X=5.25 $Y=2.435
r190 68 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.365
+ $X2=1.695 $Y2=1.2
r191 67 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.365
+ $X2=1.695 $Y2=1.2
r192 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.695
+ $Y=1.365 $X2=1.695 $Y2=1.365
r193 63 64 6.78944 $w=4.43e-07 $l=8.5e-08 $layer=LI1_cond $X=0.332 $Y=2.035
+ $X2=0.332 $Y2=1.95
r194 59 86 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.61
+ $X2=5.175 $Y2=1.775
r195 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.61 $X2=5.175 $Y2=1.61
r196 56 58 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.75 $Y=1.61
+ $X2=5.175 $Y2=1.61
r197 55 56 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.665 $Y=1.445
+ $X2=4.75 $Y2=1.61
r198 54 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=1.045
+ $X2=4.665 $Y2=0.96
r199 54 55 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.665 $Y=1.045
+ $X2=4.665 $Y2=1.445
r200 52 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.285
+ $X2=4.245 $Y2=1.12
r201 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.245
+ $Y=1.285 $X2=4.245 $Y2=1.285
r202 49 73 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.245 $Y=0.96
+ $X2=4.665 $Y2=0.96
r203 49 51 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.245 $Y=1.045
+ $X2=4.245 $Y2=1.285
r204 48 71 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0.96
+ $X2=2.625 $Y2=0.96
r205 47 49 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=0.96
+ $X2=4.245 $Y2=0.96
r206 47 48 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.08 $Y=0.96
+ $X2=2.79 $Y2=0.96
r207 45 80 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.285
+ $X2=2.625 $Y2=1.45
r208 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.285 $X2=2.625 $Y2=1.285
r209 42 71 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.045
+ $X2=2.625 $Y2=0.96
r210 42 44 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.625 $Y=1.045
+ $X2=2.625 $Y2=1.285
r211 41 71 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.545 $Y=0.875
+ $X2=2.625 $Y2=0.96
r212 40 41 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.545 $Y=0.425
+ $X2=2.545 $Y2=0.875
r213 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=0.34
+ $X2=2.545 $Y2=0.425
r214 38 39 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.46 $Y=0.34
+ $X2=1.7 $Y2=0.34
r215 36 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=1.03
+ $X2=1.615 $Y2=0.945
r216 36 69 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.615 $Y=1.03
+ $X2=1.615 $Y2=1.2
r217 35 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.86
+ $X2=1.615 $Y2=0.945
r218 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=0.425
+ $X2=1.7 $Y2=0.34
r219 34 35 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.615 $Y=0.425
+ $X2=1.615 $Y2=0.86
r220 33 61 2.79892 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.445 $Y=0.945
+ $X2=0.277 $Y2=0.945
r221 32 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=0.945
+ $X2=1.615 $Y2=0.945
r222 32 33 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=1.53 $Y=0.945
+ $X2=0.445 $Y2=0.945
r223 28 63 3.54797 $w=4.43e-07 $l=1.37e-07 $layer=LI1_cond $X=0.332 $Y=2.172
+ $X2=0.332 $Y2=2.035
r224 28 30 14.0624 $w=4.43e-07 $l=5.43e-07 $layer=LI1_cond $X=0.332 $Y=2.172
+ $X2=0.332 $Y2=2.715
r225 26 61 3.67481 $w=2.52e-07 $l=1.19143e-07 $layer=LI1_cond $X=0.195 $Y=1.03
+ $X2=0.277 $Y2=0.945
r226 26 64 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.195 $Y=1.03
+ $X2=0.195 $Y2=1.95
r227 22 61 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=0.86
+ $X2=0.277 $Y2=0.945
r228 22 24 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=0.277 $Y=0.86
+ $X2=0.277 $Y2=0.515
r229 20 86 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.25 $Y=2.435
+ $X2=5.25 $Y2=1.775
r230 17 82 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.155 $Y=0.69
+ $X2=4.155 $Y2=1.12
r231 13 80 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=2.61 $Y=2.205
+ $X2=2.61 $Y2=1.45
r232 9 76 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.635 $Y=0.69
+ $X2=1.635 $Y2=1.2
r233 2 63 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.035
r234 2 30 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.715
r235 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A1 3 7 9 10 14 15
r40 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.38
+ $X2=3.165 $Y2=1.545
r41 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.38
+ $X2=3.165 $Y2=1.215
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=1.38 $X2=3.165 $Y2=1.38
r43 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.165 $Y=1.665
+ $X2=3.165 $Y2=2.035
r44 9 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.165 $Y=1.665
+ $X2=3.165 $Y2=1.38
r45 7 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=2.205
+ $X2=3.12 $Y2=1.545
r46 3 16 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.075 $Y=0.69
+ $X2=3.075 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A2 3 7 9 10 14 15
r37 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.38
+ $X2=3.705 $Y2=1.545
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.38
+ $X2=3.705 $Y2=1.215
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.38 $X2=3.705 $Y2=1.38
r40 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.685 $Y=1.665
+ $X2=3.685 $Y2=2.035
r41 9 15 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.685 $Y=1.665
+ $X2=3.685 $Y2=1.38
r42 7 16 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.765 $Y=0.69
+ $X2=3.765 $Y2=1.215
r43 3 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.74 $Y=2.205
+ $X2=3.74 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%S0 3 8 9 10 11 14 17 18 23 24 25 27 28 30 31
+ 32 35 37 40 41
c122 40 0 1.81924e-19 $X=0.615 $Y=1.38
c123 31 0 1.25715e-19 $X=2.16 $Y=1.085
c124 28 0 1.11257e-19 $X=4.82 $Y=1.085
c125 11 0 1.37343e-19 $X=2.16 $Y=1.175
r126 40 43 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.38
+ $X2=0.6 $Y2=1.545
r127 40 42 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.38
+ $X2=0.6 $Y2=1.215
r128 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.615
+ $Y=1.38 $X2=0.615 $Y2=1.38
r129 37 41 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.635 $Y=1.665
+ $X2=0.635 $Y2=1.38
r130 33 35 48.7128 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=4.725 $Y=1.16
+ $X2=4.82 $Y2=1.16
r131 28 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.82 $Y=1.085
+ $X2=4.82 $Y2=1.16
r132 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.82 $Y=1.085
+ $X2=4.82 $Y2=0.69
r133 26 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.725 $Y=1.235
+ $X2=4.725 $Y2=1.16
r134 26 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.725 $Y=1.235
+ $X2=4.725 $Y2=1.69
r135 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.65 $Y=1.765
+ $X2=4.725 $Y2=1.69
r136 24 25 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.65 $Y=1.765
+ $X2=4.335 $Y2=1.765
r137 21 23 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=4.245 $Y=3.075
+ $X2=4.245 $Y2=2.435
r138 20 25 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.245 $Y=1.84
+ $X2=4.335 $Y2=1.765
r139 20 23 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=4.245 $Y=1.84
+ $X2=4.245 $Y2=2.435
r140 19 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.25 $Y=3.15 $X2=2.16
+ $Y2=3.15
r141 18 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.155 $Y=3.15
+ $X2=4.245 $Y2=3.075
r142 18 19 976.819 $w=1.5e-07 $l=1.905e-06 $layer=POLY_cond $X=4.155 $Y=3.15
+ $X2=2.25 $Y2=3.15
r143 17 31 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.175 $Y=0.69
+ $X2=2.175 $Y2=1.085
r144 12 32 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=3.075
+ $X2=2.16 $Y2=3.15
r145 12 14 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=2.16 $Y=3.075
+ $X2=2.16 $Y2=2.205
r146 11 31 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=1.175
+ $X2=2.16 $Y2=1.085
r147 11 14 400.371 $w=1.8e-07 $l=1.03e-06 $layer=POLY_cond $X=2.16 $Y=1.175
+ $X2=2.16 $Y2=2.205
r148 9 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.07 $Y=3.15 $X2=2.16
+ $Y2=3.15
r149 9 10 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=2.07 $Y=3.15
+ $X2=0.705 $Y2=3.15
r150 8 43 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=0.615 $Y=2.34
+ $X2=0.615 $Y2=1.545
r151 6 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.615 $Y=3.075
+ $X2=0.705 $Y2=3.15
r152 6 8 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=0.615 $Y=3.075
+ $X2=0.615 $Y2=2.34
r153 3 42 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=0.495 $Y=0.69
+ $X2=0.495 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A3 1 3 4 5 6 8 9
c42 9 0 4.73862e-20 $X=6 $Y=1.665
c43 5 0 1.11609e-19 $X=5.285 $Y=1.16
r44 11 13 41.3143 $w=5.25e-07 $l=4.5e-07 $layer=POLY_cond $X=5.88 $Y=1.16
+ $X2=5.88 $Y2=1.61
r45 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.015
+ $Y=1.61 $X2=6.015 $Y2=1.61
r46 6 13 45.6215 $w=5.25e-07 $l=3.44347e-07 $layer=POLY_cond $X=5.67 $Y=1.865
+ $X2=5.88 $Y2=1.61
r47 6 8 152.633 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=5.67 $Y=1.865 $X2=5.67
+ $Y2=2.435
r48 4 11 32.6451 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.61 $Y=1.16 $X2=5.88
+ $Y2=1.16
r49 4 5 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=5.285 $Y2=1.16
r50 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.21 $Y=1.085
+ $X2=5.285 $Y2=1.16
r51 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.21 $Y=1.085
+ $X2=5.21 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A_1396_99# 1 2 9 13 15 17 22 27 29 31 33 36
c63 13 0 2.17476e-19 $X=7.18 $Y=2.46
r64 33 35 17.4812 $w=5.43e-07 $l=5.15e-07 $layer=LI1_cond $X=8.137 $Y=0.665
+ $X2=8.137 $Y2=1.18
r65 30 31 10.4914 $w=1.83e-07 $l=1.75e-07 $layer=LI1_cond $X=7.942 $Y=1.775
+ $X2=7.942 $Y2=1.95
r66 29 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.95 $Y=1.445
+ $X2=7.95 $Y2=1.18
r67 28 36 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.795 $Y=1.61
+ $X2=7.795 $Y2=1.515
r68 27 30 8.13117 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.832 $Y=1.61
+ $X2=7.832 $Y2=1.775
r69 27 29 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.832 $Y=1.61
+ $X2=7.832 $Y2=1.445
r70 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.795
+ $Y=1.61 $X2=7.795 $Y2=1.61
r71 22 31 7.96936 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=2.115
+ $X2=8.015 $Y2=1.95
r72 16 17 6.66866 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.27 $Y=1.515
+ $X2=7.125 $Y2=1.515
r73 15 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.795 $Y2=1.515
r74 15 16 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.27 $Y2=1.515
r75 11 17 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=7.18 $Y=1.59
+ $X2=7.125 $Y2=1.515
r76 11 13 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=7.18 $Y=1.59
+ $X2=7.18 $Y2=2.46
r77 7 17 18.8402 $w=1.65e-07 $l=1.04283e-07 $layer=POLY_cond $X=7.055 $Y=1.44
+ $X2=7.125 $Y2=1.515
r78 7 9 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.055 $Y=1.44
+ $X2=7.055 $Y2=0.945
r79 2 22 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=7.87
+ $Y=1.935 $X2=8.015 $Y2=2.115
r80 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=8.1
+ $Y=0.52 $X2=8.245 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%S1 4 7 9 10 11 13 18 20 21 25
c77 20 0 4.73862e-20 $X=6.655 $Y=1.49
c78 11 0 7.34196e-20 $X=8.29 $Y=1.77
c79 4 0 1.50188e-19 $X=6.615 $Y=0.945
r80 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.37
+ $Y=1.515 $X2=8.37 $Y2=1.515
r81 21 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=8.37 $Y=1.665
+ $X2=8.37 $Y2=1.515
r82 19 20 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.655 $Y=1.34
+ $X2=6.655 $Y2=1.49
r83 16 24 38.5662 $w=2.97e-07 $l=2.06325e-07 $layer=POLY_cond $X=8.46 $Y=1.35
+ $X2=8.367 $Y2=1.515
r84 16 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=8.46 $Y=1.35
+ $X2=8.46 $Y2=0.84
r85 15 18 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=8.46 $Y=0.255
+ $X2=8.46 $Y2=0.84
r86 11 24 48.8089 $w=2.97e-07 $l=2.90964e-07 $layer=POLY_cond $X=8.29 $Y=1.77
+ $X2=8.367 $Y2=1.515
r87 11 13 258.492 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=8.29 $Y=1.77
+ $X2=8.29 $Y2=2.435
r88 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.385 $Y=0.18
+ $X2=8.46 $Y2=0.255
r89 9 10 869.138 $w=1.5e-07 $l=1.695e-06 $layer=POLY_cond $X=8.385 $Y=0.18
+ $X2=6.69 $Y2=0.18
r90 7 20 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=6.68 $Y=2.46 $X2=6.68
+ $Y2=1.49
r91 4 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.615 $Y=0.945
+ $X2=6.615 $Y2=1.34
r92 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.615 $Y=0.255
+ $X2=6.69 $Y2=0.18
r93 1 4 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.615 $Y=0.255
+ $X2=6.615 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A_1338_125# 1 2 9 13 15 18 21 22 24 25 26 28
+ 32 39
c80 25 0 7.34196e-20 $X=8.745 $Y=2.035
c81 15 0 1.50188e-19 $X=6.955 $Y=1.285
r82 38 39 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=9.03 $Y=1.515 $X2=9.08
+ $Y2=1.515
r83 33 38 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=8.91 $Y=1.515
+ $X2=9.03 $Y2=1.515
r84 32 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=1.515
+ $X2=8.91 $Y2=1.68
r85 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.91
+ $Y=1.515 $X2=8.91 $Y2=1.515
r86 28 35 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.83 $Y=1.95 $X2=8.83
+ $Y2=1.68
r87 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.83 $Y2=1.95
r88 25 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.52 $Y2=2.035
r89 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.435 $Y=2.12
+ $X2=8.52 $Y2=2.035
r90 23 24 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.435 $Y=2.12
+ $X2=8.435 $Y2=2.905
r91 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.35 $Y=2.99
+ $X2=8.435 $Y2=2.905
r92 21 22 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=8.35 $Y=2.99
+ $X2=7.12 $Y2=2.99
r93 18 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.955 $Y=2.105
+ $X2=6.955 $Y2=2.815
r94 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.955 $Y=2.905
+ $X2=7.12 $Y2=2.99
r95 16 20 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.955 $Y=2.905
+ $X2=6.955 $Y2=2.815
r96 15 30 6.41518 $w=3.3e-07 $l=1.76125e-07 $layer=LI1_cond $X=6.955 $Y=1.285
+ $X2=6.932 $Y2=1.12
r97 15 18 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=6.955 $Y=1.285
+ $X2=6.955 $Y2=2.105
r98 11 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.08 $Y=1.68
+ $X2=9.08 $Y2=1.515
r99 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.08 $Y=1.68
+ $X2=9.08 $Y2=2.4
r100 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.03 $Y=1.35
+ $X2=9.03 $Y2=1.515
r101 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.03 $Y=1.35 $X2=9.03
+ $Y2=0.79
r102 2 20 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.96 $X2=6.955 $Y2=2.815
r103 2 18 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.96 $X2=6.955 $Y2=2.105
r104 1 30 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=6.69
+ $Y=0.625 $X2=6.835 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%VPWR 1 2 3 4 15 21 25 29 32 33 35 36 37 49 56
+ 63 64 67 70
c91 25 0 1.87958e-19 $X=5.895 $Y=2.775
c92 15 0 1.81924e-19 $X=0.89 $Y=2.035
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r94 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r95 64 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r97 61 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.02 $Y=3.33
+ $X2=8.855 $Y2=3.33
r98 61 63 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.02 $Y=3.33
+ $X2=9.36 $Y2=3.33
r99 60 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r100 60 68 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33 $X2=6
+ $Y2=3.33
r101 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r102 57 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=5.895 $Y2=3.33
r103 57 59 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=8.4 $Y2=3.33
r104 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.69 $Y=3.33
+ $X2=8.855 $Y2=3.33
r105 56 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.69 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 55 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r107 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.895 $Y2=3.33
r111 49 54 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r112 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 45 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 44 47 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 41 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 37 55 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 37 52 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 35 47 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.12 $Y2=3.33
r122 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.43 $Y2=3.33
r123 34 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.43 $Y2=3.33
r125 32 40 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r127 31 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r129 27 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=3.245
+ $X2=8.855 $Y2=3.33
r130 27 29 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=8.855 $Y=3.245
+ $X2=8.855 $Y2=2.455
r131 23 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.895 $Y=3.245
+ $X2=5.895 $Y2=3.33
r132 23 25 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.895 $Y=3.245
+ $X2=5.895 $Y2=2.775
r133 19 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r134 19 21 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.84
r135 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.89 $Y=2.035
+ $X2=0.89 $Y2=2.715
r136 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r137 13 18 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.715
r138 4 29 300 $w=1.7e-07 $l=7.19305e-07 $layer=licon1_PDIFF $count=2 $X=8.38
+ $Y=1.935 $X2=8.855 $Y2=2.455
r139 3 25 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=5.76
+ $Y=1.935 $X2=5.895 $Y2=2.775
r140 2 21 600 $w=1.7e-07 $l=1.24013e-06 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.705 $X2=3.43 $Y2=2.84
r141 1 18 600 $w=1.7e-07 $l=9.63068e-07 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.84 $X2=0.89 $Y2=2.715
r142 1 15 300 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=2 $X=0.705
+ $Y=1.84 $X2=0.89 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A_342_74# 1 2 3 4 16 17 20 21 22 24 25 26 28
+ 30 33 38 42 45 46 47 51 52 54 55
c138 52 0 1.25754e-19 $X=6.455 $Y=2.42
c139 33 0 1.2171e-19 $X=6.455 $Y=2.815
c140 30 0 9.57651e-20 $X=6.455 $Y=2.115
r141 54 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.27 $Y=0.77
+ $X2=7.105 $Y2=0.77
r142 47 49 3.22021 $w=5.18e-07 $l=1.4e-07 $layer=LI1_cond $X=2.29 $Y=2.42
+ $X2=2.29 $Y2=2.56
r143 45 46 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=1.85
+ $X2=2.29 $Y2=1.685
r144 40 42 4.10641 $w=4.33e-07 $l=1.55e-07 $layer=LI1_cond $X=1.96 $Y=0.812
+ $X2=2.115 $Y2=0.812
r145 38 55 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.575 $Y=0.7
+ $X2=7.105 $Y2=0.7
r146 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.49 $Y=0.785
+ $X2=6.575 $Y2=0.7
r147 35 51 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=6.49 $Y=0.785
+ $X2=6.49 $Y2=1.95
r148 31 52 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.505
+ $X2=6.455 $Y2=2.42
r149 31 33 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.455 $Y=2.505
+ $X2=6.455 $Y2=2.815
r150 30 51 7.49019 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=2.115
+ $X2=6.455 $Y2=1.95
r151 28 52 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.335
+ $X2=6.455 $Y2=2.42
r152 28 30 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.455 $Y=2.335
+ $X2=6.455 $Y2=2.115
r153 25 52 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.29 $Y=2.42
+ $X2=6.455 $Y2=2.42
r154 25 26 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.29 $Y=2.42
+ $X2=5.55 $Y2=2.42
r155 23 26 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.45 $Y=2.505
+ $X2=5.55 $Y2=2.42
r156 23 24 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=5.45 $Y=2.505
+ $X2=5.45 $Y2=2.905
r157 21 24 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.35 $Y=2.99
+ $X2=5.45 $Y2=2.905
r158 21 22 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=5.35 $Y=2.99
+ $X2=4.02 $Y2=2.99
r159 20 22 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.907 $Y=2.905
+ $X2=4.02 $Y2=2.99
r160 19 20 20.4879 $w=2.23e-07 $l=4e-07 $layer=LI1_cond $X=3.907 $Y=2.505
+ $X2=3.907 $Y2=2.905
r161 18 47 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.55 $Y=2.42
+ $X2=2.29 $Y2=2.42
r162 17 19 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.795 $Y=2.42
+ $X2=3.907 $Y2=2.505
r163 17 18 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=3.795 $Y=2.42
+ $X2=2.55 $Y2=2.42
r164 16 47 1.95513 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.335
+ $X2=2.29 $Y2=2.42
r165 15 45 2.18514 $w=5.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.29 $Y=1.945
+ $X2=2.29 $Y2=1.85
r166 15 16 8.97059 $w=5.18e-07 $l=3.9e-07 $layer=LI1_cond $X=2.29 $Y=1.945
+ $X2=2.29 $Y2=2.335
r167 13 42 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=2.115 $Y=1.03
+ $X2=2.115 $Y2=0.812
r168 13 46 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.115 $Y=1.03
+ $X2=2.115 $Y2=1.685
r169 4 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.31
+ $Y=1.96 $X2=6.455 $Y2=2.815
r170 4 30 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=6.31
+ $Y=1.96 $X2=6.455 $Y2=2.115
r171 3 49 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.705 $X2=2.385 $Y2=2.56
r172 3 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.705 $X2=2.385 $Y2=1.85
r173 2 54 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.625 $X2=7.27 $Y2=0.77
r174 1 40 182 $w=1.7e-07 $l=5.50999e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=0.37 $X2=1.96 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%A_846_74# 1 2 3 4 13 18 19 20 21 24 25 27 30
+ 31 33 39 42 46 47 50 53 55
c122 46 0 2.43471e-20 $X=5.165 $Y=2.365
r123 51 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.375 $Y=1.19
+ $X2=7.61 $Y2=1.19
r124 44 46 10.6559 $w=7.38e-07 $l=1.4e-07 $layer=LI1_cond $X=5.025 $Y=2.365
+ $X2=5.165 $Y2=2.365
r125 42 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.61 $Y=1.105
+ $X2=7.61 $Y2=1.19
r126 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.61 $Y=0.435
+ $X2=7.61 $Y2=1.105
r127 39 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=2.11
+ $X2=7.455 $Y2=1.945
r128 35 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.375 $Y=1.275
+ $X2=7.375 $Y2=1.19
r129 35 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.375 $Y=1.275
+ $X2=7.375 $Y2=1.945
r130 33 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.525 $Y=0.35
+ $X2=7.61 $Y2=0.435
r131 33 50 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=7.525 $Y=0.35
+ $X2=6.485 $Y2=0.35
r132 32 49 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6.235 $Y=0.355
+ $X2=6.11 $Y2=0.355
r133 31 50 5.59224 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=6.395 $Y=0.355
+ $X2=6.485 $Y2=0.355
r134 31 32 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=6.395 $Y=0.355
+ $X2=6.235 $Y2=0.355
r135 28 30 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.11 $Y=1.105
+ $X2=6.11 $Y2=0.82
r136 27 49 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.11 $Y=0.445 $X2=6.11
+ $Y2=0.355
r137 27 30 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=6.11 $Y=0.445
+ $X2=6.11 $Y2=0.82
r138 26 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=1.19
+ $X2=5.595 $Y2=1.19
r139 25 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.985 $Y=1.19
+ $X2=6.11 $Y2=1.105
r140 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.985 $Y=1.19
+ $X2=5.68 $Y2=1.19
r141 23 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.275
+ $X2=5.595 $Y2=1.19
r142 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.595 $Y=1.275
+ $X2=5.595 $Y2=1.995
r143 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.51 $Y=2.08
+ $X2=5.595 $Y2=1.995
r144 21 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.51 $Y=2.08
+ $X2=5.165 $Y2=2.08
r145 19 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=1.19
+ $X2=5.595 $Y2=1.19
r146 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.51 $Y=1.19
+ $X2=5.09 $Y2=1.19
r147 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.005 $Y=1.105
+ $X2=5.09 $Y2=1.19
r148 17 18 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.005 $Y=0.705
+ $X2=5.005 $Y2=1.105
r149 13 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.92 $Y=0.54
+ $X2=5.005 $Y2=0.705
r150 13 15 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.92 $Y=0.54
+ $X2=4.485 $Y2=0.54
r151 4 39 300 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=2 $X=7.27
+ $Y=1.96 $X2=7.455 $Y2=2.11
r152 3 44 150 $w=1.7e-07 $l=7.59045e-07 $layer=licon1_PDIFF $count=4 $X=4.335
+ $Y=1.935 $X2=5.025 $Y2=2.08
r153 2 49 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=5.995
+ $Y=0.215 $X2=6.15 $Y2=0.36
r154 2 30 182 $w=1.7e-07 $l=6.78086e-07 $layer=licon1_NDIFF $count=1 $X=5.995
+ $Y=0.215 $X2=6.15 $Y2=0.82
r155 1 15 182 $w=1.7e-07 $l=3.29204e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.37 $X2=4.485 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%X 1 2 7 8 9 10 11 12 13 30
r19 22 30 1.50814 $w=4.03e-07 $l=5.3e-08 $layer=LI1_cond $X=9.282 $Y=0.978
+ $X2=9.282 $Y2=0.925
r20 13 45 7.30194 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=9.352 $Y=2.725
+ $X2=9.352 $Y2=2.56
r21 12 45 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=9.365 $Y=2.405
+ $X2=9.365 $Y2=2.56
r22 11 12 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.365 $Y=2.035
+ $X2=9.365 $Y2=2.405
r23 10 11 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.365 $Y=1.665
+ $X2=9.365 $Y2=2.035
r24 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.365 $Y=1.295
+ $X2=9.365 $Y2=1.665
r25 9 42 5.52212 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=9.365 $Y=1.295
+ $X2=9.365 $Y2=1.18
r26 8 42 7.19001 $w=4.03e-07 $l=1.86e-07 $layer=LI1_cond $X=9.282 $Y=0.994
+ $X2=9.282 $Y2=1.18
r27 8 22 0.455286 $w=4.03e-07 $l=1.6e-08 $layer=LI1_cond $X=9.282 $Y=0.994
+ $X2=9.282 $Y2=0.978
r28 8 30 0.455286 $w=4.03e-07 $l=1.6e-08 $layer=LI1_cond $X=9.282 $Y=0.909
+ $X2=9.282 $Y2=0.925
r29 8 27 9.78865 $w=4.03e-07 $l=3.44e-07 $layer=LI1_cond $X=9.282 $Y=0.909
+ $X2=9.282 $Y2=0.565
r30 7 27 0.284554 $w=4.03e-07 $l=1e-08 $layer=LI1_cond $X=9.282 $Y=0.555
+ $X2=9.282 $Y2=0.565
r31 2 13 600 $w=1.7e-07 $l=9.52431e-07 $layer=licon1_PDIFF $count=1 $X=9.17
+ $Y=1.84 $X2=9.31 $Y2=2.725
r32 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.42 $X2=9.245 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_1%VGND 1 2 3 4 17 21 25 29 32 33 34 36 44 57 58
+ 61 64 67
r83 67 68 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r84 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r87 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r88 55 68 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=5.52
+ $Y2=0
r89 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r90 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.425
+ $Y2=0
r91 52 54 183.326 $w=1.68e-07 $l=2.81e-06 $layer=LI1_cond $X=5.59 $Y=0 $X2=8.4
+ $Y2=0
r92 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r93 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r94 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r95 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r96 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r97 45 64 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.42
+ $Y2=0
r98 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=4.08
+ $Y2=0
r99 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.425
+ $Y2=0
r100 44 50 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r101 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r102 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r103 40 43 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r104 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r105 39 42 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r106 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r107 37 61 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.895
+ $Y2=0
r108 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=1.2
+ $Y2=0
r109 36 64 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.42
+ $Y2=0
r110 36 42 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.12
+ $Y2=0
r111 34 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r112 34 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.08
+ $Y2=0
r113 32 54 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.58 $Y=0 $X2=8.4
+ $Y2=0
r114 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=0 $X2=8.745
+ $Y2=0
r115 31 57 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=0 $X2=9.36
+ $Y2=0
r116 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=0 $X2=8.745
+ $Y2=0
r117 27 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=0.085
+ $X2=8.745 $Y2=0
r118 27 29 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=8.745 $Y=0.085
+ $X2=8.745 $Y2=0.665
r119 23 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0
r120 23 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0.495
r121 19 64 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r122 19 21 8.71718 $w=5.88e-07 $l=4.3e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.515
r123 15 61 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0
r124 15 17 13.7407 $w=3.88e-07 $l=4.65e-07 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0.55
r125 4 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.535
+ $Y=0.52 $X2=8.745 $Y2=0.665
r126 3 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.425 $Y2=0.495
r127 2 21 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.37 $X2=3.42 $Y2=0.515
r128 1 17 182 $w=1.7e-07 $l=4.05123e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.895 $Y2=0.55
.ends


* File: sky130_fd_sc_ms__or2b_4.spice
* Created: Fri Aug 28 18:07:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or2b_4.pex.spice"
.subckt sky130_fd_sc_ms__or2b_4  VNB VPB A B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_81_296#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_81_296#_M1010_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1010_d N_A_81_296#_M1012_g N_X_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.11285 PD=1.09 PS=1.045 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_81_296#_M1013_g N_X_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.11285 PD=1.14217 PS=1.045 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75001.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1000 N_A_81_296#_M1000_d N_A_M1000_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.144 AS=0.108058 PD=1.09 PS=0.987826 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1007 N_A_81_296#_M1000_d N_A_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.144 AS=0.112 PD=1.09 PS=0.99 NRD=18.744 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_81_296#_M1006_d N_A_676_48#_M1006_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75003.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1017 N_A_81_296#_M1006_d N_A_676_48#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1014 N_A_676_48#_M1014_d N_B_N_M1014_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.6272 AS=0.112 PD=3.24 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75004.1
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1008 N_X_M1008_d N_A_81_296#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1008_d N_A_81_296#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1011_d N_A_81_296#_M1011_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1016 N_X_M1011_d N_A_81_296#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.199381 PD=1.39 PS=1.54792 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1003 N_A_492_392#_M1003_d N_A_M1003_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.178019 PD=1.27 PS=1.38208 NRD=0 NRS=13.7703 M=1 R=5.55556
+ SA=90002.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1004 N_A_492_392#_M1003_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_81_296#_M1001_d N_A_676_48#_M1001_g N_A_492_392#_M1001_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1002 N_A_81_296#_M1001_d N_A_676_48#_M1002_g N_A_492_392#_M1002_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1015 N_A_676_48#_M1015_d N_B_N_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18 W=1
+ AD=0.27 AS=0.275 PD=2.54 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__or2b_4.pxi.spice"
*
.ends
*
*

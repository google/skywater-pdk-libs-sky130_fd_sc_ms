* File: sky130_fd_sc_ms__a222oi_2.pxi.spice
* Created: Fri Aug 28 17:02:20 2020
* 
x_PM_SKY130_FD_SC_MS__A222OI_2%C2 N_C2_M1002_g N_C2_M1008_g N_C2_M1018_g
+ N_C2_M1010_g N_C2_c_128_n N_C2_c_129_n N_C2_c_130_n N_C2_c_131_n N_C2_c_139_n
+ N_C2_c_140_n N_C2_c_132_n N_C2_c_133_n C2 N_C2_c_135_n
+ PM_SKY130_FD_SC_MS__A222OI_2%C2
x_PM_SKY130_FD_SC_MS__A222OI_2%C1 N_C1_M1003_g N_C1_M1004_g N_C1_M1016_g
+ N_C1_M1011_g N_C1_c_218_n N_C1_c_223_n C1 N_C1_c_220_n
+ PM_SKY130_FD_SC_MS__A222OI_2%C1
x_PM_SKY130_FD_SC_MS__A222OI_2%B1 N_B1_M1020_g N_B1_M1007_g N_B1_M1014_g
+ N_B1_M1023_g N_B1_c_274_n N_B1_c_282_n N_B1_c_283_n N_B1_c_322_p N_B1_c_284_n
+ N_B1_c_275_n N_B1_c_276_n B1 N_B1_c_277_n N_B1_c_278_n
+ PM_SKY130_FD_SC_MS__A222OI_2%B1
x_PM_SKY130_FD_SC_MS__A222OI_2%B2 N_B2_M1009_g N_B2_M1012_g N_B2_M1013_g
+ N_B2_c_370_n N_B2_M1015_g B2 N_B2_c_371_n N_B2_c_372_n
+ PM_SKY130_FD_SC_MS__A222OI_2%B2
x_PM_SKY130_FD_SC_MS__A222OI_2%A1 N_A1_M1017_g N_A1_M1005_g N_A1_M1006_g
+ N_A1_M1022_g N_A1_c_436_n N_A1_c_437_n N_A1_c_482_p N_A1_c_438_n N_A1_c_430_n
+ N_A1_c_431_n A1 N_A1_c_432_n N_A1_c_433_n PM_SKY130_FD_SC_MS__A222OI_2%A1
x_PM_SKY130_FD_SC_MS__A222OI_2%A2 N_A2_M1019_g N_A2_M1000_g N_A2_M1021_g
+ N_A2_M1001_g A2 N_A2_c_521_n PM_SKY130_FD_SC_MS__A222OI_2%A2
x_PM_SKY130_FD_SC_MS__A222OI_2%Y N_Y_M1004_s N_Y_M1020_s N_Y_M1023_s N_Y_M1006_s
+ N_Y_M1002_s N_Y_M1003_d N_Y_M1018_s N_Y_c_572_n N_Y_c_573_n N_Y_c_591_n
+ N_Y_c_673_p N_Y_c_596_n N_Y_c_574_n N_Y_c_575_n N_Y_c_576_n N_Y_c_577_n
+ N_Y_c_578_n N_Y_c_579_n N_Y_c_580_n N_Y_c_607_n N_Y_c_608_n N_Y_c_610_n
+ N_Y_c_583_n Y Y Y PM_SKY130_FD_SC_MS__A222OI_2%Y
x_PM_SKY130_FD_SC_MS__A222OI_2%A_119_392# N_A_119_392#_M1002_d
+ N_A_119_392#_M1016_s N_A_119_392#_M1007_d N_A_119_392#_M1013_s
+ N_A_119_392#_c_726_n N_A_119_392#_c_720_n N_A_119_392#_c_721_n
+ N_A_119_392#_c_728_n N_A_119_392#_c_722_n N_A_119_392#_c_723_n
+ N_A_119_392#_c_724_n N_A_119_392#_c_725_n
+ PM_SKY130_FD_SC_MS__A222OI_2%A_119_392#
x_PM_SKY130_FD_SC_MS__A222OI_2%A_515_392# N_A_515_392#_M1007_s
+ N_A_515_392#_M1012_d N_A_515_392#_M1014_s N_A_515_392#_M1019_d
+ N_A_515_392#_M1022_s N_A_515_392#_c_782_n N_A_515_392#_c_826_n
+ N_A_515_392#_c_784_n N_A_515_392#_c_776_n N_A_515_392#_c_803_n
+ N_A_515_392#_c_777_n N_A_515_392#_c_807_n N_A_515_392#_c_778_n
+ N_A_515_392#_c_829_n N_A_515_392#_c_779_n N_A_515_392#_c_815_n
+ N_A_515_392#_c_780_n PM_SKY130_FD_SC_MS__A222OI_2%A_515_392#
x_PM_SKY130_FD_SC_MS__A222OI_2%VPWR N_VPWR_M1017_d N_VPWR_M1021_s N_VPWR_c_856_n
+ N_VPWR_c_857_n VPWR N_VPWR_c_858_n N_VPWR_c_859_n N_VPWR_c_860_n
+ N_VPWR_c_855_n N_VPWR_c_862_n N_VPWR_c_863_n PM_SKY130_FD_SC_MS__A222OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A222OI_2%VGND N_VGND_M1008_d N_VGND_M1010_d N_VGND_M1009_d
+ N_VGND_M1000_d N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n
+ VGND N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n
+ N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n
+ PM_SKY130_FD_SC_MS__A222OI_2%VGND
x_PM_SKY130_FD_SC_MS__A222OI_2%A_137_74# N_A_137_74#_M1008_s N_A_137_74#_M1011_d
+ N_A_137_74#_c_1015_n PM_SKY130_FD_SC_MS__A222OI_2%A_137_74#
x_PM_SKY130_FD_SC_MS__A222OI_2%A_593_74# N_A_593_74#_M1020_d N_A_593_74#_M1015_s
+ N_A_593_74#_c_1030_n N_A_593_74#_c_1028_n N_A_593_74#_c_1029_n
+ PM_SKY130_FD_SC_MS__A222OI_2%A_593_74#
x_PM_SKY130_FD_SC_MS__A222OI_2%A_981_74# N_A_981_74#_M1005_d N_A_981_74#_M1001_s
+ N_A_981_74#_c_1054_n N_A_981_74#_c_1061_n N_A_981_74#_c_1057_n
+ N_A_981_74#_c_1058_n N_A_981_74#_c_1055_n
+ PM_SKY130_FD_SC_MS__A222OI_2%A_981_74#
cc_1 VNB N_C2_M1002_g 0.0104319f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_2 VNB N_C2_M1008_g 0.0214368f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_3 VNB N_C2_c_128_n 0.0207721f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.13
cc_4 VNB N_C2_c_129_n 0.0277839f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.635
cc_5 VNB N_C2_c_130_n 0.00204176f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.8
cc_6 VNB N_C2_c_131_n 0.00280946f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_7 VNB N_C2_c_132_n 0.00263864f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_8 VNB N_C2_c_133_n 0.0188881f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_9 VNB C2 0.00453826f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_C2_c_135_n 0.033161f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.33
cc_11 VNB N_C1_M1004_g 0.0197442f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_12 VNB N_C1_M1016_g 0.00871368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C1_M1011_g 0.0196961f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_14 VNB N_C1_c_218_n 0.00871426f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.635
cc_15 VNB C1 0.00139126f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.495
cc_16 VNB N_C1_c_220_n 0.0367937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1020_g 0.0415299f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_18 VNB N_B1_M1023_g 0.0345024f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_19 VNB N_B1_c_274_n 0.00340496f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.13
cc_20 VNB N_B1_c_275_n 0.00354957f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_21 VNB N_B1_c_276_n 0.0166452f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_22 VNB N_B1_c_277_n 0.0188982f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.33
cc_23 VNB N_B1_c_278_n 0.00188639f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.33
cc_24 VNB N_B2_M1009_g 0.0261081f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_25 VNB N_B2_M1012_g 0.00348647f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_26 VNB N_B2_M1013_g 0.00359827f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=2.46
cc_27 VNB N_B2_c_370_n 0.0165083f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.13
cc_28 VNB N_B2_c_371_n 0.00359946f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.75
cc_29 VNB N_B2_c_372_n 0.0730116f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.75
cc_30 VNB N_A1_M1005_g 0.0352532f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_31 VNB N_A1_M1006_g 0.0442873f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=2.46
cc_32 VNB N_A1_c_430_n 0.0159934f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_33 VNB N_A1_c_431_n 0.00360097f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_34 VNB N_A1_c_432_n 0.0204373f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.165
cc_35 VNB N_A1_c_433_n 0.0124003f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.495
cc_36 VNB N_A2_M1000_g 0.0342909f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_37 VNB N_A2_M1001_g 0.0328015f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_38 VNB A2 0.00102026f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.13
cc_39 VNB N_A2_c_521_n 0.025771f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_40 VNB N_Y_c_572_n 0.0315443f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.75
cc_41 VNB N_Y_c_573_n 0.00803133f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_42 VNB N_Y_c_574_n 0.00739598f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_43 VNB N_Y_c_575_n 0.0077195f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.33
cc_44 VNB N_Y_c_576_n 0.0166262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_577_n 0.0234737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_578_n 0.0021982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_579_n 0.0321153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_580_n 0.0318202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_855_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.33
cc_50 VNB N_VGND_c_926_n 0.01289f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.13
cc_51 VNB N_VGND_c_927_n 0.0246219f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_52 VNB N_VGND_c_928_n 0.0128186f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.8
cc_53 VNB N_VGND_c_929_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.75
cc_54 VNB N_VGND_c_930_n 0.0378216f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.295
cc_55 VNB N_VGND_c_931_n 0.0317955f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.165
cc_56 VNB N_VGND_c_932_n 0.0415162f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.33
cc_57 VNB N_VGND_c_933_n 0.0299361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_934_n 0.370389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_935_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_936_n 0.0155699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_937_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_137_74#_c_1015_n 0.00685031f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.69
cc_63 VNB N_A_593_74#_c_1028_n 0.00204804f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=2.46
cc_64 VNB N_A_593_74#_c_1029_n 0.00204804f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_65 VNB N_A_981_74#_c_1054_n 0.00284399f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.8
cc_66 VNB N_A_981_74#_c_1055_n 0.00215161f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.69
cc_67 VPB N_C2_M1002_g 0.034302f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_68 VPB N_C2_M1018_g 0.0242077f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_69 VPB N_C2_c_130_n 0.0140112f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.8
cc_70 VPB N_C2_c_139_n 0.0205246f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.75
cc_71 VPB N_C2_c_140_n 0.00387294f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.75
cc_72 VPB N_C1_M1016_g 0.0266462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_C1_c_218_n 0.00324744f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.635
cc_74 VPB N_C1_c_223_n 0.0290913f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.8
cc_75 VPB N_B1_M1007_g 0.0244628f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.69
cc_76 VPB N_B1_M1014_g 0.0243306f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_77 VPB N_B1_c_274_n 9.55489e-19 $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_78 VPB N_B1_c_282_n 0.00269414f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.635
cc_79 VPB N_B1_c_283_n 0.00962097f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.8
cc_80 VPB N_B1_c_284_n 0.00333193f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.75
cc_81 VPB N_B1_c_275_n 0.00184657f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_82 VPB N_B1_c_276_n 0.0109595f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_83 VPB N_B1_c_277_n 0.0148352f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_84 VPB N_B1_c_278_n 0.00153498f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.33
cc_85 VPB N_B2_M1012_g 0.028157f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.69
cc_86 VPB N_B2_M1013_g 0.0298842f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_87 VPB N_B2_c_371_n 0.00323444f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.75
cc_88 VPB N_A1_M1017_g 0.0228661f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_89 VPB N_A1_M1022_g 0.0302933f $X=-0.19 $Y=1.66 $X2=1.9 $Y2=0.69
cc_90 VPB N_A1_c_436_n 0.00344758f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.635
cc_91 VPB N_A1_c_437_n 0.00488508f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.8
cc_92 VPB N_A1_c_438_n 0.00354832f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.75
cc_93 VPB N_A1_c_430_n 0.0106933f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_94 VPB N_A1_c_431_n 0.00180389f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_95 VPB N_A1_c_432_n 0.0127646f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.165
cc_96 VPB N_A1_c_433_n 0.007317f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.495
cc_97 VPB N_A2_M1019_g 0.0222357f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_98 VPB N_A2_M1021_g 0.021883f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=2.46
cc_99 VPB A2 8.34758e-19 $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_100 VPB N_A2_c_521_n 0.0148892f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_101 VPB N_Y_c_572_n 0.0125731f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.75
cc_102 VPB N_Y_c_574_n 0.00742463f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_103 VPB N_Y_c_583_n 0.0106183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB Y 0.0155085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB Y 0.0334941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_119_392#_c_720_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_107 VPB N_A_119_392#_c_721_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.635
cc_108 VPB N_A_119_392#_c_722_n 0.00534149f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_109 VPB N_A_119_392#_c_723_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_110 VPB N_A_119_392#_c_724_n 0.0142686f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.33
cc_111 VPB N_A_119_392#_c_725_n 0.0019546f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_112 VPB N_A_515_392#_c_776_n 0.00399881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_515_392#_c_777_n 0.00233129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_515_392#_c_778_n 0.0169341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_515_392#_c_779_n 0.00219668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_515_392#_c_780_n 0.029936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_856_n 0.00329267f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=1.8
cc_118 VPB N_VPWR_c_857_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.9 $Y2=1.13
cc_119 VPB N_VPWR_c_858_n 0.119356f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.13
cc_120 VPB N_VPWR_c_859_n 0.0159778f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.295
cc_121 VPB N_VPWR_c_860_n 0.0177874f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.33
cc_122 VPB N_VPWR_c_855_n 0.076024f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.33
cc_123 VPB N_VPWR_c_862_n 0.00656574f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.495
cc_124 VPB N_VPWR_c_863_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 N_C2_M1008_g N_C1_M1004_g 0.0276308f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_126 N_C2_c_129_n N_C1_M1016_g 0.0433281f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_127 N_C2_c_139_n N_C1_M1016_g 0.0157037f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_128 N_C2_c_132_n N_C1_M1016_g 0.00108316f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_129 N_C2_c_128_n N_C1_M1011_g 0.0224f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_130 N_C2_c_132_n N_C1_M1011_g 0.00174486f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_131 N_C2_c_133_n N_C1_M1011_g 0.00978324f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_132 N_C2_M1002_g N_C1_c_218_n 0.0058994f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_133 N_C2_c_131_n N_C1_c_218_n 0.00312674f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_134 N_C2_c_139_n N_C1_c_218_n 0.00520968f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_135 N_C2_M1002_g N_C1_c_223_n 0.0305024f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_136 N_C2_c_139_n N_C1_c_223_n 0.00871786f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_137 N_C2_c_139_n C1 0.0243679f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_138 N_C2_c_132_n C1 0.0110236f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_139 N_C2_c_133_n C1 8.95767e-19 $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_140 C2 C1 0.0265726f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_141 N_C2_c_135_n C1 3.29091e-19 $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_142 N_C2_c_129_n N_C1_c_220_n 0.00978324f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_143 N_C2_c_139_n N_C1_c_220_n 0.0011826f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_144 C2 N_C1_c_220_n 0.00312674f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_145 N_C2_c_135_n N_C1_c_220_n 0.0213924f $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_146 N_C2_c_133_n N_B1_M1020_g 0.00335539f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_147 N_C2_c_129_n N_B1_c_277_n 0.00519886f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_148 N_C2_M1008_g N_Y_c_572_n 0.00514335f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_149 N_C2_c_131_n N_Y_c_572_n 0.00787536f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_150 N_C2_c_140_n N_Y_c_572_n 0.00866338f $X=0.835 $Y=1.75 $X2=0 $Y2=0
cc_151 C2 N_Y_c_572_n 0.0252195f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_152 N_C2_c_135_n N_Y_c_572_n 0.018006f $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_153 N_C2_M1002_g N_Y_c_591_n 0.0164355f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_154 N_C2_c_139_n N_Y_c_591_n 0.0139362f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_155 N_C2_c_140_n N_Y_c_591_n 0.0163035f $X=0.835 $Y=1.75 $X2=0 $Y2=0
cc_156 C2 N_Y_c_591_n 0.00508596f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_157 N_C2_c_135_n N_Y_c_591_n 4.50378e-19 $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_158 N_C2_M1018_g N_Y_c_596_n 0.0142101f $X=1.885 $Y=2.46 $X2=0 $Y2=0
cc_159 N_C2_c_139_n N_Y_c_596_n 0.0433701f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_160 N_C2_M1018_g N_Y_c_574_n 0.0047678f $X=1.885 $Y=2.46 $X2=0 $Y2=0
cc_161 N_C2_c_129_n N_Y_c_574_n 0.00361657f $X=1.96 $Y=1.635 $X2=0 $Y2=0
cc_162 N_C2_c_130_n N_Y_c_574_n 5.25314e-19 $X=1.96 $Y=1.8 $X2=0 $Y2=0
cc_163 N_C2_c_139_n N_Y_c_574_n 0.0137446f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_164 N_C2_c_132_n N_Y_c_574_n 0.0273195f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_165 N_C2_c_128_n N_Y_c_575_n 0.00103145f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_166 N_C2_c_128_n N_Y_c_577_n 0.00440566f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_167 N_C2_c_132_n N_Y_c_577_n 0.0140395f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_168 N_C2_c_133_n N_Y_c_577_n 0.00192034f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_169 N_C2_c_139_n N_Y_c_607_n 0.0179902f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_170 N_C2_M1008_g N_Y_c_608_n 2.14939e-19 $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_171 N_C2_c_128_n N_Y_c_608_n 4.40457e-19 $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_172 N_C2_M1008_g N_Y_c_610_n 0.0133138f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_173 N_C2_c_139_n N_Y_c_610_n 0.00497809f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_174 C2 N_Y_c_610_n 0.0270966f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_175 N_C2_c_135_n N_Y_c_610_n 0.00145942f $X=0.59 $Y=1.33 $X2=0 $Y2=0
cc_176 N_C2_c_130_n N_Y_c_583_n 8.20456e-19 $X=1.96 $Y=1.8 $X2=0 $Y2=0
cc_177 N_C2_c_139_n N_Y_c_583_n 0.0103156f $X=1.795 $Y=1.75 $X2=0 $Y2=0
cc_178 N_C2_M1002_g Y 0.0016711f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_179 N_C2_M1002_g Y 4.70646e-19 $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_180 N_C2_M1002_g N_A_119_392#_c_726_n 0.00757756f $X=0.505 $Y=2.46 $X2=0
+ $Y2=0
cc_181 N_C2_M1002_g N_A_119_392#_c_721_n 0.00694332f $X=0.505 $Y=2.46 $X2=0
+ $Y2=0
cc_182 N_C2_M1018_g N_A_119_392#_c_728_n 0.0126153f $X=1.885 $Y=2.46 $X2=0 $Y2=0
cc_183 N_C2_M1018_g N_A_119_392#_c_723_n 0.00191106f $X=1.885 $Y=2.46 $X2=0
+ $Y2=0
cc_184 N_C2_M1018_g N_A_119_392#_c_724_n 0.0137576f $X=1.885 $Y=2.46 $X2=0 $Y2=0
cc_185 N_C2_M1002_g N_VPWR_c_858_n 0.00517089f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_186 N_C2_M1018_g N_VPWR_c_858_n 0.00333896f $X=1.885 $Y=2.46 $X2=0 $Y2=0
cc_187 N_C2_M1002_g N_VPWR_c_855_n 0.00982428f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_188 N_C2_M1018_g N_VPWR_c_855_n 0.00427929f $X=1.885 $Y=2.46 $X2=0 $Y2=0
cc_189 N_C2_M1008_g N_VGND_c_927_n 0.0105743f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_190 N_C2_c_128_n N_VGND_c_928_n 0.0118294f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_191 N_C2_c_132_n N_VGND_c_928_n 0.0114324f $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_192 N_C2_c_133_n N_VGND_c_928_n 9.66467e-19 $X=1.96 $Y=1.295 $X2=0 $Y2=0
cc_193 N_C2_M1008_g N_VGND_c_930_n 0.00433162f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_194 N_C2_c_128_n N_VGND_c_930_n 0.00383152f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_195 N_C2_M1008_g N_VGND_c_934_n 0.00446997f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_196 N_C2_c_128_n N_VGND_c_934_n 0.00757637f $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_197 N_C2_M1008_g N_A_137_74#_c_1015_n 0.00366414f $X=0.61 $Y=0.69 $X2=0 $Y2=0
cc_198 N_C2_c_128_n N_A_137_74#_c_1015_n 7.20798e-19 $X=1.96 $Y=1.13 $X2=0 $Y2=0
cc_199 N_C1_c_223_n N_Y_c_591_n 0.0142175f $X=0.99 $Y=1.885 $X2=0 $Y2=0
cc_200 N_C1_M1016_g N_Y_c_596_n 0.0142175f $X=1.435 $Y=2.46 $X2=0 $Y2=0
cc_201 N_C1_c_223_n N_Y_c_607_n 0.00132091f $X=0.99 $Y=1.885 $X2=0 $Y2=0
cc_202 N_C1_M1004_g N_Y_c_608_n 0.00185091f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_203 N_C1_M1011_g N_Y_c_608_n 0.00411699f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_204 N_C1_c_220_n N_Y_c_608_n 7.12379e-19 $X=1.47 $Y=1.33 $X2=0 $Y2=0
cc_205 N_C1_M1004_g N_Y_c_610_n 0.00815093f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_206 C1 N_Y_c_610_n 0.0221715f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_207 N_C1_M1016_g N_A_119_392#_c_726_n 5.39294e-19 $X=1.435 $Y=2.46 $X2=0
+ $Y2=0
cc_208 N_C1_c_223_n N_A_119_392#_c_726_n 0.00830259f $X=0.99 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_C1_M1016_g N_A_119_392#_c_720_n 0.011817f $X=1.435 $Y=2.46 $X2=0 $Y2=0
cc_210 N_C1_c_223_n N_A_119_392#_c_720_n 0.011817f $X=0.99 $Y=1.885 $X2=0 $Y2=0
cc_211 N_C1_c_223_n N_A_119_392#_c_721_n 0.001916f $X=0.99 $Y=1.885 $X2=0 $Y2=0
cc_212 N_C1_M1016_g N_A_119_392#_c_728_n 0.00830259f $X=1.435 $Y=2.46 $X2=0
+ $Y2=0
cc_213 N_C1_c_223_n N_A_119_392#_c_728_n 5.39294e-19 $X=0.99 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_C1_M1016_g N_A_119_392#_c_723_n 0.001916f $X=1.435 $Y=2.46 $X2=0 $Y2=0
cc_215 N_C1_M1016_g N_VPWR_c_858_n 0.00333896f $X=1.435 $Y=2.46 $X2=0 $Y2=0
cc_216 N_C1_c_223_n N_VPWR_c_858_n 0.00333896f $X=0.99 $Y=1.885 $X2=0 $Y2=0
cc_217 N_C1_M1016_g N_VPWR_c_855_n 0.00423094f $X=1.435 $Y=2.46 $X2=0 $Y2=0
cc_218 N_C1_c_223_n N_VPWR_c_855_n 0.00423094f $X=0.99 $Y=1.885 $X2=0 $Y2=0
cc_219 N_C1_M1011_g N_VGND_c_928_n 9.22378e-19 $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_220 N_C1_M1004_g N_VGND_c_930_n 0.00291649f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_221 N_C1_M1011_g N_VGND_c_930_n 0.00291649f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_222 N_C1_M1004_g N_VGND_c_934_n 0.00359219f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_223 N_C1_M1011_g N_VGND_c_934_n 0.00359219f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_224 N_C1_M1004_g N_A_137_74#_c_1015_n 0.0106323f $X=1.04 $Y=0.69 $X2=0 $Y2=0
cc_225 N_C1_M1011_g N_A_137_74#_c_1015_n 0.0156912f $X=1.47 $Y=0.69 $X2=0 $Y2=0
cc_226 N_B1_M1020_g N_B2_M1009_g 0.040022f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_227 N_B1_c_274_n N_B2_M1012_g 0.00204456f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_228 N_B1_c_282_n N_B2_M1012_g 0.00347946f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_229 N_B1_c_283_n N_B2_M1012_g 0.0143336f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_230 N_B1_c_277_n N_B2_M1012_g 0.0520199f $X=2.84 $Y=1.635 $X2=0 $Y2=0
cc_231 N_B1_M1014_g N_B2_M1013_g 0.0319503f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_232 N_B1_c_283_n N_B2_M1013_g 0.0173194f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_233 N_B1_c_284_n N_B2_M1013_g 0.00366877f $X=4.19 $Y=1.95 $X2=0 $Y2=0
cc_234 N_B1_M1023_g N_B2_c_370_n 0.0286129f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_235 N_B1_M1020_g N_B2_c_371_n 8.86752e-19 $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_236 N_B1_M1023_g N_B2_c_371_n 7.75734e-19 $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_237 N_B1_c_274_n N_B2_c_371_n 0.0256873f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_238 N_B1_c_283_n N_B2_c_371_n 0.0264559f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_239 N_B1_c_275_n N_B2_c_371_n 0.0154943f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_240 N_B1_c_277_n N_B2_c_371_n 2.29946e-19 $X=2.84 $Y=1.635 $X2=0 $Y2=0
cc_241 N_B1_M1023_g N_B2_c_372_n 0.00771183f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_242 N_B1_c_274_n N_B2_c_372_n 0.00109171f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_243 N_B1_c_283_n N_B2_c_372_n 0.00243942f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_244 N_B1_c_275_n N_B2_c_372_n 0.00273929f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_245 N_B1_c_276_n N_B2_c_372_n 0.0206191f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_246 N_B1_c_277_n N_B2_c_372_n 0.00781816f $X=2.84 $Y=1.635 $X2=0 $Y2=0
cc_247 N_B1_M1014_g N_A1_M1017_g 0.0142042f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_248 N_B1_M1023_g N_A1_M1005_g 0.0266162f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_249 N_B1_c_284_n N_A1_c_436_n 0.00477427f $X=4.19 $Y=1.95 $X2=0 $Y2=0
cc_250 N_B1_c_275_n N_A1_c_430_n 4.14342e-19 $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_251 N_B1_c_276_n N_A1_c_430_n 0.0214313f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_252 N_B1_c_275_n N_A1_c_431_n 0.0215802f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_253 N_B1_c_276_n N_A1_c_431_n 4.13565e-19 $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_254 N_B1_M1020_g N_Y_c_574_n 0.00329148f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_255 N_B1_M1007_g N_Y_c_574_n 0.0030209f $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_256 N_B1_c_282_n N_Y_c_574_n 0.0046204f $X=3.15 $Y=1.95 $X2=0 $Y2=0
cc_257 N_B1_c_322_p N_Y_c_574_n 4.83753e-19 $X=3.235 $Y=2.035 $X2=0 $Y2=0
cc_258 N_B1_c_277_n N_Y_c_574_n 0.00128193f $X=2.84 $Y=1.635 $X2=0 $Y2=0
cc_259 N_B1_c_278_n N_Y_c_574_n 0.0219971f $X=3.065 $Y=1.635 $X2=0 $Y2=0
cc_260 N_B1_M1020_g N_Y_c_575_n 0.0078351f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_261 N_B1_M1020_g N_Y_c_576_n 0.0120432f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_262 N_B1_M1023_g N_Y_c_576_n 0.0197687f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_263 N_B1_c_274_n N_Y_c_576_n 0.00818622f $X=3.15 $Y=1.8 $X2=0 $Y2=0
cc_264 N_B1_c_275_n N_Y_c_576_n 0.0164207f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_265 N_B1_c_276_n N_Y_c_576_n 0.00361622f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_266 N_B1_c_277_n N_Y_c_576_n 0.00156821f $X=2.84 $Y=1.635 $X2=0 $Y2=0
cc_267 N_B1_c_278_n N_Y_c_576_n 0.00888366f $X=3.065 $Y=1.635 $X2=0 $Y2=0
cc_268 N_B1_M1020_g N_Y_c_577_n 0.0104367f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_269 N_B1_c_277_n N_Y_c_577_n 0.00326139f $X=2.84 $Y=1.635 $X2=0 $Y2=0
cc_270 N_B1_c_278_n N_Y_c_577_n 0.0138023f $X=3.065 $Y=1.635 $X2=0 $Y2=0
cc_271 N_B1_M1023_g N_Y_c_578_n 0.00756015f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_272 N_B1_M1007_g N_Y_c_583_n 4.33202e-19 $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_273 N_B1_c_322_p N_A_119_392#_M1007_d 0.00182529f $X=3.235 $Y=2.035 $X2=0
+ $Y2=0
cc_274 N_B1_c_283_n N_A_119_392#_M1013_s 0.0036552f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_275 N_B1_M1014_g N_A_119_392#_c_722_n 0.00470938f $X=4.385 $Y=2.46 $X2=0
+ $Y2=0
cc_276 N_B1_M1007_g N_A_119_392#_c_724_n 0.0106283f $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_277 N_B1_M1007_g N_A_119_392#_c_725_n 0.0117648f $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_278 N_B1_c_283_n N_A_515_392#_M1012_d 0.00166235f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_279 N_B1_c_277_n N_A_515_392#_c_782_n 0.00298686f $X=2.84 $Y=1.635 $X2=0
+ $Y2=0
cc_280 N_B1_c_278_n N_A_515_392#_c_782_n 0.0103836f $X=3.065 $Y=1.635 $X2=0
+ $Y2=0
cc_281 N_B1_M1007_g N_A_515_392#_c_784_n 0.0138414f $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_282 N_B1_M1014_g N_A_515_392#_c_784_n 0.0139923f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_283 N_B1_c_283_n N_A_515_392#_c_784_n 0.054985f $X=4.105 $Y=2.035 $X2=0 $Y2=0
cc_284 N_B1_c_322_p N_A_515_392#_c_784_n 0.0115915f $X=3.235 $Y=2.035 $X2=0
+ $Y2=0
cc_285 N_B1_c_275_n N_A_515_392#_c_784_n 0.0046953f $X=4.31 $Y=1.615 $X2=0 $Y2=0
cc_286 N_B1_c_276_n N_A_515_392#_c_784_n 3.97349e-19 $X=4.31 $Y=1.615 $X2=0
+ $Y2=0
cc_287 N_B1_c_278_n N_A_515_392#_c_784_n 0.00678712f $X=3.065 $Y=1.635 $X2=0
+ $Y2=0
cc_288 N_B1_M1014_g N_A_515_392#_c_776_n 0.00587661f $X=4.385 $Y=2.46 $X2=0
+ $Y2=0
cc_289 N_B1_c_283_n N_A_515_392#_c_776_n 0.00682866f $X=4.105 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_B1_c_275_n N_A_515_392#_c_776_n 0.00226259f $X=4.31 $Y=1.615 $X2=0
+ $Y2=0
cc_291 N_B1_M1014_g N_A_515_392#_c_779_n 0.00181298f $X=4.385 $Y=2.46 $X2=0
+ $Y2=0
cc_292 N_B1_M1014_g N_VPWR_c_856_n 6.31214e-19 $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_293 N_B1_M1007_g N_VPWR_c_858_n 0.00333926f $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_294 N_B1_M1014_g N_VPWR_c_858_n 0.00519794f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_295 N_B1_M1007_g N_VPWR_c_855_n 0.00427931f $X=2.945 $Y=2.46 $X2=0 $Y2=0
cc_296 N_B1_M1014_g N_VPWR_c_855_n 0.00980729f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_297 N_B1_M1020_g N_VGND_c_928_n 0.00380203f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_298 N_B1_M1020_g N_VGND_c_931_n 0.00434272f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_299 N_B1_M1023_g N_VGND_c_932_n 0.00434272f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_300 N_B1_M1020_g N_VGND_c_934_n 0.00826366f $X=2.89 $Y=0.69 $X2=0 $Y2=0
cc_301 N_B1_M1023_g N_VGND_c_934_n 0.00821465f $X=4.4 $Y=0.69 $X2=0 $Y2=0
cc_302 N_B2_M1009_g N_Y_c_575_n 9.56968e-19 $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_303 N_B2_M1009_g N_Y_c_576_n 0.0158888f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_304 N_B2_c_370_n N_Y_c_576_n 0.0153959f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_305 N_B2_c_371_n N_Y_c_576_n 0.0256597f $X=3.57 $Y=1.425 $X2=0 $Y2=0
cc_306 N_B2_c_372_n N_Y_c_576_n 0.0113491f $X=3.845 $Y=1.34 $X2=0 $Y2=0
cc_307 N_B2_M1009_g N_Y_c_577_n 9.79153e-19 $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_308 N_B2_c_371_n N_Y_c_577_n 0.00116356f $X=3.57 $Y=1.425 $X2=0 $Y2=0
cc_309 N_B2_c_370_n N_Y_c_578_n 9.65066e-19 $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_310 N_B2_M1012_g N_A_119_392#_c_722_n 0.0120973f $X=3.395 $Y=2.46 $X2=0 $Y2=0
cc_311 N_B2_M1013_g N_A_119_392#_c_722_n 0.0140371f $X=3.845 $Y=2.46 $X2=0 $Y2=0
cc_312 N_B2_M1012_g N_A_119_392#_c_725_n 0.00505896f $X=3.395 $Y=2.46 $X2=0
+ $Y2=0
cc_313 N_B2_M1013_g N_A_119_392#_c_725_n 5.34023e-19 $X=3.845 $Y=2.46 $X2=0
+ $Y2=0
cc_314 N_B2_M1012_g N_A_515_392#_c_784_n 0.00975857f $X=3.395 $Y=2.46 $X2=0
+ $Y2=0
cc_315 N_B2_M1013_g N_A_515_392#_c_784_n 0.0102724f $X=3.845 $Y=2.46 $X2=0 $Y2=0
cc_316 N_B2_M1013_g N_A_515_392#_c_776_n 8.9192e-19 $X=3.845 $Y=2.46 $X2=0 $Y2=0
cc_317 N_B2_M1012_g N_VPWR_c_858_n 0.00347303f $X=3.395 $Y=2.46 $X2=0 $Y2=0
cc_318 N_B2_M1013_g N_VPWR_c_858_n 0.00349978f $X=3.845 $Y=2.46 $X2=0 $Y2=0
cc_319 N_B2_M1012_g N_VPWR_c_855_n 0.00428491f $X=3.395 $Y=2.46 $X2=0 $Y2=0
cc_320 N_B2_M1013_g N_VPWR_c_855_n 0.00430421f $X=3.845 $Y=2.46 $X2=0 $Y2=0
cc_321 N_B2_M1009_g N_VGND_c_931_n 0.00316493f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_322 N_B2_c_370_n N_VGND_c_932_n 0.00316493f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_323 N_B2_M1009_g N_VGND_c_934_n 0.00393725f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_324 N_B2_c_370_n N_VGND_c_934_n 0.00393725f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_325 N_B2_M1009_g N_VGND_c_936_n 0.00381881f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_326 N_B2_c_370_n N_VGND_c_936_n 0.00381881f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_327 N_B2_M1009_g N_A_593_74#_c_1030_n 0.00966972f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_328 N_B2_c_370_n N_A_593_74#_c_1030_n 0.00966972f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_329 N_B2_M1009_g N_A_593_74#_c_1028_n 0.00590335f $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_330 N_B2_c_370_n N_A_593_74#_c_1028_n 8.35363e-19 $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_331 N_B2_M1009_g N_A_593_74#_c_1029_n 8.35363e-19 $X=3.32 $Y=0.69 $X2=0 $Y2=0
cc_332 N_B2_c_370_n N_A_593_74#_c_1029_n 0.00590335f $X=3.97 $Y=1.09 $X2=0 $Y2=0
cc_333 N_A1_M1017_g N_A2_M1019_g 0.0360637f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_334 N_A1_c_436_n N_A2_M1019_g 0.00383206f $X=5.03 $Y=1.95 $X2=0 $Y2=0
cc_335 N_A1_c_437_n N_A2_M1019_g 0.0125883f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_336 N_A1_M1005_g N_A2_M1000_g 0.0300052f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_337 N_A1_M1022_g N_A2_M1021_g 0.0282552f $X=6.215 $Y=2.46 $X2=0 $Y2=0
cc_338 N_A1_c_437_n N_A2_M1021_g 0.0138227f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_339 N_A1_c_438_n N_A2_M1021_g 0.00417136f $X=5.97 $Y=1.95 $X2=0 $Y2=0
cc_340 N_A1_M1006_g N_A2_M1001_g 0.0266095f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_341 N_A1_c_437_n A2 0.0244048f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_342 N_A1_c_430_n A2 2.99931e-19 $X=4.85 $Y=1.615 $X2=0 $Y2=0
cc_343 N_A1_c_431_n A2 0.0244979f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_344 N_A1_c_432_n A2 2.19852e-19 $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_345 N_A1_c_433_n A2 0.0204271f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_346 N_A1_c_437_n N_A2_c_521_n 6.34453e-19 $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_347 N_A1_c_430_n N_A2_c_521_n 0.0214942f $X=4.85 $Y=1.615 $X2=0 $Y2=0
cc_348 N_A1_c_431_n N_A2_c_521_n 0.00243494f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_349 N_A1_c_432_n N_A2_c_521_n 0.0282552f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_350 N_A1_c_433_n N_A2_c_521_n 0.00375221f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_351 N_A1_M1005_g N_Y_c_576_n 3.91998e-19 $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_352 N_A1_c_430_n N_Y_c_576_n 6.75574e-19 $X=4.85 $Y=1.615 $X2=0 $Y2=0
cc_353 N_A1_c_431_n N_Y_c_576_n 0.00244567f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_354 N_A1_M1005_g N_Y_c_578_n 0.00279931f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_355 N_A1_M1005_g N_Y_c_579_n 0.0135003f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_356 N_A1_M1006_g N_Y_c_579_n 0.0156502f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_357 N_A1_c_437_n N_Y_c_579_n 0.0110324f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_358 N_A1_c_430_n N_Y_c_579_n 0.00348128f $X=4.85 $Y=1.615 $X2=0 $Y2=0
cc_359 N_A1_c_431_n N_Y_c_579_n 0.0299139f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_360 N_A1_c_432_n N_Y_c_579_n 0.00426984f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_361 N_A1_c_433_n N_Y_c_579_n 0.0444698f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_362 N_A1_M1006_g N_Y_c_580_n 0.00453147f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_363 N_A1_c_437_n N_A_515_392#_M1019_d 0.00165831f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_364 N_A1_M1017_g N_A_515_392#_c_776_n 0.00570833f $X=4.835 $Y=2.46 $X2=0
+ $Y2=0
cc_365 N_A1_c_482_p N_A_515_392#_c_776_n 0.00682866f $X=5.115 $Y=2.035 $X2=0
+ $Y2=0
cc_366 N_A1_c_430_n N_A_515_392#_c_776_n 0.00139157f $X=4.85 $Y=1.615 $X2=0
+ $Y2=0
cc_367 N_A1_c_431_n N_A_515_392#_c_776_n 0.007278f $X=5.03 $Y=1.615 $X2=0 $Y2=0
cc_368 N_A1_M1017_g N_A_515_392#_c_803_n 0.0119461f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_369 N_A1_c_437_n N_A_515_392#_c_803_n 0.0161169f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_370 N_A1_c_482_p N_A_515_392#_c_803_n 0.0103235f $X=5.115 $Y=2.035 $X2=0
+ $Y2=0
cc_371 N_A1_c_431_n N_A_515_392#_c_803_n 0.00473085f $X=5.03 $Y=1.615 $X2=0
+ $Y2=0
cc_372 N_A1_M1022_g N_A_515_392#_c_807_n 0.0117491f $X=6.215 $Y=2.46 $X2=0 $Y2=0
cc_373 N_A1_c_437_n N_A_515_392#_c_807_n 0.0233707f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_374 N_A1_c_433_n N_A_515_392#_c_807_n 0.00600414f $X=6.29 $Y=1.615 $X2=0
+ $Y2=0
cc_375 N_A1_M1022_g N_A_515_392#_c_778_n 0.00589675f $X=6.215 $Y=2.46 $X2=0
+ $Y2=0
cc_376 N_A1_c_437_n N_A_515_392#_c_778_n 0.0115259f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_377 N_A1_c_432_n N_A_515_392#_c_778_n 0.00348818f $X=6.29 $Y=1.615 $X2=0
+ $Y2=0
cc_378 N_A1_c_433_n N_A_515_392#_c_778_n 0.014868f $X=6.29 $Y=1.615 $X2=0 $Y2=0
cc_379 N_A1_M1017_g N_A_515_392#_c_779_n 0.00125921f $X=4.835 $Y=2.46 $X2=0
+ $Y2=0
cc_380 N_A1_c_437_n N_A_515_392#_c_815_n 0.0127071f $X=5.885 $Y=2.035 $X2=0
+ $Y2=0
cc_381 N_A1_M1022_g N_A_515_392#_c_780_n 0.00221423f $X=6.215 $Y=2.46 $X2=0
+ $Y2=0
cc_382 N_A1_c_437_n N_VPWR_M1017_d 5.54118e-19 $X=5.885 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_383 N_A1_c_482_p N_VPWR_M1017_d 0.00196024f $X=5.115 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_384 N_A1_c_437_n N_VPWR_M1021_s 0.00321233f $X=5.885 $Y=2.035 $X2=0 $Y2=0
cc_385 N_A1_M1017_g N_VPWR_c_856_n 0.00849298f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_386 N_A1_M1022_g N_VPWR_c_857_n 0.0105392f $X=6.215 $Y=2.46 $X2=0 $Y2=0
cc_387 N_A1_M1017_g N_VPWR_c_858_n 0.00460063f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_388 N_A1_M1022_g N_VPWR_c_860_n 0.00460063f $X=6.215 $Y=2.46 $X2=0 $Y2=0
cc_389 N_A1_M1017_g N_VPWR_c_855_n 0.00463426f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_390 N_A1_M1022_g N_VPWR_c_855_n 0.00467058f $X=6.215 $Y=2.46 $X2=0 $Y2=0
cc_391 N_A1_M1005_g N_VGND_c_929_n 5.94048e-19 $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_392 N_A1_M1006_g N_VGND_c_929_n 5.48301e-19 $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_393 N_A1_M1005_g N_VGND_c_932_n 0.00439937f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_394 N_A1_M1006_g N_VGND_c_933_n 0.00433834f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_395 N_A1_M1005_g N_VGND_c_934_n 0.00840422f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_396 N_A1_M1006_g N_VGND_c_934_n 0.00824802f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_397 N_A1_M1005_g N_A_981_74#_c_1054_n 0.00450875f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_398 N_A1_M1005_g N_A_981_74#_c_1057_n 0.00192658f $X=4.83 $Y=0.69 $X2=0 $Y2=0
cc_399 N_A1_M1006_g N_A_981_74#_c_1058_n 0.00215008f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_400 N_A1_M1006_g N_A_981_74#_c_1055_n 0.00587363f $X=6.2 $Y=0.69 $X2=0 $Y2=0
cc_401 N_A2_M1000_g N_Y_c_579_n 0.0116566f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_402 N_A2_M1001_g N_Y_c_579_n 0.0127854f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_403 A2 N_Y_c_579_n 0.0244045f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_404 N_A2_c_521_n N_Y_c_579_n 0.00202495f $X=5.77 $Y=1.615 $X2=0 $Y2=0
cc_405 N_A2_M1019_g N_A_515_392#_c_776_n 9.14751e-19 $X=5.315 $Y=2.46 $X2=0
+ $Y2=0
cc_406 N_A2_M1019_g N_A_515_392#_c_803_n 0.0118989f $X=5.315 $Y=2.46 $X2=0 $Y2=0
cc_407 N_A2_M1019_g N_A_515_392#_c_777_n 3.35321e-19 $X=5.315 $Y=2.46 $X2=0
+ $Y2=0
cc_408 N_A2_M1021_g N_A_515_392#_c_777_n 3.35321e-19 $X=5.765 $Y=2.46 $X2=0
+ $Y2=0
cc_409 N_A2_M1021_g N_A_515_392#_c_807_n 0.0117019f $X=5.765 $Y=2.46 $X2=0 $Y2=0
cc_410 N_A2_M1021_g N_A_515_392#_c_778_n 9.37392e-19 $X=5.765 $Y=2.46 $X2=0
+ $Y2=0
cc_411 N_A2_M1019_g N_VPWR_c_856_n 0.00838578f $X=5.315 $Y=2.46 $X2=0 $Y2=0
cc_412 N_A2_M1021_g N_VPWR_c_856_n 4.12401e-19 $X=5.765 $Y=2.46 $X2=0 $Y2=0
cc_413 N_A2_M1019_g N_VPWR_c_857_n 4.12707e-19 $X=5.315 $Y=2.46 $X2=0 $Y2=0
cc_414 N_A2_M1021_g N_VPWR_c_857_n 0.00825058f $X=5.765 $Y=2.46 $X2=0 $Y2=0
cc_415 N_A2_M1019_g N_VPWR_c_859_n 0.00460063f $X=5.315 $Y=2.46 $X2=0 $Y2=0
cc_416 N_A2_M1021_g N_VPWR_c_859_n 0.00460063f $X=5.765 $Y=2.46 $X2=0 $Y2=0
cc_417 N_A2_M1019_g N_VPWR_c_855_n 0.00463365f $X=5.315 $Y=2.46 $X2=0 $Y2=0
cc_418 N_A2_M1021_g N_VPWR_c_855_n 0.00463365f $X=5.765 $Y=2.46 $X2=0 $Y2=0
cc_419 N_A2_M1000_g N_VGND_c_929_n 0.00681232f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_420 N_A2_M1001_g N_VGND_c_929_n 0.0066056f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_421 N_A2_M1000_g N_VGND_c_932_n 0.00398535f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_422 N_A2_M1001_g N_VGND_c_933_n 0.00398535f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_423 N_A2_M1000_g N_VGND_c_934_n 0.00384569f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_424 N_A2_M1001_g N_VGND_c_934_n 0.00383955f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_425 N_A2_M1000_g N_A_981_74#_c_1054_n 0.00227555f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_426 N_A2_M1000_g N_A_981_74#_c_1061_n 0.0119053f $X=5.33 $Y=0.69 $X2=0 $Y2=0
cc_427 N_A2_M1001_g N_A_981_74#_c_1061_n 0.00951514f $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_428 N_A2_M1001_g N_A_981_74#_c_1055_n 2.96277e-19 $X=5.77 $Y=0.69 $X2=0 $Y2=0
cc_429 N_Y_c_591_n N_A_119_392#_M1002_d 0.00319799f $X=1.065 $Y=2.09 $X2=-0.19
+ $Y2=-0.245
cc_430 N_Y_c_596_n N_A_119_392#_M1016_s 0.00332066f $X=1.995 $Y=2.09 $X2=0 $Y2=0
cc_431 N_Y_c_591_n N_A_119_392#_c_726_n 0.0170259f $X=1.065 $Y=2.09 $X2=0 $Y2=0
cc_432 N_Y_M1003_d N_A_119_392#_c_720_n 0.00197722f $X=1.045 $Y=1.96 $X2=0 $Y2=0
cc_433 N_Y_c_673_p N_A_119_392#_c_720_n 0.014157f $X=1.195 $Y=2.57 $X2=0 $Y2=0
cc_434 Y N_A_119_392#_c_721_n 0.00346205f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_435 N_Y_c_596_n N_A_119_392#_c_728_n 0.0170259f $X=1.995 $Y=2.09 $X2=0 $Y2=0
cc_436 N_Y_M1018_s N_A_119_392#_c_724_n 0.00335038f $X=1.975 $Y=1.96 $X2=0 $Y2=0
cc_437 N_Y_c_583_n N_A_119_392#_c_724_n 0.0333411f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_438 N_Y_c_574_n N_A_515_392#_c_782_n 0.00255112f $X=2.38 $Y=2.005 $X2=0 $Y2=0
cc_439 N_Y_c_577_n N_A_515_392#_c_782_n 0.0013185f $X=2.84 $Y=1.005 $X2=0 $Y2=0
cc_440 N_Y_c_583_n N_A_515_392#_c_782_n 0.0232783f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_441 N_Y_c_583_n N_A_515_392#_c_826_n 0.0220282f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_442 N_Y_c_576_n N_A_515_392#_c_776_n 0.00748381f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_443 N_Y_c_579_n N_A_515_392#_c_778_n 0.0044659f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_444 N_Y_c_583_n N_A_515_392#_c_829_n 0.0151272f $X=2.16 $Y=2.17 $X2=0 $Y2=0
cc_445 Y N_VPWR_c_858_n 0.0124046f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_446 Y N_VPWR_c_855_n 0.0102675f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_447 N_Y_c_572_n N_VGND_M1008_d 2.6293e-19 $X=0.17 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_448 N_Y_c_573_n N_VGND_M1008_d 0.00243255f $X=0.255 $Y=0.91 $X2=-0.19
+ $Y2=-0.245
cc_449 N_Y_c_610_n N_VGND_M1008_d 0.00982502f $X=1.09 $Y=0.887 $X2=-0.19
+ $Y2=-0.245
cc_450 N_Y_c_576_n N_VGND_M1009_d 0.00480292f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_451 N_Y_c_573_n N_VGND_c_927_n 0.0122781f $X=0.255 $Y=0.91 $X2=0 $Y2=0
cc_452 N_Y_c_610_n N_VGND_c_927_n 0.0176875f $X=1.09 $Y=0.887 $X2=0 $Y2=0
cc_453 N_Y_c_575_n N_VGND_c_928_n 0.0383948f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_454 N_Y_c_577_n N_VGND_c_928_n 0.00143078f $X=2.84 $Y=1.005 $X2=0 $Y2=0
cc_455 N_Y_c_608_n N_VGND_c_928_n 0.00172463f $X=1.255 $Y=0.865 $X2=0 $Y2=0
cc_456 N_Y_c_575_n N_VGND_c_931_n 0.0145639f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_457 N_Y_c_578_n N_VGND_c_932_n 0.0116636f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_458 N_Y_c_580_n N_VGND_c_933_n 0.0115122f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_459 N_Y_c_573_n N_VGND_c_934_n 0.00175584f $X=0.255 $Y=0.91 $X2=0 $Y2=0
cc_460 N_Y_c_575_n N_VGND_c_934_n 0.0119984f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_461 N_Y_c_578_n N_VGND_c_934_n 0.00959771f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_462 N_Y_c_580_n N_VGND_c_934_n 0.0095288f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_463 N_Y_c_610_n N_VGND_c_934_n 0.00688546f $X=1.09 $Y=0.887 $X2=0 $Y2=0
cc_464 N_Y_c_610_n N_A_137_74#_M1008_s 0.00441403f $X=1.09 $Y=0.887 $X2=-0.19
+ $Y2=-0.245
cc_465 N_Y_M1004_s N_A_137_74#_c_1015_n 0.0016448f $X=1.115 $Y=0.37 $X2=0 $Y2=0
cc_466 N_Y_c_608_n N_A_137_74#_c_1015_n 0.0156706f $X=1.255 $Y=0.865 $X2=0 $Y2=0
cc_467 N_Y_c_610_n N_A_137_74#_c_1015_n 0.0181933f $X=1.09 $Y=0.887 $X2=0 $Y2=0
cc_468 N_Y_c_576_n N_A_593_74#_M1020_d 0.00176461f $X=4.45 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_469 N_Y_c_576_n N_A_593_74#_M1015_s 0.00176461f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_470 N_Y_c_576_n N_A_593_74#_c_1030_n 0.0449815f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_471 N_Y_c_575_n N_A_593_74#_c_1028_n 0.0150645f $X=2.675 $Y=0.515 $X2=0 $Y2=0
cc_472 N_Y_c_576_n N_A_593_74#_c_1028_n 0.0146914f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_473 N_Y_c_576_n N_A_593_74#_c_1029_n 0.0146914f $X=4.45 $Y=1.005 $X2=0 $Y2=0
cc_474 N_Y_c_578_n N_A_593_74#_c_1029_n 0.0145907f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_475 N_Y_c_578_n N_A_981_74#_c_1054_n 0.0164865f $X=4.615 $Y=0.515 $X2=0 $Y2=0
cc_476 N_Y_c_579_n N_A_981_74#_c_1061_n 0.0411874f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_477 N_Y_c_579_n N_A_981_74#_c_1057_n 0.023557f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_478 N_Y_c_579_n N_A_981_74#_c_1058_n 0.0176844f $X=6.32 $Y=1.195 $X2=0 $Y2=0
cc_479 N_Y_c_580_n N_A_981_74#_c_1055_n 0.0158295f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_480 N_A_119_392#_c_724_n N_A_515_392#_M1007_s 0.00434847f $X=3.005 $Y=2.852
+ $X2=-0.19 $Y2=1.66
cc_481 N_A_119_392#_c_722_n N_A_515_392#_M1012_d 0.00177865f $X=4.115 $Y=2.815
+ $X2=0 $Y2=0
cc_482 N_A_119_392#_c_724_n N_A_515_392#_c_826_n 0.0123303f $X=3.005 $Y=2.852
+ $X2=0 $Y2=0
cc_483 N_A_119_392#_M1007_d N_A_515_392#_c_784_n 0.003321f $X=3.035 $Y=1.96
+ $X2=0 $Y2=0
cc_484 N_A_119_392#_M1013_s N_A_515_392#_c_784_n 0.00525856f $X=3.935 $Y=1.96
+ $X2=0 $Y2=0
cc_485 N_A_119_392#_c_722_n N_A_515_392#_c_784_n 0.0516394f $X=4.115 $Y=2.815
+ $X2=0 $Y2=0
cc_486 N_A_119_392#_c_724_n N_A_515_392#_c_784_n 0.0046334f $X=3.005 $Y=2.852
+ $X2=0 $Y2=0
cc_487 N_A_119_392#_c_725_n N_A_515_392#_c_784_n 0.0165186f $X=3.335 $Y=2.852
+ $X2=0 $Y2=0
cc_488 N_A_119_392#_c_722_n N_A_515_392#_c_779_n 0.0141875f $X=4.115 $Y=2.815
+ $X2=0 $Y2=0
cc_489 N_A_119_392#_c_720_n N_VPWR_c_858_n 0.0377252f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_490 N_A_119_392#_c_721_n N_VPWR_c_858_n 0.0234458f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_491 N_A_119_392#_c_722_n N_VPWR_c_858_n 0.0407895f $X=4.115 $Y=2.815 $X2=0
+ $Y2=0
cc_492 N_A_119_392#_c_723_n N_VPWR_c_858_n 0.0234131f $X=1.66 $Y=2.99 $X2=0
+ $Y2=0
cc_493 N_A_119_392#_c_724_n N_VPWR_c_858_n 0.0976566f $X=3.005 $Y=2.852 $X2=0
+ $Y2=0
cc_494 N_A_119_392#_c_720_n N_VPWR_c_855_n 0.0211866f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_495 N_A_119_392#_c_721_n N_VPWR_c_855_n 0.0125551f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_496 N_A_119_392#_c_722_n N_VPWR_c_855_n 0.0339574f $X=4.115 $Y=2.815 $X2=0
+ $Y2=0
cc_497 N_A_119_392#_c_723_n N_VPWR_c_855_n 0.0125504f $X=1.66 $Y=2.99 $X2=0
+ $Y2=0
cc_498 N_A_119_392#_c_724_n N_VPWR_c_855_n 0.0554027f $X=3.005 $Y=2.852 $X2=0
+ $Y2=0
cc_499 N_A_515_392#_c_803_n N_VPWR_M1017_d 0.0039058f $X=5.425 $Y=2.385
+ $X2=-0.19 $Y2=1.66
cc_500 N_A_515_392#_c_807_n N_VPWR_M1021_s 0.00340622f $X=6.275 $Y=2.385 $X2=0
+ $Y2=0
cc_501 N_A_515_392#_c_803_n N_VPWR_c_856_n 0.0191959f $X=5.425 $Y=2.385 $X2=0
+ $Y2=0
cc_502 N_A_515_392#_c_777_n N_VPWR_c_856_n 0.0132968f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_503 N_A_515_392#_c_779_n N_VPWR_c_856_n 0.0126977f $X=4.61 $Y=2.465 $X2=0
+ $Y2=0
cc_504 N_A_515_392#_c_777_n N_VPWR_c_857_n 0.0131308f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_505 N_A_515_392#_c_807_n N_VPWR_c_857_n 0.016789f $X=6.275 $Y=2.385 $X2=0
+ $Y2=0
cc_506 N_A_515_392#_c_780_n N_VPWR_c_857_n 0.0140562f $X=6.44 $Y=2.455 $X2=0
+ $Y2=0
cc_507 N_A_515_392#_c_779_n N_VPWR_c_858_n 0.00950426f $X=4.61 $Y=2.465 $X2=0
+ $Y2=0
cc_508 N_A_515_392#_c_777_n N_VPWR_c_859_n 0.0101844f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_509 N_A_515_392#_c_780_n N_VPWR_c_860_n 0.0129995f $X=6.44 $Y=2.455 $X2=0
+ $Y2=0
cc_510 N_A_515_392#_c_803_n N_VPWR_c_855_n 0.00921423f $X=5.425 $Y=2.385 $X2=0
+ $Y2=0
cc_511 N_A_515_392#_c_777_n N_VPWR_c_855_n 0.00842501f $X=5.54 $Y=2.815 $X2=0
+ $Y2=0
cc_512 N_A_515_392#_c_807_n N_VPWR_c_855_n 0.00911854f $X=6.275 $Y=2.385 $X2=0
+ $Y2=0
cc_513 N_A_515_392#_c_779_n N_VPWR_c_855_n 0.00989327f $X=4.61 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_515_392#_c_780_n N_VPWR_c_855_n 0.012042f $X=6.44 $Y=2.455 $X2=0
+ $Y2=0
cc_515 N_VGND_c_927_n N_A_137_74#_c_1015_n 0.0111115f $X=0.295 $Y=0.49 $X2=0
+ $Y2=0
cc_516 N_VGND_c_928_n N_A_137_74#_c_1015_n 0.0106879f $X=2.115 $Y=0.515 $X2=0
+ $Y2=0
cc_517 N_VGND_c_930_n N_A_137_74#_c_1015_n 0.0460738f $X=1.95 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_934_n N_A_137_74#_c_1015_n 0.0386873f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_M1009_d N_A_593_74#_c_1030_n 0.00883733f $X=3.395 $Y=0.37 $X2=0
+ $Y2=0
cc_520 N_VGND_c_931_n N_A_593_74#_c_1030_n 0.0029521f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_932_n N_A_593_74#_c_1030_n 0.0029521f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_934_n N_A_593_74#_c_1030_n 0.0115024f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_936_n N_A_593_74#_c_1030_n 0.0288883f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_931_n N_A_593_74#_c_1028_n 0.0105866f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_934_n N_A_593_74#_c_1028_n 0.00888607f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_936_n N_A_593_74#_c_1028_n 0.00283955f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_932_n N_A_593_74#_c_1029_n 0.0105866f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_934_n N_A_593_74#_c_1029_n 0.00888607f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_936_n N_A_593_74#_c_1029_n 0.00283955f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_929_n N_A_981_74#_c_1054_n 0.0101711f $X=5.55 $Y=0.515 $X2=0
+ $Y2=0
cc_531 N_VGND_c_932_n N_A_981_74#_c_1054_n 0.0144296f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_934_n N_A_981_74#_c_1054_n 0.0119645f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_M1000_d N_A_981_74#_c_1061_n 0.00353971f $X=5.405 $Y=0.37 $X2=0
+ $Y2=0
cc_534 N_VGND_c_929_n N_A_981_74#_c_1061_n 0.0166493f $X=5.55 $Y=0.515 $X2=0
+ $Y2=0
cc_535 N_VGND_c_934_n N_A_981_74#_c_1061_n 0.0123108f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_929_n N_A_981_74#_c_1055_n 0.0109329f $X=5.55 $Y=0.515 $X2=0
+ $Y2=0
cc_537 N_VGND_c_933_n N_A_981_74#_c_1055_n 0.0118609f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_934_n N_A_981_74#_c_1055_n 0.00912082f $X=6.48 $Y=0 $X2=0 $Y2=0

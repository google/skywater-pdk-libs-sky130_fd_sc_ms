* NGSPICE file created from sky130_fd_sc_ms__dlrbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR RESET_B a_889_92# VPB pshort w=1.12e+06u l=180000u
+  ad=2.18775e+12p pd=1.595e+07u as=3.136e+11p ps=2.8e+06u
M1001 a_608_74# a_27_424# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.4043e+12p ps=1.104e+07u
M1002 a_686_74# a_231_74# a_608_74# VNB nlowvt w=640000u l=150000u
+  ad=3.835e+11p pd=2.53e+06u as=0p ps=0u
M1003 a_231_74# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 a_805_508# a_231_74# a_686_74# VPB pshort w=420000u l=180000u
+  ad=2.121e+11p pd=1.85e+06u as=3.115e+11p ps=2.71e+06u
M1005 VGND RESET_B a_1133_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1006 a_686_74# a_373_74# a_614_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1007 a_231_74# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 VGND D a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 Q_N a_1437_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1010 VGND a_889_92# a_1437_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.925e+11p ps=1.8e+06u
M1011 VPWR a_889_92# a_805_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR D a_27_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 a_889_92# a_686_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_841_118# a_373_74# a_686_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 VGND a_231_74# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 Q a_889_92# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1017 a_1133_74# a_686_74# a_889_92# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 Q a_889_92# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 a_614_392# a_27_424# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_1437_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 VPWR a_889_92# a_1437_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1022 VPWR a_231_74# a_373_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=3.704e+11p ps=2.85e+06u
M1023 VGND a_889_92# a_841_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__dlxbn_2.pxi.spice
* Created: Wed Sep  2 12:06:10 2020
* 
x_PM_SKY130_FD_SC_MS__DLXBN_2%D N_D_M1018_g N_D_M1020_g D N_D_c_169_n
+ PM_SKY130_FD_SC_MS__DLXBN_2%D
x_PM_SKY130_FD_SC_MS__DLXBN_2%GATE_N N_GATE_N_M1019_g N_GATE_N_M1001_g GATE_N
+ N_GATE_N_c_203_n N_GATE_N_c_206_n PM_SKY130_FD_SC_MS__DLXBN_2%GATE_N
x_PM_SKY130_FD_SC_MS__DLXBN_2%A_232_98# N_A_232_98#_M1001_d N_A_232_98#_M1019_d
+ N_A_232_98#_c_239_n N_A_232_98#_M1004_g N_A_232_98#_c_253_n
+ N_A_232_98#_M1023_g N_A_232_98#_c_241_n N_A_232_98#_M1013_g
+ N_A_232_98#_c_242_n N_A_232_98#_c_243_n N_A_232_98#_c_244_n
+ N_A_232_98#_M1006_g N_A_232_98#_c_245_n N_A_232_98#_c_246_n
+ N_A_232_98#_c_247_n N_A_232_98#_c_256_n N_A_232_98#_c_248_n
+ N_A_232_98#_c_258_n N_A_232_98#_c_259_n N_A_232_98#_c_249_n
+ N_A_232_98#_c_260_n N_A_232_98#_c_250_n N_A_232_98#_c_251_n
+ N_A_232_98#_c_252_n PM_SKY130_FD_SC_MS__DLXBN_2%A_232_98#
x_PM_SKY130_FD_SC_MS__DLXBN_2%A_27_136# N_A_27_136#_M1018_s N_A_27_136#_M1020_s
+ N_A_27_136#_M1011_g N_A_27_136#_M1012_g N_A_27_136#_c_389_n
+ N_A_27_136#_c_390_n N_A_27_136#_c_391_n N_A_27_136#_c_392_n
+ N_A_27_136#_c_393_n N_A_27_136#_c_394_n N_A_27_136#_c_397_n
+ N_A_27_136#_c_395_n PM_SKY130_FD_SC_MS__DLXBN_2%A_27_136#
x_PM_SKY130_FD_SC_MS__DLXBN_2%A_343_74# N_A_343_74#_M1004_s N_A_343_74#_M1023_s
+ N_A_343_74#_M1017_g N_A_343_74#_c_466_n N_A_343_74#_M1025_g
+ N_A_343_74#_c_467_n N_A_343_74#_c_476_n N_A_343_74#_c_468_n
+ N_A_343_74#_c_478_n N_A_343_74#_c_469_n N_A_343_74#_c_470_n
+ N_A_343_74#_c_471_n N_A_343_74#_c_479_n N_A_343_74#_c_472_n
+ N_A_343_74#_c_473_n N_A_343_74#_c_474_n PM_SKY130_FD_SC_MS__DLXBN_2%A_343_74#
x_PM_SKY130_FD_SC_MS__DLXBN_2%A_887_270# N_A_887_270#_M1015_d
+ N_A_887_270#_M1009_d N_A_887_270#_M1021_g N_A_887_270#_M1022_g
+ N_A_887_270#_M1002_g N_A_887_270#_M1000_g N_A_887_270#_M1008_g
+ N_A_887_270#_M1024_g N_A_887_270#_M1016_g N_A_887_270#_M1010_g
+ N_A_887_270#_c_593_n N_A_887_270#_c_583_n N_A_887_270#_c_595_n
+ N_A_887_270#_c_596_n N_A_887_270#_c_597_n N_A_887_270#_c_598_n
+ N_A_887_270#_c_584_n N_A_887_270#_c_600_n N_A_887_270#_c_585_n
+ N_A_887_270#_c_586_n N_A_887_270#_c_587_n N_A_887_270#_c_602_n
+ N_A_887_270#_c_603_n N_A_887_270#_c_701_p N_A_887_270#_c_588_n
+ PM_SKY130_FD_SC_MS__DLXBN_2%A_887_270#
x_PM_SKY130_FD_SC_MS__DLXBN_2%A_647_79# N_A_647_79#_M1013_d N_A_647_79#_M1017_d
+ N_A_647_79#_M1015_g N_A_647_79#_M1009_g N_A_647_79#_c_750_n
+ N_A_647_79#_c_741_n N_A_647_79#_c_742_n N_A_647_79#_c_743_n
+ N_A_647_79#_c_744_n N_A_647_79#_c_745_n N_A_647_79#_c_763_n
+ N_A_647_79#_c_746_n PM_SKY130_FD_SC_MS__DLXBN_2%A_647_79#
x_PM_SKY130_FD_SC_MS__DLXBN_2%A_1442_94# N_A_1442_94#_M1016_d
+ N_A_1442_94#_M1010_d N_A_1442_94#_M1003_g N_A_1442_94#_M1007_g
+ N_A_1442_94#_c_831_n N_A_1442_94#_M1005_g N_A_1442_94#_M1014_g
+ N_A_1442_94#_c_834_n N_A_1442_94#_c_835_n N_A_1442_94#_c_836_n
+ N_A_1442_94#_c_841_n N_A_1442_94#_c_861_p N_A_1442_94#_c_837_n
+ N_A_1442_94#_c_838_n PM_SKY130_FD_SC_MS__DLXBN_2%A_1442_94#
x_PM_SKY130_FD_SC_MS__DLXBN_2%VPWR N_VPWR_M1020_d N_VPWR_M1023_d N_VPWR_M1021_d
+ N_VPWR_M1000_d N_VPWR_M1024_d N_VPWR_M1003_s N_VPWR_M1005_s N_VPWR_c_895_n
+ N_VPWR_c_896_n N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_900_n
+ N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n
+ N_VPWR_c_906_n VPWR N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n
+ N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n N_VPWR_c_914_n
+ N_VPWR_c_894_n PM_SKY130_FD_SC_MS__DLXBN_2%VPWR
x_PM_SKY130_FD_SC_MS__DLXBN_2%Q N_Q_M1002_d N_Q_M1000_s N_Q_c_998_n N_Q_c_999_n
+ N_Q_c_995_n N_Q_c_996_n Q Q PM_SKY130_FD_SC_MS__DLXBN_2%Q
x_PM_SKY130_FD_SC_MS__DLXBN_2%Q_N N_Q_N_M1007_d N_Q_N_M1003_d N_Q_N_c_1039_n
+ N_Q_N_c_1040_n Q_N Q_N Q_N Q_N N_Q_N_c_1041_n PM_SKY130_FD_SC_MS__DLXBN_2%Q_N
x_PM_SKY130_FD_SC_MS__DLXBN_2%VGND N_VGND_M1018_d N_VGND_M1004_d N_VGND_M1022_d
+ N_VGND_M1002_s N_VGND_M1008_s N_VGND_M1007_s N_VGND_M1014_s N_VGND_c_1063_n
+ N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n N_VGND_c_1067_n
+ N_VGND_c_1068_n N_VGND_c_1069_n N_VGND_c_1070_n N_VGND_c_1071_n
+ N_VGND_c_1072_n N_VGND_c_1073_n N_VGND_c_1074_n N_VGND_c_1075_n VGND
+ N_VGND_c_1076_n N_VGND_c_1077_n N_VGND_c_1078_n N_VGND_c_1079_n
+ N_VGND_c_1080_n N_VGND_c_1081_n PM_SKY130_FD_SC_MS__DLXBN_2%VGND
cc_1 VNB N_D_M1018_g 0.0287808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_2 VNB D 0.00360823f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_c_169_n 0.0259122f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_4 VNB N_GATE_N_M1001_g 0.039987f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.54
cc_5 VNB N_GATE_N_c_203_n 0.00726573f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_6 VNB N_A_232_98#_c_239_n 0.0122688f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.54
cc_7 VNB N_A_232_98#_M1004_g 0.0264819f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.615
cc_8 VNB N_A_232_98#_c_241_n 0.0136955f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_9 VNB N_A_232_98#_c_242_n 0.0395632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_232_98#_c_243_n 0.00597718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_232_98#_c_244_n 0.0118988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_232_98#_c_245_n 0.00862749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_232_98#_c_246_n 0.0129672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_232_98#_c_247_n 0.00460145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_232_98#_c_248_n 0.00230542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_232_98#_c_249_n 0.0105749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_232_98#_c_250_n 0.0306934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_98#_c_251_n 0.00196916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_232_98#_c_252_n 0.0414802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_136#_M1011_g 0.00637675f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_21 VNB N_A_27_136#_M1012_g 0.0211101f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_22 VNB N_A_27_136#_c_389_n 0.0126258f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_23 VNB N_A_27_136#_c_390_n 0.00888898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_136#_c_391_n 0.0114703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_136#_c_392_n 0.00142827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_136#_c_393_n 0.033354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_136#_c_394_n 0.0128373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_136#_c_395_n 0.0193092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_343_74#_c_466_n 0.0443862f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_30 VNB N_A_343_74#_c_467_n 0.00179953f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_31 VNB N_A_343_74#_c_468_n 0.00446714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_343_74#_c_469_n 0.00242174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_343_74#_c_470_n 0.00692449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_343_74#_c_471_n 0.0500834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_343_74#_c_472_n 0.00381535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_343_74#_c_473_n 0.0161126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_343_74#_c_474_n 0.00455507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_887_270#_M1022_g 0.0300984f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_39 VNB N_A_887_270#_M1002_g 0.0244965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_887_270#_M1000_g 0.00187765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_887_270#_M1008_g 0.0227093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_887_270#_M1024_g 0.00159345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_887_270#_M1016_g 0.0242938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_887_270#_M1010_g 0.00158006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_887_270#_c_583_n 0.0276879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_887_270#_c_584_n 0.0151601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_887_270#_c_585_n 0.00159323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_887_270#_c_586_n 4.70257e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_887_270#_c_587_n 0.0112925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_887_270#_c_588_n 0.0733926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_647_79#_M1009_g 0.00687504f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_52 VNB N_A_647_79#_c_741_n 0.00377565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_647_79#_c_742_n 0.0120605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_647_79#_c_743_n 0.00476855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_647_79#_c_744_n 0.00210366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_647_79#_c_745_n 0.0349638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_647_79#_c_746_n 0.0205599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1442_94#_M1003_g 5.87138e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_59 VNB N_A_1442_94#_M1007_g 0.0251049f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_60 VNB N_A_1442_94#_c_831_n 0.0527129f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.78
cc_61 VNB N_A_1442_94#_M1005_g 9.14676e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1442_94#_M1014_g 0.0292907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1442_94#_c_834_n 0.0664837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1442_94#_c_835_n 0.0078387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1442_94#_c_836_n 0.00449706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1442_94#_c_837_n 0.00162453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1442_94#_c_838_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VPWR_c_894_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_995_n 0.00211954f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_70 VNB N_Q_c_996_n 0.00341266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB Q 0.00492273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_Q_N_c_1039_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_73 VNB N_Q_N_c_1040_n 0.00238514f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_74 VNB N_Q_N_c_1041_n 0.00367433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1063_n 0.0108989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1064_n 0.00557196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1065_n 0.0163546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1066_n 0.0214178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1067_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1068_n 0.050535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1069_n 0.0509137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1070_n 0.0502315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1071_n 0.00740538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1072_n 0.0220478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1073_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1074_n 0.0168757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1075_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1076_n 0.0194574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1077_n 0.0213793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1078_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1079_n 0.023189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1080_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1081_n 0.511181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VPB N_D_M1020_g 0.0385062f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.54
cc_95 VPB D 0.0015504f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_96 VPB N_D_c_169_n 0.0152032f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_97 VPB N_GATE_N_M1019_g 0.0268663f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.955
cc_98 VPB N_GATE_N_c_203_n 0.0276884f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_99 VPB N_GATE_N_c_206_n 0.00330344f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_100 VPB N_A_232_98#_c_253_n 0.0266405f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.78
cc_101 VPB N_A_232_98#_M1006_g 0.0271639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_232_98#_c_246_n 0.00822477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_232_98#_c_256_n 0.0107841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_232_98#_c_248_n 0.0140995f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_232_98#_c_258_n 0.0296065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_232_98#_c_259_n 0.00354838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_232_98#_c_260_n 0.00701033f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_232_98#_c_250_n 0.0184768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_232_98#_c_251_n 6.7826e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_136#_M1011_g 0.0299183f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_111 VPB N_A_27_136#_c_397_n 0.0441474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_136#_c_395_n 0.0214398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_343_74#_M1017_g 0.0265628f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_114 VPB N_A_343_74#_c_476_n 0.00329195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_343_74#_c_468_n 6.37444e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_343_74#_c_478_n 0.0230163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_343_74#_c_479_n 0.00392418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_343_74#_c_472_n 0.00357223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_343_74#_c_473_n 0.0136449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_887_270#_M1021_g 0.0330344f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_121 VPB N_A_887_270#_M1000_g 0.0256956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_887_270#_M1024_g 0.0222385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_887_270#_M1010_g 0.0347837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_887_270#_c_593_n 4.61567e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_887_270#_c_583_n 0.00602384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_887_270#_c_595_n 0.00456729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_887_270#_c_596_n 0.00319544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_887_270#_c_597_n 0.00492787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_887_270#_c_598_n 0.0107396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_887_270#_c_584_n 0.0013859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_887_270#_c_600_n 0.0130362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_887_270#_c_586_n 0.00295505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_887_270#_c_602_n 0.00954478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_887_270#_c_603_n 5.97334e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_647_79#_M1009_g 0.0274363f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_136 VPB N_A_647_79#_c_741_n 0.00405049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_1442_94#_M1003_g 0.0250694f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_138 VPB N_A_1442_94#_M1005_g 0.0280436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1442_94#_c_841_n 0.0156401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_895_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_896_n 0.012439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_897_n 0.0316603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_898_n 0.00548364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_899_n 0.0057229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_900_n 0.0211595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_901_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_902_n 0.0645583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_903_n 0.0627859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_904_n 0.00786036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_905_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_906_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_907_n 0.0412238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_908_n 0.0224872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_909_n 0.0207632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_910_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_911_n 0.0261175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_912_n 0.00612764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_913_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_914_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_894_n 0.137463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_Q_c_998_n 3.97757e-19 $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.54
cc_162 VPB N_Q_c_999_n 0.0022119f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_163 VPB Q 0.00138605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB Q_N 0.0034565f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.45
cc_165 VPB N_Q_N_c_1041_n 0.00288708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 N_D_M1020_g N_GATE_N_M1019_g 0.014313f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_167 N_D_M1018_g N_GATE_N_M1001_g 0.0235236f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_168 D N_GATE_N_M1001_g 0.0016953f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_169 N_D_c_169_n N_GATE_N_M1001_g 0.00900297f $X=0.605 $Y=1.615 $X2=0 $Y2=0
cc_170 N_D_M1020_g N_GATE_N_c_203_n 0.00791719f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_171 D N_GATE_N_c_203_n 0.00124643f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_172 N_D_c_169_n N_GATE_N_c_203_n 0.009114f $X=0.605 $Y=1.615 $X2=0 $Y2=0
cc_173 N_D_M1020_g N_GATE_N_c_206_n 0.00425511f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_174 D N_GATE_N_c_206_n 0.00674868f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_175 N_D_M1018_g N_A_232_98#_c_247_n 0.00153513f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_176 D N_A_232_98#_c_248_n 0.00516007f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_177 N_D_M1018_g N_A_232_98#_c_249_n 8.44735e-19 $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_178 D N_A_232_98#_c_249_n 0.00386002f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_179 N_D_M1018_g N_A_27_136#_c_389_n 0.00695111f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_180 N_D_M1018_g N_A_27_136#_c_390_n 0.0118249f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_181 N_D_M1018_g N_A_27_136#_c_391_n 0.00418997f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_182 N_D_M1018_g N_A_27_136#_c_394_n 0.00679591f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_183 N_D_M1020_g N_A_27_136#_c_397_n 0.0178136f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_184 N_D_c_169_n N_A_27_136#_c_397_n 9.89549e-19 $X=0.605 $Y=1.615 $X2=0 $Y2=0
cc_185 N_D_M1018_g N_A_27_136#_c_395_n 0.012924f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_186 N_D_M1020_g N_A_27_136#_c_395_n 0.00883162f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_187 D N_A_27_136#_c_395_n 0.0250154f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_188 N_D_M1020_g N_VPWR_c_895_n 0.0161576f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_189 D N_VPWR_c_895_n 0.00451046f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_190 N_D_c_169_n N_VPWR_c_895_n 0.00138384f $X=0.605 $Y=1.615 $X2=0 $Y2=0
cc_191 N_D_M1020_g N_VPWR_c_911_n 0.00460063f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_192 N_D_M1020_g N_VPWR_c_894_n 0.00912557f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_193 N_D_M1018_g N_VGND_c_1076_n 0.00297615f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_194 N_D_M1018_g N_VGND_c_1081_n 0.00454494f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_195 N_GATE_N_c_206_n N_A_232_98#_M1019_d 0.00117007f $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_196 N_GATE_N_M1001_g N_A_232_98#_c_247_n 0.00801187f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_197 N_GATE_N_M1019_g N_A_232_98#_c_256_n 0.00589806f $X=1.09 $Y=2.54 $X2=0
+ $Y2=0
cc_198 N_GATE_N_M1019_g N_A_232_98#_c_248_n 0.0044318f $X=1.09 $Y=2.54 $X2=0
+ $Y2=0
cc_199 N_GATE_N_M1001_g N_A_232_98#_c_248_n 0.00134619f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_200 N_GATE_N_c_203_n N_A_232_98#_c_248_n 0.00771834f $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_201 N_GATE_N_c_206_n N_A_232_98#_c_248_n 0.0349338f $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_202 N_GATE_N_M1001_g N_A_232_98#_c_249_n 0.00964542f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_203 N_GATE_N_c_203_n N_A_232_98#_c_249_n 0.00389431f $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_204 N_GATE_N_c_206_n N_A_232_98#_c_249_n 0.014229f $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_205 N_GATE_N_M1019_g N_A_232_98#_c_260_n 0.00326002f $X=1.09 $Y=2.54 $X2=0
+ $Y2=0
cc_206 N_GATE_N_c_203_n N_A_232_98#_c_260_n 5.25096e-19 $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_207 N_GATE_N_c_206_n N_A_232_98#_c_260_n 0.00844358f $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_208 N_GATE_N_M1001_g N_A_232_98#_c_252_n 0.0092413f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_209 N_GATE_N_M1001_g N_A_27_136#_c_389_n 0.00225232f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_210 N_GATE_N_M1001_g N_A_27_136#_c_390_n 0.0176665f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_211 N_GATE_N_c_206_n N_A_27_136#_c_397_n 7.06413e-19 $X=1.15 $Y=1.795 $X2=0
+ $Y2=0
cc_212 N_GATE_N_M1019_g N_VPWR_c_895_n 0.00345319f $X=1.09 $Y=2.54 $X2=0 $Y2=0
cc_213 N_GATE_N_M1019_g N_VPWR_c_907_n 0.005209f $X=1.09 $Y=2.54 $X2=0 $Y2=0
cc_214 N_GATE_N_M1019_g N_VPWR_c_894_n 0.00982678f $X=1.09 $Y=2.54 $X2=0 $Y2=0
cc_215 N_GATE_N_M1001_g N_VGND_c_1069_n 0.00374721f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_216 N_GATE_N_M1001_g N_VGND_c_1079_n 0.00210264f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_217 N_GATE_N_M1001_g N_VGND_c_1081_n 0.00508379f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_218 N_A_232_98#_c_253_n N_A_27_136#_M1011_g 0.0356864f $X=2.215 $Y=1.88 $X2=0
+ $Y2=0
cc_219 N_A_232_98#_c_246_n N_A_27_136#_M1011_g 0.00755691f $X=2.215 $Y=1.79
+ $X2=0 $Y2=0
cc_220 N_A_232_98#_c_258_n N_A_27_136#_M1011_g 0.0150769f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_221 N_A_232_98#_M1004_g N_A_27_136#_M1012_g 0.0208763f $X=2.155 $Y=0.74 $X2=0
+ $Y2=0
cc_222 N_A_232_98#_c_241_n N_A_27_136#_M1012_g 0.0251774f $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_223 N_A_232_98#_M1001_d N_A_27_136#_c_390_n 0.00711247f $X=1.16 $Y=0.49 $X2=0
+ $Y2=0
cc_224 N_A_232_98#_M1004_g N_A_27_136#_c_390_n 0.0143931f $X=2.155 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_232_98#_c_247_n N_A_27_136#_c_390_n 0.0207561f $X=1.3 $Y=1.085 $X2=0
+ $Y2=0
cc_226 N_A_232_98#_c_249_n N_A_27_136#_c_390_n 0.00787715f $X=1.72 $Y=1.425
+ $X2=0 $Y2=0
cc_227 N_A_232_98#_c_252_n N_A_27_136#_c_390_n 0.00282316f $X=1.72 $Y=1.335
+ $X2=0 $Y2=0
cc_228 N_A_232_98#_M1004_g N_A_27_136#_c_392_n 0.00611624f $X=2.155 $Y=0.74
+ $X2=0 $Y2=0
cc_229 N_A_232_98#_c_241_n N_A_27_136#_c_392_n 5.65676e-19 $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_230 N_A_232_98#_c_245_n N_A_27_136#_c_392_n 0.0010854f $X=2.177 $Y=1.335
+ $X2=0 $Y2=0
cc_231 N_A_232_98#_M1004_g N_A_27_136#_c_393_n 0.00156579f $X=2.155 $Y=0.74
+ $X2=0 $Y2=0
cc_232 N_A_232_98#_c_243_n N_A_27_136#_c_393_n 0.0251774f $X=3.235 $Y=1.185
+ $X2=0 $Y2=0
cc_233 N_A_232_98#_c_245_n N_A_27_136#_c_393_n 0.0152915f $X=2.177 $Y=1.335
+ $X2=0 $Y2=0
cc_234 N_A_232_98#_c_258_n N_A_343_74#_M1023_s 0.00751229f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_235 N_A_232_98#_M1006_g N_A_343_74#_M1017_g 0.00457063f $X=3.995 $Y=2.17
+ $X2=0 $Y2=0
cc_236 N_A_232_98#_c_258_n N_A_343_74#_M1017_g 0.0161603f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_237 N_A_232_98#_c_242_n N_A_343_74#_c_466_n 0.00302518f $X=3.655 $Y=1.185
+ $X2=0 $Y2=0
cc_238 N_A_232_98#_c_250_n N_A_343_74#_c_466_n 0.00755032f $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_239 N_A_232_98#_M1004_g N_A_343_74#_c_467_n 0.00926159f $X=2.155 $Y=0.74
+ $X2=0 $Y2=0
cc_240 N_A_232_98#_c_247_n N_A_343_74#_c_467_n 0.0117856f $X=1.3 $Y=1.085 $X2=0
+ $Y2=0
cc_241 N_A_232_98#_c_249_n N_A_343_74#_c_467_n 0.0138199f $X=1.72 $Y=1.425 $X2=0
+ $Y2=0
cc_242 N_A_232_98#_c_252_n N_A_343_74#_c_467_n 0.0080401f $X=1.72 $Y=1.335 $X2=0
+ $Y2=0
cc_243 N_A_232_98#_c_253_n N_A_343_74#_c_476_n 0.00888376f $X=2.215 $Y=1.88
+ $X2=0 $Y2=0
cc_244 N_A_232_98#_c_248_n N_A_343_74#_c_476_n 0.0269151f $X=1.57 $Y=2.32 $X2=0
+ $Y2=0
cc_245 N_A_232_98#_c_258_n N_A_343_74#_c_476_n 0.0214834f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_246 N_A_232_98#_c_239_n N_A_343_74#_c_468_n 0.0033888f $X=2.08 $Y=1.335 $X2=0
+ $Y2=0
cc_247 N_A_232_98#_M1004_g N_A_343_74#_c_468_n 0.00594454f $X=2.155 $Y=0.74
+ $X2=0 $Y2=0
cc_248 N_A_232_98#_c_245_n N_A_343_74#_c_468_n 0.00443569f $X=2.177 $Y=1.335
+ $X2=0 $Y2=0
cc_249 N_A_232_98#_c_246_n N_A_343_74#_c_468_n 0.00896731f $X=2.215 $Y=1.79
+ $X2=0 $Y2=0
cc_250 N_A_232_98#_c_247_n N_A_343_74#_c_468_n 0.00534234f $X=1.3 $Y=1.085 $X2=0
+ $Y2=0
cc_251 N_A_232_98#_c_248_n N_A_343_74#_c_468_n 0.00743655f $X=1.57 $Y=2.32 $X2=0
+ $Y2=0
cc_252 N_A_232_98#_c_249_n N_A_343_74#_c_468_n 0.0204605f $X=1.72 $Y=1.425 $X2=0
+ $Y2=0
cc_253 N_A_232_98#_c_252_n N_A_343_74#_c_468_n 8.96662e-19 $X=1.72 $Y=1.335
+ $X2=0 $Y2=0
cc_254 N_A_232_98#_c_253_n N_A_343_74#_c_478_n 0.00436771f $X=2.215 $Y=1.88
+ $X2=0 $Y2=0
cc_255 N_A_232_98#_c_246_n N_A_343_74#_c_478_n 0.00338494f $X=2.215 $Y=1.79
+ $X2=0 $Y2=0
cc_256 N_A_232_98#_c_258_n N_A_343_74#_c_478_n 0.0222768f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_257 N_A_232_98#_c_241_n N_A_343_74#_c_469_n 0.00467657f $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_258 N_A_232_98#_c_241_n N_A_343_74#_c_470_n 0.00745016f $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_259 N_A_232_98#_c_242_n N_A_343_74#_c_470_n 0.00261047f $X=3.655 $Y=1.185
+ $X2=0 $Y2=0
cc_260 N_A_232_98#_c_241_n N_A_343_74#_c_471_n 0.00781125f $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_261 N_A_232_98#_c_242_n N_A_343_74#_c_471_n 0.0027429f $X=3.655 $Y=1.185
+ $X2=0 $Y2=0
cc_262 N_A_232_98#_c_239_n N_A_343_74#_c_479_n 0.00365223f $X=2.08 $Y=1.335
+ $X2=0 $Y2=0
cc_263 N_A_232_98#_c_253_n N_A_343_74#_c_479_n 0.00452394f $X=2.215 $Y=1.88
+ $X2=0 $Y2=0
cc_264 N_A_232_98#_c_246_n N_A_343_74#_c_479_n 0.00233389f $X=2.215 $Y=1.79
+ $X2=0 $Y2=0
cc_265 N_A_232_98#_c_248_n N_A_343_74#_c_479_n 0.014358f $X=1.57 $Y=2.32 $X2=0
+ $Y2=0
cc_266 N_A_232_98#_c_258_n N_A_343_74#_c_479_n 0.00216797f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_267 N_A_232_98#_c_249_n N_A_343_74#_c_479_n 0.00456809f $X=1.72 $Y=1.425
+ $X2=0 $Y2=0
cc_268 N_A_232_98#_c_252_n N_A_343_74#_c_479_n 0.00148506f $X=1.72 $Y=1.335
+ $X2=0 $Y2=0
cc_269 N_A_232_98#_c_243_n N_A_343_74#_c_472_n 0.00128368f $X=3.235 $Y=1.185
+ $X2=0 $Y2=0
cc_270 N_A_232_98#_c_258_n N_A_343_74#_c_472_n 0.00609329f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_271 N_A_232_98#_c_250_n N_A_343_74#_c_472_n 2.95224e-19 $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_272 N_A_232_98#_c_243_n N_A_343_74#_c_473_n 0.018811f $X=3.235 $Y=1.185 $X2=0
+ $Y2=0
cc_273 N_A_232_98#_M1006_g N_A_343_74#_c_473_n 7.53672e-19 $X=3.995 $Y=2.17
+ $X2=0 $Y2=0
cc_274 N_A_232_98#_c_250_n N_A_343_74#_c_473_n 0.0126885f $X=4.06 $Y=1.585 $X2=0
+ $Y2=0
cc_275 N_A_232_98#_c_241_n N_A_343_74#_c_474_n 0.0190136f $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_276 N_A_232_98#_c_243_n N_A_343_74#_c_474_n 0.00607852f $X=3.235 $Y=1.185
+ $X2=0 $Y2=0
cc_277 N_A_232_98#_c_244_n N_A_343_74#_c_474_n 0.00104113f $X=3.73 $Y=1.42 $X2=0
+ $Y2=0
cc_278 N_A_232_98#_M1006_g N_A_887_270#_M1021_g 0.0204185f $X=3.995 $Y=2.17
+ $X2=0 $Y2=0
cc_279 N_A_232_98#_c_258_n N_A_887_270#_M1021_g 0.0013122f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_280 N_A_232_98#_c_259_n N_A_887_270#_M1021_g 0.00774455f $X=4.19 $Y=2.39
+ $X2=0 $Y2=0
cc_281 N_A_232_98#_c_242_n N_A_887_270#_M1022_g 0.00397576f $X=3.655 $Y=1.185
+ $X2=0 $Y2=0
cc_282 N_A_232_98#_c_244_n N_A_887_270#_c_593_n 3.09175e-19 $X=3.73 $Y=1.42
+ $X2=0 $Y2=0
cc_283 N_A_232_98#_c_250_n N_A_887_270#_c_593_n 3.27874e-19 $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_284 N_A_232_98#_c_251_n N_A_887_270#_c_593_n 0.0239718f $X=4.19 $Y=1.585
+ $X2=0 $Y2=0
cc_285 N_A_232_98#_c_244_n N_A_887_270#_c_583_n 0.00147634f $X=3.73 $Y=1.42
+ $X2=0 $Y2=0
cc_286 N_A_232_98#_c_250_n N_A_887_270#_c_583_n 0.0205099f $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_287 N_A_232_98#_c_251_n N_A_887_270#_c_583_n 0.001888f $X=4.19 $Y=1.585 $X2=0
+ $Y2=0
cc_288 N_A_232_98#_c_259_n N_A_887_270#_c_596_n 0.0111881f $X=4.19 $Y=2.39 $X2=0
+ $Y2=0
cc_289 N_A_232_98#_c_251_n N_A_887_270#_c_596_n 0.00247167f $X=4.19 $Y=1.585
+ $X2=0 $Y2=0
cc_290 N_A_232_98#_c_258_n N_A_647_79#_M1017_d 0.00629f $X=4.105 $Y=2.475 $X2=0
+ $Y2=0
cc_291 N_A_232_98#_c_258_n N_A_647_79#_c_750_n 0.0450916f $X=4.105 $Y=2.475
+ $X2=0 $Y2=0
cc_292 N_A_232_98#_c_242_n N_A_647_79#_c_741_n 0.00785202f $X=3.655 $Y=1.185
+ $X2=0 $Y2=0
cc_293 N_A_232_98#_c_244_n N_A_647_79#_c_741_n 0.00951903f $X=3.73 $Y=1.42 $X2=0
+ $Y2=0
cc_294 N_A_232_98#_M1006_g N_A_647_79#_c_741_n 0.0027097f $X=3.995 $Y=2.17 $X2=0
+ $Y2=0
cc_295 N_A_232_98#_c_259_n N_A_647_79#_c_741_n 0.0108171f $X=4.19 $Y=2.39 $X2=0
+ $Y2=0
cc_296 N_A_232_98#_c_250_n N_A_647_79#_c_741_n 0.0104544f $X=4.06 $Y=1.585 $X2=0
+ $Y2=0
cc_297 N_A_232_98#_c_251_n N_A_647_79#_c_741_n 0.0238146f $X=4.19 $Y=1.585 $X2=0
+ $Y2=0
cc_298 N_A_232_98#_c_250_n N_A_647_79#_c_742_n 0.00138087f $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_299 N_A_232_98#_c_251_n N_A_647_79#_c_742_n 0.0122748f $X=4.19 $Y=1.585 $X2=0
+ $Y2=0
cc_300 N_A_232_98#_c_241_n N_A_647_79#_c_743_n 0.0080375f $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_301 N_A_232_98#_c_242_n N_A_647_79#_c_743_n 0.0205903f $X=3.655 $Y=1.185
+ $X2=0 $Y2=0
cc_302 N_A_232_98#_c_250_n N_A_647_79#_c_743_n 0.00754817f $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_303 N_A_232_98#_c_251_n N_A_647_79#_c_743_n 0.0112164f $X=4.19 $Y=1.585 $X2=0
+ $Y2=0
cc_304 N_A_232_98#_M1006_g N_A_647_79#_c_763_n 0.00284565f $X=3.995 $Y=2.17
+ $X2=0 $Y2=0
cc_305 N_A_232_98#_c_250_n N_A_647_79#_c_763_n 0.00552112f $X=4.06 $Y=1.585
+ $X2=0 $Y2=0
cc_306 N_A_232_98#_c_251_n N_A_647_79#_c_763_n 0.00157703f $X=4.19 $Y=1.585
+ $X2=0 $Y2=0
cc_307 N_A_232_98#_c_258_n N_VPWR_M1023_d 0.00691066f $X=4.105 $Y=2.475 $X2=0
+ $Y2=0
cc_308 N_A_232_98#_c_256_n N_VPWR_c_895_n 0.0165862f $X=1.317 $Y=2.56 $X2=0
+ $Y2=0
cc_309 N_A_232_98#_c_253_n N_VPWR_c_896_n 0.00403165f $X=2.215 $Y=1.88 $X2=0
+ $Y2=0
cc_310 N_A_232_98#_c_258_n N_VPWR_c_896_n 0.0211657f $X=4.105 $Y=2.475 $X2=0
+ $Y2=0
cc_311 N_A_232_98#_c_258_n N_VPWR_c_897_n 0.00848257f $X=4.105 $Y=2.475 $X2=0
+ $Y2=0
cc_312 N_A_232_98#_c_259_n N_VPWR_c_897_n 0.00644887f $X=4.19 $Y=2.39 $X2=0
+ $Y2=0
cc_313 N_A_232_98#_c_253_n N_VPWR_c_907_n 0.00562877f $X=2.215 $Y=1.88 $X2=0
+ $Y2=0
cc_314 N_A_232_98#_c_256_n N_VPWR_c_907_n 0.0142726f $X=1.317 $Y=2.56 $X2=0
+ $Y2=0
cc_315 N_A_232_98#_c_253_n N_VPWR_c_894_n 0.00595788f $X=2.215 $Y=1.88 $X2=0
+ $Y2=0
cc_316 N_A_232_98#_c_256_n N_VPWR_c_894_n 0.0119658f $X=1.317 $Y=2.56 $X2=0
+ $Y2=0
cc_317 N_A_232_98#_c_258_n N_VPWR_c_894_n 0.0579251f $X=4.105 $Y=2.475 $X2=0
+ $Y2=0
cc_318 N_A_232_98#_c_260_n N_VPWR_c_894_n 0.0318218f $X=1.655 $Y=2.44 $X2=0
+ $Y2=0
cc_319 N_A_232_98#_c_258_n A_568_392# 0.00466147f $X=4.105 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_320 N_A_232_98#_c_259_n A_817_392# 0.00679946f $X=4.19 $Y=2.39 $X2=-0.19
+ $Y2=-0.245
cc_321 N_A_232_98#_M1004_g N_VGND_c_1069_n 0.00758354f $X=2.155 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_232_98#_c_241_n N_VGND_c_1070_n 9.62872e-19 $X=3.16 $Y=1.11 $X2=0
+ $Y2=0
cc_323 N_A_232_98#_M1004_g N_VGND_c_1081_n 0.00409717f $X=2.155 $Y=0.74 $X2=0
+ $Y2=0
cc_324 N_A_27_136#_c_390_n N_A_343_74#_M1004_s 0.00966132f $X=2.515 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_325 N_A_27_136#_M1011_g N_A_343_74#_M1017_g 0.0735542f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_326 N_A_27_136#_c_390_n N_A_343_74#_c_467_n 0.0349225f $X=2.515 $Y=0.665
+ $X2=0 $Y2=0
cc_327 N_A_27_136#_c_392_n N_A_343_74#_c_467_n 0.00919669f $X=2.68 $Y=1.385
+ $X2=0 $Y2=0
cc_328 N_A_27_136#_M1011_g N_A_343_74#_c_476_n 0.00156565f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_329 N_A_27_136#_M1011_g N_A_343_74#_c_468_n 8.67244e-19 $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_330 N_A_27_136#_c_392_n N_A_343_74#_c_468_n 0.0214523f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_331 N_A_27_136#_c_393_n N_A_343_74#_c_468_n 0.0011754f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_332 N_A_27_136#_M1011_g N_A_343_74#_c_478_n 0.0133699f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_333 N_A_27_136#_c_392_n N_A_343_74#_c_478_n 0.025539f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_334 N_A_27_136#_c_393_n N_A_343_74#_c_478_n 0.00345141f $X=2.68 $Y=1.385
+ $X2=0 $Y2=0
cc_335 N_A_27_136#_M1012_g N_A_343_74#_c_469_n 0.00389603f $X=2.77 $Y=0.715
+ $X2=0 $Y2=0
cc_336 N_A_27_136#_M1011_g N_A_343_74#_c_472_n 0.00389005f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_337 N_A_27_136#_c_393_n N_A_343_74#_c_472_n 0.00398233f $X=2.68 $Y=1.385
+ $X2=0 $Y2=0
cc_338 N_A_27_136#_M1011_g N_A_343_74#_c_473_n 0.0149276f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_339 N_A_27_136#_c_393_n N_A_343_74#_c_473_n 0.00500108f $X=2.68 $Y=1.385
+ $X2=0 $Y2=0
cc_340 N_A_27_136#_M1012_g N_A_343_74#_c_474_n 0.00599955f $X=2.77 $Y=0.715
+ $X2=0 $Y2=0
cc_341 N_A_27_136#_c_390_n N_A_343_74#_c_474_n 0.0133619f $X=2.515 $Y=0.665
+ $X2=0 $Y2=0
cc_342 N_A_27_136#_c_392_n N_A_343_74#_c_474_n 0.0592147f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_343 N_A_27_136#_M1011_g N_A_647_79#_c_750_n 7.99808e-19 $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_344 N_A_27_136#_c_397_n N_VPWR_c_895_n 0.0220172f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_345 N_A_27_136#_M1011_g N_VPWR_c_896_n 0.0103389f $X=2.75 $Y=2.46 $X2=0 $Y2=0
cc_346 N_A_27_136#_M1011_g N_VPWR_c_903_n 0.00460063f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_347 N_A_27_136#_c_397_n N_VPWR_c_911_n 0.015305f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_348 N_A_27_136#_M1011_g N_VPWR_c_894_n 0.00443063f $X=2.75 $Y=2.46 $X2=0
+ $Y2=0
cc_349 N_A_27_136#_c_397_n N_VPWR_c_894_n 0.0126681f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_350 N_A_27_136#_c_390_n N_VGND_M1018_d 0.0162931f $X=2.515 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_351 N_A_27_136#_c_390_n N_VGND_M1004_d 0.0132139f $X=2.515 $Y=0.665 $X2=0
+ $Y2=0
cc_352 N_A_27_136#_c_392_n N_VGND_M1004_d 0.00360055f $X=2.68 $Y=1.385 $X2=0
+ $Y2=0
cc_353 N_A_27_136#_M1012_g N_VGND_c_1069_n 0.001789f $X=2.77 $Y=0.715 $X2=0
+ $Y2=0
cc_354 N_A_27_136#_c_390_n N_VGND_c_1069_n 0.0514958f $X=2.515 $Y=0.665 $X2=0
+ $Y2=0
cc_355 N_A_27_136#_M1012_g N_VGND_c_1070_n 0.00423046f $X=2.77 $Y=0.715 $X2=0
+ $Y2=0
cc_356 N_A_27_136#_c_390_n N_VGND_c_1070_n 0.00368689f $X=2.515 $Y=0.665 $X2=0
+ $Y2=0
cc_357 N_A_27_136#_c_390_n N_VGND_c_1076_n 0.00345394f $X=2.515 $Y=0.665 $X2=0
+ $Y2=0
cc_358 N_A_27_136#_c_391_n N_VGND_c_1076_n 0.00780247f $X=0.445 $Y=0.665 $X2=0
+ $Y2=0
cc_359 N_A_27_136#_c_390_n N_VGND_c_1079_n 0.0246008f $X=2.515 $Y=0.665 $X2=0
+ $Y2=0
cc_360 N_A_27_136#_M1012_g N_VGND_c_1081_n 0.00537853f $X=2.77 $Y=0.715 $X2=0
+ $Y2=0
cc_361 N_A_27_136#_c_390_n N_VGND_c_1081_n 0.0539352f $X=2.515 $Y=0.665 $X2=0
+ $Y2=0
cc_362 N_A_27_136#_c_391_n N_VGND_c_1081_n 0.0108671f $X=0.445 $Y=0.665 $X2=0
+ $Y2=0
cc_363 N_A_343_74#_c_466_n N_A_887_270#_M1022_g 0.0272682f $X=4.12 $Y=0.505
+ $X2=0 $Y2=0
cc_364 N_A_343_74#_c_470_n N_A_647_79#_M1013_d 0.00253551f $X=4.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_365 N_A_343_74#_M1017_g N_A_647_79#_c_750_n 0.00418839f $X=3.17 $Y=2.46 $X2=0
+ $Y2=0
cc_366 N_A_343_74#_c_472_n N_A_647_79#_c_750_n 0.00996264f $X=3.22 $Y=1.635
+ $X2=0 $Y2=0
cc_367 N_A_343_74#_c_473_n N_A_647_79#_c_750_n 6.00906e-19 $X=3.22 $Y=1.635
+ $X2=0 $Y2=0
cc_368 N_A_343_74#_M1017_g N_A_647_79#_c_741_n 0.00326542f $X=3.17 $Y=2.46 $X2=0
+ $Y2=0
cc_369 N_A_343_74#_c_472_n N_A_647_79#_c_741_n 0.0314209f $X=3.22 $Y=1.635 $X2=0
+ $Y2=0
cc_370 N_A_343_74#_c_473_n N_A_647_79#_c_741_n 0.00214697f $X=3.22 $Y=1.635
+ $X2=0 $Y2=0
cc_371 N_A_343_74#_c_474_n N_A_647_79#_c_741_n 0.0119182f $X=3.2 $Y=1.47 $X2=0
+ $Y2=0
cc_372 N_A_343_74#_c_466_n N_A_647_79#_c_742_n 0.0081273f $X=4.12 $Y=0.505 $X2=0
+ $Y2=0
cc_373 N_A_343_74#_c_470_n N_A_647_79#_c_742_n 0.00478234f $X=4.1 $Y=0.34 $X2=0
+ $Y2=0
cc_374 N_A_343_74#_c_466_n N_A_647_79#_c_743_n 0.00869586f $X=4.12 $Y=0.505
+ $X2=0 $Y2=0
cc_375 N_A_343_74#_c_470_n N_A_647_79#_c_743_n 0.0415775f $X=4.1 $Y=0.34 $X2=0
+ $Y2=0
cc_376 N_A_343_74#_c_471_n N_A_647_79#_c_743_n 0.00734404f $X=4.1 $Y=0.34 $X2=0
+ $Y2=0
cc_377 N_A_343_74#_c_472_n N_A_647_79#_c_743_n 0.00120024f $X=3.22 $Y=1.635
+ $X2=0 $Y2=0
cc_378 N_A_343_74#_c_474_n N_A_647_79#_c_743_n 0.0317057f $X=3.2 $Y=1.47 $X2=0
+ $Y2=0
cc_379 N_A_343_74#_M1017_g N_VPWR_c_896_n 0.00174454f $X=3.17 $Y=2.46 $X2=0
+ $Y2=0
cc_380 N_A_343_74#_M1017_g N_VPWR_c_903_n 0.00553757f $X=3.17 $Y=2.46 $X2=0
+ $Y2=0
cc_381 N_A_343_74#_M1017_g N_VPWR_c_894_n 0.00540034f $X=3.17 $Y=2.46 $X2=0
+ $Y2=0
cc_382 N_A_343_74#_c_466_n N_VGND_c_1063_n 0.00488592f $X=4.12 $Y=0.505 $X2=0
+ $Y2=0
cc_383 N_A_343_74#_c_470_n N_VGND_c_1063_n 0.0117986f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_384 N_A_343_74#_c_469_n N_VGND_c_1069_n 0.00751318f $X=3.185 $Y=0.38 $X2=0
+ $Y2=0
cc_385 N_A_343_74#_c_469_n N_VGND_c_1070_n 0.0121867f $X=3.185 $Y=0.38 $X2=0
+ $Y2=0
cc_386 N_A_343_74#_c_470_n N_VGND_c_1070_n 0.0693566f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_387 N_A_343_74#_c_471_n N_VGND_c_1070_n 0.0131137f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_388 N_A_343_74#_c_466_n N_VGND_c_1081_n 0.00664082f $X=4.12 $Y=0.505 $X2=0
+ $Y2=0
cc_389 N_A_343_74#_c_469_n N_VGND_c_1081_n 0.00660921f $X=3.185 $Y=0.38 $X2=0
+ $Y2=0
cc_390 N_A_343_74#_c_470_n N_VGND_c_1081_n 0.0378549f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_391 N_A_343_74#_c_471_n N_VGND_c_1081_n 0.0119786f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_392 N_A_343_74#_c_469_n A_569_79# 0.00148387f $X=3.185 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_393 N_A_343_74#_c_474_n A_569_79# 0.0046631f $X=3.2 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_394 N_A_887_270#_M1021_g N_A_647_79#_M1009_g 0.0158644f $X=4.525 $Y=2.17
+ $X2=0 $Y2=0
cc_395 N_A_887_270#_c_593_n N_A_647_79#_M1009_g 0.00163644f $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_396 N_A_887_270#_c_583_n N_A_647_79#_M1009_g 0.0053658f $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_397 N_A_887_270#_c_595_n N_A_647_79#_M1009_g 0.01389f $X=5.25 $Y=1.805 $X2=0
+ $Y2=0
cc_398 N_A_887_270#_c_597_n N_A_647_79#_M1009_g 0.00655648f $X=5.415 $Y=1.985
+ $X2=0 $Y2=0
cc_399 N_A_887_270#_c_598_n N_A_647_79#_M1009_g 0.0078776f $X=5.415 $Y=2.815
+ $X2=0 $Y2=0
cc_400 N_A_887_270#_c_584_n N_A_647_79#_M1009_g 0.00568868f $X=5.57 $Y=1.72
+ $X2=0 $Y2=0
cc_401 N_A_887_270#_c_602_n N_A_647_79#_M1009_g 0.00342996f $X=5.452 $Y=1.805
+ $X2=0 $Y2=0
cc_402 N_A_887_270#_c_603_n N_A_647_79#_M1009_g 0.00195991f $X=5.452 $Y=2.325
+ $X2=0 $Y2=0
cc_403 N_A_887_270#_M1015_d N_A_647_79#_c_742_n 0.00157147f $X=5.21 $Y=0.37
+ $X2=0 $Y2=0
cc_404 N_A_887_270#_M1022_g N_A_647_79#_c_742_n 0.0149129f $X=4.58 $Y=0.825
+ $X2=0 $Y2=0
cc_405 N_A_887_270#_c_593_n N_A_647_79#_c_742_n 0.0251561f $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_406 N_A_887_270#_c_583_n N_A_647_79#_c_742_n 0.00474267f $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_407 N_A_887_270#_c_595_n N_A_647_79#_c_742_n 0.007112f $X=5.25 $Y=1.805 $X2=0
+ $Y2=0
cc_408 N_A_887_270#_c_584_n N_A_647_79#_c_742_n 0.014063f $X=5.57 $Y=1.72 $X2=0
+ $Y2=0
cc_409 N_A_887_270#_c_587_n N_A_647_79#_c_742_n 0.00615278f $X=5.57 $Y=0.597
+ $X2=0 $Y2=0
cc_410 N_A_887_270#_M1022_g N_A_647_79#_c_743_n 0.00117111f $X=4.58 $Y=0.825
+ $X2=0 $Y2=0
cc_411 N_A_887_270#_M1022_g N_A_647_79#_c_744_n 0.00148093f $X=4.58 $Y=0.825
+ $X2=0 $Y2=0
cc_412 N_A_887_270#_c_593_n N_A_647_79#_c_744_n 0.0123578f $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_413 N_A_887_270#_c_583_n N_A_647_79#_c_744_n 7.18735e-19 $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_414 N_A_887_270#_c_595_n N_A_647_79#_c_744_n 0.0201041f $X=5.25 $Y=1.805
+ $X2=0 $Y2=0
cc_415 N_A_887_270#_c_584_n N_A_647_79#_c_744_n 0.0275348f $X=5.57 $Y=1.72 $X2=0
+ $Y2=0
cc_416 N_A_887_270#_c_602_n N_A_647_79#_c_744_n 0.0054737f $X=5.452 $Y=1.805
+ $X2=0 $Y2=0
cc_417 N_A_887_270#_M1022_g N_A_647_79#_c_745_n 0.00521165f $X=4.58 $Y=0.825
+ $X2=0 $Y2=0
cc_418 N_A_887_270#_c_593_n N_A_647_79#_c_745_n 6.79167e-19 $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_419 N_A_887_270#_c_583_n N_A_647_79#_c_745_n 0.0122491f $X=4.61 $Y=1.515
+ $X2=0 $Y2=0
cc_420 N_A_887_270#_c_595_n N_A_647_79#_c_745_n 7.99874e-19 $X=5.25 $Y=1.805
+ $X2=0 $Y2=0
cc_421 N_A_887_270#_c_584_n N_A_647_79#_c_745_n 0.00739878f $X=5.57 $Y=1.72
+ $X2=0 $Y2=0
cc_422 N_A_887_270#_c_587_n N_A_647_79#_c_745_n 3.84739e-19 $X=5.57 $Y=0.597
+ $X2=0 $Y2=0
cc_423 N_A_887_270#_c_602_n N_A_647_79#_c_745_n 2.69101e-19 $X=5.452 $Y=1.805
+ $X2=0 $Y2=0
cc_424 N_A_887_270#_M1022_g N_A_647_79#_c_746_n 0.015054f $X=4.58 $Y=0.825 $X2=0
+ $Y2=0
cc_425 N_A_887_270#_c_584_n N_A_647_79#_c_746_n 0.00632728f $X=5.57 $Y=1.72
+ $X2=0 $Y2=0
cc_426 N_A_887_270#_c_587_n N_A_647_79#_c_746_n 0.00802501f $X=5.57 $Y=0.597
+ $X2=0 $Y2=0
cc_427 N_A_887_270#_c_588_n N_A_1442_94#_c_834_n 0.0182623f $X=7.135 $Y=1.465
+ $X2=0 $Y2=0
cc_428 N_A_887_270#_M1016_g N_A_1442_94#_c_835_n 0.00611061f $X=7.135 $Y=0.79
+ $X2=0 $Y2=0
cc_429 N_A_887_270#_M1016_g N_A_1442_94#_c_836_n 0.00742201f $X=7.135 $Y=0.79
+ $X2=0 $Y2=0
cc_430 N_A_887_270#_c_585_n N_A_1442_94#_c_836_n 0.00109962f $X=6.87 $Y=1.63
+ $X2=0 $Y2=0
cc_431 N_A_887_270#_c_588_n N_A_1442_94#_c_836_n 0.00148793f $X=7.135 $Y=1.465
+ $X2=0 $Y2=0
cc_432 N_A_887_270#_M1024_g N_A_1442_94#_c_841_n 0.00124359f $X=6.65 $Y=2.4
+ $X2=0 $Y2=0
cc_433 N_A_887_270#_M1010_g N_A_1442_94#_c_841_n 0.024961f $X=7.155 $Y=2.46
+ $X2=0 $Y2=0
cc_434 N_A_887_270#_c_600_n N_A_1442_94#_c_841_n 0.0101259f $X=6.785 $Y=2.325
+ $X2=0 $Y2=0
cc_435 N_A_887_270#_c_586_n N_A_1442_94#_c_841_n 0.0316465f $X=6.87 $Y=2.24
+ $X2=0 $Y2=0
cc_436 N_A_887_270#_M1016_g N_A_1442_94#_c_837_n 0.00337479f $X=7.135 $Y=0.79
+ $X2=0 $Y2=0
cc_437 N_A_887_270#_c_588_n N_A_1442_94#_c_837_n 2.4036e-19 $X=7.135 $Y=1.465
+ $X2=0 $Y2=0
cc_438 N_A_887_270#_M1010_g N_A_1442_94#_c_838_n 4.50765e-19 $X=7.155 $Y=2.46
+ $X2=0 $Y2=0
cc_439 N_A_887_270#_c_585_n N_A_1442_94#_c_838_n 0.0186054f $X=6.87 $Y=1.63
+ $X2=0 $Y2=0
cc_440 N_A_887_270#_c_586_n N_A_1442_94#_c_838_n 0.00110185f $X=6.87 $Y=2.24
+ $X2=0 $Y2=0
cc_441 N_A_887_270#_c_588_n N_A_1442_94#_c_838_n 0.00974945f $X=7.135 $Y=1.465
+ $X2=0 $Y2=0
cc_442 N_A_887_270#_c_595_n N_VPWR_M1021_d 0.0022138f $X=5.25 $Y=1.805 $X2=0
+ $Y2=0
cc_443 N_A_887_270#_c_600_n N_VPWR_M1000_d 0.00886389f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_444 N_A_887_270#_c_600_n N_VPWR_M1024_d 0.00379308f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_445 N_A_887_270#_c_586_n N_VPWR_M1024_d 0.00614027f $X=6.87 $Y=2.24 $X2=0
+ $Y2=0
cc_446 N_A_887_270#_M1021_g N_VPWR_c_897_n 0.00398805f $X=4.525 $Y=2.17 $X2=0
+ $Y2=0
cc_447 N_A_887_270#_c_583_n N_VPWR_c_897_n 5.03772e-19 $X=4.61 $Y=1.515 $X2=0
+ $Y2=0
cc_448 N_A_887_270#_c_595_n N_VPWR_c_897_n 0.0209569f $X=5.25 $Y=1.805 $X2=0
+ $Y2=0
cc_449 N_A_887_270#_c_596_n N_VPWR_c_897_n 0.00896127f $X=4.775 $Y=1.805 $X2=0
+ $Y2=0
cc_450 N_A_887_270#_c_598_n N_VPWR_c_897_n 0.0228467f $X=5.415 $Y=2.815 $X2=0
+ $Y2=0
cc_451 N_A_887_270#_M1000_g N_VPWR_c_898_n 0.0132135f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_452 N_A_887_270#_M1024_g N_VPWR_c_898_n 0.00149457f $X=6.65 $Y=2.4 $X2=0
+ $Y2=0
cc_453 N_A_887_270#_c_598_n N_VPWR_c_898_n 0.0258522f $X=5.415 $Y=2.815 $X2=0
+ $Y2=0
cc_454 N_A_887_270#_c_600_n N_VPWR_c_898_n 0.0153892f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_455 N_A_887_270#_M1000_g N_VPWR_c_899_n 0.00149196f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_456 N_A_887_270#_M1024_g N_VPWR_c_899_n 0.012302f $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_457 N_A_887_270#_M1010_g N_VPWR_c_899_n 0.00336208f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_458 N_A_887_270#_c_600_n N_VPWR_c_899_n 0.0164096f $X=6.785 $Y=2.325 $X2=0
+ $Y2=0
cc_459 N_A_887_270#_M1010_g N_VPWR_c_900_n 0.00496623f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_460 N_A_887_270#_M1000_g N_VPWR_c_905_n 0.00460063f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_461 N_A_887_270#_M1024_g N_VPWR_c_905_n 0.00460063f $X=6.65 $Y=2.4 $X2=0
+ $Y2=0
cc_462 N_A_887_270#_c_598_n N_VPWR_c_908_n 0.0178955f $X=5.415 $Y=2.815 $X2=0
+ $Y2=0
cc_463 N_A_887_270#_M1010_g N_VPWR_c_909_n 0.005209f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_464 N_A_887_270#_M1021_g N_VPWR_c_894_n 0.00465911f $X=4.525 $Y=2.17 $X2=0
+ $Y2=0
cc_465 N_A_887_270#_M1000_g N_VPWR_c_894_n 0.00908554f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A_887_270#_M1024_g N_VPWR_c_894_n 0.00908554f $X=6.65 $Y=2.4 $X2=0
+ $Y2=0
cc_467 N_A_887_270#_M1010_g N_VPWR_c_894_n 0.00987373f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_468 N_A_887_270#_c_598_n N_VPWR_c_894_n 0.0147443f $X=5.415 $Y=2.815 $X2=0
+ $Y2=0
cc_469 N_A_887_270#_c_600_n N_Q_M1000_s 0.0075347f $X=6.785 $Y=2.325 $X2=0 $Y2=0
cc_470 N_A_887_270#_M1000_g N_Q_c_998_n 0.00521827f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A_887_270#_c_597_n N_Q_c_998_n 0.0127317f $X=5.415 $Y=1.985 $X2=0 $Y2=0
cc_472 N_A_887_270#_c_600_n N_Q_c_998_n 0.014007f $X=6.785 $Y=2.325 $X2=0 $Y2=0
cc_473 N_A_887_270#_c_602_n N_Q_c_998_n 0.00673592f $X=5.452 $Y=1.805 $X2=0
+ $Y2=0
cc_474 N_A_887_270#_M1000_g N_Q_c_999_n 0.0121f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_475 N_A_887_270#_M1024_g N_Q_c_999_n 0.00445056f $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_476 N_A_887_270#_c_600_n N_Q_c_999_n 0.0260347f $X=6.785 $Y=2.325 $X2=0 $Y2=0
cc_477 N_A_887_270#_c_586_n N_Q_c_999_n 0.0114667f $X=6.87 $Y=2.24 $X2=0 $Y2=0
cc_478 N_A_887_270#_c_701_p N_Q_c_999_n 0.0236214f $X=6.79 $Y=1.465 $X2=0 $Y2=0
cc_479 N_A_887_270#_c_588_n N_Q_c_999_n 0.00235524f $X=7.135 $Y=1.465 $X2=0
+ $Y2=0
cc_480 N_A_887_270#_M1002_g N_Q_c_995_n 2.80152e-19 $X=6.125 $Y=0.74 $X2=0 $Y2=0
cc_481 N_A_887_270#_M1008_g N_Q_c_995_n 0.00593075f $X=6.555 $Y=0.74 $X2=0 $Y2=0
cc_482 N_A_887_270#_M1002_g N_Q_c_996_n 0.015065f $X=6.125 $Y=0.74 $X2=0 $Y2=0
cc_483 N_A_887_270#_M1008_g N_Q_c_996_n 0.00358118f $X=6.555 $Y=0.74 $X2=0 $Y2=0
cc_484 N_A_887_270#_c_584_n N_Q_c_996_n 0.0183676f $X=5.57 $Y=1.72 $X2=0 $Y2=0
cc_485 N_A_887_270#_c_701_p N_Q_c_996_n 0.0170873f $X=6.79 $Y=1.465 $X2=0 $Y2=0
cc_486 N_A_887_270#_c_588_n N_Q_c_996_n 0.00262336f $X=7.135 $Y=1.465 $X2=0
+ $Y2=0
cc_487 N_A_887_270#_M1002_g Q 0.0066884f $X=6.125 $Y=0.74 $X2=0 $Y2=0
cc_488 N_A_887_270#_M1000_g Q 0.00635149f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_489 N_A_887_270#_M1008_g Q 8.9393e-19 $X=6.555 $Y=0.74 $X2=0 $Y2=0
cc_490 N_A_887_270#_M1024_g Q 4.8868e-19 $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_491 N_A_887_270#_c_584_n Q 0.0367836f $X=5.57 $Y=1.72 $X2=0 $Y2=0
cc_492 N_A_887_270#_c_586_n Q 0.00428129f $X=6.87 $Y=2.24 $X2=0 $Y2=0
cc_493 N_A_887_270#_c_602_n Q 0.00554709f $X=5.452 $Y=1.805 $X2=0 $Y2=0
cc_494 N_A_887_270#_c_701_p Q 0.0254856f $X=6.79 $Y=1.465 $X2=0 $Y2=0
cc_495 N_A_887_270#_c_588_n Q 0.0129504f $X=7.135 $Y=1.465 $X2=0 $Y2=0
cc_496 N_A_887_270#_M1022_g N_VGND_c_1063_n 0.00931115f $X=4.58 $Y=0.825 $X2=0
+ $Y2=0
cc_497 N_A_887_270#_c_587_n N_VGND_c_1063_n 0.0204019f $X=5.57 $Y=0.597 $X2=0
+ $Y2=0
cc_498 N_A_887_270#_M1002_g N_VGND_c_1064_n 0.00866236f $X=6.125 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_887_270#_M1008_g N_VGND_c_1064_n 4.50236e-19 $X=6.555 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_887_270#_c_587_n N_VGND_c_1064_n 0.0272606f $X=5.57 $Y=0.597 $X2=0
+ $Y2=0
cc_501 N_A_887_270#_M1008_g N_VGND_c_1065_n 0.00804415f $X=6.555 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_A_887_270#_M1016_g N_VGND_c_1065_n 0.00744268f $X=7.135 $Y=0.79 $X2=0
+ $Y2=0
cc_503 N_A_887_270#_c_585_n N_VGND_c_1065_n 0.0151563f $X=6.87 $Y=1.63 $X2=0
+ $Y2=0
cc_504 N_A_887_270#_c_701_p N_VGND_c_1065_n 0.00915551f $X=6.79 $Y=1.465 $X2=0
+ $Y2=0
cc_505 N_A_887_270#_c_588_n N_VGND_c_1065_n 0.00377846f $X=7.135 $Y=1.465 $X2=0
+ $Y2=0
cc_506 N_A_887_270#_M1016_g N_VGND_c_1066_n 0.00405453f $X=7.135 $Y=0.79 $X2=0
+ $Y2=0
cc_507 N_A_887_270#_M1022_g N_VGND_c_1070_n 0.00349617f $X=4.58 $Y=0.825 $X2=0
+ $Y2=0
cc_508 N_A_887_270#_c_587_n N_VGND_c_1072_n 0.0203373f $X=5.57 $Y=0.597 $X2=0
+ $Y2=0
cc_509 N_A_887_270#_M1002_g N_VGND_c_1074_n 0.00383152f $X=6.125 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_887_270#_M1008_g N_VGND_c_1074_n 0.0043438f $X=6.555 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_887_270#_M1016_g N_VGND_c_1077_n 0.00485498f $X=7.135 $Y=0.79 $X2=0
+ $Y2=0
cc_512 N_A_887_270#_M1022_g N_VGND_c_1081_n 0.00396651f $X=4.58 $Y=0.825 $X2=0
+ $Y2=0
cc_513 N_A_887_270#_M1002_g N_VGND_c_1081_n 0.00386058f $X=6.125 $Y=0.74 $X2=0
+ $Y2=0
cc_514 N_A_887_270#_M1008_g N_VGND_c_1081_n 0.0082053f $X=6.555 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_887_270#_M1016_g N_VGND_c_1081_n 0.00514438f $X=7.135 $Y=0.79 $X2=0
+ $Y2=0
cc_516 N_A_887_270#_c_587_n N_VGND_c_1081_n 0.0170424f $X=5.57 $Y=0.597 $X2=0
+ $Y2=0
cc_517 N_A_647_79#_M1009_g N_VPWR_c_897_n 0.0181104f $X=5.19 $Y=2.4 $X2=0 $Y2=0
cc_518 N_A_647_79#_M1009_g N_VPWR_c_898_n 0.00317114f $X=5.19 $Y=2.4 $X2=0 $Y2=0
cc_519 N_A_647_79#_M1009_g N_VPWR_c_908_n 0.005209f $X=5.19 $Y=2.4 $X2=0 $Y2=0
cc_520 N_A_647_79#_M1009_g N_VPWR_c_894_n 0.0099186f $X=5.19 $Y=2.4 $X2=0 $Y2=0
cc_521 N_A_647_79#_M1009_g N_Q_c_998_n 5.72896e-19 $X=5.19 $Y=2.4 $X2=0 $Y2=0
cc_522 N_A_647_79#_M1009_g Q 2.67281e-19 $X=5.19 $Y=2.4 $X2=0 $Y2=0
cc_523 N_A_647_79#_c_742_n N_VGND_M1022_d 0.00313795f $X=4.985 $Y=1.1 $X2=0
+ $Y2=0
cc_524 N_A_647_79#_c_742_n N_VGND_c_1063_n 0.0255566f $X=4.985 $Y=1.1 $X2=0
+ $Y2=0
cc_525 N_A_647_79#_c_743_n N_VGND_c_1063_n 0.00363658f $X=4.07 $Y=1.1 $X2=0
+ $Y2=0
cc_526 N_A_647_79#_c_746_n N_VGND_c_1063_n 0.00955147f $X=5.15 $Y=1.22 $X2=0
+ $Y2=0
cc_527 N_A_647_79#_c_746_n N_VGND_c_1064_n 0.00290507f $X=5.15 $Y=1.22 $X2=0
+ $Y2=0
cc_528 N_A_647_79#_c_746_n N_VGND_c_1072_n 0.00433162f $X=5.15 $Y=1.22 $X2=0
+ $Y2=0
cc_529 N_A_647_79#_c_746_n N_VGND_c_1081_n 0.00826407f $X=5.15 $Y=1.22 $X2=0
+ $Y2=0
cc_530 N_A_647_79#_c_742_n A_839_123# 0.00718311f $X=4.985 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_531 N_A_1442_94#_c_841_n N_VPWR_c_899_n 0.0154383f $X=7.38 $Y=2.105 $X2=0
+ $Y2=0
cc_532 N_A_1442_94#_M1003_g N_VPWR_c_900_n 0.00649215f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_533 N_A_1442_94#_c_834_n N_VPWR_c_900_n 0.00577732f $X=8.075 $Y=1.485 $X2=0
+ $Y2=0
cc_534 N_A_1442_94#_c_841_n N_VPWR_c_900_n 0.0765956f $X=7.38 $Y=2.105 $X2=0
+ $Y2=0
cc_535 N_A_1442_94#_c_861_p N_VPWR_c_900_n 0.0209147f $X=7.99 $Y=1.485 $X2=0
+ $Y2=0
cc_536 N_A_1442_94#_M1005_g N_VPWR_c_902_n 0.00649215f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_537 N_A_1442_94#_c_841_n N_VPWR_c_909_n 0.014549f $X=7.38 $Y=2.105 $X2=0
+ $Y2=0
cc_538 N_A_1442_94#_M1003_g N_VPWR_c_910_n 0.005209f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_539 N_A_1442_94#_M1005_g N_VPWR_c_910_n 0.005209f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_540 N_A_1442_94#_M1003_g N_VPWR_c_894_n 0.00987399f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_541 N_A_1442_94#_M1005_g N_VPWR_c_894_n 0.00986008f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_542 N_A_1442_94#_c_841_n N_VPWR_c_894_n 0.0119743f $X=7.38 $Y=2.105 $X2=0
+ $Y2=0
cc_543 N_A_1442_94#_M1007_g N_Q_N_c_1039_n 0.00792614f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_A_1442_94#_M1014_g N_Q_N_c_1039_n 0.00505299f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_545 N_A_1442_94#_M1007_g N_Q_N_c_1040_n 0.00270721f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_A_1442_94#_M1003_g Q_N 0.0173318f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_547 N_A_1442_94#_c_831_n Q_N 0.00481639f $X=8.615 $Y=1.645 $X2=0 $Y2=0
cc_548 N_A_1442_94#_M1005_g Q_N 0.0173318f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_549 N_A_1442_94#_M1003_g N_Q_N_c_1041_n 0.00396377f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_550 N_A_1442_94#_M1007_g N_Q_N_c_1041_n 0.00451055f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_551 N_A_1442_94#_c_831_n N_Q_N_c_1041_n 0.0289506f $X=8.615 $Y=1.645 $X2=0
+ $Y2=0
cc_552 N_A_1442_94#_M1005_g N_Q_N_c_1041_n 0.00429389f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_553 N_A_1442_94#_c_861_p N_Q_N_c_1041_n 0.0250004f $X=7.99 $Y=1.485 $X2=0
+ $Y2=0
cc_554 N_A_1442_94#_c_835_n N_VGND_c_1065_n 0.0258547f $X=7.35 $Y=0.615 $X2=0
+ $Y2=0
cc_555 N_A_1442_94#_M1007_g N_VGND_c_1066_n 0.0184013f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_556 N_A_1442_94#_c_834_n N_VGND_c_1066_n 0.0075646f $X=8.075 $Y=1.485 $X2=0
+ $Y2=0
cc_557 N_A_1442_94#_c_835_n N_VGND_c_1066_n 0.0458112f $X=7.35 $Y=0.615 $X2=0
+ $Y2=0
cc_558 N_A_1442_94#_c_861_p N_VGND_c_1066_n 0.0254428f $X=7.99 $Y=1.485 $X2=0
+ $Y2=0
cc_559 N_A_1442_94#_M1007_g N_VGND_c_1068_n 6.13445e-19 $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_560 N_A_1442_94#_c_831_n N_VGND_c_1068_n 2.01871e-19 $X=8.615 $Y=1.645 $X2=0
+ $Y2=0
cc_561 N_A_1442_94#_M1014_g N_VGND_c_1068_n 0.0160357f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_562 N_A_1442_94#_c_835_n N_VGND_c_1077_n 0.0103491f $X=7.35 $Y=0.615 $X2=0
+ $Y2=0
cc_563 N_A_1442_94#_M1007_g N_VGND_c_1078_n 0.00434272f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_564 N_A_1442_94#_M1014_g N_VGND_c_1078_n 0.00383152f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_565 N_A_1442_94#_M1007_g N_VGND_c_1081_n 0.00825059f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_566 N_A_1442_94#_M1014_g N_VGND_c_1081_n 0.0075754f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_567 N_A_1442_94#_c_835_n N_VGND_c_1081_n 0.0113354f $X=7.35 $Y=0.615 $X2=0
+ $Y2=0
cc_568 N_VPWR_M1000_d N_Q_c_998_n 0.00507725f $X=5.83 $Y=1.84 $X2=0 $Y2=0
cc_569 N_VPWR_c_900_n Q_N 0.0395357f $X=7.94 $Y=1.985 $X2=0 $Y2=0
cc_570 N_VPWR_c_902_n Q_N 0.0395357f $X=8.84 $Y=1.985 $X2=0 $Y2=0
cc_571 N_VPWR_c_910_n Q_N 0.0144623f $X=8.755 $Y=3.33 $X2=0 $Y2=0
cc_572 N_VPWR_c_894_n Q_N 0.0118344f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_573 N_Q_c_996_n N_VGND_M1002_s 0.00417801f $X=6.375 $Y=0.99 $X2=0 $Y2=0
cc_574 N_Q_c_995_n N_VGND_c_1064_n 0.0122486f $X=6.34 $Y=0.52 $X2=0 $Y2=0
cc_575 N_Q_c_996_n N_VGND_c_1064_n 0.0107023f $X=6.375 $Y=0.99 $X2=0 $Y2=0
cc_576 N_Q_c_995_n N_VGND_c_1065_n 0.0184898f $X=6.34 $Y=0.52 $X2=0 $Y2=0
cc_577 N_Q_c_996_n N_VGND_c_1065_n 0.0122991f $X=6.375 $Y=0.99 $X2=0 $Y2=0
cc_578 N_Q_c_995_n N_VGND_c_1074_n 0.0109621f $X=6.34 $Y=0.52 $X2=0 $Y2=0
cc_579 N_Q_c_995_n N_VGND_c_1081_n 0.00928322f $X=6.34 $Y=0.52 $X2=0 $Y2=0
cc_580 N_Q_c_996_n N_VGND_c_1081_n 0.00585568f $X=6.375 $Y=0.99 $X2=0 $Y2=0
cc_581 N_Q_N_c_1039_n N_VGND_c_1066_n 0.0295934f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_582 N_Q_N_c_1039_n N_VGND_c_1068_n 0.0294122f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_583 N_Q_N_c_1039_n N_VGND_c_1078_n 0.0109942f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_584 N_Q_N_c_1039_n N_VGND_c_1081_n 0.00904371f $X=8.41 $Y=0.515 $X2=0 $Y2=0

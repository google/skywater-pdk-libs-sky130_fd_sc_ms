* NGSPICE file created from sky130_fd_sc_ms__a221oi_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_117_368# B1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.8144e+12p pd=1.668e+07u as=2.6992e+12p ps=2.498e+07u
M1001 VGND A2 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=1.2432e+12p pd=1.224e+07u as=1.0138e+12p ps=1.014e+07u
M1002 VPWR A2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.4672e+12p pd=1.158e+07u as=0p ps=0u
M1003 a_531_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1326_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0138e+12p pd=1.014e+07u as=0p ps=0u
M1005 VGND A2 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B2 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_531_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_117_368# B1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1326_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.4282e+12p ps=1.422e+07u
M1010 a_534_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_531_368# B1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1326_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_531_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_117_368# B2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_534_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_531_368# B2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_534_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1326_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B2 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_117_368# B2 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A1 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y B1 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_531_368# B2 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_531_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A1 a_531_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=8.848e+11p ps=8.3e+06u
M1032 Y C1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y A1 a_534_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_534_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_117_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y B1 a_1326_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y C1 a_117_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_531_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


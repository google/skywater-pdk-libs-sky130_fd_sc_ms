* File: sky130_fd_sc_ms__nand3_4.pex.spice
* Created: Fri Aug 28 17:43:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND3_4%A 1 3 6 8 10 11 13 16 18 20 21 22 34 35
r61 33 35 12.8452 $w=3.94e-07 $l=1.05e-07 $layer=POLY_cond $X=1.37 $Y=1.452
+ $X2=1.475 $Y2=1.452
r62 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.515 $X2=1.37 $Y2=1.515
r63 31 33 3.05838 $w=3.94e-07 $l=2.5e-08 $layer=POLY_cond $X=1.345 $Y=1.452
+ $X2=1.37 $Y2=1.452
r64 30 31 52.6041 $w=3.94e-07 $l=4.3e-07 $layer=POLY_cond $X=0.915 $Y=1.452
+ $X2=1.345 $Y2=1.452
r65 28 30 27.5254 $w=3.94e-07 $l=2.25e-07 $layer=POLY_cond $X=0.69 $Y=1.452
+ $X2=0.915 $Y2=1.452
r66 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.515 $X2=0.69 $Y2=1.515
r67 26 28 22.632 $w=3.94e-07 $l=1.85e-07 $layer=POLY_cond $X=0.505 $Y=1.452
+ $X2=0.69 $Y2=1.452
r68 25 26 2.4467 $w=3.94e-07 $l=2e-08 $layer=POLY_cond $X=0.485 $Y=1.452
+ $X2=0.505 $Y2=1.452
r69 22 34 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.37 $Y2=1.565
r70 21 22 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r71 21 29 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.69
+ $Y2=1.565
r72 18 35 36.7005 $w=3.94e-07 $l=3.97618e-07 $layer=POLY_cond $X=1.775 $Y=1.225
+ $X2=1.475 $Y2=1.452
r73 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.775 $Y=1.225
+ $X2=1.775 $Y2=0.78
r74 14 35 21.1025 $w=1.8e-07 $l=2.28e-07 $layer=POLY_cond $X=1.475 $Y=1.68
+ $X2=1.475 $Y2=1.452
r75 14 16 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.475 $Y=1.68
+ $X2=1.475 $Y2=2.4
r76 11 31 25.4929 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=1.345 $Y=1.225
+ $X2=1.345 $Y2=1.452
r77 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.345 $Y=1.225
+ $X2=1.345 $Y2=0.78
r78 8 30 25.4929 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=0.915 $Y=1.225
+ $X2=0.915 $Y2=1.452
r79 8 10 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.915 $Y=1.225
+ $X2=0.915 $Y2=0.78
r80 4 26 21.1025 $w=1.8e-07 $l=2.28e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.452
r81 4 6 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
r82 1 25 25.4929 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=0.485 $Y=1.225
+ $X2=0.485 $Y2=1.452
r83 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.485 $Y=1.225
+ $X2=0.485 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%B 1 3 6 8 10 13 17 21 28 32 33 34 45
c66 45 0 1.88335e-19 $X=3.405 $Y=1.515
c67 21 0 4.53359e-20 $X=3.495 $Y=0.78
c68 17 0 1.20944e-20 $X=3.065 $Y=0.78
c69 6 0 1.07122e-19 $X=2.205 $Y=0.78
r70 45 47 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=3.405 $Y=1.557
+ $X2=3.495 $Y2=1.557
r71 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.405
+ $Y=1.515 $X2=3.405 $Y2=1.515
r72 43 45 43.5851 $w=3.76e-07 $l=3.4e-07 $layer=POLY_cond $X=3.065 $Y=1.557
+ $X2=3.405 $Y2=1.557
r73 40 41 26.9202 $w=3.76e-07 $l=2.1e-07 $layer=POLY_cond $X=2.425 $Y=1.557
+ $X2=2.635 $Y2=1.557
r74 34 46 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.405 $Y2=1.565
r75 33 46 7.63829 $w=4.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.405 $Y2=1.565
r76 31 43 43.5851 $w=3.76e-07 $l=3.4e-07 $layer=POLY_cond $X=2.725 $Y=1.557
+ $X2=3.065 $Y2=1.557
r77 31 41 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=2.725 $Y=1.557
+ $X2=2.635 $Y2=1.557
r78 30 32 5.82291 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.565
+ $X2=2.56 $Y2=1.565
r79 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.725
+ $Y=1.515 $X2=2.725 $Y2=1.515
r80 28 33 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.99 $Y=1.565
+ $X2=3.12 $Y2=1.565
r81 28 30 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.99 $Y=1.565
+ $X2=2.725 $Y2=1.565
r82 26 40 16.6649 $w=3.76e-07 $l=1.3e-07 $layer=POLY_cond $X=2.295 $Y=1.557
+ $X2=2.425 $Y2=1.557
r83 26 38 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=2.295 $Y=1.557
+ $X2=2.205 $Y2=1.557
r84 25 32 10.9071 $w=2.78e-07 $l=2.65e-07 $layer=LI1_cond $X=2.295 $Y=1.49
+ $X2=2.56 $Y2=1.49
r85 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.515 $X2=2.295 $Y2=1.515
r86 19 47 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=1.557
r87 19 21 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=0.78
r88 15 43 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=1.557
r89 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=0.78
r90 11 41 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=1.557
r91 11 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=0.78
r92 8 40 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.425 $Y=1.765
+ $X2=2.425 $Y2=1.557
r93 8 10 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=2.425 $Y=1.765
+ $X2=2.425 $Y2=2.4
r94 4 38 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=1.557
r95 4 6 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=0.78
r96 1 38 29.484 $w=3.76e-07 $l=3.17396e-07 $layer=POLY_cond $X=1.975 $Y=1.765
+ $X2=2.205 $Y2=1.557
r97 1 3 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=1.975 $Y=1.765
+ $X2=1.975 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%C 3 7 11 15 19 23 30 34 35 36 37 55
c63 34 0 2.21572e-19 $X=4.495 $Y=1.56
c64 23 0 1.6164e-19 $X=5.755 $Y=0.78
r65 53 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.665 $Y=1.505
+ $X2=5.755 $Y2=1.505
r66 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.665
+ $Y=1.505 $X2=5.665 $Y2=1.505
r67 51 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.325 $Y=1.505
+ $X2=5.665 $Y2=1.505
r68 49 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.985 $Y=1.505
+ $X2=5.325 $Y2=1.505
r69 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.505 $X2=4.985 $Y2=1.505
r70 47 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.895 $Y=1.505
+ $X2=4.985 $Y2=1.505
r71 44 45 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.35 $Y=1.505
+ $X2=4.465 $Y2=1.505
r72 37 54 8.77428 $w=4.38e-07 $l=3.35e-07 $layer=LI1_cond $X=6 $Y=1.56 $X2=5.665
+ $Y2=1.56
r73 36 54 3.79782 $w=4.38e-07 $l=1.45e-07 $layer=LI1_cond $X=5.52 $Y=1.56
+ $X2=5.665 $Y2=1.56
r74 35 36 12.5721 $w=4.38e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.56
+ $X2=5.52 $Y2=1.56
r75 35 50 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=5.04 $Y=1.56
+ $X2=4.985 $Y2=1.56
r76 33 47 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.645 $Y=1.505
+ $X2=4.895 $Y2=1.505
r77 33 45 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.645 $Y=1.505
+ $X2=4.465 $Y2=1.505
r78 32 34 5.26886 $w=4.38e-07 $l=1.5e-07 $layer=LI1_cond $X=4.645 $Y=1.56
+ $X2=4.495 $Y2=1.56
r79 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.645
+ $Y=1.505 $X2=4.645 $Y2=1.505
r80 30 50 1.30959 $w=4.38e-07 $l=5e-08 $layer=LI1_cond $X=4.935 $Y=1.56
+ $X2=4.985 $Y2=1.56
r81 30 32 7.59565 $w=4.38e-07 $l=2.9e-07 $layer=LI1_cond $X=4.935 $Y=1.56
+ $X2=4.645 $Y2=1.56
r82 28 44 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=4.305 $Y=1.505
+ $X2=4.35 $Y2=1.505
r83 28 41 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=4.305 $Y=1.505
+ $X2=3.9 $Y2=1.505
r84 27 34 7.55049 $w=2.88e-07 $l=1.9e-07 $layer=LI1_cond $X=4.305 $Y=1.485
+ $X2=4.495 $Y2=1.485
r85 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=1.505 $X2=4.305 $Y2=1.505
r86 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=1.34
+ $X2=5.755 $Y2=1.505
r87 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.755 $Y=1.34
+ $X2=5.755 $Y2=0.78
r88 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.34
+ $X2=5.325 $Y2=1.505
r89 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.325 $Y=1.34
+ $X2=5.325 $Y2=0.78
r90 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=1.34
+ $X2=4.895 $Y2=1.505
r91 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.895 $Y=1.34
+ $X2=4.895 $Y2=0.78
r92 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=1.34
+ $X2=4.465 $Y2=1.505
r93 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.465 $Y=1.34
+ $X2=4.465 $Y2=0.78
r94 5 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.67
+ $X2=4.35 $Y2=1.505
r95 5 7 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=4.35 $Y=1.67 $X2=4.35
+ $Y2=2.4
r96 1 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.67 $X2=3.9
+ $Y2=1.505
r97 1 3 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=3.9 $Y=1.67 $X2=3.9
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%VPWR 1 2 3 4 13 15 19 21 23 33 40 41 47 52
+ 60 62
r52 71 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r53 65 68 3.36552 $w=1.303e-06 $l=3.6e-07 $layer=LI1_cond $X=5.112 $Y=2.455
+ $X2=5.112 $Y2=2.815
r54 62 65 3.17854 $w=1.303e-06 $l=3.4e-07 $layer=LI1_cond $X=5.112 $Y=2.115
+ $X2=5.112 $Y2=2.455
r55 59 60 13.0375 $w=1.123e-06 $l=1.2e-07 $layer=LI1_cond $X=3.67 $Y=2.852
+ $X2=3.79 $Y2=2.852
r56 56 59 0.759111 $w=1.123e-06 $l=7e-08 $layer=LI1_cond $X=3.6 $Y=2.852
+ $X2=3.67 $Y2=2.852
r57 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 54 56 10.248 $w=1.123e-06 $l=9.45e-07 $layer=LI1_cond $X=2.655 $Y=2.852
+ $X2=3.6 $Y2=2.852
r59 50 54 0.162667 $w=1.123e-06 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=2.655 $Y2=2.852
r60 50 52 12.8748 $w=1.123e-06 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=2.535 $Y2=2.852
r61 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 41 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r65 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r66 38 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33 $X2=6
+ $Y2=3.33
r67 37 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r68 37 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 36 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.79 $Y2=3.33
r70 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 33 38 13.5804 $w=1.7e-07 $l=6.53e-07 $layer=LI1_cond $X=5.112 $Y=3.33
+ $X2=5.765 $Y2=3.33
r72 33 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 33 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 33 68 4.81456 $w=1.303e-06 $l=5.15e-07 $layer=LI1_cond $X=5.112 $Y=3.33
+ $X2=5.112 $Y2=2.815
r75 33 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 31 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.535 $Y2=3.33
r79 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 29 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.7 $Y2=3.33
r81 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 27 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 27 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 24 44 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r86 24 26 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r87 23 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.7 $Y2=3.33
r88 23 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.2 $Y2=3.33
r89 21 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r90 21 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r91 17 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=3.245 $X2=1.7
+ $Y2=3.33
r92 17 19 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.7 $Y=3.245 $X2=1.7
+ $Y2=2.455
r93 13 44 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r94 13 15 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.395
r95 4 68 200 $w=1.7e-07 $l=1.19106e-06 $layer=licon1_PDIFF $count=3 $X=4.44
+ $Y=1.84 $X2=4.92 $Y2=2.815
r96 4 65 200 $w=1.7e-07 $l=1.43492e-06 $layer=licon1_PDIFF $count=3 $X=4.44
+ $Y=1.84 $X2=5.6 $Y2=2.455
r97 4 65 200 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=3 $X=4.44
+ $Y=1.84 $X2=4.58 $Y2=2.455
r98 4 62 200 $w=1.7e-07 $l=6.01997e-07 $layer=licon1_PDIFF $count=3 $X=4.44
+ $Y=1.84 $X2=4.92 $Y2=2.115
r99 3 59 200 $w=1.7e-07 $l=1.42981e-06 $layer=licon1_PDIFF $count=3 $X=2.515
+ $Y=1.84 $X2=3.67 $Y2=2.455
r100 3 54 200 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=3 $X=2.515
+ $Y=1.84 $X2=2.655 $Y2=2.455
r101 2 19 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.84 $X2=1.7 $Y2=2.455
r102 1 15 300 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%Y 1 2 3 4 5 16 17 18 19 22 26 28 30 34 38 40
+ 42 44 48 50 52 55 56
c95 28 0 9.50231e-20 $X=1.395 $Y=1.095
r96 55 56 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r97 47 56 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.95
+ $X2=0.24 $Y2=1.665
r98 46 55 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r99 42 54 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.125 $Y=2.12
+ $X2=4.125 $Y2=1.97
r100 42 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.125 $Y=2.12
+ $X2=4.125 $Y2=2.815
r101 41 52 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.365 $Y=2.035
+ $X2=2.2 $Y2=1.97
r102 40 54 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=4.125 $Y2=1.97
r103 40 41 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=2.365 $Y2=2.035
r104 36 52 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=2.2 $Y=2.12 $X2=2.2
+ $Y2=1.97
r105 36 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.2 $Y=2.12
+ $X2=2.2 $Y2=2.815
r106 32 34 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.56 $Y=1.01
+ $X2=1.56 $Y2=0.68
r107 31 50 14.1623 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=1.365 $Y=2.035
+ $X2=0.99 $Y2=2.035
r108 30 52 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=2.2 $Y2=1.97
r109 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=1.365 $Y2=2.035
r110 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=1.095
+ $X2=0.7 $Y2=1.095
r111 28 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.395 $Y=1.095
+ $X2=1.56 $Y2=1.01
r112 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.395 $Y=1.095
+ $X2=0.865 $Y2=1.095
r113 24 50 3.00456 $w=7.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=2.12
+ $X2=0.99 $Y2=2.035
r114 24 26 11.0837 $w=7.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.99 $Y=2.12
+ $X2=0.99 $Y2=2.815
r115 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.01 $X2=0.7
+ $Y2=1.095
r116 20 22 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.7 $Y=1.01 $X2=0.7
+ $Y2=0.68
r117 19 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.035
+ $X2=0.24 $Y2=1.95
r118 18 50 14.1623 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.99 $Y2=2.035
r119 18 19 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.355 $Y2=2.035
r120 17 46 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.095
+ $X2=0.24 $Y2=1.18
r121 16 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=1.095
+ $X2=0.7 $Y2=1.095
r122 16 17 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.535 $Y=1.095
+ $X2=0.355 $Y2=1.095
r123 5 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.125 $Y2=1.985
r124 5 44 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.125 $Y2=2.815
r125 4 52 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.84 $X2=2.2 $Y2=1.985
r126 4 38 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.84 $X2=2.2 $Y2=2.815
r127 3 50 200 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=3 $X=0.595
+ $Y=1.84 $X2=0.735 $Y2=2.115
r128 3 26 200 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=3 $X=0.595
+ $Y=1.84 $X2=0.735 $Y2=2.815
r129 2 34 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.41 $X2=1.56 $Y2=0.68
r130 1 22 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.41 $X2=0.7 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%A_27_82# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 45 46
r66 40 42 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=3.745 $Y=0.425
+ $X2=3.745 $Y2=0.57
r67 39 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.85 $Y2=0.34
r68 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.615 $Y=0.34
+ $X2=3.745 $Y2=0.425
r69 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.615 $Y=0.34
+ $X2=2.945 $Y2=0.34
r70 34 46 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=0.425
+ $X2=2.85 $Y2=0.34
r71 34 36 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.85 $Y=0.425
+ $X2=2.85 $Y2=0.57
r72 33 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.34
+ $X2=1.99 $Y2=0.34
r73 32 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.755 $Y=0.34
+ $X2=2.85 $Y2=0.34
r74 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.755 $Y=0.34
+ $X2=2.075 $Y2=0.34
r75 28 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.425
+ $X2=1.99 $Y2=0.34
r76 28 30 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.99 $Y=0.425
+ $X2=1.99 $Y2=0.555
r77 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.34
+ $X2=1.13 $Y2=0.34
r78 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=0.34
+ $X2=1.99 $Y2=0.34
r79 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.905 $Y=0.34
+ $X2=1.215 $Y2=0.34
r80 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.13 $Y2=0.34
r81 22 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.13 $Y2=0.615
r82 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.13 $Y2=0.34
r83 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.355 $Y2=0.34
r84 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=0.425
+ $X2=0.355 $Y2=0.34
r85 16 18 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.23 $Y=0.425
+ $X2=0.23 $Y2=0.615
r86 5 42 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.41 $X2=3.71 $Y2=0.57
r87 4 36 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.41 $X2=2.85 $Y2=0.57
r88 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.85
+ $Y=0.41 $X2=1.99 $Y2=0.555
r89 2 24 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.41 $X2=1.13 $Y2=0.615
r90 1 18 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.41 $X2=0.27 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%A_456_82# 1 2 3 4 13 15 19 21 23 25 28 33 38
c66 23 0 1.6164e-19 $X=5.54 $Y=0.92
c67 15 0 1.20944e-20 $X=4.585 $Y=1.045
c68 13 0 2.41975e-20 $X=3.115 $Y=1.045
r69 33 35 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.28 $Y=0.68
+ $X2=3.28 $Y2=1.045
r70 28 30 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.42 $Y=0.68
+ $X2=2.42 $Y2=1.045
r71 23 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.54 $Y=0.92
+ $X2=5.54 $Y2=1.045
r72 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.54 $Y=0.92
+ $X2=5.54 $Y2=0.555
r73 22 38 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.775 $Y=1.045
+ $X2=4.68 $Y2=1.045
r74 21 40 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.455 $Y=1.045
+ $X2=5.54 $Y2=1.045
r75 21 22 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=5.455 $Y=1.045
+ $X2=4.775 $Y2=1.045
r76 17 38 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.68 $Y=0.92
+ $X2=4.68 $Y2=1.045
r77 17 19 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=4.68 $Y=0.92
+ $X2=4.68 $Y2=0.555
r78 16 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=1.045
+ $X2=3.28 $Y2=1.045
r79 15 38 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.585 $Y=1.045
+ $X2=4.68 $Y2=1.045
r80 15 16 52.5514 $w=2.48e-07 $l=1.14e-06 $layer=LI1_cond $X=4.585 $Y=1.045
+ $X2=3.445 $Y2=1.045
r81 14 30 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=1.045
+ $X2=2.42 $Y2=1.045
r82 13 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=1.045
+ $X2=3.28 $Y2=1.045
r83 13 14 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=3.115 $Y=1.045
+ $X2=2.585 $Y2=1.045
r84 4 40 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.41 $X2=5.54 $Y2=1.005
r85 4 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.41 $X2=5.54 $Y2=0.555
r86 3 38 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.54
+ $Y=0.41 $X2=4.68 $Y2=1.005
r87 3 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.54
+ $Y=0.41 $X2=4.68 $Y2=0.555
r88 2 33 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.41 $X2=3.28 $Y2=0.68
r89 1 28 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=2.28
+ $Y=0.41 $X2=2.42 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3_4%VGND 1 2 3 12 16 18 20 23 24 25 34 38 44 48
r67 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r68 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r69 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r70 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r71 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r72 39 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.11
+ $Y2=0
r73 39 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.52
+ $Y2=0
r74 38 47 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=5.805 $Y=0 $X2=6.022
+ $Y2=0
r75 38 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.805 $Y=0 $X2=5.52
+ $Y2=0
r76 37 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r77 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 34 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.11
+ $Y2=0
r79 34 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=4.56
+ $Y2=0
r80 33 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r81 32 33 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r82 28 32 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r83 28 29 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r84 25 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r85 25 29 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=0.24
+ $Y2=0
r86 23 32 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.08
+ $Y2=0
r87 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.25
+ $Y2=0
r88 22 36 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.415 $Y=0 $X2=4.56
+ $Y2=0
r89 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=0 $X2=4.25
+ $Y2=0
r90 18 47 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=6.022 $Y2=0
r91 18 20 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.555
r92 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=0.085
+ $X2=5.11 $Y2=0
r93 14 16 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=5.11 $Y=0.085 $X2=5.11
+ $Y2=0.585
r94 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0.085
+ $X2=4.25 $Y2=0
r95 10 12 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.25 $Y=0.085 $X2=4.25
+ $Y2=0.585
r96 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.83
+ $Y=0.41 $X2=5.97 $Y2=0.555
r97 2 16 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.41 $X2=5.11 $Y2=0.585
r98 1 12 182 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_NDIFF $count=1 $X=4.115
+ $Y=0.41 $X2=4.25 $Y2=0.585
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__clkinv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  5.040000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.985000 1.180000 10.935000 1.410000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  5.040000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575000 1.920000 10.935000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.115000  0.085000  0.445000 0.840000 ;
      RECT  0.115000  1.900000  0.445000 3.245000 ;
      RECT  0.615000  0.380000  0.805000 0.775000 ;
      RECT  0.625000  0.775000  0.805000 1.820000 ;
      RECT  0.625000  1.820000  0.815000 2.980000 ;
      RECT  0.975000  0.085000  1.260000 0.840000 ;
      RECT  0.975000  1.150000  1.295000 1.650000 ;
      RECT  1.015000  1.820000  1.265000 3.245000 ;
      RECT  1.440000  0.380000  1.700000 0.775000 ;
      RECT  1.465000  0.775000  1.695000 1.885000 ;
      RECT  1.465000  1.885000  1.795000 2.980000 ;
      RECT  1.865000  1.150000  2.195000 1.650000 ;
      RECT  1.885000  0.085000  2.165000 0.840000 ;
      RECT  1.995000  1.820000  2.165000 3.245000 ;
      RECT  2.350000  0.380000  2.665000 0.775000 ;
      RECT  2.365000  0.775000  2.665000 1.885000 ;
      RECT  2.365000  1.885000  2.695000 2.980000 ;
      RECT  2.835000  1.150000  3.165000 1.650000 ;
      RECT  2.845000  0.085000  3.095000 0.840000 ;
      RECT  2.895000  1.820000  3.065000 3.245000 ;
      RECT  3.300000  0.380000  3.595000 0.775000 ;
      RECT  3.335000  0.775000  3.595000 2.980000 ;
      RECT  3.765000  0.085000  4.095000 0.840000 ;
      RECT  3.765000  1.150000  4.095000 1.650000 ;
      RECT  3.795000  1.820000  3.965000 3.245000 ;
      RECT  4.165000  1.850000  4.525000 1.900000 ;
      RECT  4.165000  1.900000  4.495000 2.980000 ;
      RECT  4.265000  0.380000  4.525000 1.850000 ;
      RECT  4.695000  1.820000  4.865000 3.245000 ;
      RECT  4.755000  1.150000  5.085000 1.650000 ;
      RECT  4.765000  0.085000  5.085000 0.840000 ;
      RECT  5.065000  1.850000  5.425000 2.010000 ;
      RECT  5.065000  2.010000  5.395000 2.980000 ;
      RECT  5.255000  0.380000  5.525000 0.775000 ;
      RECT  5.255000  0.775000  5.425000 1.850000 ;
      RECT  5.595000  1.150000  5.925000 1.650000 ;
      RECT  5.595000  1.820000  5.845000 3.245000 ;
      RECT  5.695000  0.085000  5.980000 0.840000 ;
      RECT  6.015000  1.820000  6.330000 2.980000 ;
      RECT  6.095000  1.010000  6.340000 1.760000 ;
      RECT  6.095000  1.760000  6.330000 1.820000 ;
      RECT  6.160000  0.380000  6.385000 0.785000 ;
      RECT  6.160000  0.785000  6.340000 1.010000 ;
      RECT  6.510000  1.820000  6.795000 3.245000 ;
      RECT  6.545000  1.150000  6.875000 1.650000 ;
      RECT  6.555000  0.085000  6.875000 0.840000 ;
      RECT  7.045000  0.380000  7.290000 2.980000 ;
      RECT  7.475000  1.820000  7.805000 3.245000 ;
      RECT  7.485000  0.085000  9.825000 0.710000 ;
      RECT  7.525000  1.150000 10.915000 1.650000 ;
      RECT  8.005000  1.820000  8.175000 2.980000 ;
      RECT  8.375000  1.820000  8.625000 3.245000 ;
      RECT  8.905000  1.820000  9.075000 2.980000 ;
      RECT  9.275000  1.820000  9.605000 3.245000 ;
      RECT  9.805000  1.820000  9.975000 2.980000 ;
      RECT 10.175000  1.820000 10.505000 3.245000 ;
      RECT 10.705000  1.820000 10.875000 2.980000 ;
      RECT 11.075000  1.820000 11.405000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  1.950000  0.805000 2.120000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.045000  1.210000  1.215000 1.380000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.545000  1.950000  1.715000 2.120000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  1.945000  1.210000  2.115000 1.380000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.445000  1.950000  2.615000 2.120000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  2.915000  1.210000  3.085000 1.380000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.375000  1.950000  3.545000 2.120000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.845000  1.210000  4.015000 1.380000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.245000  1.950000  4.415000 2.120000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.835000  1.210000  5.005000 1.380000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.145000  1.950000  5.315000 2.120000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.675000  1.210000  5.845000 1.380000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.095000  1.950000  6.265000 2.120000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.625000  1.210000  6.795000 1.380000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.075000  1.950000  7.245000 2.120000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.745000  1.210000  7.915000 1.380000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.005000  1.950000  8.175000 2.120000 ;
      RECT  8.105000  1.210000  8.275000 1.380000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.465000  1.210000  8.635000 1.380000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  8.825000  1.210000  8.995000 1.380000 ;
      RECT  8.905000  1.950000  9.075000 2.120000 ;
      RECT  9.185000  1.210000  9.355000 1.380000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.545000  1.210000  9.715000 1.380000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.805000  1.950000  9.975000 2.120000 ;
      RECT  9.905000  1.210000 10.075000 1.380000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.265000  1.210000 10.435000 1.380000 ;
      RECT 10.625000  1.210000 10.795000 1.380000 ;
      RECT 10.705000  1.950000 10.875000 2.120000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
  END
END sky130_fd_sc_ms__clkinv_16
END LIBRARY

* File: sky130_fd_sc_ms__a211o_4.spice
* Created: Fri Aug 28 16:56:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a211o_4.pex.spice"
.subckt sky130_fd_sc_ms__a211o_4  VNB VPB B1 C1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_105_280#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1001_d N_A_105_280#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1008_d N_A_105_280#_M1008_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1019 N_X_M1008_d N_A_105_280#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_105_280#_M1005_d N_B1_M1005_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.113206 PD=0.92 PS=1.00174 NRD=0 NRS=11.712 M=1 R=4.26667
+ SA=75002 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1020 N_A_105_280#_M1005_d N_C1_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.114925 PD=0.92 PS=1.05 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.4
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1021 N_A_105_280#_M1021_d N_C1_M1021_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.110562 AS=0.114925 PD=1.04 PS=1.05 NRD=4.68 NRS=12.18 M=1 R=4.26667
+ SA=75002.6 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1013 N_A_105_280#_M1021_d N_B1_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.110562 AS=0.2304 PD=1.04 PS=1.36 NRD=3.744 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1000 N_A_1064_123#_M1000_d N_A2_M1000_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2304 PD=0.92 PS=1.36 NRD=0 NRS=82.5 M=1 R=4.26667
+ SA=75003.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_105_280#_M1002_d N_A1_M1002_g N_A_1064_123#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1017 N_A_105_280#_M1002_d N_A1_M1017_g N_A_1064_123#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.4 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_1064_123#_M1017_s N_A2_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_X_M1006_d N_A_105_280#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1006_d N_A_105_280#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1015 N_X_M1015_d N_A_105_280#_M1015_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1016 N_X_M1015_d N_A_105_280#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1010 N_A_605_392#_M1010_d N_B1_M1010_g N_A_517_392#_M1010_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.26 PD=1.32 PS=2.52 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90003.8 A=0.18 P=2.36 MULT=1
MM1009 N_A_105_280#_M1009_d N_C1_M1009_g N_A_605_392#_M1010_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1012 N_A_105_280#_M1009_d N_C1_M1012_g N_A_605_392#_M1012_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.1475 PD=1.27 PS=1.295 NRD=0 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1018 N_A_605_392#_M1012_s N_B1_M1018_g N_A_517_392#_M1018_s VPB PSHORT L=0.18
+ W=1 AD=0.1475 AS=0.1375 PD=1.295 PS=1.275 NRD=1.9503 NRS=0 M=1 R=5.55556
+ SA=90001.6 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1004 N_A_517_392#_M1018_s N_A2_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1
+ AD=0.1375 AS=0.3125 PD=1.275 PS=1.625 NRD=0 NRS=0 M=1 R=5.55556 SA=90002
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1004_s N_A1_M1003_g N_A_517_392#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.3125 AS=0.135 PD=1.625 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.9
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1022_d N_A1_M1022_g N_A_517_392#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90003.3
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1014 N_A_517_392#_M1014_d N_A2_M1014_g N_VPWR_M1022_d VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90003.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ms__a211o_4.pxi.spice"
*
.ends
*
*

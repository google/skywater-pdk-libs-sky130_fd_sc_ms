* File: sky130_fd_sc_ms__sdfrbp_1.spice
* Created: Wed Sep  2 12:30:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfrbp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfrbp_1  VNB VPB SCE D SCD CLK RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1038 N_VGND_M1038_d N_SCE_M1038_g N_A_27_74#_M1038_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 noxref_26 N_A_27_74#_M1023_g N_noxref_25_M1023_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.07455 AS=0.1197 PD=0.775 PS=1.41 NRD=34.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_413_90#_M1002_d N_D_M1002_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.107537 AS=0.07455 PD=0.965 PS=0.775 NRD=65.712 NRS=34.992 M=1 R=2.8
+ SA=75000.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1032 noxref_27 N_SCE_M1032_g N_A_413_90#_M1002_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.107537 PD=0.63 PS=0.965 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1022 N_noxref_25_M1022_d N_SCD_M1022_g noxref_27 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0721875 AS=0.0441 PD=0.79 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_RESET_B_M1028_g N_noxref_25_M1022_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0721875 PD=1.37 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75002 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_CLK_M1013_g N_A_819_119#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.179025 AS=0.254 PD=1.335 PS=2.22 NRD=12.156 NRS=2.424 M=1
+ R=4.93333 SA=75000.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_1037_119#_M1014_d N_A_819_119#_M1014_g N_VGND_M1013_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1998 AS=0.179025 PD=2.02 PS=1.335 NRD=0 NRS=12.156 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_1235_119#_M1031_d N_A_819_119#_M1031_g N_A_413_90#_M1031_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1036 A_1321_119# N_A_1037_119#_M1036_g N_A_1235_119#_M1031_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1004 A_1399_119# N_A_1369_93#_M1004_g A_1321_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_RESET_B_M1034_g A_1399_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.209713 AS=0.0504 PD=1.26 PS=0.66 NRD=126.936 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1041 N_A_1369_93#_M1041_d N_A_1235_119#_M1041_g N_VGND_M1034_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.319562 PD=0.92 PS=1.92 NRD=0 NRS=83.304 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1029 N_A_1747_74#_M1029_d N_A_1037_119#_M1029_g N_A_1369_93#_M1041_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.272845 AS=0.0896 PD=1.91396 PS=0.92 NRD=92.808 NRS=0
+ M=1 R=4.26667 SA=75002.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1016 A_1966_74# N_A_819_119#_M1016_g N_A_1747_74#_M1029_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.179055 PD=0.63 PS=1.25604 NRD=14.28 NRS=48.564 M=1 R=2.8
+ SA=75002.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_2008_48#_M1005_g A_1966_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1009 A_2124_74# N_RESET_B_M1009_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_2008_48#_M1012_d N_A_1747_74#_M1012_g A_2124_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_Q_N_M1010_d N_A_1747_74#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.3159 PD=2.04 PS=2.57 NRD=0 NRS=60.3 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_1747_74#_M1003_g N_A_2513_424#_M1003_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.101196 AS=0.14575 PD=0.92093 PS=1.63 NRD=13.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1037 N_Q_M1037_d N_A_2513_424#_M1037_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.136154 PD=2.05 PS=1.23907 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_VPWR_M1018_d N_SCE_M1018_g N_A_27_74#_M1018_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.5696 PD=0.96 PS=3.06 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.8
+ SB=90002.7 A=0.1152 P=1.64 MULT=1
MM1017 A_341_464# N_SCE_M1017_g N_VPWR_M1018_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90001.3
+ SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1027 N_A_413_90#_M1027_d N_D_M1027_g A_341_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.7
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1030 A_515_464# N_A_27_74#_M1030_g N_A_413_90#_M1027_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1152 AS=0.0864 PD=1 PS=0.91 NRD=38.4741 NRS=0 M=1 R=3.55556
+ SA=90002.2 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1001 N_VPWR_M1001_d N_SCD_M1001_g A_515_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1248 AS=0.1152 PD=1.03 PS=1 NRD=3.0732 NRS=38.4741 M=1 R=3.55556
+ SA=90002.7 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1011 N_A_413_90#_M1011_d N_RESET_B_M1011_g N_VPWR_M1001_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.1248 PD=1.84 PS=1.03 NRD=0 NRS=30.7714 M=1 R=3.55556
+ SA=90003.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1025 N_VPWR_M1025_d N_CLK_M1025_g N_A_819_119#_M1025_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1035 N_A_1037_119#_M1035_d N_A_819_119#_M1035_g N_VPWR_M1025_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1019 N_A_1235_119#_M1019_d N_A_1037_119#_M1019_g N_A_413_90#_M1019_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.0567 AS=0.1134 PD=0.69 PS=1.38 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1024 A_1331_463# N_A_819_119#_M1024_g N_A_1235_119#_M1019_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_1369_93#_M1006_g A_1331_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.119925 AS=0.0441 PD=1.075 PS=0.63 NRD=108.114 NRS=23.443 M=1 R=2.33333
+ SA=90001 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1040 N_A_1235_119#_M1040_d N_RESET_B_M1040_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1134 AS=0.119925 PD=1.38 PS=1.075 NRD=0 NRS=108.114 M=1 R=2.33333
+ SA=90001.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1007 N_A_1369_93#_M1007_d N_A_1235_119#_M1007_g N_VPWR_M1007_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1015 N_A_1747_74#_M1015_d N_A_819_119#_M1015_g N_A_1369_93#_M1007_d VPB PSHORT
+ L=0.18 W=1 AD=0.277148 AS=0.135 PD=2.42958 PS=1.27 NRD=20.3501 NRS=0 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1033 A_1972_489# N_A_1037_119#_M1033_g N_A_1747_74#_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.116402 PD=0.63 PS=1.02042 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90001 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1039 N_VPWR_M1039_d N_A_2008_48#_M1039_g A_1972_489# VPB PSHORT L=0.18 W=0.42
+ AD=0.111562 AS=0.0441 PD=0.98 PS=0.63 NRD=42.1974 NRS=23.443 M=1 R=2.33333
+ SA=90001.4 SB=90002 A=0.0756 P=1.2 MULT=1
MM1020 N_A_2008_48#_M1020_d N_RESET_B_M1020_g N_VPWR_M1039_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.111562 PD=0.69 PS=0.98 NRD=0 NRS=44.5417 M=1 R=2.33333
+ SA=90002.1 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1021 N_VPWR_M1021_d N_A_1747_74#_M1021_g N_A_2008_48#_M1020_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.115309 AS=0.0567 PD=0.883636 PS=0.69 NRD=68.0044 NRS=0 M=1
+ R=2.33333 SA=90002.5 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1026 N_Q_N_M1026_d N_A_1747_74#_M1026_g N_VPWR_M1021_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.307491 PD=2.8 PS=2.35636 NRD=0 NRS=9.3772 M=1 R=6.22222
+ SA=90001.3 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A_1747_74#_M1008_g N_A_2513_424#_M1008_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1536 AS=0.2184 PD=1.25143 PS=2.2 NRD=7.0329 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1000 N_Q_M1000_d N_A_2513_424#_M1000_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2048 PD=2.76 PS=1.66857 NRD=0 NRS=3.2111 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX42_noxref VNB VPB NWDIODE A=26.7791 P=32.56
*
.include "sky130_fd_sc_ms__sdfrbp_1.pxi.spice"
*
.ends
*
*

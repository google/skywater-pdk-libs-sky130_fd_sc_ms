* File: sky130_fd_sc_ms__nand3b_4.pxi.spice
* Created: Wed Sep  2 12:14:03 2020
* 
x_PM_SKY130_FD_SC_MS__NAND3B_4%A_N N_A_N_M1000_g N_A_N_c_104_n N_A_N_M1017_g
+ N_A_N_c_101_n N_A_N_c_106_n N_A_N_M1020_g A_N N_A_N_c_102_n N_A_N_c_103_n
+ PM_SKY130_FD_SC_MS__NAND3B_4%A_N
x_PM_SKY130_FD_SC_MS__NAND3B_4%C N_C_c_151_n N_C_M1006_g N_C_c_152_n N_C_c_153_n
+ N_C_c_154_n N_C_M1010_g N_C_c_155_n N_C_M1011_g N_C_M1001_g N_C_M1018_g
+ N_C_c_156_n N_C_M1012_g N_C_c_157_n C C C N_C_c_159_n
+ PM_SKY130_FD_SC_MS__NAND3B_4%C
x_PM_SKY130_FD_SC_MS__NAND3B_4%A_89_172# N_A_89_172#_M1000_s N_A_89_172#_M1017_d
+ N_A_89_172#_M1008_g N_A_89_172#_c_230_n N_A_89_172#_M1005_g
+ N_A_89_172#_M1009_g N_A_89_172#_c_232_n N_A_89_172#_M1013_g
+ N_A_89_172#_c_233_n N_A_89_172#_c_234_n N_A_89_172#_M1014_g
+ N_A_89_172#_c_235_n N_A_89_172#_c_236_n N_A_89_172#_M1019_g
+ N_A_89_172#_c_237_n N_A_89_172#_c_238_n N_A_89_172#_c_251_n
+ N_A_89_172#_c_239_n N_A_89_172#_c_240_n N_A_89_172#_c_241_n
+ N_A_89_172#_c_242_n N_A_89_172#_c_278_n N_A_89_172#_c_243_n
+ N_A_89_172#_c_244_n PM_SKY130_FD_SC_MS__NAND3B_4%A_89_172#
x_PM_SKY130_FD_SC_MS__NAND3B_4%B N_B_c_364_n N_B_M1002_g N_B_c_356_n N_B_c_357_n
+ N_B_M1003_g N_B_c_367_n N_B_M1004_g N_B_M1007_g N_B_M1015_g N_B_M1016_g B B B
+ N_B_c_362_n N_B_c_363_n PM_SKY130_FD_SC_MS__NAND3B_4%B
x_PM_SKY130_FD_SC_MS__NAND3B_4%VPWR N_VPWR_M1017_s N_VPWR_M1020_s N_VPWR_M1018_d
+ N_VPWR_M1009_d N_VPWR_M1004_s N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n
+ N_VPWR_c_427_n VPWR N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_430_n
+ N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_423_n
+ PM_SKY130_FD_SC_MS__NAND3B_4%VPWR
x_PM_SKY130_FD_SC_MS__NAND3B_4%Y N_Y_M1005_s N_Y_M1014_s N_Y_M1001_s N_Y_M1008_s
+ N_Y_M1002_d N_Y_c_495_n N_Y_c_496_n N_Y_c_492_n N_Y_c_497_n N_Y_c_500_n
+ N_Y_c_541_n Y Y Y N_Y_c_494_n PM_SKY130_FD_SC_MS__NAND3B_4%Y
x_PM_SKY130_FD_SC_MS__NAND3B_4%VGND N_VGND_M1000_d N_VGND_M1010_s N_VGND_M1012_s
+ N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n N_VGND_c_560_n VGND
+ N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n
+ PM_SKY130_FD_SC_MS__NAND3B_4%VGND
x_PM_SKY130_FD_SC_MS__NAND3B_4%A_297_82# N_A_297_82#_M1006_d N_A_297_82#_M1011_d
+ N_A_297_82#_M1003_s N_A_297_82#_M1015_s N_A_297_82#_c_624_n
+ N_A_297_82#_c_625_n N_A_297_82#_c_639_n N_A_297_82#_c_631_n
+ N_A_297_82#_c_696_n N_A_297_82#_c_641_n N_A_297_82#_c_707_n
+ N_A_297_82#_c_650_n N_A_297_82#_c_664_n N_A_297_82#_c_681_n
+ N_A_297_82#_c_632_n N_A_297_82#_c_633_n N_A_297_82#_c_626_n
+ N_A_297_82#_c_627_n N_A_297_82#_c_628_n N_A_297_82#_c_629_n
+ PM_SKY130_FD_SC_MS__NAND3B_4%A_297_82#
x_PM_SKY130_FD_SC_MS__NAND3B_4%A_744_74# N_A_744_74#_M1005_d N_A_744_74#_M1013_d
+ N_A_744_74#_M1019_d N_A_744_74#_M1007_d N_A_744_74#_M1016_d
+ N_A_744_74#_c_749_n N_A_744_74#_c_750_n N_A_744_74#_c_751_n
+ N_A_744_74#_c_752_n PM_SKY130_FD_SC_MS__NAND3B_4%A_744_74#
cc_1 VNB N_A_N_M1000_g 0.0287326f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.78
cc_2 VNB N_A_N_c_101_n 0.0107003f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.69
cc_3 VNB N_A_N_c_102_n 0.00482071f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_4 VNB N_A_N_c_103_n 0.0526828f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.557
cc_5 VNB N_C_c_151_n 0.0150735f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.35
cc_6 VNB N_C_c_152_n 0.0210958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C_c_153_n 0.00896832f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.765
cc_8 VNB N_C_c_154_n 0.0158871f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.26
cc_9 VNB N_C_c_155_n 0.0164552f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.69
cc_10 VNB N_C_c_156_n 0.059874f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_11 VNB N_C_c_157_n 0.0132043f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.665
cc_12 VNB C 0.00633246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_159_n 0.0375955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_89_172#_M1008_g 0.00211793f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.69
cc_15 VNB N_A_89_172#_c_230_n 0.0173647f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.26
cc_16 VNB N_A_89_172#_M1009_g 0.00213854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_89_172#_c_232_n 0.0152147f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.557
cc_18 VNB N_A_89_172#_c_233_n 0.015184f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.557
cc_19 VNB N_A_89_172#_c_234_n 0.014791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_89_172#_c_235_n 0.0241507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_89_172#_c_236_n 0.015888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_89_172#_c_237_n 0.00678911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_89_172#_c_238_n 0.00339641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_89_172#_c_239_n 0.00551243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_89_172#_c_240_n 0.03265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_89_172#_c_241_n 0.00351706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_89_172#_c_242_n 0.00467773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_89_172#_c_243_n 0.00586556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_89_172#_c_244_n 0.0953027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_356_n 0.0113503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_c_357_n 0.0101726f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.765
cc_32 VNB N_B_M1003_g 0.0220707f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=1.69
cc_33 VNB N_B_M1007_g 0.0209473f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.557
cc_34 VNB N_B_M1015_g 0.0209424f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_35 VNB N_B_M1016_g 0.0278788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_c_362_n 0.0850853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_363_n 0.00991188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_423_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_492_n 0.0100981f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.665
cc_40 VNB Y 0.00834423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_494_n 0.00413956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_557_n 0.0145618f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.26
cc_43 VNB N_VGND_c_558_n 0.0450868f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.557
cc_44 VNB N_VGND_c_559_n 0.0184795f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.515
cc_45 VNB N_VGND_c_560_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_561_n 0.0179406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_562_n 0.10598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_563_n 0.422046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_564_n 0.0209864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_297_82#_c_624_n 0.0446775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_297_82#_c_625_n 0.0100851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_297_82#_c_626_n 0.0200968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_297_82#_c_627_n 0.0103159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_297_82#_c_628_n 0.00255379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_297_82#_c_629_n 0.00296506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_744_74#_c_749_n 0.00258449f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_57 VNB N_A_744_74#_c_750_n 0.0237054f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.665
cc_58 VNB N_A_744_74#_c_751_n 0.00534237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_744_74#_c_752_n 0.00766753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_A_N_c_104_n 0.0185567f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.765
cc_61 VPB N_A_N_c_101_n 0.00823689f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=1.69
cc_62 VPB N_A_N_c_106_n 0.0190716f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.765
cc_63 VPB N_A_N_c_102_n 0.00488844f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_64 VPB N_A_N_c_103_n 0.0215841f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.557
cc_65 VPB N_C_M1001_g 0.0253908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_C_M1018_g 0.0216595f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.557
cc_67 VPB N_C_c_156_n 0.00489206f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_68 VPB N_C_c_157_n 0.00490368f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.665
cc_69 VPB C 0.0174982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_C_c_159_n 0.0183479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_89_172#_M1008_g 0.0276387f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.69
cc_72 VPB N_A_89_172#_M1009_g 0.0290702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_B_c_364_n 0.0210416f $X=-0.19 $Y=1.66 $X2=0.805 $Y2=1.35
cc_74 VPB N_B_c_356_n 0.0032339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_B_c_357_n 0.00299068f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.765
cc_76 VPB N_B_c_367_n 0.0232721f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.765
cc_77 VPB N_B_c_362_n 0.0407356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_424_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_425_n 0.0528544f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.557
cc_80 VPB N_VPWR_c_426_n 0.00408418f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.515
cc_81 VPB N_VPWR_c_427_n 0.0165163f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.665
cc_82 VPB N_VPWR_c_428_n 0.017758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_429_n 0.0331904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_430_n 0.0457448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_431_n 0.00910695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_432_n 0.0298504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_433_n 0.0228918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_434_n 0.0934196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_423_n 0.0811708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_Y_c_495_n 0.00818226f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_91 VPB N_Y_c_496_n 0.00112215f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.557
cc_92 VPB N_Y_c_497_n 0.0105296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB Y 0.00476158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_297_82#_c_624_n 0.0127365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_297_82#_c_631_n 0.00866242f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.557
cc_96 VPB N_A_297_82#_c_632_n 0.0080099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_297_82#_c_633_n 0.00120381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_297_82#_c_626_n 0.0102237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 N_A_N_M1000_g N_C_c_151_n 0.0258441f $X=0.805 $Y=0.78 $X2=-0.19 $Y2=-0.245
cc_100 N_A_N_c_101_n N_C_c_153_n 0.00556329f $X=1.255 $Y=1.69 $X2=0 $Y2=0
cc_101 N_A_N_c_103_n N_C_c_153_n 0.00139393f $X=1.095 $Y=1.557 $X2=0 $Y2=0
cc_102 N_A_N_c_101_n N_C_c_157_n 0.00248024f $X=1.255 $Y=1.69 $X2=0 $Y2=0
cc_103 N_A_N_c_103_n N_C_c_157_n 0.00268185f $X=1.095 $Y=1.557 $X2=0 $Y2=0
cc_104 N_A_N_c_101_n C 0.00264236f $X=1.255 $Y=1.69 $X2=0 $Y2=0
cc_105 N_A_N_M1000_g N_A_89_172#_c_238_n 0.00915372f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_106 N_A_N_c_101_n N_A_89_172#_c_238_n 0.00490597f $X=1.255 $Y=1.69 $X2=0
+ $Y2=0
cc_107 N_A_N_c_102_n N_A_89_172#_c_238_n 0.0256619f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_N_c_103_n N_A_89_172#_c_238_n 0.0014897f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_109 N_A_N_c_104_n N_A_89_172#_c_251_n 0.00300824f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_N_c_106_n N_A_89_172#_c_251_n 0.00872631f $X=1.345 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_N_c_102_n N_A_89_172#_c_251_n 0.00885832f $X=0.93 $Y=1.515 $X2=0
+ $Y2=0
cc_112 N_A_N_c_103_n N_A_89_172#_c_251_n 0.00253974f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_113 N_A_N_M1000_g N_A_89_172#_c_239_n 0.00291514f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_114 N_A_N_c_104_n N_A_89_172#_c_239_n 8.17481e-19 $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_N_c_101_n N_A_89_172#_c_239_n 0.00834478f $X=1.255 $Y=1.69 $X2=0
+ $Y2=0
cc_116 N_A_N_c_106_n N_A_89_172#_c_239_n 0.0114333f $X=1.345 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_N_c_102_n N_A_89_172#_c_239_n 0.0335776f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_N_c_103_n N_A_89_172#_c_239_n 0.00302054f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_119 N_A_N_M1000_g N_A_89_172#_c_242_n 0.0040074f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_120 N_A_N_c_102_n N_A_89_172#_c_242_n 0.0261451f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A_N_c_103_n N_A_89_172#_c_242_n 0.00220658f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_122 N_A_N_c_104_n N_VPWR_c_425_n 0.0110695f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_N_c_104_n N_VPWR_c_429_n 0.00482866f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_N_c_106_n N_VPWR_c_429_n 0.00482866f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_N_c_106_n N_VPWR_c_430_n 0.00671647f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_N_c_104_n N_VPWR_c_423_n 0.00555093f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_N_c_106_n N_VPWR_c_423_n 0.00555093f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_N_M1000_g N_VGND_c_558_n 0.00798327f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_129 N_A_N_M1000_g N_VGND_c_563_n 0.00533081f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_130 N_A_N_M1000_g N_A_297_82#_c_624_n 0.00747069f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_131 N_A_N_c_104_n N_A_297_82#_c_624_n 0.0040318f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_N_c_102_n N_A_297_82#_c_624_n 0.0342298f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_N_c_103_n N_A_297_82#_c_624_n 0.0108353f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_134 N_A_N_c_102_n N_A_297_82#_c_639_n 0.0282995f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A_N_c_103_n N_A_297_82#_c_639_n 0.00241497f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_136 N_A_N_c_104_n N_A_297_82#_c_641_n 0.0160698f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_N_c_106_n N_A_297_82#_c_641_n 0.01521f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_N_c_102_n N_A_297_82#_c_641_n 0.00471811f $X=0.93 $Y=1.515 $X2=0
+ $Y2=0
cc_139 N_A_N_M1000_g N_A_297_82#_c_627_n 0.0144512f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_140 N_A_N_M1000_g N_A_297_82#_c_628_n 0.00116196f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_141 N_C_c_156_n N_A_89_172#_M1008_g 0.0265873f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_142 N_C_c_151_n N_A_89_172#_c_239_n 0.00135568f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_143 N_C_c_153_n N_A_89_172#_c_239_n 0.00965829f $X=1.485 $Y=1.3 $X2=0 $Y2=0
cc_144 N_C_c_154_n N_A_89_172#_c_239_n 2.47368e-19 $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_145 N_C_c_157_n N_A_89_172#_c_239_n 0.00106338f $X=1.84 $Y=1.452 $X2=0 $Y2=0
cc_146 C N_A_89_172#_c_239_n 0.0204898f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_147 N_C_c_151_n N_A_89_172#_c_240_n 0.00544416f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_148 N_C_c_152_n N_A_89_172#_c_240_n 0.00392416f $X=1.765 $Y=1.3 $X2=0 $Y2=0
cc_149 N_C_c_154_n N_A_89_172#_c_240_n 0.0118156f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_150 N_C_c_155_n N_A_89_172#_c_240_n 0.0121942f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_151 N_C_c_156_n N_A_89_172#_c_240_n 0.0213471f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_152 C N_A_89_172#_c_240_n 0.111296f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_153 N_C_c_159_n N_A_89_172#_c_240_n 0.0116694f $X=2.515 $Y=1.452 $X2=0 $Y2=0
cc_154 N_C_c_151_n N_A_89_172#_c_242_n 4.85079e-19 $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_155 N_C_c_151_n N_A_89_172#_c_278_n 0.00624968f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_156 N_C_c_156_n N_A_89_172#_c_243_n 0.00201075f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_157 C N_A_89_172#_c_243_n 0.0127818f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_158 N_C_c_156_n N_A_89_172#_c_244_n 0.0265873f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_159 C N_A_89_172#_c_244_n 0.00601111f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_160 N_C_M1001_g N_VPWR_c_426_n 0.00128552f $X=2.625 $Y=2.4 $X2=0 $Y2=0
cc_161 N_C_M1018_g N_VPWR_c_426_n 0.0165714f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_162 N_C_M1001_g N_VPWR_c_428_n 0.00460063f $X=2.625 $Y=2.4 $X2=0 $Y2=0
cc_163 N_C_M1018_g N_VPWR_c_428_n 0.00460063f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_164 N_C_M1001_g N_VPWR_c_430_n 0.0125814f $X=2.625 $Y=2.4 $X2=0 $Y2=0
cc_165 N_C_M1018_g N_VPWR_c_430_n 0.00128042f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_166 N_C_M1001_g N_VPWR_c_423_n 0.00461676f $X=2.625 $Y=2.4 $X2=0 $Y2=0
cc_167 N_C_M1018_g N_VPWR_c_423_n 0.00463365f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_168 N_C_M1018_g N_Y_c_496_n 5.69669e-19 $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_169 N_C_M1001_g N_Y_c_500_n 0.00980014f $X=2.625 $Y=2.4 $X2=0 $Y2=0
cc_170 N_C_M1018_g N_Y_c_500_n 0.0111406f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_171 N_C_c_156_n N_Y_c_500_n 4.92363e-19 $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_172 C N_Y_c_500_n 0.0363507f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_173 N_C_c_155_n N_VGND_c_557_n 6.53784e-19 $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_174 N_C_c_156_n N_VGND_c_557_n 0.0110145f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_175 N_C_c_151_n N_VGND_c_558_n 0.00345905f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_176 N_C_c_155_n N_VGND_c_559_n 0.00419934f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_177 N_C_c_156_n N_VGND_c_559_n 0.00455951f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_178 N_C_c_151_n N_VGND_c_561_n 0.00411482f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_179 N_C_c_154_n N_VGND_c_561_n 0.00418922f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_180 N_C_c_151_n N_VGND_c_563_n 0.00533081f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_181 N_C_c_154_n N_VGND_c_563_n 0.00533081f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_182 N_C_c_155_n N_VGND_c_563_n 0.00533081f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_183 N_C_c_156_n N_VGND_c_563_n 0.00447788f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_184 N_C_c_154_n N_VGND_c_564_n 0.00458735f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_185 N_C_c_155_n N_VGND_c_564_n 0.00456635f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_186 N_C_M1001_g N_A_297_82#_c_641_n 0.0170116f $X=2.625 $Y=2.4 $X2=0 $Y2=0
cc_187 N_C_M1018_g N_A_297_82#_c_641_n 0.0138959f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_188 N_C_c_157_n N_A_297_82#_c_641_n 0.00331897f $X=1.84 $Y=1.452 $X2=0 $Y2=0
cc_189 C N_A_297_82#_c_641_n 0.030624f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_190 N_C_c_154_n N_A_297_82#_c_650_n 0.00974223f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_191 N_C_c_155_n N_A_297_82#_c_650_n 0.0102985f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_192 N_C_c_151_n N_A_297_82#_c_627_n 0.00922607f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_193 N_C_c_151_n N_A_297_82#_c_628_n 0.00749188f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_194 N_C_c_154_n N_A_297_82#_c_628_n 0.0106036f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_195 N_C_c_155_n N_A_297_82#_c_629_n 0.0108343f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_196 N_C_c_156_n N_A_297_82#_c_629_n 0.00240868f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_197 N_C_c_156_n N_A_744_74#_c_751_n 7.1746e-19 $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_198 N_A_89_172#_c_235_n N_B_c_357_n 0.00692021f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_199 N_A_89_172#_c_236_n N_B_M1003_g 0.0315164f $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_200 N_A_89_172#_c_235_n N_B_c_362_n 8.25902e-19 $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_201 N_A_89_172#_c_236_n N_B_c_363_n 7.20156e-19 $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_202 N_A_89_172#_M1008_g N_VPWR_c_426_n 0.0283726f $X=3.69 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_89_172#_M1008_g N_VPWR_c_432_n 0.00460063f $X=3.69 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_89_172#_M1009_g N_VPWR_c_432_n 0.00460063f $X=4.52 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_89_172#_M1009_g N_VPWR_c_433_n 0.0250658f $X=4.52 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_89_172#_M1008_g N_VPWR_c_423_n 0.00466128f $X=3.69 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_89_172#_M1009_g N_VPWR_c_423_n 0.00464439f $X=4.52 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_89_172#_M1009_g N_Y_c_495_n 0.0186322f $X=4.52 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_89_172#_c_233_n N_Y_c_495_n 0.00943567f $X=4.89 $Y=1.26 $X2=0 $Y2=0
cc_210 N_A_89_172#_M1008_g N_Y_c_496_n 0.0047366f $X=3.69 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A_89_172#_c_241_n N_Y_c_496_n 0.0601856f $X=4.445 $Y=1.465 $X2=0 $Y2=0
cc_212 N_A_89_172#_c_243_n N_Y_c_496_n 0.00137336f $X=3.685 $Y=1.095 $X2=0 $Y2=0
cc_213 N_A_89_172#_c_244_n N_Y_c_496_n 0.0118177f $X=4.61 $Y=1.407 $X2=0 $Y2=0
cc_214 N_A_89_172#_c_230_n N_Y_c_492_n 0.011661f $X=4.08 $Y=1.185 $X2=0 $Y2=0
cc_215 N_A_89_172#_c_232_n N_Y_c_492_n 0.0131408f $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A_89_172#_c_233_n N_Y_c_492_n 0.00420528f $X=4.89 $Y=1.26 $X2=0 $Y2=0
cc_217 N_A_89_172#_c_234_n N_Y_c_492_n 0.0069204f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_218 N_A_89_172#_c_241_n N_Y_c_492_n 0.0372722f $X=4.445 $Y=1.465 $X2=0 $Y2=0
cc_219 N_A_89_172#_c_243_n N_Y_c_492_n 0.00525886f $X=3.685 $Y=1.095 $X2=0 $Y2=0
cc_220 N_A_89_172#_c_244_n N_Y_c_492_n 0.00355854f $X=4.61 $Y=1.407 $X2=0 $Y2=0
cc_221 N_A_89_172#_c_235_n N_Y_c_497_n 0.00687428f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_222 N_A_89_172#_M1008_g N_Y_c_500_n 0.0106011f $X=3.69 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_89_172#_c_243_n N_Y_c_500_n 0.00680492f $X=3.685 $Y=1.095 $X2=0 $Y2=0
cc_224 N_A_89_172#_c_232_n Y 3.1248e-19 $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_225 N_A_89_172#_c_234_n Y 0.00164483f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_226 N_A_89_172#_c_235_n Y 0.00822151f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_227 N_A_89_172#_c_236_n Y 0.00114729f $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_228 N_A_89_172#_c_237_n Y 0.0104475f $X=4.965 $Y=1.26 $X2=0 $Y2=0
cc_229 N_A_89_172#_c_241_n Y 0.0167252f $X=4.445 $Y=1.465 $X2=0 $Y2=0
cc_230 N_A_89_172#_c_244_n Y 0.00775966f $X=4.61 $Y=1.407 $X2=0 $Y2=0
cc_231 N_A_89_172#_c_234_n N_Y_c_494_n 0.00625476f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_232 N_A_89_172#_c_235_n N_Y_c_494_n 0.00319434f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_233 N_A_89_172#_c_236_n N_Y_c_494_n 0.0088709f $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_234 N_A_89_172#_c_238_n N_VGND_M1000_d 0.00489649f $X=1.265 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_235 N_A_89_172#_c_240_n N_VGND_M1010_s 0.00702535f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_236 N_A_89_172#_c_240_n N_VGND_M1012_s 0.00259019f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_237 N_A_89_172#_c_230_n N_VGND_c_557_n 0.00715259f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_238 N_A_89_172#_c_240_n N_VGND_c_557_n 0.0220913f $X=3.6 $Y=1.095 $X2=0 $Y2=0
cc_239 N_A_89_172#_c_230_n N_VGND_c_562_n 0.00291649f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_240 N_A_89_172#_c_232_n N_VGND_c_562_n 0.00291649f $X=4.535 $Y=1.185 $X2=0
+ $Y2=0
cc_241 N_A_89_172#_c_234_n N_VGND_c_562_n 0.00291649f $X=4.965 $Y=1.185 $X2=0
+ $Y2=0
cc_242 N_A_89_172#_c_236_n N_VGND_c_562_n 0.00291649f $X=5.395 $Y=1.185 $X2=0
+ $Y2=0
cc_243 N_A_89_172#_c_230_n N_VGND_c_563_n 0.00364365f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_244 N_A_89_172#_c_232_n N_VGND_c_563_n 0.00359366f $X=4.535 $Y=1.185 $X2=0
+ $Y2=0
cc_245 N_A_89_172#_c_234_n N_VGND_c_563_n 0.00359121f $X=4.965 $Y=1.185 $X2=0
+ $Y2=0
cc_246 N_A_89_172#_c_236_n N_VGND_c_563_n 0.00359833f $X=5.395 $Y=1.185 $X2=0
+ $Y2=0
cc_247 N_A_89_172#_c_240_n N_A_297_82#_M1006_d 0.00176891f $X=3.6 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_248 N_A_89_172#_c_240_n N_A_297_82#_M1011_d 0.00250873f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_249 N_A_89_172#_c_242_n N_A_297_82#_c_624_n 0.020614f $X=0.59 $Y=1.005 $X2=0
+ $Y2=0
cc_250 N_A_89_172#_M1017_d N_A_297_82#_c_641_n 0.00473027f $X=0.985 $Y=1.84
+ $X2=0 $Y2=0
cc_251 N_A_89_172#_M1008_g N_A_297_82#_c_641_n 0.0154035f $X=3.69 $Y=2.4 $X2=0
+ $Y2=0
cc_252 N_A_89_172#_M1009_g N_A_297_82#_c_641_n 0.0167389f $X=4.52 $Y=2.4 $X2=0
+ $Y2=0
cc_253 N_A_89_172#_c_251_n N_A_297_82#_c_641_n 0.0268888f $X=1.265 $Y=2.045
+ $X2=0 $Y2=0
cc_254 N_A_89_172#_c_236_n N_A_297_82#_c_664_n 5.14228e-19 $X=5.395 $Y=1.185
+ $X2=0 $Y2=0
cc_255 N_A_89_172#_M1000_s N_A_297_82#_c_627_n 0.00566964f $X=0.445 $Y=0.86
+ $X2=0 $Y2=0
cc_256 N_A_89_172#_c_238_n N_A_297_82#_c_627_n 0.0234296f $X=1.265 $Y=1.095
+ $X2=0 $Y2=0
cc_257 N_A_89_172#_c_240_n N_A_297_82#_c_627_n 0.0011585f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_258 N_A_89_172#_c_242_n N_A_297_82#_c_627_n 0.0203761f $X=0.59 $Y=1.005 $X2=0
+ $Y2=0
cc_259 N_A_89_172#_c_278_n N_A_297_82#_c_627_n 0.00618821f $X=1.35 $Y=1.095
+ $X2=0 $Y2=0
cc_260 N_A_89_172#_c_240_n N_A_297_82#_c_628_n 0.0688738f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_261 N_A_89_172#_c_240_n N_A_297_82#_c_629_n 0.0203381f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_262 N_A_89_172#_c_243_n N_A_744_74#_M1005_d 0.00139751f $X=3.685 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_263 N_A_89_172#_c_230_n N_A_744_74#_c_751_n 0.0024281f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_264 N_A_89_172#_c_241_n N_A_744_74#_c_751_n 0.00585628f $X=4.445 $Y=1.465
+ $X2=0 $Y2=0
cc_265 N_A_89_172#_c_243_n N_A_744_74#_c_751_n 0.00332029f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_266 N_A_89_172#_c_244_n N_A_744_74#_c_751_n 0.00465854f $X=4.61 $Y=1.407
+ $X2=0 $Y2=0
cc_267 N_A_89_172#_c_230_n N_A_744_74#_c_752_n 0.0122631f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_268 N_A_89_172#_c_232_n N_A_744_74#_c_752_n 0.0106216f $X=4.535 $Y=1.185
+ $X2=0 $Y2=0
cc_269 N_A_89_172#_c_234_n N_A_744_74#_c_752_n 0.0102551f $X=4.965 $Y=1.185
+ $X2=0 $Y2=0
cc_270 N_A_89_172#_c_236_n N_A_744_74#_c_752_n 0.0175315f $X=5.395 $Y=1.185
+ $X2=0 $Y2=0
cc_271 N_B_c_364_n N_VPWR_c_427_n 0.00307643f $X=5.46 $Y=1.725 $X2=0 $Y2=0
cc_272 N_B_c_367_n N_VPWR_c_427_n 0.00307643f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_273 N_B_c_364_n N_VPWR_c_433_n 0.0125746f $X=5.46 $Y=1.725 $X2=0 $Y2=0
cc_274 N_B_c_367_n N_VPWR_c_433_n 0.00127991f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_275 N_B_c_364_n N_VPWR_c_434_n 0.00128463f $X=5.46 $Y=1.725 $X2=0 $Y2=0
cc_276 N_B_c_367_n N_VPWR_c_434_n 0.0188613f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_277 N_B_c_364_n N_VPWR_c_423_n 0.00461676f $X=5.46 $Y=1.725 $X2=0 $Y2=0
cc_278 N_B_c_367_n N_VPWR_c_423_n 0.00461676f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_279 N_B_c_364_n N_Y_c_497_n 0.0209674f $X=5.46 $Y=1.725 $X2=0 $Y2=0
cc_280 N_B_c_356_n N_Y_c_497_n 0.00360837f $X=5.74 $Y=1.65 $X2=0 $Y2=0
cc_281 N_B_c_367_n N_Y_c_497_n 0.00511506f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_282 N_B_c_363_n N_Y_c_497_n 0.00230862f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_283 N_B_c_357_n Y 0.00855912f $X=5.55 $Y=1.65 $X2=0 $Y2=0
cc_284 N_B_c_362_n Y 0.00471144f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_285 N_B_c_363_n Y 0.0127966f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_286 N_B_M1003_g N_Y_c_494_n 0.00141517f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_287 N_B_M1003_g N_VGND_c_562_n 0.00291649f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_288 N_B_M1007_g N_VGND_c_562_n 0.00291649f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_289 N_B_M1015_g N_VGND_c_562_n 0.00291649f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_290 N_B_M1016_g N_VGND_c_562_n 0.00291649f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_291 N_B_M1003_g N_VGND_c_563_n 0.00359833f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_292 N_B_M1007_g N_VGND_c_563_n 0.00359121f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_293 N_B_M1015_g N_VGND_c_563_n 0.00359121f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_294 N_B_M1016_g N_VGND_c_563_n 0.00362779f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_295 N_B_c_364_n N_A_297_82#_c_641_n 0.0151925f $X=5.46 $Y=1.725 $X2=0 $Y2=0
cc_296 N_B_c_367_n N_A_297_82#_c_641_n 0.0165919f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_297 N_B_c_363_n N_A_297_82#_c_641_n 0.00431983f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_298 N_B_M1003_g N_A_297_82#_c_664_n 0.00384298f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_299 N_B_M1007_g N_A_297_82#_c_664_n 0.00843705f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B_M1015_g N_A_297_82#_c_664_n 0.00843705f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_301 N_B_M1016_g N_A_297_82#_c_664_n 0.0129826f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B_c_362_n N_A_297_82#_c_664_n 0.00149218f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_303 N_B_c_363_n N_A_297_82#_c_664_n 0.0772269f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_304 N_B_c_367_n N_A_297_82#_c_681_n 0.0101691f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_305 N_B_c_362_n N_A_297_82#_c_632_n 0.0303401f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_306 N_B_c_363_n N_A_297_82#_c_632_n 0.0652259f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_307 N_B_c_367_n N_A_297_82#_c_633_n 0.00418654f $X=5.91 $Y=1.725 $X2=0 $Y2=0
cc_308 N_B_c_362_n N_A_297_82#_c_633_n 0.00473088f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_309 N_B_c_363_n N_A_297_82#_c_633_n 0.0146559f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_310 N_B_M1015_g N_A_297_82#_c_626_n 7.10626e-19 $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_311 N_B_M1016_g N_A_297_82#_c_626_n 0.00947193f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_312 N_B_c_362_n N_A_297_82#_c_626_n 0.0137996f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_313 N_B_c_363_n N_A_297_82#_c_626_n 0.036909f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_314 N_B_M1003_g N_A_744_74#_c_749_n 0.00118092f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_315 N_B_c_362_n N_A_744_74#_c_749_n 0.00145872f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_316 N_B_c_363_n N_A_744_74#_c_749_n 0.00389228f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_317 N_B_M1003_g N_A_744_74#_c_750_n 0.0122981f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_318 N_B_M1007_g N_A_744_74#_c_750_n 0.0120586f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_319 N_B_M1015_g N_A_744_74#_c_750_n 0.0120586f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_320 N_B_M1016_g N_A_744_74#_c_750_n 0.0122066f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_321 N_VPWR_M1009_d N_Y_c_495_n 0.00501014f $X=4.61 $Y=1.84 $X2=0 $Y2=0
cc_322 N_VPWR_M1009_d N_Y_c_497_n 0.0022686f $X=4.61 $Y=1.84 $X2=0 $Y2=0
cc_323 N_VPWR_M1018_d N_Y_c_500_n 0.0162631f $X=3.165 $Y=1.84 $X2=0 $Y2=0
cc_324 N_VPWR_M1009_d N_Y_c_541_n 0.00637067f $X=4.61 $Y=1.84 $X2=0 $Y2=0
cc_325 N_VPWR_M1017_s N_A_297_82#_c_624_n 0.00242459f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_326 N_VPWR_M1017_s N_A_297_82#_c_639_n 0.0222151f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_425_n N_A_297_82#_c_639_n 0.0153403f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_328 N_VPWR_M1017_s N_A_297_82#_c_631_n 0.00244603f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_425_n N_A_297_82#_c_631_n 0.0125546f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_330 N_VPWR_M1017_s N_A_297_82#_c_696_n 0.00681249f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_425_n N_A_297_82#_c_696_n 0.00149212f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_332 N_VPWR_M1020_s N_A_297_82#_c_641_n 0.0393528f $X=1.435 $Y=1.84 $X2=0
+ $Y2=0
cc_333 N_VPWR_M1018_d N_A_297_82#_c_641_n 0.00748652f $X=3.165 $Y=1.84 $X2=0
+ $Y2=0
cc_334 N_VPWR_M1009_d N_A_297_82#_c_641_n 0.0173926f $X=4.61 $Y=1.84 $X2=0 $Y2=0
cc_335 N_VPWR_M1004_s N_A_297_82#_c_641_n 0.00420712f $X=6 $Y=1.84 $X2=0 $Y2=0
cc_336 N_VPWR_c_426_n N_A_297_82#_c_641_n 0.0298907f $X=3.38 $Y=2.815 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_430_n N_A_297_82#_c_641_n 0.0803372f $X=2.565 $Y=3.032 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_433_n N_A_297_82#_c_641_n 0.0555716f $X=5.4 $Y=3.032 $X2=0 $Y2=0
cc_339 N_VPWR_c_434_n N_A_297_82#_c_641_n 0.032597f $X=7.4 $Y=2.325 $X2=0 $Y2=0
cc_340 N_VPWR_c_423_n N_A_297_82#_c_641_n 0.0965196f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_341 N_VPWR_M1017_s N_A_297_82#_c_707_n 0.00507182f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_425_n N_A_297_82#_c_707_n 0.0144778f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_423_n N_A_297_82#_c_707_n 0.00648262f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_344 N_VPWR_M1004_s N_A_297_82#_c_681_n 0.0129914f $X=6 $Y=1.84 $X2=0 $Y2=0
cc_345 N_VPWR_c_434_n N_A_297_82#_c_681_n 0.0121673f $X=7.4 $Y=2.325 $X2=0 $Y2=0
cc_346 N_VPWR_M1004_s N_A_297_82#_c_632_n 0.0309213f $X=6 $Y=1.84 $X2=0 $Y2=0
cc_347 N_VPWR_c_434_n N_A_297_82#_c_632_n 0.0889948f $X=7.4 $Y=2.325 $X2=0 $Y2=0
cc_348 N_VPWR_M1004_s N_A_297_82#_c_633_n 0.00278928f $X=6 $Y=1.84 $X2=0 $Y2=0
cc_349 N_Y_c_492_n N_VGND_c_557_n 0.00115716f $X=4.925 $Y=0.965 $X2=0 $Y2=0
cc_350 N_Y_M1001_s N_A_297_82#_c_641_n 0.00474966f $X=2.715 $Y=1.84 $X2=0 $Y2=0
cc_351 N_Y_M1008_s N_A_297_82#_c_641_n 0.0189322f $X=3.78 $Y=1.84 $X2=0 $Y2=0
cc_352 N_Y_M1002_d N_A_297_82#_c_641_n 0.00473982f $X=5.55 $Y=1.84 $X2=0 $Y2=0
cc_353 N_Y_c_497_n N_A_297_82#_c_641_n 0.0387838f $X=5.685 $Y=2.02 $X2=0 $Y2=0
cc_354 N_Y_c_500_n N_A_297_82#_c_641_n 0.134784f $X=3.75 $Y=1.98 $X2=0 $Y2=0
cc_355 N_Y_c_541_n N_A_297_82#_c_641_n 0.0187125f $X=5.04 $Y=1.98 $X2=0 $Y2=0
cc_356 N_Y_c_494_n N_A_297_82#_c_664_n 0.00497712f $X=5.04 $Y=1.13 $X2=0 $Y2=0
cc_357 N_Y_c_497_n N_A_297_82#_c_681_n 0.00990768f $X=5.685 $Y=2.02 $X2=0 $Y2=0
cc_358 N_Y_c_497_n N_A_297_82#_c_633_n 0.0125668f $X=5.685 $Y=2.02 $X2=0 $Y2=0
cc_359 N_Y_c_492_n N_A_744_74#_M1013_d 0.00189973f $X=4.925 $Y=0.965 $X2=0 $Y2=0
cc_360 N_Y_M1005_s N_A_744_74#_c_752_n 0.00207408f $X=4.155 $Y=0.37 $X2=0 $Y2=0
cc_361 N_Y_M1014_s N_A_744_74#_c_752_n 0.00168993f $X=5.04 $Y=0.37 $X2=0 $Y2=0
cc_362 N_Y_c_492_n N_A_744_74#_c_752_n 0.0365346f $X=4.925 $Y=0.965 $X2=0 $Y2=0
cc_363 N_Y_c_494_n N_A_744_74#_c_752_n 0.0233947f $X=5.04 $Y=1.13 $X2=0 $Y2=0
cc_364 N_VGND_c_558_n N_A_297_82#_c_625_n 0.00387622f $X=0.935 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_563_n N_A_297_82#_c_625_n 0.00537088f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_M1010_s N_A_297_82#_c_650_n 0.0117523f $X=1.915 $Y=0.41 $X2=0
+ $Y2=0
cc_367 N_VGND_c_559_n N_A_297_82#_c_650_n 0.00237563f $X=3.14 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_561_n N_A_297_82#_c_650_n 0.00236949f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_563_n N_A_297_82#_c_650_n 0.011866f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_564_n N_A_297_82#_c_650_n 0.0374471f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_M1000_d N_A_297_82#_c_627_n 0.00852962f $X=0.88 $Y=0.41 $X2=0
+ $Y2=0
cc_372 N_VGND_c_558_n N_A_297_82#_c_627_n 0.0381142f $X=0.935 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_c_561_n N_A_297_82#_c_627_n 0.00294479f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_374 N_VGND_c_563_n N_A_297_82#_c_627_n 0.0271405f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_558_n N_A_297_82#_c_628_n 0.00145202f $X=0.935 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_c_561_n N_A_297_82#_c_628_n 0.0121348f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_377 N_VGND_c_563_n N_A_297_82#_c_628_n 0.0116628f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_564_n N_A_297_82#_c_628_n 0.00469436f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_557_n N_A_297_82#_c_629_n 0.0176756f $X=3.305 $Y=0.615 $X2=0
+ $Y2=0
cc_380 N_VGND_c_559_n N_A_297_82#_c_629_n 0.0121755f $X=3.14 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_563_n N_A_297_82#_c_629_n 0.0116241f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_564_n N_A_297_82#_c_629_n 0.00474851f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_557_n N_A_744_74#_c_751_n 0.0197752f $X=3.305 $Y=0.615 $X2=0
+ $Y2=0
cc_384 N_VGND_c_562_n N_A_744_74#_c_751_n 0.158354f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_563_n N_A_744_74#_c_751_n 0.132997f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_386 N_A_297_82#_c_664_n N_A_744_74#_M1007_d 0.00333133f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0
cc_387 N_A_297_82#_c_664_n N_A_744_74#_M1016_d 0.00874113f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0
cc_388 N_A_297_82#_c_626_n N_A_744_74#_M1016_d 0.0037774f $X=7.33 $Y=1.82 $X2=0
+ $Y2=0
cc_389 N_A_297_82#_M1003_s N_A_744_74#_c_750_n 0.00172259f $X=5.97 $Y=0.37 $X2=0
+ $Y2=0
cc_390 N_A_297_82#_M1015_s N_A_744_74#_c_750_n 0.00172259f $X=6.83 $Y=0.37 $X2=0
+ $Y2=0
cc_391 N_A_297_82#_c_664_n N_A_744_74#_c_750_n 0.0780631f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0

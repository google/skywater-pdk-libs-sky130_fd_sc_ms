# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__xnor3_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__xnor3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.915000 1.375000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.771000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.940000 1.350000 4.270000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.780000 1.350000 7.110000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.280000 1.840000 8.640000 2.980000 ;
        RECT 8.345000 0.470000 8.675000 1.170000 ;
        RECT 8.470000 1.170000 8.675000 1.420000 ;
        RECT 8.470000 1.420000 9.535000 1.625000 ;
        RECT 8.470000 1.625000 8.640000 1.840000 ;
        RECT 9.180000 1.625000 9.535000 2.980000 ;
        RECT 9.205000 0.440000 9.535000 1.420000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.665000  0.085000  0.995000 0.865000 ;
        RECT 4.270000  0.085000  4.600000 0.445000 ;
        RECT 6.900000  0.085000  8.165000 0.490000 ;
        RECT 7.230000  0.490000  8.165000 0.840000 ;
        RECT 7.915000  0.840000  8.165000 1.170000 ;
        RECT 8.855000  0.085000  9.025000 1.250000 ;
        RECT 9.715000  0.085000  9.965000 1.250000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.565000 2.290000  0.895000 3.245000 ;
        RECT 4.390000 2.730000  4.720000 3.245000 ;
        RECT 7.485000 2.290000  8.110000 3.245000 ;
        RECT 7.685000 1.840000  8.110000 2.290000 ;
        RECT 8.810000 1.820000  8.980000 3.245000 ;
        RECT 9.710000 1.820000  9.960000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.365000 0.495000 0.865000 ;
      RECT 0.085000 0.865000 0.285000 1.845000 ;
      RECT 0.085000 1.845000 0.365000 2.885000 ;
      RECT 0.455000 1.035000 1.425000 1.205000 ;
      RECT 0.455000 1.205000 0.705000 1.465000 ;
      RECT 0.535000 1.465000 0.705000 1.950000 ;
      RECT 0.535000 1.950000 1.395000 2.120000 ;
      RECT 1.065000 2.120000 1.395000 2.905000 ;
      RECT 1.065000 2.905000 3.680000 3.075000 ;
      RECT 1.175000 0.255000 3.530000 0.425000 ;
      RECT 1.175000 0.425000 1.425000 1.035000 ;
      RECT 1.565000 1.375000 1.765000 2.565000 ;
      RECT 1.565000 2.565000 2.725000 2.735000 ;
      RECT 1.595000 1.165000 2.385000 1.335000 ;
      RECT 1.595000 1.335000 1.765000 1.375000 ;
      RECT 1.625000 0.595000 2.725000 0.615000 ;
      RECT 1.625000 0.615000 5.160000 0.765000 ;
      RECT 1.625000 0.765000 1.955000 0.995000 ;
      RECT 1.935000 1.505000 2.755000 1.675000 ;
      RECT 1.935000 1.675000 2.245000 2.120000 ;
      RECT 1.935000 2.120000 2.135000 2.155000 ;
      RECT 2.135000 0.935000 2.385000 1.165000 ;
      RECT 2.305000 2.290000 2.725000 2.565000 ;
      RECT 2.555000 0.765000 5.160000 0.785000 ;
      RECT 2.555000 0.955000 3.020000 1.205000 ;
      RECT 2.555000 1.205000 2.755000 1.505000 ;
      RECT 2.895000 1.875000 3.145000 2.370000 ;
      RECT 2.895000 2.370000 4.610000 2.390000 ;
      RECT 2.895000 2.390000 6.270000 2.540000 ;
      RECT 2.895000 2.540000 3.145000 2.545000 ;
      RECT 2.995000 1.375000 3.770000 1.705000 ;
      RECT 3.200000 0.425000 3.530000 0.445000 ;
      RECT 3.350000 2.710000 3.680000 2.905000 ;
      RECT 3.600000 0.955000 4.090000 1.125000 ;
      RECT 3.600000 1.125000 3.770000 1.375000 ;
      RECT 3.600000 1.705000 3.770000 1.950000 ;
      RECT 3.600000 1.950000 4.270000 2.200000 ;
      RECT 4.440000 0.785000 5.160000 1.030000 ;
      RECT 4.440000 1.030000 4.610000 2.370000 ;
      RECT 4.440000 2.540000 6.270000 2.560000 ;
      RECT 4.780000 1.210000 6.160000 1.380000 ;
      RECT 4.780000 1.380000 4.950000 1.950000 ;
      RECT 4.780000 1.950000 5.280000 2.220000 ;
      RECT 4.830000 0.350000 5.160000 0.615000 ;
      RECT 5.120000 1.550000 6.610000 1.720000 ;
      RECT 5.120000 1.720000 5.450000 1.780000 ;
      RECT 5.330000 0.255000 6.500000 0.425000 ;
      RECT 5.330000 0.425000 5.660000 1.010000 ;
      RECT 5.405000 1.180000 6.160000 1.210000 ;
      RECT 5.485000 2.730000 5.815000 2.905000 ;
      RECT 5.485000 2.905000 7.315000 3.075000 ;
      RECT 5.830000 0.595000 6.160000 1.180000 ;
      RECT 6.020000 1.970000 6.270000 2.390000 ;
      RECT 6.020000 2.560000 6.270000 2.735000 ;
      RECT 6.330000 0.425000 6.500000 0.660000 ;
      RECT 6.330000 0.660000 7.060000 0.830000 ;
      RECT 6.390000 1.000000 6.720000 1.170000 ;
      RECT 6.390000 1.170000 6.610000 1.550000 ;
      RECT 6.440000 1.720000 6.610000 1.990000 ;
      RECT 6.440000 1.990000 6.960000 2.500000 ;
      RECT 6.890000 0.830000 7.060000 1.010000 ;
      RECT 6.890000 1.010000 7.490000 1.180000 ;
      RECT 7.130000 1.950000 7.490000 2.120000 ;
      RECT 7.130000 2.120000 7.315000 2.905000 ;
      RECT 7.320000 1.180000 7.490000 1.340000 ;
      RECT 7.320000 1.340000 8.300000 1.670000 ;
      RECT 7.320000 1.670000 7.490000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 1.950000 0.325000 2.120000 ;
      RECT 1.595000 1.950000 1.765000 2.120000 ;
      RECT 2.075000 1.950000 2.245000 2.120000 ;
      RECT 4.955000 1.950000 5.125000 2.120000 ;
    LAYER met1 ;
      RECT 0.095000 1.920000 0.385000 1.965000 ;
      RECT 0.095000 1.965000 1.825000 2.105000 ;
      RECT 0.095000 2.105000 0.385000 2.150000 ;
      RECT 1.535000 1.920000 1.825000 1.965000 ;
      RECT 1.535000 2.105000 1.825000 2.150000 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 1.965000 5.185000 2.105000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 4.895000 1.920000 5.185000 1.965000 ;
      RECT 4.895000 2.105000 5.185000 2.150000 ;
  END
END sky130_fd_sc_ms__xnor3_4

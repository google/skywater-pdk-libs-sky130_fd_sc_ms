* File: sky130_fd_sc_ms__dlxtn_4.pex.spice
* Created: Fri Aug 28 17:29:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLXTN_4%D 3 7 9 13 16
c28 3 0 1.04866e-19 $X=0.495 $Y=0.85
r29 15 16 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.525 $Y2=1.465
r30 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.495 $Y2=1.465
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r32 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r33 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.63
+ $X2=0.525 $Y2=1.465
r34 5 7 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.525 $Y=1.63
+ $X2=0.525 $Y2=2.54
r35 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r36 1 3 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%GATE_N 3 7 9 12
c40 3 0 1.68883e-19 $X=1.075 $Y=2.54
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.83
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.5
r43 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.665 $X2=1.15 $Y2=1.665
r44 7 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.085 $Y=0.94
+ $X2=1.085 $Y2=1.5
r45 3 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.075 $Y=2.54
+ $X2=1.075 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%A_232_114# 1 2 9 11 13 14 16 18 21 25 27 31
+ 32 35 39 40 42 44 45 50 52 56 57 64
c145 38 0 5.47968e-20 $X=3.075 $Y=2.905
c146 27 0 1.04866e-19 $X=1.485 $Y=1.165
c147 25 0 6.91456e-20 $X=3.855 $Y=1.185
r148 66 68 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.855 $Y=1.57
+ $X2=3.87 $Y2=1.57
r149 57 68 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=4.215 $Y=1.57
+ $X2=3.87 $Y2=1.57
r150 56 59 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=1.57
+ $X2=4.215 $Y2=1.735
r151 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.215
+ $Y=1.57 $X2=4.215 $Y2=1.57
r152 53 64 45.7069 $w=5.22e-07 $l=4.95e-07 $layer=POLY_cond $X=1.72 $Y=1.477
+ $X2=2.215 $Y2=1.477
r153 53 60 13.513 $w=3.3e-07 $l=2.92e-07 $layer=POLY_cond $X=1.72 $Y=1.477
+ $X2=1.72 $Y2=1.185
r154 52 54 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.605
+ $X2=1.685 $Y2=1.77
r155 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.605 $X2=1.72 $Y2=1.605
r156 50 60 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.72 $Y=0.925
+ $X2=1.72 $Y2=1.185
r157 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=0.925 $X2=1.72 $Y2=0.925
r158 45 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.57 $Y=2.1
+ $X2=1.57 $Y2=1.77
r159 44 46 4.83032 $w=5.18e-07 $l=2.1e-07 $layer=LI1_cond $X=1.395 $Y=2.265
+ $X2=1.395 $Y2=2.475
r160 44 45 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.265
+ $X2=1.395 $Y2=2.1
r161 42 59 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.135 $Y=2.905
+ $X2=4.135 $Y2=1.735
r162 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.05 $Y=2.99
+ $X2=4.135 $Y2=2.905
r163 39 40 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.05 $Y=2.99
+ $X2=3.16 $Y2=2.99
r164 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.905
+ $X2=3.16 $Y2=2.99
r165 37 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.075 $Y=2.56
+ $X2=3.075 $Y2=2.905
r166 36 46 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.655 $Y=2.475
+ $X2=1.395 $Y2=2.475
r167 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=3.075 $Y2=2.56
r168 35 36 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=1.655 $Y2=2.475
r169 32 52 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.685 $Y=1.57
+ $X2=1.685 $Y2=1.605
r170 31 49 3.24963 $w=4e-07 $l=2.85e-07 $layer=LI1_cond $X=1.685 $Y=1.33
+ $X2=1.685 $Y2=1.045
r171 31 32 6.91466 $w=3.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.685 $Y=1.33
+ $X2=1.685 $Y2=1.57
r172 27 49 3.6487 $w=3.3e-07 $l=2.52982e-07 $layer=LI1_cond $X=1.485 $Y=1.165
+ $X2=1.685 $Y2=1.045
r173 27 29 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.485 $Y=1.165
+ $X2=1.3 $Y2=1.165
r174 23 25 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.605 $Y=1.185
+ $X2=3.855 $Y2=1.185
r175 19 68 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.87 $Y=1.735
+ $X2=3.87 $Y2=1.57
r176 19 21 394.54 $w=1.8e-07 $l=1.015e-06 $layer=POLY_cond $X=3.87 $Y=1.735
+ $X2=3.87 $Y2=2.75
r177 18 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.405
+ $X2=3.855 $Y2=1.57
r178 17 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.855 $Y=1.26
+ $X2=3.855 $Y2=1.185
r179 17 18 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.855 $Y=1.26
+ $X2=3.855 $Y2=1.405
r180 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.605 $Y=1.11
+ $X2=3.605 $Y2=1.185
r181 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=1.11
+ $X2=3.605 $Y2=0.715
r182 11 64 12.9272 $w=5.22e-07 $l=3.55168e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.215 $Y2=1.477
r183 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.74
r184 7 64 27.9254 $w=1.8e-07 $l=2.93e-07 $layer=POLY_cond $X=2.215 $Y=1.77
+ $X2=2.215 $Y2=1.477
r185 7 9 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=2.215 $Y=1.77
+ $X2=2.215 $Y2=2.38
r186 2 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.165
+ $Y=2.12 $X2=1.3 $Y2=2.265
r187 1 29 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.57 $X2=1.3 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%A_27_115# 1 2 9 11 13 16 19 20 21 23 24 25
+ 27 33 38 42
r110 39 42 7.97426 $w=2.72e-07 $l=4.5e-08 $layer=POLY_cond $X=2.835 $Y=1.33
+ $X2=2.88 $Y2=1.33
r111 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.835
+ $Y=1.385 $X2=2.835 $Y2=1.385
r112 35 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.56 $Y=1.385
+ $X2=2.835 $Y2=1.385
r113 29 30 10.0885 $w=5.2e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.842
+ $X2=0.71 $Y2=0.842
r114 27 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=1.22
+ $X2=2.56 $Y2=1.385
r115 26 27 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=1.22
r116 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=2.56 $Y2=0.425
r117 24 25 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=1.315 $Y2=0.34
r118 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.315 $Y2=0.34
r119 22 23 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.66
r120 21 30 7.9572 $w=5.2e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.795 $Y=0.745
+ $X2=0.71 $Y2=0.842
r121 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=0.745
+ $X2=1.23 $Y2=0.66
r122 20 21 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.145 $Y=0.745
+ $X2=0.795 $Y2=0.745
r123 19 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.71 $Y2=2.035
r124 18 30 7.40362 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=0.842
r125 18 19 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r126 14 33 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.3 $Y=2.035
+ $X2=0.71 $Y2=2.035
r127 14 16 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.3 $Y=2.12
+ $X2=0.3 $Y2=2.265
r128 11 42 59.364 $w=2.72e-07 $l=4.3119e-07 $layer=POLY_cond $X=3.215 $Y=1.11
+ $X2=2.88 $Y2=1.33
r129 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.215 $Y=1.11
+ $X2=3.215 $Y2=0.715
r130 7 42 12.4592 $w=1.8e-07 $l=2.2e-07 $layer=POLY_cond $X=2.88 $Y=1.55
+ $X2=2.88 $Y2=1.33
r131 7 9 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=2.88 $Y=1.55 $X2=2.88
+ $Y2=2.46
r132 2 16 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.12 $X2=0.3 $Y2=2.265
r133 1 29 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.575 $X2=0.28 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%A_369_392# 1 2 9 11 13 16 18 22 24 27 31 32
+ 33 41
c94 31 0 6.91456e-20 $X=3.375 $Y=1.635
c95 27 0 1.68883e-19 $X=2.065 $Y=1.805
c96 24 0 6.33553e-20 $X=4.28 $Y=0.34
c97 22 0 1.82656e-20 $X=3.485 $Y=0.38
r98 32 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.635
+ $X2=3.375 $Y2=1.8
r99 31 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.375 $Y=1.635
+ $X2=3.375 $Y2=1.805
r100 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=1.635
+ $X2=3.375 $Y2=1.47
r101 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.375
+ $Y=1.635 $X2=3.375 $Y2=1.635
r102 27 29 11.7883 $w=3.26e-07 $l=3.15e-07 $layer=LI1_cond $X=2.065 $Y=1.805
+ $X2=2.065 $Y2=2.12
r103 25 41 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.28 $Y=0.34
+ $X2=4.4 $Y2=0.34
r104 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=0.34 $X2=4.28 $Y2=0.34
r105 22 24 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=3.485 $Y=0.38
+ $X2=4.28 $Y2=0.38
r106 20 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.4 $Y=0.505
+ $X2=3.485 $Y2=0.38
r107 20 33 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.4 $Y=0.505
+ $X2=3.4 $Y2=1.47
r108 19 27 4.55145 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=2.305 $Y=1.805
+ $X2=2.065 $Y2=1.805
r109 18 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=1.805
+ $X2=3.375 $Y2=1.805
r110 18 19 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=3.21 $Y=1.805
+ $X2=2.305 $Y2=1.805
r111 14 27 3.87481 $w=3.26e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.18 $Y=1.72
+ $X2=2.065 $Y2=1.805
r112 14 16 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=2.18 $Y=1.72
+ $X2=2.18 $Y2=0.86
r113 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=0.505
+ $X2=4.4 $Y2=0.34
r114 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.4 $Y=0.505
+ $X2=4.4 $Y2=0.825
r115 9 38 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.3 $Y=2.46 $X2=3.3
+ $Y2=1.8
r116 2 29 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.12
r117 1 16 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.37 $X2=2.14 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%A_840_395# 1 2 9 13 17 21 23 27 31 35 39 43
+ 47 49 52 58 61 63 67 69 73 77 79 89
c154 67 0 1.4938e-19 $X=6.305 $Y=1.485
c155 63 0 9.68457e-20 $X=5.745 $Y=1.82
c156 58 0 1.44963e-19 $X=5.485 $Y=0.54
c157 13 0 6.33553e-20 $X=4.76 $Y=0.825
r158 89 90 2.22462 $w=3.25e-07 $l=1.5e-08 $layer=POLY_cond $X=7.64 $Y=1.485
+ $X2=7.655 $Y2=1.485
r159 86 87 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=7.165 $Y=1.485
+ $X2=7.205 $Y2=1.485
r160 85 86 60.8062 $w=3.25e-07 $l=4.1e-07 $layer=POLY_cond $X=6.755 $Y=1.485
+ $X2=7.165 $Y2=1.485
r161 84 85 2.96615 $w=3.25e-07 $l=2e-08 $layer=POLY_cond $X=6.735 $Y=1.485
+ $X2=6.755 $Y2=1.485
r162 70 89 46.7169 $w=3.25e-07 $l=3.15e-07 $layer=POLY_cond $X=7.325 $Y=1.485
+ $X2=7.64 $Y2=1.485
r163 70 87 17.7969 $w=3.25e-07 $l=1.2e-07 $layer=POLY_cond $X=7.325 $Y=1.485
+ $X2=7.205 $Y2=1.485
r164 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.325
+ $Y=1.485 $X2=7.325 $Y2=1.485
r165 66 69 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.305 $Y=1.485
+ $X2=7.325 $Y2=1.485
r166 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.305
+ $Y=1.485 $X2=6.305 $Y2=1.485
r167 64 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=1.485
+ $X2=5.745 $Y2=1.485
r168 64 66 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.83 $Y=1.485
+ $X2=6.305 $Y2=1.485
r169 63 73 8.71429 $w=3.71e-07 $l=3.66545e-07 $layer=LI1_cond $X=5.745 $Y=1.82
+ $X2=5.48 $Y2=2.062
r170 62 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=1.65
+ $X2=5.745 $Y2=1.485
r171 62 63 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.745 $Y=1.65
+ $X2=5.745 $Y2=1.82
r172 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=1.32
+ $X2=5.745 $Y2=1.485
r173 60 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=1.15
+ $X2=5.745 $Y2=1.065
r174 60 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.745 $Y=1.15
+ $X2=5.745 $Y2=1.32
r175 56 77 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.445 $Y=1.065
+ $X2=5.745 $Y2=1.065
r176 56 58 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=5.445 $Y=0.98
+ $X2=5.445 $Y2=0.54
r177 52 82 27.2956 $w=3.62e-07 $l=2.05e-07 $layer=POLY_cond $X=4.555 $Y=2.032
+ $X2=4.76 $Y2=2.032
r178 52 80 35.2845 $w=3.62e-07 $l=2.65e-07 $layer=POLY_cond $X=4.555 $Y=2.032
+ $X2=4.29 $Y2=2.032
r179 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.555
+ $Y=2.14 $X2=4.555 $Y2=2.14
r180 49 73 5.60386 $w=3.71e-07 $l=2.00237e-07 $layer=LI1_cond $X=5.315 $Y=2.14
+ $X2=5.48 $Y2=2.062
r181 49 51 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.315 $Y=2.14
+ $X2=4.555 $Y2=2.14
r182 45 90 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.65
+ $X2=7.655 $Y2=1.485
r183 45 47 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.655 $Y=1.65
+ $X2=7.655 $Y2=2.4
r184 41 89 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.64 $Y=1.32
+ $X2=7.64 $Y2=1.485
r185 41 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.64 $Y=1.32
+ $X2=7.64 $Y2=0.74
r186 37 87 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=1.65
+ $X2=7.205 $Y2=1.485
r187 37 39 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.205 $Y=1.65
+ $X2=7.205 $Y2=2.4
r188 33 86 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.32
+ $X2=7.165 $Y2=1.485
r189 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.165 $Y=1.32
+ $X2=7.165 $Y2=0.74
r190 29 85 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.755 $Y=1.65
+ $X2=6.755 $Y2=1.485
r191 29 31 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.755 $Y=1.65
+ $X2=6.755 $Y2=2.4
r192 25 84 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.32
+ $X2=6.735 $Y2=1.485
r193 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.735 $Y=1.32
+ $X2=6.735 $Y2=0.74
r194 24 67 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.32 $Y=1.485
+ $X2=6.23 $Y2=1.485
r195 23 84 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=1.485
+ $X2=6.735 $Y2=1.485
r196 23 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.66 $Y=1.485
+ $X2=6.32 $Y2=1.485
r197 19 67 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.65
+ $X2=6.23 $Y2=1.485
r198 19 21 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.23 $Y=1.65
+ $X2=6.23 $Y2=2.4
r199 15 67 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=6.215 $Y=1.32
+ $X2=6.23 $Y2=1.485
r200 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.215 $Y=1.32
+ $X2=6.215 $Y2=0.74
r201 11 82 23.4391 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.76 $Y=1.76
+ $X2=4.76 $Y2=2.032
r202 11 13 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=4.76 $Y=1.76
+ $X2=4.76 $Y2=0.825
r203 7 80 19.0988 $w=1.8e-07 $l=2.73e-07 $layer=POLY_cond $X=4.29 $Y=2.305
+ $X2=4.29 $Y2=2.032
r204 7 9 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=4.29 $Y=2.305
+ $X2=4.29 $Y2=2.75
r205 2 73 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=5.31
+ $Y=2.12 $X2=5.48 $Y2=2.265
r206 1 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.345
+ $Y=0.395 $X2=5.485 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%A_678_392# 1 2 9 13 17 21 25 26 30 31 33 37
+ 38 43
c103 33 0 1.4938e-19 $X=5.325 $Y=1.485
c104 21 0 1.64715e-19 $X=5.725 $Y=2.54
c105 17 0 3.11092e-19 $X=5.7 $Y=0.715
r106 43 44 3.46264 $w=3.48e-07 $l=2.5e-08 $layer=POLY_cond $X=5.7 $Y=1.53
+ $X2=5.725 $Y2=1.53
r107 40 41 6.92529 $w=3.48e-07 $l=5e-08 $layer=POLY_cond $X=5.22 $Y=1.53
+ $X2=5.27 $Y2=1.53
r108 37 38 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=2.225
+ $X2=3.62 $Y2=2.06
r109 34 43 51.9397 $w=3.48e-07 $l=3.75e-07 $layer=POLY_cond $X=5.325 $Y=1.53
+ $X2=5.7 $Y2=1.53
r110 34 41 7.61782 $w=3.48e-07 $l=5.5e-08 $layer=POLY_cond $X=5.325 $Y=1.53
+ $X2=5.27 $Y2=1.53
r111 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.325
+ $Y=1.485 $X2=5.325 $Y2=1.485
r112 31 33 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=4.72 $Y=1.485
+ $X2=5.325 $Y2=1.485
r113 30 31 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.635 $Y=1.32
+ $X2=4.72 $Y2=1.485
r114 29 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.635 $Y=1.055
+ $X2=4.635 $Y2=1.32
r115 26 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.88 $Y=0.89
+ $X2=4.185 $Y2=0.89
r116 25 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.55 $Y=0.89
+ $X2=4.635 $Y2=1.055
r117 25 28 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.55 $Y=0.89
+ $X2=4.185 $Y2=0.89
r118 23 26 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.795 $Y=1.055
+ $X2=3.88 $Y2=0.89
r119 23 38 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=3.795 $Y=1.055
+ $X2=3.795 $Y2=2.06
r120 19 44 18.1727 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.725 $Y=1.74
+ $X2=5.725 $Y2=1.53
r121 19 21 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=5.725 $Y=1.74
+ $X2=5.725 $Y2=2.54
r122 15 43 22.4912 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.7 $Y=1.32 $X2=5.7
+ $Y2=1.53
r123 15 17 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=5.7 $Y=1.32
+ $X2=5.7 $Y2=0.715
r124 11 41 22.4912 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.27 $Y=1.32
+ $X2=5.27 $Y2=1.53
r125 11 13 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=5.27 $Y=1.32
+ $X2=5.27 $Y2=0.715
r126 7 40 18.1727 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.22 $Y=1.74
+ $X2=5.22 $Y2=1.53
r127 7 9 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=5.22 $Y=1.74 $X2=5.22
+ $Y2=2.54
r128 2 37 300 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=2 $X=3.39
+ $Y=1.96 $X2=3.525 $Y2=2.225
r129 1 28 91 $w=1.7e-07 $l=7.10634e-07 $layer=licon1_NDIFF $count=2 $X=3.68
+ $Y=0.395 $X2=4.185 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%VPWR 1 2 3 4 5 6 21 25 29 33 35 37 39 41 46
+ 62 67 72 78 81 85 89 91 94 98
r98 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r99 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r100 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r101 87 89 10.7168 $w=8.23e-07 $l=1.05e-07 $layer=LI1_cond $X=5.04 $Y=3.002
+ $X2=5.145 $Y2=3.002
r102 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 84 87 0.869875 $w=8.23e-07 $l=6e-08 $layer=LI1_cond $X=4.98 $Y=3.002
+ $X2=5.04 $Y2=3.002
r104 84 85 17.7483 $w=8.23e-07 $l=5.9e-07 $layer=LI1_cond $X=4.98 $Y=3.002
+ $X2=4.39 $Y2=3.002
r105 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 76 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 76 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 73 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=3.33
+ $X2=6.98 $Y2=3.33
r111 73 75 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.145 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 72 97 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.937 $Y2=3.33
r113 72 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 71 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r116 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r117 68 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=3.33
+ $X2=5.98 $Y2=3.33
r118 68 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.145 $Y=3.33
+ $X2=6.48 $Y2=3.33
r119 67 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.815 $Y=3.33
+ $X2=6.98 $Y2=3.33
r120 67 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r122 66 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 65 89 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=5.145 $Y2=3.33
r124 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r125 62 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.98 $Y2=3.33
r126 62 65 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.52 $Y2=3.33
r127 60 85 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=4.39 $Y2=3.33
r128 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 55 81 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.59 $Y2=3.33
r132 55 57 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=3.33 $X2=3.12
+ $Y2=3.33
r133 53 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r135 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 50 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r138 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 47 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r140 47 49 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r141 46 81 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.59 $Y2=3.33
r142 46 52 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r143 44 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r145 41 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r146 41 43 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r147 39 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r148 39 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r149 39 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 35 97 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.937 $Y2=3.33
r151 35 37 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.405
r152 31 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=3.245
+ $X2=6.98 $Y2=3.33
r153 31 33 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=6.98 $Y=3.245
+ $X2=6.98 $Y2=2.265
r154 27 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=3.245
+ $X2=5.98 $Y2=3.33
r155 27 29 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=5.98 $Y=3.245
+ $X2=5.98 $Y2=2.325
r156 23 81 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=3.245
+ $X2=2.59 $Y2=3.33
r157 23 25 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=2.59 $Y=3.245
+ $X2=2.59 $Y2=2.815
r158 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r159 19 21 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.455
r160 6 37 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=2.405
r161 5 33 300 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_PDIFF $count=2 $X=6.845
+ $Y=1.84 $X2=6.98 $Y2=2.265
r162 4 29 300 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_PDIFF $count=2 $X=5.815
+ $Y=2.12 $X2=5.98 $Y2=2.325
r163 3 84 300 $w=1.7e-07 $l=6.99285e-07 $layer=licon1_PDIFF $count=2 $X=4.38
+ $Y=2.54 $X2=4.98 $Y2=2.755
r164 2 25 600 $w=1.7e-07 $l=9.87269e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.96 $X2=2.59 $Y2=2.815
r165 1 21 300 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_PDIFF $count=2 $X=0.615
+ $Y=2.12 $X2=0.8 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%Q 1 2 3 4 15 17 19 21 22 27 31 33 37 39 40
+ 41 52
c73 22 0 1.66129e-19 $X=6.615 $Y=1.065
c74 17 0 1.64715e-19 $X=6.48 $Y=1.99
r75 51 52 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.43 $Y=1.985
+ $X2=7.315 $Y2=1.985
r76 41 51 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=7.92 $Y=1.985
+ $X2=7.43 $Y2=1.985
r77 41 45 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.985
+ $X2=7.92 $Y2=1.82
r78 40 45 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.82
r79 39 40 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.665
r80 38 39 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.92 $Y=1.15
+ $X2=7.92 $Y2=1.295
r81 34 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.545 $Y=1.065
+ $X2=7.42 $Y2=1.065
r82 33 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.065
+ $X2=7.92 $Y2=1.15
r83 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.805 $Y=1.065
+ $X2=7.545 $Y2=1.065
r84 29 51 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=2.15
+ $X2=7.43 $Y2=1.985
r85 29 31 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.43 $Y=2.15
+ $X2=7.43 $Y2=2.4
r86 25 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.42 $Y=0.98
+ $X2=7.42 $Y2=1.065
r87 25 27 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=7.42 $Y=0.98
+ $X2=7.42 $Y2=0.515
r88 24 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=1.905
+ $X2=6.48 $Y2=1.905
r89 24 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.645 $Y=1.905
+ $X2=7.315 $Y2=1.905
r90 21 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=1.065
+ $X2=7.42 $Y2=1.065
r91 21 22 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.295 $Y=1.065
+ $X2=6.615 $Y2=1.065
r92 17 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=1.99 $X2=6.48
+ $Y2=1.905
r93 17 19 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=6.48 $Y=1.99
+ $X2=6.48 $Y2=2.815
r94 13 22 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=6.44 $Y=0.98
+ $X2=6.615 $Y2=1.065
r95 13 15 15.311 $w=3.48e-07 $l=4.65e-07 $layer=LI1_cond $X=6.44 $Y=0.98
+ $X2=6.44 $Y2=0.515
r96 4 51 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.43 $Y2=1.985
r97 4 31 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=7.295
+ $Y=1.84 $X2=7.43 $Y2=2.4
r98 3 36 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.84 $X2=6.48 $Y2=1.985
r99 3 19 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.84 $X2=6.48 $Y2=2.815
r100 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.37 $X2=7.38 $Y2=0.515
r101 1 15 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=6.29
+ $Y=0.37 $X2=6.44 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 46 48 53 61 70 74 80 83 86 89 93
r112 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r113 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r114 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r115 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r116 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r118 78 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r119 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r120 75 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=6.95
+ $Y2=0
r121 75 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=0
+ $X2=7.44 $Y2=0
r122 74 92 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.937 $Y2=0
r123 74 77 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.44 $Y2=0
r124 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r125 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r126 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=0 $X2=6.95
+ $Y2=0
r127 70 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.785 $Y=0
+ $X2=6.48 $Y2=0
r128 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r129 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r130 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r131 66 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.015
+ $Y2=0
r132 66 68 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.52
+ $Y2=0
r133 65 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r134 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r135 62 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=2.98
+ $Y2=0
r136 62 64 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.145 $Y=0
+ $X2=4.56 $Y2=0
r137 61 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.89 $Y=0 $X2=5.015
+ $Y2=0
r138 61 64 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.89 $Y=0 $X2=4.56
+ $Y2=0
r139 60 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r140 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r141 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r142 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r143 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r144 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r145 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r146 54 56 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r147 53 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.98
+ $Y2=0
r148 53 59 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=0
+ $X2=2.64 $Y2=0
r149 51 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r150 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r151 48 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r152 48 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r153 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r154 46 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r155 44 68 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.52
+ $Y2=0
r156 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.915
+ $Y2=0
r157 43 72 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=6.48
+ $Y2=0
r158 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=5.915
+ $Y2=0
r159 39 92 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.937 $Y2=0
r160 39 41 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.62
r161 35 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=0.085
+ $X2=6.95 $Y2=0
r162 35 37 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=6.95 $Y=0.085
+ $X2=6.95 $Y2=0.62
r163 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=0.085
+ $X2=5.915 $Y2=0
r164 31 33 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=5.915 $Y=0.085
+ $X2=5.915 $Y2=0.59
r165 27 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.015 $Y=0.085
+ $X2=5.015 $Y2=0
r166 27 29 34.1123 $w=2.48e-07 $l=7.4e-07 $layer=LI1_cond $X=5.015 $Y=0.085
+ $X2=5.015 $Y2=0.825
r167 23 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0
r168 23 25 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0.54
r169 19 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r170 19 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r171 6 41 182 $w=1.7e-07 $l=3.22102e-07 $layer=licon1_NDIFF $count=1 $X=7.715
+ $Y=0.37 $X2=7.88 $Y2=0.62
r172 5 37 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.37 $X2=6.95 $Y2=0.62
r173 4 33 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=5.775
+ $Y=0.395 $X2=5.915 $Y2=0.59
r174 3 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.835
+ $Y=0.615 $X2=4.975 $Y2=0.825
r175 2 25 91 $w=1.7e-07 $l=6.29285e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.37 $X2=2.98 $Y2=0.54
r176 1 21 182 $w=1.7e-07 $l=3.42783e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.575 $X2=0.79 $Y2=0.325
.ends


* File: sky130_fd_sc_ms__sdfstp_2.spice
* Created: Wed Sep  2 12:31:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfstp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfstp_2  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1043 N_VGND_M1043_d N_SCE_M1043_g N_A_27_74#_M1043_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.09975 AS=0.1197 PD=0.895 PS=1.41 NRD=37.14 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1038 A_239_74# N_A_27_74#_M1038_g N_VGND_M1043_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.09975 PD=0.66 PS=0.895 NRD=18.564 NRS=18.564 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1028 N_A_293_464#_M1028_d N_D_M1028_g A_239_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1039 A_403_74# N_SCE_M1039_g N_A_293_464#_M1028_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_SCD_M1035_g A_403_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0672 PD=1.41 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75002.1 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_CLK_M1012_g N_A_608_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1006 N_A_795_74#_M1006_d N_A_608_74#_M1006_g N_VGND_M1012_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.1295 PD=2.04 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_991_81#_M1024_d N_A_608_74#_M1024_g N_A_293_464#_M1024_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1176 PD=1.03 PS=1.4 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1031 A_1143_81# N_A_795_74#_M1031_g N_A_991_81#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1281 PD=0.63 PS=1.03 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1185_55#_M1020_g A_1143_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.2316 AS=0.0441 PD=2.11 PS=0.63 NRD=141.828 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1026 A_1429_74# N_A_991_81#_M1026_g N_A_1185_55#_M1026_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_SET_B_M1027_g A_1429_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.108328 AS=0.0504 PD=0.919245 PS=0.66 NRD=24.276 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1029 N_A_1641_74#_M1029_d N_A_991_81#_M1029_g N_VGND_M1027_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.165072 PD=0.92 PS=1.40075 NRD=0 NRS=29.052 M=1 R=4.26667
+ SA=75000.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1033 N_A_1641_74#_M1029_d N_A_991_81#_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2336 PD=0.92 PS=2.01 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.3 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1001 N_A_1804_424#_M1001_d N_A_795_74#_M1001_g N_A_1641_74#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2272 AS=0.0896 PD=1.99 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1036 N_A_1804_424#_M1036_d N_A_795_74#_M1036_g N_A_1641_74#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.121962 AS=0.0896 PD=1.19547 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.7 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1044 A_2141_74# N_A_608_74#_M1044_g N_A_1804_424#_M1036_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0800377 PD=0.66 PS=0.784528 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1041 A_2219_74# N_A_2186_367#_M1041_g A_2141_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_SET_B_M1025_g A_2219_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.14385 AS=0.0882 PD=1.105 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75002.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1030 N_A_2186_367#_M1030_d N_A_1804_424#_M1030_g N_VGND_M1025_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.14385 PD=1.41 PS=1.105 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75003 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1804_424#_M1022_g N_A_2611_98#_M1022_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.124754 AS=0.1824 PD=1.0342 PS=1.85 NRD=17.34 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1014 N_Q_M1014_d N_A_2611_98#_M1014_g N_VGND_M1022_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.144246 PD=1.02 PS=1.1958 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1037 N_Q_M1014_d N_A_2611_98#_M1037_g N_VGND_M1037_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.222 PD=1.02 PS=2.08 NRD=0 NRS=2.424 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_SCE_M1015_g N_A_27_74#_M1015_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.1792 PD=0.91 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1016 A_209_464# N_SCE_M1016_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.0864 PD=0.88 PS=0.91 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.6
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1023 N_A_293_464#_M1023_d N_D_M1023_g A_209_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.144 AS=0.0768 PD=1.09 PS=0.88 NRD=26.1616 NRS=19.9955 M=1 R=3.55556
+ SA=90001.1 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1005 A_419_464# N_A_27_74#_M1005_g N_A_293_464#_M1023_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.144 PD=0.88 PS=1.09 NRD=19.9955 NRS=26.1616 M=1
+ R=3.55556 SA=90001.7 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1017 N_VPWR_M1017_d N_SCD_M1017_g A_419_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.2653 AS=0.0768 PD=2.32 PS=0.88 NRD=23.0687 NRS=19.9955 M=1 R=3.55556
+ SA=90002.1 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1032 N_VPWR_M1032_d N_CLK_M1032_g N_A_608_74#_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1040 N_A_795_74#_M1040_d N_A_608_74#_M1040_g N_VPWR_M1032_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2908 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1034 N_A_991_81#_M1034_d N_A_795_74#_M1034_g N_A_293_464#_M1034_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.085925 AS=0.1176 PD=0.905 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1018 A_1120_483# N_A_608_74#_M1018_g N_A_991_81#_M1034_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0794 AS=0.085925 PD=0.86 PS=0.905 NRD=62.8627 NRS=39.8531 M=1
+ R=2.33333 SA=90000.6 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1042 N_VPWR_M1042_d N_A_1185_55#_M1042_g A_1120_483# VPB PSHORT L=0.18 W=0.42
+ AD=0.10605 AS=0.0794 PD=0.925 PS=0.86 NRD=0 NRS=62.8627 M=1 R=2.33333
+ SA=90000.9 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1011 N_A_1185_55#_M1011_d N_A_991_81#_M1011_g N_VPWR_M1042_d VPB PSHORT L=0.18
+ W=0.42 AD=0.06615 AS=0.10605 PD=0.735 PS=0.925 NRD=0 NRS=105.533 M=1 R=2.33333
+ SA=90001.6 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1021 N_VPWR_M1021_d N_SET_B_M1021_g N_A_1185_55#_M1011_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1029 AS=0.06615 PD=0.863333 PS=0.735 NRD=84.4145 NRS=18.7544 M=1
+ R=2.33333 SA=90002.1 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1000 N_A_1587_379#_M1000_d N_A_991_81#_M1000_g N_VPWR_M1021_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.2058 PD=1.11 PS=1.72667 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90001.5 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1007 N_A_1587_379#_M1000_d N_A_991_81#_M1007_g N_VPWR_M1007_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.2226 PD=1.11 PS=2.21 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90001.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1003 N_A_1587_379#_M1003_d N_A_608_74#_M1003_g N_A_1804_424#_M1003_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.2772 PD=1.11 PS=2.34 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90000.2 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1010 N_A_1587_379#_M1003_d N_A_608_74#_M1010_g N_A_1804_424#_M1010_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.2268 PD=1.11 PS=1.86667 NRD=0 NRS=35.1645
+ M=1 R=4.66667 SA=90000.7 SB=90001 A=0.1512 P=2.04 MULT=1
MM1019 A_2144_508# N_A_795_74#_M1019_g N_A_1804_424#_M1010_s VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.1134 PD=0.63 PS=0.933333 NRD=23.443 NRS=60.9715 M=1
+ R=2.33333 SA=90001.4 SB=90001 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_A_2186_367#_M1008_g A_2144_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333 SA=90001.8
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1013 N_A_1804_424#_M1013_d N_SET_B_M1013_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.0567 PD=1.37 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90002.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_A_1804_424#_M1009_g N_A_2186_367#_M1009_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_1804_424#_M1002_g N_A_2611_98#_M1002_s VPB PSHORT
+ L=0.18 W=1 AD=0.167453 AS=0.265 PD=1.36321 PS=2.53 NRD=8.8453 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1002_d N_A_2611_98#_M1004_g N_Q_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.187547 AS=0.1512 PD=1.52679 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1045 N_VPWR_M1045_d N_A_2611_98#_M1045_g N_Q_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX46_noxref VNB VPB NWDIODE A=28.3836 P=34.24
c_166 VNB 0 7.29682e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sdfstp_2.pxi.spice"
*
.ends
*
*

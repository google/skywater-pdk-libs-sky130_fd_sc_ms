* File: sky130_fd_sc_ms__or4_1.spice
* Created: Fri Aug 28 18:08:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4_1.pex.spice"
.subckt sky130_fd_sc_ms__or4_1  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1003 N_A_44_392#_M1003_d N_D_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.19525 PD=0.83 PS=1.81 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.3
+ SB=75002.5 A=0.0825 P=1.4 MULT=1
MM1002 N_VGND_M1002_d N_C_M1002_g N_A_44_392#_M1003_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.1674 AS=0.077 PD=1.165 PS=0.83 NRD=32.724 NRS=0 M=1 R=3.66667 SA=75000.7
+ SB=75002 A=0.0825 P=1.4 MULT=1
MM1006 N_A_44_392#_M1006_d N_B_M1006_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.121 AS=0.1674 PD=0.99 PS=1.165 NRD=17.448 NRS=33.816 M=1 R=3.66667
+ SA=75001.4 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_44_392#_M1006_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.107506 AS=0.121 PD=0.937984 PS=0.99 NRD=17.448 NRS=17.448 M=1 R=3.66667
+ SA=75002 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1007 N_X_M1007_d N_A_44_392#_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.144644 PD=2.05 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_136_392# N_D_M1001_g N_A_44_392#_M1001_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90002.4
+ A=0.18 P=2.36 MULT=1
MM1008 A_220_392# N_C_M1008_g A_136_392# VPB PSHORT L=0.18 W=1 AD=0.195 AS=0.12
+ PD=1.39 PS=1.24 NRD=27.5603 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90002
+ A=0.18 P=2.36 MULT=1
MM1005 A_334_392# N_B_M1005_g A_220_392# VPB PSHORT L=0.18 W=1 AD=0.195 AS=0.195
+ PD=1.39 PS=1.39 NRD=27.5603 NRS=27.5603 M=1 R=5.55556 SA=90001.2 SB=90001.4
+ A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g A_334_392# VPB PSHORT L=0.18 W=1 AD=0.254717
+ AS=0.195 PD=1.53774 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90001.7
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_44_392#_M1000_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.285283 PD=2.8 PS=1.72226 NRD=0 NRS=41.3306 M=1 R=6.22222
+ SA=90002.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__or4_1.pxi.spice"
*
.ends
*
*

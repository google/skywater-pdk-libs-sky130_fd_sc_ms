* File: sky130_fd_sc_ms__nand2b_1.pex.spice
* Created: Wed Sep  2 12:13:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND2B_1%A_N 3 7 9 10 17
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.465 $X2=0.61 $Y2=1.465
r36 15 17 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.61 $Y2=1.465
r37 13 15 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r38 10 18 2.74101 $w=4.78e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.61 $Y2=1.54
r39 9 18 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.54 $X2=0.61
+ $Y2=1.54
r40 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r41 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.835
r42 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r43 1 3 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_1%B 3 7 9 12 13
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.515
+ $X2=1.18 $Y2=1.68
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.515
+ $X2=1.18 $Y2=1.35
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.515 $X2=1.18 $Y2=1.515
r45 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.515
r46 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.27 $Y=0.74 $X2=1.27
+ $Y2=1.35
r47 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.175 $Y=2.4
+ $X2=1.175 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_1%A_27_112# 1 2 9 13 17 21 22 23 28 30 32 33
+ 34
c74 28 0 1.74227e-19 $X=1.6 $Y=1.95
c75 13 0 1.78244e-19 $X=1.675 $Y=2.4
r76 33 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.465
+ $X2=1.75 $Y2=1.63
r77 33 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.465
+ $X2=1.75 $Y2=1.3
r78 32 35 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.465
+ $X2=1.715 $Y2=1.63
r79 32 34 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.465
+ $X2=1.715 $Y2=1.3
r80 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.465 $X2=1.75 $Y2=1.465
r81 28 35 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.6 $Y=1.95 $X2=1.6
+ $Y2=1.63
r82 25 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.6 $Y=1.13 $X2=1.6
+ $Y2=1.3
r83 24 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r84 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=1.6 $Y2=1.95
r85 23 24 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=0.445 $Y2=2.035
r86 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.045
+ $X2=1.6 $Y2=1.13
r87 21 22 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=1.515 $Y=1.045
+ $X2=0.38 $Y2=1.045
r88 15 22 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.247 $Y=0.96
+ $X2=0.38 $Y2=1.045
r89 15 17 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=0.247 $Y=0.96
+ $X2=0.247 $Y2=0.835
r90 13 38 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.675 $Y=2.4
+ $X2=1.675 $Y2=1.63
r91 9 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.66 $Y=0.74 $X2=1.66
+ $Y2=1.3
r92 2 30 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r93 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_1%VPWR 1 2 11 17 20 21 22 29 30 33
r30 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 24 33 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.782 $Y2=3.33
r35 24 26 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 20 26 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 20 21 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.902 $Y2=3.33
r40 19 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=3.33 $X2=2.16
+ $Y2=3.33
r41 19 21 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.902 $Y2=3.33
r42 15 21 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.902 $Y=3.245
+ $X2=1.902 $Y2=3.33
r43 15 17 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=1.902 $Y=3.245
+ $X2=1.902 $Y2=2.815
r44 11 14 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=0.782 $Y=2.455
+ $X2=0.782 $Y2=2.795
r45 9 33 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=3.245
+ $X2=0.782 $Y2=3.33
r46 9 14 19.5698 $w=2.63e-07 $l=4.5e-07 $layer=LI1_cond $X=0.782 $Y=3.245
+ $X2=0.782 $Y2=2.795
r47 2 17 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.84 $X2=1.9 $Y2=2.815
r48 1 14 600 $w=1.7e-07 $l=1.06156e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.82 $Y2=2.795
r49 1 11 600 $w=1.7e-07 $l=7.18749e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.82 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_1%Y 1 2 7 11 14 15 16 17 21
c36 16 0 1.78244e-19 $X=1.2 $Y=2.405
r37 16 21 2.36995 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=2.375
+ $X2=1.325 $Y2=2.46
r38 16 17 7.47549 $w=4.78e-07 $l=3e-07 $layer=LI1_cond $X=1.325 $Y=2.475
+ $X2=1.325 $Y2=2.775
r39 16 21 0.373774 $w=4.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.325 $Y=2.475
+ $X2=1.325 $Y2=2.46
r40 14 15 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.17 $Y=2.29
+ $X2=2.17 $Y2=1.13
r41 9 15 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=2.055 $Y=0.93 $X2=2.055
+ $Y2=1.13
r42 9 11 11.9566 $w=3.98e-07 $l=4.15e-07 $layer=LI1_cond $X=2.055 $Y=0.93
+ $X2=2.055 $Y2=0.515
r43 8 16 6.69163 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.565 $Y=2.375
+ $X2=1.325 $Y2=2.375
r44 7 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=2.375
+ $X2=2.17 $Y2=2.29
r45 7 8 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.085 $Y=2.375
+ $X2=1.565 $Y2=2.375
r46 2 16 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.265
+ $Y=1.84 $X2=1.4 $Y2=2.455
r47 1 11 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=1.735
+ $Y=0.37 $X2=1.94 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_1%VGND 1 6 8 10 17 18 21
r22 21 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r23 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r24 15 21 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=0.885
+ $Y2=0
r25 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=2.16
+ $Y2=0
r26 13 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r27 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 10 21 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.885
+ $Y2=0
r29 10 12 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r30 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r31 8 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r32 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 4 21 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0.085
+ $X2=0.885 $Y2=0
r34 4 6 11.0682 $w=6.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.885 $Y=0.085
+ $X2=0.885 $Y2=0.705
r35 1 6 91 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.56 $X2=1.055 $Y2=0.705
.ends


* File: sky130_fd_sc_ms__o221ai_2.pxi.spice
* Created: Fri Aug 28 17:57:32 2020
* 
x_PM_SKY130_FD_SC_MS__O221AI_2%C1 N_C1_M1017_g N_C1_M1013_g N_C1_M1018_g
+ N_C1_M1014_g C1 N_C1_c_101_n N_C1_c_102_n PM_SKY130_FD_SC_MS__O221AI_2%C1
x_PM_SKY130_FD_SC_MS__O221AI_2%B1 N_B1_c_140_n N_B1_M1008_g N_B1_c_141_n
+ N_B1_M1012_g N_B1_M1010_g N_B1_M1016_g N_B1_c_156_p N_B1_c_143_n N_B1_c_144_n
+ B1 B1 B1 N_B1_c_145_n PM_SKY130_FD_SC_MS__O221AI_2%B1
x_PM_SKY130_FD_SC_MS__O221AI_2%B2 N_B2_c_235_n N_B2_M1002_g N_B2_M1000_g
+ N_B2_c_232_n N_B2_M1009_g N_B2_M1004_g B2 N_B2_c_234_n
+ PM_SKY130_FD_SC_MS__O221AI_2%B2
x_PM_SKY130_FD_SC_MS__O221AI_2%A1 N_A1_M1003_g N_A1_M1006_g N_A1_M1015_g
+ N_A1_M1019_g N_A1_c_285_n N_A1_c_286_n N_A1_c_309_p N_A1_c_304_n A1
+ N_A1_c_287_n N_A1_c_288_n PM_SKY130_FD_SC_MS__O221AI_2%A1
x_PM_SKY130_FD_SC_MS__O221AI_2%A2 N_A2_M1001_g N_A2_M1005_g N_A2_M1007_g
+ N_A2_M1011_g A2 N_A2_c_372_n N_A2_c_373_n PM_SKY130_FD_SC_MS__O221AI_2%A2
x_PM_SKY130_FD_SC_MS__O221AI_2%VPWR N_VPWR_M1013_s N_VPWR_M1014_s N_VPWR_M1010_s
+ N_VPWR_M1015_s N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n
+ N_VPWR_c_427_n VPWR N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_430_n
+ N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_422_n PM_SKY130_FD_SC_MS__O221AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O221AI_2%Y N_Y_M1017_d N_Y_M1013_d N_Y_M1002_d N_Y_M1005_d
+ N_Y_c_506_n N_Y_c_525_n N_Y_c_496_n N_Y_c_512_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_MS__O221AI_2%Y
x_PM_SKY130_FD_SC_MS__O221AI_2%A_379_368# N_A_379_368#_M1008_d
+ N_A_379_368#_M1009_s N_A_379_368#_c_553_n N_A_379_368#_c_554_n
+ N_A_379_368#_c_555_n PM_SKY130_FD_SC_MS__O221AI_2%A_379_368#
x_PM_SKY130_FD_SC_MS__O221AI_2%A_779_368# N_A_779_368#_M1006_d
+ N_A_779_368#_M1007_s N_A_779_368#_c_581_n N_A_779_368#_c_589_n
+ N_A_779_368#_c_582_n PM_SKY130_FD_SC_MS__O221AI_2%A_779_368#
x_PM_SKY130_FD_SC_MS__O221AI_2%A_27_74# N_A_27_74#_M1017_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1012_d N_A_27_74#_M1004_s N_A_27_74#_c_609_n N_A_27_74#_c_610_n
+ N_A_27_74#_c_611_n N_A_27_74#_c_612_n N_A_27_74#_c_613_n N_A_27_74#_c_614_n
+ N_A_27_74#_c_649_p N_A_27_74#_c_615_n N_A_27_74#_c_634_n N_A_27_74#_c_616_n
+ PM_SKY130_FD_SC_MS__O221AI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O221AI_2%A_311_85# N_A_311_85#_M1012_s N_A_311_85#_M1000_d
+ N_A_311_85#_M1016_s N_A_311_85#_M1001_d N_A_311_85#_M1019_s
+ N_A_311_85#_c_660_n N_A_311_85#_c_661_n N_A_311_85#_c_662_n
+ N_A_311_85#_c_675_n N_A_311_85#_c_663_n N_A_311_85#_c_686_n
+ N_A_311_85#_c_664_n N_A_311_85#_c_665_n N_A_311_85#_c_666_n
+ N_A_311_85#_c_667_n N_A_311_85#_c_668_n N_A_311_85#_c_669_n
+ N_A_311_85#_c_670_n PM_SKY130_FD_SC_MS__O221AI_2%A_311_85#
x_PM_SKY130_FD_SC_MS__O221AI_2%VGND N_VGND_M1003_d N_VGND_M1011_s N_VGND_c_739_n
+ N_VGND_c_740_n VGND N_VGND_c_741_n N_VGND_c_742_n N_VGND_c_743_n
+ N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n PM_SKY130_FD_SC_MS__O221AI_2%VGND
cc_1 VNB N_C1_M1017_g 0.0274728f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_C1_M1013_g 0.00155225f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_3 VNB N_C1_M1018_g 0.025282f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_C1_M1014_g 0.00393622f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_5 VNB N_C1_c_101_n 0.00617983f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_6 VNB N_C1_c_102_n 0.0863785f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_7 VNB N_B1_c_140_n 0.0331484f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_8 VNB N_B1_c_141_n 0.0215291f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.63
cc_9 VNB N_B1_M1016_g 0.021044f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_10 VNB N_B1_c_143_n 0.00167757f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_11 VNB N_B1_c_144_n 0.0268438f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_12 VNB N_B1_c_145_n 0.0119268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B2_M1000_g 0.0192446f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_14 VNB N_B2_c_232_n 0.0331801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_M1004_g 0.0206166f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_16 VNB N_B2_c_234_n 8.29228e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_17 VNB N_A1_M1003_g 0.0211602f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_18 VNB N_A1_M1019_g 0.0288546f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_19 VNB N_A1_c_285_n 0.00167078f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_20 VNB N_A1_c_286_n 0.0270321f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_21 VNB N_A1_c_287_n 0.0288655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_288_n 0.0202222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1001_g 0.0219922f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_24 VNB N_A2_M1011_g 0.0214811f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_25 VNB N_A2_c_372_n 0.00139482f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_26 VNB N_A2_c_373_n 0.036614f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_27 VNB N_VPWR_c_422_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.00220761f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_29 VNB N_A_27_74#_c_609_n 0.0275751f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_30 VNB N_A_27_74#_c_610_n 0.00664238f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_A_27_74#_c_611_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_612_n 0.0062256f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_33 VNB N_A_27_74#_c_613_n 0.0143267f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.465
cc_34 VNB N_A_27_74#_c_614_n 0.00353358f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_35 VNB N_A_27_74#_c_615_n 0.0147249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_616_n 0.00154467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_311_85#_c_660_n 0.00367062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_311_85#_c_661_n 0.00702435f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_39 VNB N_A_311_85#_c_662_n 0.00454744f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_40 VNB N_A_311_85#_c_663_n 0.0135463f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_41 VNB N_A_311_85#_c_664_n 0.00924121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_311_85#_c_665_n 0.00789247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_311_85#_c_666_n 0.00316307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_311_85#_c_667_n 0.0148853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_311_85#_c_668_n 0.0249008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_311_85#_c_669_n 0.00238018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_311_85#_c_670_n 0.00312418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_739_n 0.0108406f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_49 VNB N_VGND_c_740_n 0.00891632f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.59
cc_50 VNB N_VGND_c_741_n 0.0937136f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_51 VNB N_VGND_c_742_n 0.0189057f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.465
cc_52 VNB N_VGND_c_743_n 0.0178712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_744_n 0.34449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_745_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_746_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_C1_M1013_g 0.0247757f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_57 VPB N_C1_M1014_g 0.0240263f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_58 VPB N_C1_c_101_n 0.0106052f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_59 VPB N_B1_c_140_n 0.00566622f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_60 VPB N_B1_M1008_g 0.0230334f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_61 VPB N_B1_M1010_g 0.0214037f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_62 VPB N_B1_c_143_n 0.0025087f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_63 VPB N_B1_c_144_n 0.0056302f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_64 VPB N_B1_c_145_n 0.00242791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B2_c_235_n 0.0157946f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_66 VPB N_B2_c_232_n 0.0103032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_B2_M1009_g 0.0205f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_68 VPB N_B2_c_234_n 0.0027336f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_69 VPB N_A1_M1006_g 0.0214037f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_70 VPB N_A1_M1015_g 0.0227838f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_71 VPB N_A1_c_285_n 0.00264918f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_72 VPB N_A1_c_286_n 0.00564554f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_73 VPB N_A1_c_287_n 0.00581685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A1_c_288_n 0.0205668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A2_M1005_g 0.0208757f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_76 VPB N_A2_M1007_g 0.0203097f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_77 VPB N_A2_c_372_n 0.00251564f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_78 VPB N_A2_c_373_n 0.00465871f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_79 VPB N_VPWR_c_423_n 0.011928f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.59
cc_80 VPB N_VPWR_c_424_n 0.0488269f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_81 VPB N_VPWR_c_425_n 0.00888209f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_82 VPB N_VPWR_c_426_n 0.0121872f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.465
cc_83 VPB N_VPWR_c_427_n 0.0387956f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.465
cc_84 VPB N_VPWR_c_428_n 0.0185562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_429_n 0.0401011f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_430_n 0.0389457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_431_n 0.0207863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_432_n 0.00631492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_422_n 0.0685364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB Y 0.00126143f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_91 VPB Y 0.00202354f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_92 VPB N_A_379_368#_c_553_n 0.00267435f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_93 VPB N_A_379_368#_c_554_n 0.00237125f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_94 VPB N_A_379_368#_c_555_n 0.00237138f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_95 VPB N_A_779_368#_c_581_n 0.0042639f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_96 VPB N_A_779_368#_c_582_n 0.00237138f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_97 N_C1_M1018_g N_B1_c_140_n 2.45528e-19 $X=0.925 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_98 N_C1_c_102_n N_B1_c_140_n 0.00714113f $X=0.925 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_99 N_C1_M1014_g N_B1_M1008_g 0.0166303f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_100 N_C1_c_102_n N_B1_c_145_n 0.0120372f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_101 N_C1_M1013_g N_VPWR_c_424_n 0.00370078f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_102 N_C1_c_101_n N_VPWR_c_424_n 0.0219687f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_103 N_C1_c_102_n N_VPWR_c_424_n 0.00135527f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_104 N_C1_M1013_g N_VPWR_c_428_n 0.005209f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_105 N_C1_M1014_g N_VPWR_c_428_n 0.00461464f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_106 N_C1_M1013_g N_VPWR_c_431_n 4.49936e-19 $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_107 N_C1_M1014_g N_VPWR_c_431_n 0.00989081f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_108 N_C1_M1013_g N_VPWR_c_422_n 0.00986139f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_109 N_C1_M1014_g N_VPWR_c_422_n 0.00908554f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_110 N_C1_M1014_g N_Y_c_496_n 0.0208715f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_111 N_C1_M1017_g Y 0.00526147f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_112 N_C1_M1013_g Y 0.0154776f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_113 N_C1_M1018_g Y 0.0147581f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_114 N_C1_M1014_g Y 0.00220545f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_115 N_C1_c_101_n Y 0.0360521f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_116 N_C1_c_102_n Y 0.0228477f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_117 N_C1_M1013_g Y 0.00930908f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_118 N_C1_M1014_g Y 2.60789e-19 $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_119 N_C1_M1017_g N_A_27_74#_c_609_n 0.00161118f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_120 N_C1_c_101_n N_A_27_74#_c_609_n 0.0215684f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_121 N_C1_c_102_n N_A_27_74#_c_609_n 0.00196285f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_122 N_C1_M1017_g N_A_27_74#_c_610_n 0.0139957f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_123 N_C1_M1018_g N_A_27_74#_c_610_n 0.0132617f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_124 N_C1_M1018_g N_A_27_74#_c_614_n 0.00162302f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_125 N_C1_c_102_n N_A_27_74#_c_614_n 0.0015325f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_126 N_C1_M1018_g N_A_311_85#_c_662_n 5.96586e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_127 N_C1_M1017_g N_VGND_c_741_n 0.00278271f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_128 N_C1_M1018_g N_VGND_c_741_n 0.00278271f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_129 N_C1_M1017_g N_VGND_c_744_n 0.00357086f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_C1_M1018_g N_VGND_c_744_n 0.00358427f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B1_c_156_p N_B2_c_235_n 0.00970587f $X=3.075 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_132 N_B1_c_145_n N_B2_c_235_n 0.0109186f $X=2.275 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_133 N_B1_c_141_n N_B2_M1000_g 0.0167366f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_134 N_B1_c_140_n N_B2_c_232_n 0.0274805f $X=1.805 $Y=1.68 $X2=0 $Y2=0
cc_135 N_B1_M1008_g N_B2_c_232_n 0.044666f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_136 N_B1_c_156_p N_B2_c_232_n 0.00215676f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_137 N_B1_c_143_n N_B2_c_232_n 0.00132505f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B1_c_144_n N_B2_c_232_n 0.019357f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_139 N_B1_c_145_n N_B2_c_232_n 0.0144766f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_140 N_B1_M1010_g N_B2_M1009_g 0.0416294f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_141 N_B1_c_156_p N_B2_M1009_g 0.0119965f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_142 N_B1_c_143_n N_B2_M1009_g 0.00417437f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B1_c_145_n N_B2_M1009_g 9.55047e-19 $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_144 N_B1_M1016_g N_B2_M1004_g 0.0194733f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_145 N_B1_M1010_g N_B2_c_234_n 3.1567e-19 $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_146 N_B1_c_156_p N_B2_c_234_n 0.022819f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_147 N_B1_c_143_n N_B2_c_234_n 0.0266358f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B1_c_144_n N_B2_c_234_n 0.00118382f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_149 N_B1_c_145_n N_B2_c_234_n 0.0259253f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_150 N_B1_M1016_g N_A1_M1003_g 0.0172352f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_151 N_B1_M1010_g N_A1_M1006_g 0.0350668f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_152 N_B1_c_156_p N_A1_M1006_g 6.71906e-19 $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_153 N_B1_c_143_n N_A1_M1006_g 9.28507e-19 $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_154 N_B1_M1010_g N_A1_c_285_n 9.48357e-19 $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_155 N_B1_c_143_n N_A1_c_285_n 0.0360501f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_156 N_B1_c_144_n N_A1_c_285_n 0.00121489f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_157 N_B1_c_143_n N_A1_c_286_n 0.00121489f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_158 N_B1_c_144_n N_A1_c_286_n 0.017083f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_159 N_B1_M1010_g N_A1_c_304_n 6.86064e-19 $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_160 N_B1_c_156_p N_A1_c_304_n 0.0118526f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_161 N_B1_c_145_n N_VPWR_M1014_s 0.0116587f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_162 N_B1_c_156_p N_VPWR_M1010_s 0.0017942f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_163 N_B1_c_143_n N_VPWR_M1010_s 0.00112896f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_164 N_B1_M1010_g N_VPWR_c_425_n 0.00150765f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B1_M1008_g N_VPWR_c_429_n 0.00518311f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_166 N_B1_M1010_g N_VPWR_c_429_n 0.00518311f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_167 N_B1_M1008_g N_VPWR_c_431_n 0.00202669f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_168 N_B1_M1008_g N_VPWR_c_422_n 0.00983575f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_169 N_B1_M1010_g N_VPWR_c_422_n 0.0098206f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B1_c_156_p N_Y_M1002_d 0.00453933f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_171 N_B1_M1010_g N_Y_c_506_n 0.0167741f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_172 N_B1_c_156_p N_Y_c_506_n 0.016388f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_173 N_B1_c_144_n N_Y_c_506_n 2.00421e-19 $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_174 N_B1_c_140_n N_Y_c_496_n 3.17242e-19 $X=1.805 $Y=1.68 $X2=0 $Y2=0
cc_175 N_B1_M1008_g N_Y_c_496_n 0.0175862f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_176 N_B1_c_145_n N_Y_c_496_n 0.0609847f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_177 N_B1_M1008_g N_Y_c_512_n 7.36225e-19 $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B1_M1010_g N_Y_c_512_n 7.50787e-19 $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B1_c_156_p N_Y_c_512_n 0.0609847f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_180 N_B1_c_145_n Y 0.0433228f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_181 N_B1_c_145_n N_A_379_368#_M1008_d 0.00212405f $X=2.275 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_182 N_B1_c_156_p N_A_379_368#_M1009_s 0.0087506f $X=3.075 $Y=2.035 $X2=0
+ $Y2=0
cc_183 N_B1_c_143_n N_A_379_368#_M1009_s 0.00143139f $X=3.24 $Y=1.515 $X2=0
+ $Y2=0
cc_184 N_B1_M1008_g N_A_379_368#_c_554_n 0.00701668f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_185 N_B1_M1010_g N_A_379_368#_c_555_n 0.00687709f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_186 N_B1_c_141_n N_A_27_74#_c_610_n 5.53247e-19 $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_187 N_B1_c_141_n N_A_27_74#_c_612_n 0.00501983f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_188 N_B1_c_140_n N_A_27_74#_c_613_n 0.00565069f $X=1.805 $Y=1.68 $X2=0 $Y2=0
cc_189 N_B1_c_141_n N_A_27_74#_c_613_n 0.0133087f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_190 N_B1_c_145_n N_A_27_74#_c_613_n 0.0599647f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_191 N_B1_c_145_n N_A_27_74#_c_614_n 0.0205272f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_192 N_B1_M1016_g N_A_27_74#_c_615_n 0.00232271f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_193 N_B1_c_143_n N_A_27_74#_c_615_n 0.0178644f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_194 N_B1_c_144_n N_A_27_74#_c_615_n 0.00138314f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_195 N_B1_c_145_n N_A_27_74#_c_615_n 0.00496728f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_196 N_B1_M1016_g N_A_27_74#_c_634_n 0.0046047f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_197 N_B1_c_145_n N_A_27_74#_c_616_n 0.0156866f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_198 N_B1_c_141_n N_A_311_85#_c_660_n 0.00631411f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_199 N_B1_c_141_n N_A_311_85#_c_661_n 0.00817976f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_200 N_B1_c_141_n N_A_311_85#_c_662_n 0.0032816f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_201 N_B1_c_141_n N_A_311_85#_c_675_n 5.66812e-19 $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_202 N_B1_M1016_g N_A_311_85#_c_675_n 5.11849e-19 $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_203 N_B1_M1016_g N_A_311_85#_c_663_n 0.01343f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_204 N_B1_c_141_n N_VGND_c_741_n 8.82278e-19 $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_205 N_B1_M1016_g N_VGND_c_741_n 8.63546e-19 $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_206 N_B2_c_235_n N_VPWR_c_429_n 0.00333926f $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_207 N_B2_M1009_g N_VPWR_c_429_n 0.00333926f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_208 N_B2_c_235_n N_VPWR_c_422_n 0.00423273f $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_209 N_B2_M1009_g N_VPWR_c_422_n 0.00423405f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_210 N_B2_M1009_g N_Y_c_506_n 0.010049f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B2_c_235_n N_Y_c_496_n 0.0107581f $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_212 N_B2_c_235_n N_Y_c_512_n 0.00551896f $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_213 N_B2_M1009_g N_Y_c_512_n 0.00652147f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B2_c_235_n N_A_379_368#_c_553_n 0.0101522f $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_215 N_B2_M1009_g N_A_379_368#_c_553_n 0.0101083f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_216 N_B2_c_235_n N_A_379_368#_c_554_n 7.00934e-19 $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_217 N_B2_M1009_g N_A_379_368#_c_555_n 4.1224e-19 $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_218 N_B2_M1000_g N_A_27_74#_c_615_n 0.0156966f $X=2.345 $Y=0.795 $X2=0 $Y2=0
cc_219 N_B2_c_232_n N_A_27_74#_c_615_n 0.00126891f $X=2.755 $Y=1.68 $X2=0 $Y2=0
cc_220 N_B2_M1004_g N_A_27_74#_c_615_n 0.0127188f $X=2.775 $Y=0.795 $X2=0 $Y2=0
cc_221 N_B2_c_234_n N_A_27_74#_c_615_n 0.0247257f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_222 N_B2_M1000_g N_A_311_85#_c_660_n 5.66812e-19 $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_223 N_B2_M1000_g N_A_311_85#_c_661_n 0.00817976f $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_224 N_B2_M1000_g N_A_311_85#_c_675_n 0.00603381f $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_225 N_B2_M1004_g N_A_311_85#_c_675_n 0.00647806f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_226 N_B2_M1004_g N_A_311_85#_c_663_n 0.00866507f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_227 N_B2_M1000_g N_A_311_85#_c_669_n 0.00221614f $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_228 N_B2_M1004_g N_A_311_85#_c_669_n 0.00221614f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_229 N_B2_M1000_g N_VGND_c_741_n 8.82278e-19 $X=2.345 $Y=0.795 $X2=0 $Y2=0
cc_230 N_B2_M1004_g N_VGND_c_741_n 8.82278e-19 $X=2.775 $Y=0.795 $X2=0 $Y2=0
cc_231 N_A1_M1003_g N_A2_M1001_g 0.0242339f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_232 N_A1_M1006_g N_A2_M1005_g 0.0413385f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A1_c_285_n N_A2_M1005_g 0.00453755f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_234 N_A1_c_309_p N_A2_M1005_g 0.0158698f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_235 N_A1_M1015_g N_A2_M1007_g 0.0243267f $X=5.205 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A1_c_309_p N_A2_M1007_g 0.0204393f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_237 N_A1_c_288_n N_A2_M1007_g 2.62404e-19 $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A1_M1019_g N_A2_M1011_g 0.0286785f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_239 N_A1_c_285_n N_A2_c_372_n 0.0176717f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A1_c_286_n N_A2_c_372_n 9.97094e-19 $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A1_c_309_p N_A2_c_372_n 0.0217013f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_242 N_A1_c_287_n N_A2_c_372_n 3.27266e-19 $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_243 N_A1_c_288_n N_A2_c_372_n 0.027167f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A1_c_285_n N_A2_c_373_n 0.00147358f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_245 N_A1_c_286_n N_A2_c_373_n 0.0184457f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A1_c_309_p N_A2_c_373_n 4.89879e-19 $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_247 N_A1_c_287_n N_A2_c_373_n 0.0243267f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A1_c_288_n N_A2_c_373_n 0.00963203f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A1_c_285_n N_VPWR_M1010_s 0.00112423f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_250 N_A1_c_304_n N_VPWR_M1010_s 0.0019198f $X=3.975 $Y=2.035 $X2=0 $Y2=0
cc_251 N_A1_c_288_n N_VPWR_M1015_s 0.00517975f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_252 N_A1_M1006_g N_VPWR_c_425_n 0.00150765f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A1_M1015_g N_VPWR_c_427_n 0.00341401f $X=5.205 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A1_c_287_n N_VPWR_c_427_n 3.71773e-19 $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_255 N_A1_c_288_n N_VPWR_c_427_n 0.0254574f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A1_M1006_g N_VPWR_c_430_n 0.00518311f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A1_M1015_g N_VPWR_c_430_n 0.00517089f $X=5.205 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A1_M1006_g N_VPWR_c_422_n 0.0098206f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A1_M1015_g N_VPWR_c_422_n 0.00980819f $X=5.205 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A1_c_309_p N_Y_M1005_d 0.00314031f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_261 N_A1_M1006_g N_Y_c_506_n 0.0167741f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A1_c_286_n N_Y_c_506_n 3.13234e-19 $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_263 N_A1_c_309_p N_Y_c_506_n 0.0378628f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_264 N_A1_c_304_n N_Y_c_506_n 0.0165507f $X=3.975 $Y=2.035 $X2=0 $Y2=0
cc_265 N_A1_M1006_g N_Y_c_525_n 7.49979e-19 $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_266 N_A1_c_285_n N_A_779_368#_M1006_d 0.00144296f $X=3.81 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A1_c_309_p N_A_779_368#_M1006_d 0.00888372f $X=4.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A1_c_304_n N_A_779_368#_M1006_d 2.44056e-19 $X=3.975 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A1_c_309_p N_A_779_368#_M1007_s 0.00153059f $X=4.925 $Y=2.035 $X2=0
+ $Y2=0
cc_270 N_A1_c_288_n N_A_779_368#_M1007_s 0.0033177f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_271 N_A1_M1015_g N_A_779_368#_c_581_n 0.00345561f $X=5.205 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A1_M1015_g N_A_779_368#_c_589_n 0.00761488f $X=5.205 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A1_c_309_p N_A_779_368#_c_589_n 0.00403821f $X=4.925 $Y=2.035 $X2=0
+ $Y2=0
cc_274 N_A1_c_288_n N_A_779_368#_c_589_n 0.0143139f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_275 N_A1_M1006_g N_A_779_368#_c_582_n 0.00687709f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A1_M1003_g N_A_311_85#_c_663_n 0.00322639f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_277 N_A1_M1003_g N_A_311_85#_c_686_n 0.0083539f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_278 N_A1_M1003_g N_A_311_85#_c_664_n 0.0116199f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_279 N_A1_c_285_n N_A_311_85#_c_664_n 0.0205962f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_280 N_A1_c_286_n N_A_311_85#_c_664_n 9.74228e-19 $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_281 N_A1_M1003_g N_A_311_85#_c_665_n 8.73939e-19 $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_282 N_A1_c_285_n N_A_311_85#_c_665_n 0.0055933f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_283 N_A1_c_286_n N_A_311_85#_c_665_n 3.08675e-19 $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_284 N_A1_M1019_g N_A_311_85#_c_666_n 9.38284e-19 $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_285 N_A1_M1019_g N_A_311_85#_c_667_n 0.012834f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_286 N_A1_c_287_n N_A_311_85#_c_667_n 0.00130772f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_287 N_A1_c_288_n N_A_311_85#_c_667_n 0.0599533f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_288 N_A1_M1019_g N_A_311_85#_c_668_n 0.0014977f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_289 N_A1_M1003_g N_VGND_c_739_n 0.00335812f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_290 N_A1_M1019_g N_VGND_c_740_n 0.0121211f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_291 N_A1_M1003_g N_VGND_c_741_n 0.00462669f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_292 N_A1_M1019_g N_VGND_c_743_n 0.00447026f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_293 N_A1_M1003_g N_VGND_c_744_n 0.00440294f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_294 N_A1_M1019_g N_VGND_c_744_n 0.00443817f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_295 N_A2_M1005_g N_VPWR_c_430_n 0.00333926f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A2_M1007_g N_VPWR_c_430_n 0.00333896f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A2_M1005_g N_VPWR_c_422_n 0.00423254f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A2_M1007_g N_VPWR_c_422_n 0.00422796f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A2_M1005_g N_Y_c_506_n 0.0111468f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A2_M1005_g N_Y_c_525_n 0.00511267f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_301 N_A2_M1005_g N_A_779_368#_c_581_n 0.0100424f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_302 N_A2_M1007_g N_A_779_368#_c_581_n 0.0135118f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A2_M1005_g N_A_779_368#_c_589_n 6.69226e-19 $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A2_M1007_g N_A_779_368#_c_589_n 0.00904087f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A2_M1005_g N_A_779_368#_c_582_n 4.1224e-19 $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A2_M1001_g N_A_311_85#_c_686_n 6.11774e-19 $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_307 N_A2_M1001_g N_A_311_85#_c_664_n 0.0176612f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_308 N_A2_c_372_n N_A_311_85#_c_664_n 0.00251202f $X=4.51 $Y=1.515 $X2=0 $Y2=0
cc_309 N_A2_M1001_g N_A_311_85#_c_666_n 4.62671e-19 $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_310 N_A2_M1011_g N_A_311_85#_c_666_n 0.00846178f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_311 N_A2_M1011_g N_A_311_85#_c_667_n 0.0162625f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_312 N_A2_M1011_g N_A_311_85#_c_670_n 0.0011955f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_313 N_A2_c_372_n N_A_311_85#_c_670_n 0.025376f $X=4.51 $Y=1.515 $X2=0 $Y2=0
cc_314 N_A2_c_373_n N_A_311_85#_c_670_n 0.00118154f $X=4.77 $Y=1.515 $X2=0 $Y2=0
cc_315 N_A2_M1001_g N_VGND_c_739_n 0.00231397f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_316 N_A2_M1011_g N_VGND_c_740_n 0.0039639f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_317 N_A2_M1001_g N_VGND_c_742_n 0.00537957f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_318 N_A2_M1011_g N_VGND_c_742_n 0.00523995f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_319 N_A2_M1001_g N_VGND_c_744_n 0.00528353f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_320 N_A2_M1011_g N_VGND_c_744_n 0.00528353f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_321 N_VPWR_M1010_s N_Y_c_506_n 0.0120673f $X=3.345 $Y=1.84 $X2=0 $Y2=0
cc_322 N_VPWR_c_425_n N_Y_c_506_n 0.0206651f $X=3.53 $Y=2.805 $X2=0 $Y2=0
cc_323 N_VPWR_M1014_s N_Y_c_496_n 0.0134696f $X=1.085 $Y=1.84 $X2=0 $Y2=0
cc_324 N_VPWR_c_431_n N_Y_c_496_n 0.044148f $X=1.58 $Y=2.795 $X2=0 $Y2=0
cc_325 N_VPWR_c_424_n Y 0.0170624f $X=0.32 $Y=2.115 $X2=0 $Y2=0
cc_326 N_VPWR_c_428_n Y 0.0109793f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_431_n Y 0.0134355f $X=1.58 $Y=2.795 $X2=0 $Y2=0
cc_328 N_VPWR_c_422_n Y 0.00901959f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_329 N_VPWR_c_429_n N_A_379_368#_c_553_n 0.0421123f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_422_n N_A_379_368#_c_553_n 0.0235523f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_429_n N_A_379_368#_c_554_n 0.0226835f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_431_n N_A_379_368#_c_554_n 0.0219393f $X=1.58 $Y=2.795 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_422_n N_A_379_368#_c_554_n 0.0124822f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_425_n N_A_379_368#_c_555_n 0.0214403f $X=3.53 $Y=2.805 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_429_n N_A_379_368#_c_555_n 0.0226835f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_422_n N_A_379_368#_c_555_n 0.0124822f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_427_n N_A_779_368#_c_581_n 0.0119238f $X=5.48 $Y=2.455 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_430_n N_A_779_368#_c_581_n 0.0623983f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_422_n N_A_779_368#_c_581_n 0.0343606f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_425_n N_A_779_368#_c_582_n 0.0214403f $X=3.53 $Y=2.805 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_430_n N_A_779_368#_c_582_n 0.0226835f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_422_n N_A_779_368#_c_582_n 0.0124822f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_343 N_Y_c_496_n N_A_379_368#_M1008_d 0.00405858f $X=2.365 $Y=2.512 $X2=-0.19
+ $Y2=-0.245
cc_344 N_Y_c_506_n N_A_379_368#_M1009_s 0.00434519f $X=4.365 $Y=2.375 $X2=0
+ $Y2=0
cc_345 N_Y_M1002_d N_A_379_368#_c_553_n 0.00182219f $X=2.38 $Y=1.84 $X2=0 $Y2=0
cc_346 N_Y_c_506_n N_A_379_368#_c_553_n 0.0046334f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_347 N_Y_c_496_n N_A_379_368#_c_553_n 0.00509985f $X=2.365 $Y=2.512 $X2=0
+ $Y2=0
cc_348 N_Y_c_512_n N_A_379_368#_c_553_n 0.0156189f $X=2.695 $Y=2.512 $X2=0 $Y2=0
cc_349 N_Y_c_496_n N_A_379_368#_c_554_n 0.0171102f $X=2.365 $Y=2.512 $X2=0 $Y2=0
cc_350 N_Y_c_506_n N_A_379_368#_c_555_n 0.0182896f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_351 N_Y_c_506_n N_A_779_368#_M1006_d 0.00435429f $X=4.365 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_352 N_Y_M1005_d N_A_779_368#_c_581_n 0.00165831f $X=4.395 $Y=1.84 $X2=0 $Y2=0
cc_353 N_Y_c_506_n N_A_779_368#_c_581_n 0.0046334f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_354 N_Y_c_525_n N_A_779_368#_c_581_n 0.0134956f $X=4.49 $Y=2.46 $X2=0 $Y2=0
cc_355 N_Y_c_506_n N_A_779_368#_c_582_n 0.0182896f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_356 Y N_A_27_74#_c_609_n 0.00119776f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_357 N_Y_M1017_d N_A_27_74#_c_610_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_358 Y N_A_27_74#_c_610_n 0.0143448f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_359 Y N_A_27_74#_c_614_n 0.00902371f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_613_n N_A_311_85#_M1012_s 0.00343588f $X=2.045 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_361 N_A_27_74#_c_615_n N_A_311_85#_M1000_d 0.00184993f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_c_612_n N_A_311_85#_c_660_n 0.0260161f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_613_n N_A_311_85#_c_660_n 0.0198855f $X=2.045 $Y=1.095 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_613_n N_A_311_85#_c_661_n 0.00390898f $X=2.045 $Y=1.095
+ $X2=0 $Y2=0
cc_365 N_A_27_74#_c_649_p N_A_311_85#_c_661_n 0.0127861f $X=2.13 $Y=0.885 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_615_n N_A_311_85#_c_661_n 0.00390898f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_367 N_A_27_74#_c_610_n N_A_311_85#_c_662_n 0.0128665f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_615_n N_A_311_85#_c_675_n 0.0154602f $X=2.895 $Y=1.095 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_615_n N_A_311_85#_c_663_n 0.00376163f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_370 N_A_27_74#_c_634_n N_A_311_85#_c_663_n 0.0265061f $X=3.085 $Y=0.68 $X2=0
+ $Y2=0
cc_371 N_A_27_74#_c_615_n N_A_311_85#_c_665_n 0.00749835f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_c_610_n N_VGND_c_741_n 0.0614387f $X=1.055 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_611_n N_VGND_c_741_n 0.0179217f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_610_n N_VGND_c_744_n 0.0342887f $X=1.055 $Y=0.34 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_611_n N_VGND_c_744_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_376 N_A_311_85#_c_664_n N_VGND_M1003_d 0.00313482f $X=4.38 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_377 N_A_311_85#_c_667_n N_VGND_M1011_s 0.00251857f $X=5.39 $Y=1.095 $X2=0
+ $Y2=0
cc_378 N_A_311_85#_c_663_n N_VGND_c_739_n 0.0144041f $X=3.46 $Y=0.34 $X2=0 $Y2=0
cc_379 N_A_311_85#_c_664_n N_VGND_c_739_n 0.0199169f $X=4.38 $Y=1.095 $X2=0
+ $Y2=0
cc_380 N_A_311_85#_c_666_n N_VGND_c_739_n 0.00158095f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_381 N_A_311_85#_c_666_n N_VGND_c_740_n 0.0163623f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_382 N_A_311_85#_c_667_n N_VGND_c_740_n 0.0185548f $X=5.39 $Y=1.095 $X2=0
+ $Y2=0
cc_383 N_A_311_85#_c_668_n N_VGND_c_740_n 0.0156043f $X=5.475 $Y=0.57 $X2=0
+ $Y2=0
cc_384 N_A_311_85#_c_661_n N_VGND_c_741_n 0.0340834f $X=2.395 $Y=0.34 $X2=0
+ $Y2=0
cc_385 N_A_311_85#_c_662_n N_VGND_c_741_n 0.0233304f $X=1.865 $Y=0.34 $X2=0
+ $Y2=0
cc_386 N_A_311_85#_c_663_n N_VGND_c_741_n 0.0652108f $X=3.46 $Y=0.34 $X2=0 $Y2=0
cc_387 N_A_311_85#_c_669_n N_VGND_c_741_n 0.0233304f $X=2.56 $Y=0.34 $X2=0 $Y2=0
cc_388 N_A_311_85#_c_666_n N_VGND_c_742_n 0.0119397f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_389 N_A_311_85#_c_668_n N_VGND_c_743_n 0.0092394f $X=5.475 $Y=0.57 $X2=0
+ $Y2=0
cc_390 N_A_311_85#_c_661_n N_VGND_c_744_n 0.0199188f $X=2.395 $Y=0.34 $X2=0
+ $Y2=0
cc_391 N_A_311_85#_c_662_n N_VGND_c_744_n 0.0127683f $X=1.865 $Y=0.34 $X2=0
+ $Y2=0
cc_392 N_A_311_85#_c_663_n N_VGND_c_744_n 0.0373458f $X=3.46 $Y=0.34 $X2=0 $Y2=0
cc_393 N_A_311_85#_c_666_n N_VGND_c_744_n 0.0116912f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_394 N_A_311_85#_c_668_n N_VGND_c_744_n 0.0090278f $X=5.475 $Y=0.57 $X2=0
+ $Y2=0
cc_395 N_A_311_85#_c_669_n N_VGND_c_744_n 0.0127683f $X=2.56 $Y=0.34 $X2=0 $Y2=0

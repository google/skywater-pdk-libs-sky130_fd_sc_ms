* File: sky130_fd_sc_ms__nor2b_2.pxi.spice
* Created: Fri Aug 28 17:47:30 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2B_2%B_N N_B_N_M1004_g N_B_N_M1005_g B_N N_B_N_c_63_n
+ PM_SKY130_FD_SC_MS__NOR2B_2%B_N
x_PM_SKY130_FD_SC_MS__NOR2B_2%A_27_392# N_A_27_392#_M1005_s N_A_27_392#_M1004_s
+ N_A_27_392#_c_93_n N_A_27_392#_M1003_g N_A_27_392#_c_102_n N_A_27_392#_M1000_g
+ N_A_27_392#_c_94_n N_A_27_392#_M1006_g N_A_27_392#_M1009_g N_A_27_392#_c_96_n
+ N_A_27_392#_c_97_n N_A_27_392#_c_98_n N_A_27_392#_c_99_n N_A_27_392#_c_100_n
+ N_A_27_392#_c_101_n PM_SKY130_FD_SC_MS__NOR2B_2%A_27_392#
x_PM_SKY130_FD_SC_MS__NOR2B_2%A N_A_M1007_g N_A_M1001_g N_A_M1008_g N_A_M1002_g
+ A A N_A_c_175_n PM_SKY130_FD_SC_MS__NOR2B_2%A
x_PM_SKY130_FD_SC_MS__NOR2B_2%VPWR N_VPWR_M1004_d N_VPWR_M1001_d N_VPWR_c_225_n
+ N_VPWR_c_226_n VPWR N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_224_n N_VPWR_c_231_n N_VPWR_c_232_n PM_SKY130_FD_SC_MS__NOR2B_2%VPWR
x_PM_SKY130_FD_SC_MS__NOR2B_2%A_228_368# N_A_228_368#_M1000_d
+ N_A_228_368#_M1009_d N_A_228_368#_M1002_s N_A_228_368#_c_265_n
+ N_A_228_368#_c_266_n N_A_228_368#_c_267_n N_A_228_368#_c_280_n
+ N_A_228_368#_c_281_n N_A_228_368#_c_288_n N_A_228_368#_c_268_n
+ N_A_228_368#_c_269_n PM_SKY130_FD_SC_MS__NOR2B_2%A_228_368#
x_PM_SKY130_FD_SC_MS__NOR2B_2%Y N_Y_M1003_d N_Y_M1007_d N_Y_M1000_s N_Y_c_310_n
+ N_Y_c_311_n N_Y_c_312_n N_Y_c_313_n N_Y_c_314_n N_Y_c_315_n N_Y_c_316_n Y
+ N_Y_c_317_n PM_SKY130_FD_SC_MS__NOR2B_2%Y
x_PM_SKY130_FD_SC_MS__NOR2B_2%VGND N_VGND_M1005_d N_VGND_M1006_s N_VGND_M1008_s
+ N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n VGND
+ N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n
+ N_VGND_c_370_n PM_SKY130_FD_SC_MS__NOR2B_2%VGND
cc_1 VNB N_B_N_M1005_g 0.0367247f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.79
cc_2 VNB B_N 0.00207353f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_B_N_c_63_n 0.0284219f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.635
cc_4 VNB N_A_27_392#_c_93_n 0.018486f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.79
cc_5 VNB N_A_27_392#_c_94_n 0.016567f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.635
cc_6 VNB N_A_27_392#_M1009_g 0.00232647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_392#_c_96_n 0.0432843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_392#_c_97_n 0.0192881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_392#_c_98_n 0.0121892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_392#_c_99_n 0.0145497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_100_n 0.00587637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_392#_c_101_n 0.0724696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1007_g 0.023477f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_14 VNB N_A_M1008_g 0.0269184f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.635
cc_15 VNB A 0.00224035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_c_175_n 0.0445892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_224_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_310_n 0.00280126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_311_n 5.19053e-19 $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.635
cc_20 VNB N_Y_c_312_n 0.00135442f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.635
cc_21 VNB N_Y_c_313_n 0.00392956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_314_n 0.00252696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_315_n 0.00292043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_316_n 0.00186002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_317_n 0.0212378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_361_n 0.0127511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_362_n 0.00277973f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.635
cc_28 VNB N_VGND_c_363_n 0.0120457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_364_n 0.0279043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_365_n 0.0292002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_366_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_367_n 0.0167762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_368_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_369_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_370_n 0.210833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B_N_M1004_g 0.029246f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.46
cc_37 VPB B_N 0.00249009f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_38 VPB N_B_N_c_63_n 0.0237944f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.635
cc_39 VPB N_A_27_392#_c_102_n 0.0194019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_392#_M1009_g 0.0211437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_392#_c_97_n 0.0558534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_392#_c_101_n 0.00825727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_M1001_g 0.0202484f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=0.79
cc_44 VPB N_A_M1002_g 0.028529f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.635
cc_45 VPB A 0.00596021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_c_175_n 0.00615722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_225_n 0.0152809f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_48 VPB N_VPWR_c_226_n 0.00522117f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.635
cc_49 VPB N_VPWR_c_227_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_228_n 0.0407783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_229_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_224_n 0.0706674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_231_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_232_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_228_368#_c_265_n 0.0129601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_228_368#_c_266_n 0.00388794f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.635
cc_57 VPB N_A_228_368#_c_267_n 0.00413156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_228_368#_c_268_n 0.0159566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_228_368#_c_269_n 0.0341141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_Y_c_312_n 0.00318572f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=1.635
cc_61 N_B_N_M1005_g N_A_27_392#_c_93_n 0.0171333f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_62 N_B_N_c_63_n N_A_27_392#_c_102_n 0.00107404f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_63 N_B_N_M1005_g N_A_27_392#_c_96_n 0.0106849f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_64 N_B_N_M1005_g N_A_27_392#_c_97_n 0.00477364f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_65 B_N N_A_27_392#_c_97_n 0.025547f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_N_c_63_n N_A_27_392#_c_97_n 0.016455f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_67 N_B_N_M1005_g N_A_27_392#_c_98_n 0.0118985f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_68 B_N N_A_27_392#_c_98_n 0.00563709f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B_N_M1005_g N_A_27_392#_c_99_n 0.00476166f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_70 B_N N_A_27_392#_c_99_n 0.0209889f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_71 N_B_N_c_63_n N_A_27_392#_c_99_n 0.00762197f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_72 N_B_N_M1005_g N_A_27_392#_c_100_n 0.00158684f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_73 B_N N_A_27_392#_c_100_n 0.00397231f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B_N_M1005_g N_A_27_392#_c_101_n 0.0191582f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_75 B_N N_A_27_392#_c_101_n 0.00151118f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_76 N_B_N_c_63_n N_A_27_392#_c_101_n 0.00667987f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_77 N_B_N_M1004_g N_VPWR_c_225_n 0.020999f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_78 B_N N_VPWR_c_225_n 0.0220408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_79 N_B_N_c_63_n N_VPWR_c_225_n 0.00297012f $X=0.83 $Y=1.635 $X2=0 $Y2=0
cc_80 N_B_N_M1004_g N_VPWR_c_227_n 0.00460063f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_81 N_B_N_M1004_g N_VPWR_c_224_n 0.00912278f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_82 N_B_N_M1004_g N_A_228_368#_c_265_n 0.00377212f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_83 N_B_N_M1004_g N_A_228_368#_c_267_n 6.08298e-19 $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_84 N_B_N_M1005_g N_VGND_c_361_n 0.0080577f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_85 N_B_N_M1005_g N_VGND_c_365_n 0.00485498f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_86 N_B_N_M1005_g N_VGND_c_370_n 0.00514438f $X=0.83 $Y=0.79 $X2=0 $Y2=0
cc_87 N_A_27_392#_c_94_n N_A_M1007_g 0.0239839f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_88 N_A_27_392#_c_101_n N_A_M1007_g 0.0131574f $X=1.915 $Y=1.49 $X2=0 $Y2=0
cc_89 N_A_27_392#_M1009_g N_A_M1001_g 0.0143437f $X=1.96 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_27_392#_M1009_g A 0.00371905f $X=1.96 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_27_392#_c_101_n A 0.00723344f $X=1.915 $Y=1.49 $X2=0 $Y2=0
cc_92 N_A_27_392#_M1009_g N_A_c_175_n 0.0131574f $X=1.96 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A_27_392#_c_102_n N_VPWR_c_225_n 0.00263089f $X=1.51 $Y=1.76 $X2=0 $Y2=0
cc_94 N_A_27_392#_c_97_n N_VPWR_c_225_n 0.0339508f $X=0.275 $Y=2.105 $X2=0 $Y2=0
cc_95 N_A_27_392#_c_98_n N_VPWR_c_225_n 8.30447e-19 $X=1.145 $Y=1.215 $X2=0
+ $Y2=0
cc_96 N_A_27_392#_c_97_n N_VPWR_c_227_n 0.011066f $X=0.275 $Y=2.105 $X2=0 $Y2=0
cc_97 N_A_27_392#_c_102_n N_VPWR_c_228_n 0.00333896f $X=1.51 $Y=1.76 $X2=0 $Y2=0
cc_98 N_A_27_392#_M1009_g N_VPWR_c_228_n 0.00333896f $X=1.96 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_27_392#_c_102_n N_VPWR_c_224_n 0.00427818f $X=1.51 $Y=1.76 $X2=0 $Y2=0
cc_100 N_A_27_392#_M1009_g N_VPWR_c_224_n 0.00422796f $X=1.96 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_27_392#_c_97_n N_VPWR_c_224_n 0.00915947f $X=0.275 $Y=2.105 $X2=0
+ $Y2=0
cc_102 N_A_27_392#_c_102_n N_A_228_368#_c_265_n 0.0159301f $X=1.51 $Y=1.76 $X2=0
+ $Y2=0
cc_103 N_A_27_392#_M1009_g N_A_228_368#_c_265_n 7.14937e-19 $X=1.96 $Y=2.4 $X2=0
+ $Y2=0
cc_104 N_A_27_392#_c_98_n N_A_228_368#_c_265_n 9.32104e-19 $X=1.145 $Y=1.215
+ $X2=0 $Y2=0
cc_105 N_A_27_392#_c_100_n N_A_228_368#_c_265_n 0.0183181f $X=1.31 $Y=1.215
+ $X2=0 $Y2=0
cc_106 N_A_27_392#_c_101_n N_A_228_368#_c_265_n 0.0035845f $X=1.915 $Y=1.49
+ $X2=0 $Y2=0
cc_107 N_A_27_392#_c_102_n N_A_228_368#_c_266_n 0.0116345f $X=1.51 $Y=1.76 $X2=0
+ $Y2=0
cc_108 N_A_27_392#_M1009_g N_A_228_368#_c_266_n 0.0135505f $X=1.96 $Y=2.4 $X2=0
+ $Y2=0
cc_109 N_A_27_392#_c_102_n N_A_228_368#_c_267_n 0.00291744f $X=1.51 $Y=1.76
+ $X2=0 $Y2=0
cc_110 N_A_27_392#_M1009_g N_A_228_368#_c_280_n 0.00332448f $X=1.96 $Y=2.4 $X2=0
+ $Y2=0
cc_111 N_A_27_392#_c_102_n N_A_228_368#_c_281_n 6.26485e-19 $X=1.51 $Y=1.76
+ $X2=0 $Y2=0
cc_112 N_A_27_392#_M1009_g N_A_228_368#_c_281_n 0.0106426f $X=1.96 $Y=2.4 $X2=0
+ $Y2=0
cc_113 N_A_27_392#_c_93_n N_Y_c_310_n 0.00505604f $X=1.435 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A_27_392#_c_93_n N_Y_c_311_n 0.00778619f $X=1.435 $Y=1.22 $X2=0 $Y2=0
cc_115 N_A_27_392#_c_100_n N_Y_c_311_n 0.00421645f $X=1.31 $Y=1.215 $X2=0 $Y2=0
cc_116 N_A_27_392#_c_101_n N_Y_c_311_n 0.00194033f $X=1.915 $Y=1.49 $X2=0 $Y2=0
cc_117 N_A_27_392#_c_93_n N_Y_c_312_n 2.53709e-19 $X=1.435 $Y=1.22 $X2=0 $Y2=0
cc_118 N_A_27_392#_c_94_n N_Y_c_312_n 0.00100575f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_119 N_A_27_392#_M1009_g N_Y_c_312_n 0.00362743f $X=1.96 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_27_392#_c_100_n N_Y_c_312_n 0.0265536f $X=1.31 $Y=1.215 $X2=0 $Y2=0
cc_121 N_A_27_392#_c_101_n N_Y_c_312_n 0.0302586f $X=1.915 $Y=1.49 $X2=0 $Y2=0
cc_122 N_A_27_392#_c_94_n N_Y_c_313_n 0.0200565f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A_27_392#_c_101_n N_Y_c_313_n 0.00285281f $X=1.915 $Y=1.49 $X2=0 $Y2=0
cc_124 N_A_27_392#_c_93_n N_VGND_c_361_n 0.00714781f $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_125 N_A_27_392#_c_96_n N_VGND_c_361_n 0.036192f $X=0.615 $Y=0.615 $X2=0 $Y2=0
cc_126 N_A_27_392#_c_98_n N_VGND_c_361_n 0.0131477f $X=1.145 $Y=1.215 $X2=0
+ $Y2=0
cc_127 N_A_27_392#_c_100_n N_VGND_c_361_n 0.0143981f $X=1.31 $Y=1.215 $X2=0
+ $Y2=0
cc_128 N_A_27_392#_c_101_n N_VGND_c_361_n 0.00102906f $X=1.915 $Y=1.49 $X2=0
+ $Y2=0
cc_129 N_A_27_392#_c_93_n N_VGND_c_362_n 4.45911e-19 $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_130 N_A_27_392#_c_94_n N_VGND_c_362_n 0.00825039f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_131 N_A_27_392#_c_96_n N_VGND_c_365_n 0.0211421f $X=0.615 $Y=0.615 $X2=0
+ $Y2=0
cc_132 N_A_27_392#_c_93_n N_VGND_c_366_n 0.00434272f $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_133 N_A_27_392#_c_94_n N_VGND_c_366_n 0.00444681f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_134 N_A_27_392#_c_93_n N_VGND_c_370_n 0.00825538f $X=1.435 $Y=1.22 $X2=0
+ $Y2=0
cc_135 N_A_27_392#_c_94_n N_VGND_c_370_n 0.00877997f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_136 N_A_27_392#_c_96_n N_VGND_c_370_n 0.0231103f $X=0.615 $Y=0.615 $X2=0
+ $Y2=0
cc_137 N_A_M1001_g N_VPWR_c_226_n 0.00126302f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_M1002_g N_VPWR_c_226_n 0.0153844f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_M1001_g N_VPWR_c_228_n 0.00517089f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_M1002_g N_VPWR_c_229_n 0.00460063f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VPWR_c_224_n 0.00977588f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_VPWR_c_224_n 0.00912278f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_A_228_368#_c_266_n 0.00347836f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_A_228_368#_c_280_n 8.84614e-19 $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_145 A N_A_228_368#_c_280_n 0.0215149f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A_M1001_g N_A_228_368#_c_281_n 0.010841f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_M1002_g N_A_228_368#_c_281_n 4.47651e-19 $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_M1001_g N_A_228_368#_c_288_n 0.012931f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_M1002_g N_A_228_368#_c_288_n 0.0196406f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_150 A N_A_228_368#_c_288_n 0.0276263f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A_c_175_n N_A_228_368#_c_288_n 4.90767e-19 $X=2.845 $Y=1.515 $X2=0
+ $Y2=0
cc_152 N_A_M1002_g N_A_228_368#_c_268_n 8.13654e-19 $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_A_228_368#_c_269_n 0.00147311f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_M1007_g N_Y_c_312_n 5.38267e-19 $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_155 A N_Y_c_312_n 0.0267892f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A_M1007_g N_Y_c_313_n 0.0147681f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_157 A N_Y_c_313_n 0.0356018f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_M1007_g N_Y_c_314_n 4.49298e-19 $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_M1008_g N_Y_c_314_n 4.7485e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_M1008_g N_Y_c_315_n 0.0188325f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_161 A N_Y_c_315_n 7.29585e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A_c_175_n N_Y_c_315_n 0.0010611f $X=2.845 $Y=1.515 $X2=0 $Y2=0
cc_163 A N_Y_c_316_n 0.0214748f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A_c_175_n N_Y_c_316_n 0.003731f $X=2.845 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A_M1008_g N_Y_c_317_n 0.00964993f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_166 A N_Y_c_317_n 0.00361538f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A_M1007_g N_VGND_c_362_n 0.00982302f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_M1008_g N_VGND_c_362_n 4.5319e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_M1007_g N_VGND_c_364_n 4.40885e-19 $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_M1008_g N_VGND_c_364_n 0.0111523f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_M1007_g N_VGND_c_367_n 0.00383152f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_M1008_g N_VGND_c_367_n 0.00444681f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_M1007_g N_VGND_c_370_n 0.00758019f $X=2.365 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_M1008_g N_VGND_c_370_n 0.00877997f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_175 N_VPWR_c_225_n N_A_228_368#_c_265_n 0.0630024f $X=0.725 $Y=2.135 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_226_n N_A_228_368#_c_266_n 0.0103534f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_228_n N_A_228_368#_c_266_n 0.0592384f $X=2.55 $Y=3.33 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_224_n N_A_228_368#_c_266_n 0.0326137f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_225_n N_A_228_368#_c_267_n 0.0121616f $X=0.725 $Y=2.135 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_228_n N_A_228_368#_c_267_n 0.0235512f $X=2.55 $Y=3.33 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_224_n N_A_228_368#_c_267_n 0.0126924f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_182 N_VPWR_M1001_d N_A_228_368#_c_288_n 0.00314376f $X=2.5 $Y=1.84 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_226_n N_A_228_368#_c_288_n 0.0148589f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_226_n N_A_228_368#_c_269_n 0.0224614f $X=2.635 $Y=2.455 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_229_n N_A_228_368#_c_269_n 0.011066f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_224_n N_A_228_368#_c_269_n 0.00915947f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_187 N_A_228_368#_c_266_n N_Y_M1000_s 0.00165831f $X=2.02 $Y=2.99 $X2=0 $Y2=0
cc_188 N_A_228_368#_c_265_n N_Y_c_312_n 0.0314126f $X=1.285 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_228_368#_c_266_n N_Y_c_312_n 0.0118736f $X=2.02 $Y=2.99 $X2=0 $Y2=0
cc_190 N_A_228_368#_c_268_n N_Y_c_317_n 0.0111281f $X=3.125 $Y=2.12 $X2=0 $Y2=0
cc_191 N_Y_c_313_n N_VGND_M1006_s 0.001993f $X=2.495 $Y=1.07 $X2=0 $Y2=0
cc_192 N_Y_c_315_n N_VGND_M1008_s 5.90379e-19 $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_193 N_Y_c_317_n N_VGND_M1008_s 0.0033108f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_194 N_Y_c_310_n N_VGND_c_361_n 0.0174504f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_195 N_Y_c_310_n N_VGND_c_362_n 0.0173003f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_196 N_Y_c_313_n N_VGND_c_362_n 0.0174872f $X=2.495 $Y=1.07 $X2=0 $Y2=0
cc_197 N_Y_c_314_n N_VGND_c_362_n 0.0164981f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_198 N_Y_c_314_n N_VGND_c_364_n 0.0191439f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_199 N_Y_c_315_n N_VGND_c_364_n 0.00254062f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_200 N_Y_c_317_n N_VGND_c_364_n 0.0198092f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_201 N_Y_c_310_n N_VGND_c_366_n 0.0145091f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_202 N_Y_c_314_n N_VGND_c_367_n 0.011066f $X=2.58 $Y=0.515 $X2=0 $Y2=0
cc_203 N_Y_c_310_n N_VGND_c_370_n 0.0119768f $X=1.65 $Y=0.515 $X2=0 $Y2=0
cc_204 N_Y_c_314_n N_VGND_c_370_n 0.00915947f $X=2.58 $Y=0.515 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__sedfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1549_74# a_1351_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=2.80005e+12p ps=2.337e+07u
M1001 a_1747_118# a_1351_74# a_697_113# VNB nlowvt w=420000u l=150000u
+  ad=2.478e+11p pd=2.02e+06u as=3.885e+11p ps=4.37e+06u
M1002 a_1895_118# a_1549_74# a_1747_118# VNB nlowvt w=420000u l=150000u
+  ad=1.617e+11p pd=1.61e+06u as=0p ps=0u
M1003 a_575_305# a_2463_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1004 Q_N a_575_305# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.2449e+12p ps=1.863e+07u
M1005 VPWR DE a_161_394# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 a_27_90# a_575_305# a_533_113# VNB nlowvt w=420000u l=150000u
+  ad=3.276e+11p pd=3.24e+06u as=1.008e+11p ps=1.32e+06u
M1007 a_2650_508# a_1549_74# a_2463_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=3.115e+11p ps=2.71e+06u
M1008 a_1071_462# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1009 a_1934_508# a_1351_74# a_1747_118# VPB pshort w=420000u l=180000u
+  ad=1.05e+11p pd=1.34e+06u as=1.344e+11p ps=1.48e+06u
M1010 a_1747_118# a_1549_74# a_697_113# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=4.823e+11p ps=5.11e+06u
M1011 a_1549_74# a_1351_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_119_464# D a_27_90# VPB pshort w=640000u l=180000u
+  ad=1.344e+11p pd=1.7e+06u as=3.52e+11p ps=3.66e+06u
M1013 VPWR a_1972_92# a_1934_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q_N a_575_305# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 VPWR a_2463_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1016 a_1351_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1017 a_533_113# a_161_394# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_697_113# SCE a_1075_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 VGND DE a_161_394# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1020 VPWR a_575_305# a_2650_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_157_90# D a_27_90# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 VGND DE a_157_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1351_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 a_2391_74# a_1972_92# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1025 a_2463_74# a_1549_74# a_2391_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1026 a_559_464# DE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1027 VGND a_1972_92# a_1895_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1075_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_161_394# a_119_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_90# a_575_305# a_559_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_575_305# a_2463_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1032 a_697_113# a_667_87# a_1071_462# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_697_113# a_667_87# a_27_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2463_74# a_1351_74# a_2348_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.95e+11p ps=3.59e+06u
M1035 a_1972_92# a_1747_118# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1036 a_2565_74# a_1351_74# a_2463_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1037 VGND a_575_305# a_2565_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR SCE a_667_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.208e+11p ps=1.97e+06u
M1039 a_697_113# SCE a_27_90# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1972_92# a_1747_118# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1041 VGND a_2463_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1042 VGND SCE a_667_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1043 a_2348_392# a_1972_92# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


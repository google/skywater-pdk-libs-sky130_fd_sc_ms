* File: sky130_fd_sc_ms__a21o_1.pex.spice
* Created: Fri Aug 28 16:59:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21O_1%A_81_264# 1 2 9 11 13 15 16 25 27 31 33 35 36
+ 40
c65 36 0 1.84796e-19 $X=1.425 $Y=1.95
c66 11 0 8.11701e-20 $X=1.13 $Y=1.47
r67 35 36 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.115
+ $X2=1.425 $Y2=1.95
r68 29 31 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.97 $Y=1.11
+ $X2=1.97 $Y2=0.805
r69 28 33 3.70735 $w=2.5e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.415 $Y=1.195
+ $X2=1.33 $Y2=1.38
r70 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.805 $Y=1.195
+ $X2=1.97 $Y2=1.11
r71 27 28 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.805 $Y=1.195
+ $X2=1.415 $Y2=1.195
r72 23 35 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.425 $Y=2.13
+ $X2=1.425 $Y2=2.115
r73 23 25 21.9284 $w=3.58e-07 $l=6.85e-07 $layer=LI1_cond $X=1.425 $Y=2.13
+ $X2=1.425 $Y2=2.815
r74 21 33 2.76166 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.33 $Y=1.65 $X2=1.33
+ $Y2=1.38
r75 21 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.33 $Y=1.65 $X2=1.33
+ $Y2=1.95
r76 19 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.485
+ $X2=0.755 $Y2=1.485
r77 19 37 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.59 $Y=1.485
+ $X2=0.495 $Y2=1.485
r78 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.485 $X2=0.59 $Y2=1.485
r79 16 33 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.245 $Y=1.485
+ $X2=1.33 $Y2=1.38
r80 16 18 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.245 $Y=1.485
+ $X2=0.59 $Y2=1.485
r81 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.205 $Y=1.395
+ $X2=1.205 $Y2=0.95
r82 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.13 $Y=1.47
+ $X2=1.205 $Y2=1.395
r83 11 40 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.13 $Y=1.47
+ $X2=0.755 $Y2=1.47
r84 7 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.65
+ $X2=0.495 $Y2=1.485
r85 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.495 $Y=1.65
+ $X2=0.495 $Y2=2.4
r86 2 35 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.115
r87 2 25 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.815
r88 1 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.83
+ $Y=0.68 $X2=1.97 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%B1 3 7 9 12
c35 9 0 8.11701e-20 $X=1.68 $Y=1.665
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.615
+ $X2=1.67 $Y2=1.78
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.615
+ $X2=1.67 $Y2=1.45
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.615 $X2=1.67 $Y2=1.615
r39 7 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.755 $Y=1 $X2=1.755
+ $Y2=1.45
r40 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.745 $Y=2.46
+ $X2=1.745 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%A1 3 7 9 12
c37 3 0 4.71918e-20 $X=2.195 $Y=2.46
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.615
+ $X2=2.21 $Y2=1.78
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.615
+ $X2=2.21 $Y2=1.45
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.615 $X2=2.21 $Y2=1.615
r41 7 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.185 $Y=1 $X2=2.185
+ $Y2=1.45
r42 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.195 $Y=2.46
+ $X2=2.195 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%A2 4 5 7 13 15 22
r34 15 22 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=0.462
+ $X2=3.005 $Y2=0.462
r35 13 17 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.81 $Y=0.405
+ $X2=2.66 $Y2=0.405
r36 12 22 7.13417 $w=3.13e-07 $l=1.95e-07 $layer=LI1_cond $X=2.81 $Y=0.412
+ $X2=3.005 $Y2=0.412
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=0.405 $X2=2.81 $Y2=0.405
r38 5 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.675 $Y=1.485 $X2=2.675
+ $Y2=1.395
r39 5 7 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=2.675 $Y=1.485
+ $X2=2.675 $Y2=2.46
r40 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.66 $Y=1 $X2=2.66
+ $Y2=1.395
r41 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=0.57
+ $X2=2.66 $Y2=0.405
r42 1 4 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.66 $Y=0.57 $X2=2.66
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%X 1 2 9 10 13 15 16 17 24 33
r20 22 24 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.26 $Y=1.995 $X2=0.26
+ $Y2=2.035
r21 16 17 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r22 15 22 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.995
r23 15 33 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.82
r24 15 16 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.405
r25 15 24 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.035
r26 11 13 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.95 $Y=0.98
+ $X2=0.95 $Y2=0.885
r27 9 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.825 $Y=1.065
+ $X2=0.95 $Y2=0.98
r28 9 10 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.825 $Y=1.065
+ $X2=0.255 $Y2=1.065
r29 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.15
+ $X2=0.255 $Y2=1.065
r30 7 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.15 $X2=0.17
+ $Y2=1.82
r31 2 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r32 2 17 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r33 1 13 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=0.865
+ $Y=0.58 $X2=0.99 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r37 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r43 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 27 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.76 $Y2=3.33
r45 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 22 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.76 $Y2=3.33
r49 22 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 18 32 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 18 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.335 $Y=3.33 $X2=2.435
+ $Y2=3.33
r54 17 35 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 17 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.535 $Y=3.33 $X2=2.435
+ $Y2=3.33
r56 13 19 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=3.33
r57 13 15 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=2.435 $Y=3.245
+ $X2=2.435 $Y2=2.455
r58 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.76 $Y=1.985
+ $X2=0.76 $Y2=2.815
r59 7 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r60 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=2.815
r61 2 15 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=2.285
+ $Y=1.96 $X2=2.435 $Y2=2.455
r62 1 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.815
r63 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%A_367_392# 1 2 7 9 11 13 15
c33 13 0 4.71918e-20 $X=2.9 $Y=2.12
r34 13 20 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.9 $Y=2.12 $X2=2.9
+ $Y2=2.03
r35 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.9 $Y=2.12 $X2=2.9
+ $Y2=2.815
r36 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=2.035
+ $X2=1.97 $Y2=2.035
r37 11 20 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.735 $Y=2.035
+ $X2=2.9 $Y2=2.03
r38 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.735 $Y=2.035
+ $X2=2.135 $Y2=2.035
r39 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=2.12 $X2=1.97
+ $Y2=2.035
r40 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.97 $Y=2.12 $X2=1.97
+ $Y2=2.815
r41 2 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.96 $X2=2.9 $Y2=2.105
r42 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.96 $X2=2.9 $Y2=2.815
r43 1 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.96 $X2=1.97 $Y2=2.115
r44 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.96 $X2=1.97 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_1%VGND 1 2 9 12 13 14 16 17 19 20 21 26 39 40
r52 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r54 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r55 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r57 29 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r58 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r60 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r61 21 24 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0.925
+ $X2=2.875 $Y2=1.09
r62 19 36 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.16
+ $Y2=0
r63 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.39
+ $Y2=0
r64 18 39 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=3.12
+ $Y2=0
r65 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.39
+ $Y2=0
r66 16 33 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r67 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.42
+ $Y2=0
r68 15 36 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=2.16
+ $Y2=0
r69 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.42
+ $Y2=0
r70 13 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.925
+ $X2=2.875 $Y2=0.925
r71 13 14 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.71 $Y=0.925
+ $X2=2.475 $Y2=0.925
r72 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.39 $Y=0.84
+ $X2=2.475 $Y2=0.925
r73 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0
r74 11 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0.84
r75 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=0.085 $X2=1.42
+ $Y2=0
r76 7 9 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.42 $Y=0.085 $X2=1.42
+ $Y2=0.775
r77 2 24 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.68 $X2=2.875 $Y2=1.09
r78 1 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.58 $X2=1.42 $Y2=0.775
.ends


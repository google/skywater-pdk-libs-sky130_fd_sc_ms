* File: sky130_fd_sc_ms__o41a_2.pxi.spice
* Created: Wed Sep  2 12:26:57 2020
* 
x_PM_SKY130_FD_SC_MS__O41A_2%A1 N_A1_M1002_g N_A1_M1011_g A1 N_A1_c_79_n
+ N_A1_c_80_n PM_SKY130_FD_SC_MS__O41A_2%A1
x_PM_SKY130_FD_SC_MS__O41A_2%A2 N_A2_M1005_g N_A2_M1013_g N_A2_c_108_n
+ N_A2_c_109_n A2 A2 A2 PM_SKY130_FD_SC_MS__O41A_2%A2
x_PM_SKY130_FD_SC_MS__O41A_2%A3 N_A3_M1008_g N_A3_M1003_g A3 A3 A3 A3
+ N_A3_c_151_n PM_SKY130_FD_SC_MS__O41A_2%A3
x_PM_SKY130_FD_SC_MS__O41A_2%A4 N_A4_M1006_g N_A4_M1000_g A4 N_A4_c_191_n
+ N_A4_c_192_n PM_SKY130_FD_SC_MS__O41A_2%A4
x_PM_SKY130_FD_SC_MS__O41A_2%B1 N_B1_M1004_g N_B1_M1009_g B1 B1 N_B1_c_227_n
+ PM_SKY130_FD_SC_MS__O41A_2%B1
x_PM_SKY130_FD_SC_MS__O41A_2%A_431_368# N_A_431_368#_M1009_d
+ N_A_431_368#_M1006_d N_A_431_368#_M1001_g N_A_431_368#_M1010_g
+ N_A_431_368#_M1007_g N_A_431_368#_M1012_g N_A_431_368#_c_280_n
+ N_A_431_368#_c_278_n N_A_431_368#_c_288_n N_A_431_368#_c_270_n
+ N_A_431_368#_c_271_n N_A_431_368#_c_272_n N_A_431_368#_c_273_n
+ N_A_431_368#_c_274_n N_A_431_368#_c_275_n
+ PM_SKY130_FD_SC_MS__O41A_2%A_431_368#
x_PM_SKY130_FD_SC_MS__O41A_2%VPWR N_VPWR_M1002_s N_VPWR_M1004_d N_VPWR_M1012_s
+ N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n VPWR
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_347_n
+ PM_SKY130_FD_SC_MS__O41A_2%VPWR
x_PM_SKY130_FD_SC_MS__O41A_2%X N_X_M1001_d N_X_M1010_d N_X_c_400_n N_X_c_401_n
+ N_X_c_402_n X PM_SKY130_FD_SC_MS__O41A_2%X
x_PM_SKY130_FD_SC_MS__O41A_2%A_27_74# N_A_27_74#_M1011_s N_A_27_74#_M1013_d
+ N_A_27_74#_M1000_d N_A_27_74#_c_423_n N_A_27_74#_c_424_n N_A_27_74#_c_425_n
+ N_A_27_74#_c_426_n N_A_27_74#_c_427_n N_A_27_74#_c_428_n N_A_27_74#_c_429_n
+ PM_SKY130_FD_SC_MS__O41A_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O41A_2%VGND N_VGND_M1011_d N_VGND_M1003_d N_VGND_M1001_s
+ N_VGND_M1007_s N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n
+ N_VGND_c_480_n N_VGND_c_481_n VGND N_VGND_c_482_n N_VGND_c_483_n
+ N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n
+ PM_SKY130_FD_SC_MS__O41A_2%VGND
cc_1 VNB N_A1_M1011_g 0.0348798f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_c_79_n 0.027683f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_3 VNB N_A1_c_80_n 0.0155193f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_4 VNB N_A2_M1013_g 0.0257807f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_5 VNB N_A2_c_108_n 0.00167106f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_6 VNB N_A2_c_109_n 0.0269673f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_7 VNB N_A3_M1003_g 0.0273614f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB A3 0.00465445f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A3_c_151_n 0.022435f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.565
cc_10 VNB N_A4_M1000_g 0.0275785f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_A4_c_191_n 0.0269767f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_12 VNB N_A4_c_192_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_13 VNB N_B1_M1009_g 0.0281622f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_14 VNB B1 0.00953293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_227_n 0.0267841f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.35
cc_16 VNB N_A_431_368#_M1001_g 0.0224767f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_A_431_368#_M1010_g 0.00166497f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_18 VNB N_A_431_368#_M1007_g 0.0265448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_431_368#_M1012_g 0.00243112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_431_368#_c_270_n 0.0104431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_431_368#_c_271_n 0.01612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_431_368#_c_272_n 0.00406491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_431_368#_c_273_n 4.08426e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_431_368#_c_274_n 0.00840116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_431_368#_c_275_n 0.0874472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_347_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_400_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_X_c_401_n 0.00415351f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_29 VNB N_X_c_402_n 4.65031e-19 $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_30 VNB N_A_27_74#_c_423_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_31 VNB N_A_27_74#_c_424_n 0.00948616f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.35
cc_32 VNB N_A_27_74#_c_425_n 0.00995328f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.68
cc_33 VNB N_A_27_74#_c_426_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_427_n 0.0188114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_428_n 0.00253059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_429_n 0.0100545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_476_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.68
cc_38 VNB N_VGND_c_477_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_478_n 0.0109596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_479_n 0.0139769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_480_n 0.0131032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_481_n 0.0117082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_482_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_483_n 0.0339528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_484_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_485_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_486_n 0.00980973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_487_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_488_n 0.285003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_A1_M1002_g 0.0253535f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_51 VPB N_A1_c_79_n 0.00579252f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_52 VPB N_A1_c_80_n 0.00816907f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_53 VPB N_A2_M1005_g 0.0223905f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_54 VPB N_A2_c_108_n 0.00136305f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_55 VPB N_A2_c_109_n 0.00564997f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_56 VPB N_A3_M1008_g 0.023977f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_57 VPB A3 0.00180784f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_58 VPB N_A3_c_151_n 0.00542952f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.565
cc_59 VPB N_A4_M1006_g 0.0250429f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_60 VPB N_A4_c_191_n 0.00564765f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_61 VPB N_A4_c_192_n 0.00206052f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_62 VPB N_B1_M1004_g 0.0250641f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_63 VPB B1 0.00745351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B1_c_227_n 0.00579128f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.35
cc_65 VPB N_A_431_368#_M1010_g 0.0246498f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_66 VPB N_A_431_368#_M1012_g 0.0289588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_431_368#_c_278_n 0.00369941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_431_368#_c_273_n 0.00339407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_348_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_349_n 0.0487491f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_71 VPB N_VPWR_c_350_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_72 VPB N_VPWR_c_351_n 0.0648097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_352_n 0.0642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_353_n 0.0163631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_354_n 0.0362502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_347_n 0.0827108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_X_c_402_n 0.00504759f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_78 N_A1_M1002_g N_A2_M1005_g 0.0443527f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A1_M1011_g N_A2_M1013_g 0.0260254f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A1_M1002_g N_A2_c_108_n 0.00452759f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A1_c_79_n N_A2_c_108_n 5.47053e-19 $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A1_c_80_n N_A2_c_108_n 0.0250943f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A1_c_79_n N_A2_c_109_n 0.0443527f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A1_c_80_n N_A2_c_109_n 0.00153341f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A1_M1002_g N_VPWR_c_349_n 0.0222166f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A1_c_79_n N_VPWR_c_349_n 7.81657e-19 $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A1_c_80_n N_VPWR_c_349_n 0.0254126f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A1_M1002_g N_VPWR_c_352_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A1_M1002_g N_VPWR_c_347_n 0.00908371f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A1_M1011_g N_A_27_74#_c_423_n 0.0103339f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_91 N_A1_M1011_g N_A_27_74#_c_424_n 0.0117984f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A1_c_79_n N_A_27_74#_c_424_n 6.59012e-19 $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_93 N_A1_c_80_n N_A_27_74#_c_424_n 0.0110042f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A1_M1011_g N_A_27_74#_c_425_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A1_c_79_n N_A_27_74#_c_425_n 0.00363055f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A1_c_80_n N_A_27_74#_c_425_n 0.0279713f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A1_M1011_g N_A_27_74#_c_426_n 6.28869e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A1_M1011_g N_VGND_c_476_n 0.00622602f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A1_M1011_g N_VGND_c_482_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A1_M1011_g N_VGND_c_488_n 0.0082497f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A2_M1005_g N_A3_M1008_g 0.0386756f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A2_c_108_n N_A3_M1008_g 0.00212152f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_103 A2 N_A3_M1008_g 0.00977703f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A2_M1013_g N_A3_M1003_g 0.019972f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A2_M1005_g A3 8.9819e-19 $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A2_c_108_n A3 0.0286217f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A2_c_109_n A3 0.00120846f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_108 A2 A3 0.0562229f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_109 N_A2_c_108_n N_A3_c_151_n 4.19484e-19 $X=1 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A2_c_109_n N_A3_c_151_n 0.0176384f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A2_M1005_g N_VPWR_c_349_n 0.00345211f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_112 A2 N_VPWR_c_349_n 0.0371956f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A2_M1005_g N_VPWR_c_352_n 0.00365007f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_114 A2 N_VPWR_c_352_n 0.0139969f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_115 N_A2_M1005_g N_VPWR_c_347_n 0.00444515f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_116 A2 N_VPWR_c_347_n 0.0157743f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_117 N_A2_c_108_n A_203_368# 9.92688e-19 $X=1 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_118 A2 A_203_368# 0.0106665f $X=1.115 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_119 A2 A_203_368# 0.0153441f $X=1.115 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_120 N_A2_M1013_g N_A_27_74#_c_423_n 6.28869e-19 $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A2_M1013_g N_A_27_74#_c_424_n 0.0117933f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A2_c_108_n N_A_27_74#_c_424_n 0.0217949f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A2_c_109_n N_A_27_74#_c_424_n 0.00107112f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A2_M1013_g N_A_27_74#_c_426_n 0.00966073f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A2_M1013_g N_A_27_74#_c_429_n 0.0015571f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A2_c_108_n N_A_27_74#_c_429_n 0.00425598f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A2_M1013_g N_VGND_c_476_n 0.00484409f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A2_M1013_g N_VGND_c_477_n 0.00434272f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A2_M1013_g N_VGND_c_488_n 0.0082141f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A3_M1008_g N_A4_M1006_g 0.0385316f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_131 A3 N_A4_M1006_g 0.0128255f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_132 N_A3_M1003_g N_A4_M1000_g 0.018224f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_133 A3 N_A4_c_191_n 0.00201946f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A3_c_151_n N_A4_c_191_n 0.0174403f $X=1.57 $Y=1.515 $X2=0 $Y2=0
cc_135 A3 N_A4_c_192_n 0.032651f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A3_c_151_n N_A4_c_192_n 3.70595e-19 $X=1.57 $Y=1.515 $X2=0 $Y2=0
cc_137 A3 N_A_431_368#_c_280_n 0.0081741f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A3_M1008_g N_A_431_368#_c_278_n 0.00102986f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_139 A3 N_A_431_368#_c_278_n 0.0349219f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A3_M1008_g N_VPWR_c_352_n 0.00533722f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_141 A3 N_VPWR_c_352_n 0.00634296f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A3_M1008_g N_VPWR_c_347_n 0.0102393f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_143 A3 N_VPWR_c_347_n 0.00785491f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_144 A3 A_317_368# 0.0155623f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_145 N_A3_M1003_g N_A_27_74#_c_426_n 0.0145272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A3_M1003_g N_A_27_74#_c_427_n 0.0122944f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_147 A3 N_A_27_74#_c_427_n 0.0260507f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A3_c_151_n N_A_27_74#_c_427_n 0.00375849f $X=1.57 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A3_M1003_g N_A_27_74#_c_429_n 0.00155819f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_150 A3 N_A_27_74#_c_429_n 0.00326062f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A3_c_151_n N_A_27_74#_c_429_n 4.08598e-19 $X=1.57 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A3_M1003_g N_VGND_c_477_n 0.00434272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A3_M1003_g N_VGND_c_478_n 0.00586574f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A3_M1003_g N_VGND_c_488_n 0.00822442f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A4_M1006_g N_B1_M1004_g 0.0208492f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A4_c_192_n N_B1_M1004_g 3.76336e-19 $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_157 N_A4_M1000_g N_B1_M1009_g 0.0193383f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A4_M1006_g B1 3.27214e-19 $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A4_c_191_n B1 0.00218973f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A4_c_192_n B1 0.0302881f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A4_c_191_n N_B1_c_227_n 0.0175566f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A4_c_192_n N_B1_c_227_n 4.04657e-19 $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A4_M1006_g N_A_431_368#_c_280_n 0.00299512f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A4_c_191_n N_A_431_368#_c_280_n 7.63688e-19 $X=2.14 $Y=1.515 $X2=0
+ $Y2=0
cc_165 N_A4_c_192_n N_A_431_368#_c_280_n 0.0130747f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_166 N_A4_M1006_g N_A_431_368#_c_278_n 0.0140998f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A4_M1006_g N_VPWR_c_352_n 0.005209f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A4_M1006_g N_VPWR_c_354_n 0.00329175f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A4_M1006_g N_VPWR_c_347_n 0.00989635f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A4_M1000_g N_A_27_74#_c_427_n 0.0145711f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A4_c_191_n N_A_27_74#_c_427_n 0.001245f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A4_c_192_n N_A_27_74#_c_427_n 0.0247664f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A4_M1000_g N_A_27_74#_c_428_n 0.013702f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A4_M1000_g N_VGND_c_478_n 0.00757529f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A4_M1000_g N_VGND_c_483_n 0.00451267f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A4_M1000_g N_VGND_c_488_n 0.00877274f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B1_M1004_g N_A_431_368#_c_278_n 0.0111422f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_178 N_B1_M1004_g N_A_431_368#_c_288_n 0.018987f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_179 B1 N_A_431_368#_c_288_n 0.0525521f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_180 N_B1_c_227_n N_A_431_368#_c_288_n 7.13232e-19 $X=2.71 $Y=1.515 $X2=0
+ $Y2=0
cc_181 N_B1_M1009_g N_A_431_368#_c_270_n 0.00161219f $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_182 B1 N_A_431_368#_c_271_n 0.00887071f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_183 N_B1_M1009_g N_A_431_368#_c_272_n 0.00162779f $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_184 B1 N_A_431_368#_c_272_n 0.0294134f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_185 N_B1_c_227_n N_A_431_368#_c_272_n 0.00186365f $X=2.71 $Y=1.515 $X2=0
+ $Y2=0
cc_186 N_B1_M1004_g N_A_431_368#_c_273_n 0.00408407f $X=2.635 $Y=2.34 $X2=0
+ $Y2=0
cc_187 B1 N_A_431_368#_c_273_n 0.0271533f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B1_c_227_n N_A_431_368#_c_273_n 3.02201e-19 $X=2.71 $Y=1.515 $X2=0
+ $Y2=0
cc_189 N_B1_M1009_g N_A_431_368#_c_274_n 0.00273312f $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_190 B1 N_A_431_368#_c_274_n 0.00969568f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_191 N_B1_M1009_g N_A_431_368#_c_275_n 6.21883e-19 $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_192 B1 N_A_431_368#_c_275_n 0.00239357f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B1_c_227_n N_A_431_368#_c_275_n 0.00488449f $X=2.71 $Y=1.515 $X2=0
+ $Y2=0
cc_194 N_B1_M1004_g N_VPWR_c_352_n 0.0049405f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_195 N_B1_M1004_g N_VPWR_c_354_n 0.0130481f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_196 N_B1_M1004_g N_VPWR_c_347_n 0.00511769f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_197 N_B1_M1009_g N_A_27_74#_c_427_n 0.00302367f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_198 B1 N_A_27_74#_c_427_n 0.00856196f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_199 N_B1_c_227_n N_A_27_74#_c_427_n 0.00149819f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_200 N_B1_M1009_g N_A_27_74#_c_428_n 0.0082268f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B1_M1009_g N_VGND_c_479_n 0.00327253f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B1_M1009_g N_VGND_c_483_n 0.00434272f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B1_M1009_g N_VGND_c_488_n 0.00826504f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_431_368#_c_288_n N_VPWR_M1004_d 0.0282656f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_205 N_A_431_368#_c_273_n N_VPWR_M1004_d 0.00386963f $X=3.57 $Y=1.95 $X2=0
+ $Y2=0
cc_206 N_A_431_368#_M1010_g N_VPWR_c_351_n 6.90496e-19 $X=3.845 $Y=2.4 $X2=0
+ $Y2=0
cc_207 N_A_431_368#_M1012_g N_VPWR_c_351_n 0.0218366f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_208 N_A_431_368#_c_278_n N_VPWR_c_352_n 0.014549f $X=2.29 $Y=2.815 $X2=0
+ $Y2=0
cc_209 N_A_431_368#_M1010_g N_VPWR_c_353_n 0.00476846f $X=3.845 $Y=2.4 $X2=0
+ $Y2=0
cc_210 N_A_431_368#_M1012_g N_VPWR_c_353_n 0.00460063f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_431_368#_M1010_g N_VPWR_c_354_n 0.0155907f $X=3.845 $Y=2.4 $X2=0
+ $Y2=0
cc_212 N_A_431_368#_M1012_g N_VPWR_c_354_n 5.00985e-19 $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_213 N_A_431_368#_c_278_n N_VPWR_c_354_n 0.0436844f $X=2.29 $Y=2.815 $X2=0
+ $Y2=0
cc_214 N_A_431_368#_c_288_n N_VPWR_c_354_n 0.0791892f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_215 N_A_431_368#_c_275_n N_VPWR_c_354_n 9.44791e-19 $X=4.235 $Y=1.465 $X2=0
+ $Y2=0
cc_216 N_A_431_368#_M1010_g N_VPWR_c_347_n 0.00938661f $X=3.845 $Y=2.4 $X2=0
+ $Y2=0
cc_217 N_A_431_368#_M1012_g N_VPWR_c_347_n 0.00908554f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_218 N_A_431_368#_c_278_n N_VPWR_c_347_n 0.0119743f $X=2.29 $Y=2.815 $X2=0
+ $Y2=0
cc_219 N_A_431_368#_M1001_g N_X_c_400_n 0.0124354f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_431_368#_M1007_g N_X_c_400_n 0.00772833f $X=4.235 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_431_368#_M1001_g N_X_c_401_n 0.006795f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_431_368#_M1007_g N_X_c_401_n 0.0150748f $X=4.235 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_431_368#_c_274_n N_X_c_401_n 0.0214332f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_224 N_A_431_368#_c_275_n N_X_c_401_n 0.0131297f $X=4.235 $Y=1.465 $X2=0 $Y2=0
cc_225 N_A_431_368#_M1010_g N_X_c_402_n 0.002166f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A_431_368#_M1012_g N_X_c_402_n 0.00524799f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_431_368#_c_273_n N_X_c_402_n 0.024103f $X=3.57 $Y=1.95 $X2=0 $Y2=0
cc_228 N_A_431_368#_c_274_n N_X_c_402_n 0.0032852f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_229 N_A_431_368#_c_275_n N_X_c_402_n 0.0185823f $X=4.235 $Y=1.465 $X2=0 $Y2=0
cc_230 N_A_431_368#_c_272_n N_A_27_74#_c_427_n 0.0104256f $X=3.125 $Y=1.095
+ $X2=0 $Y2=0
cc_231 N_A_431_368#_c_270_n N_A_27_74#_c_428_n 0.0255177f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_232 N_A_431_368#_c_271_n N_VGND_M1001_s 4.82091e-19 $X=3.405 $Y=1.095 $X2=0
+ $Y2=0
cc_233 N_A_431_368#_c_274_n N_VGND_M1001_s 0.00397467f $X=3.57 $Y=1.465 $X2=0
+ $Y2=0
cc_234 N_A_431_368#_M1001_g N_VGND_c_479_n 0.00545191f $X=3.805 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_431_368#_c_270_n N_VGND_c_479_n 0.0316872f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_A_431_368#_c_271_n N_VGND_c_479_n 0.00369599f $X=3.405 $Y=1.095 $X2=0
+ $Y2=0
cc_237 N_A_431_368#_c_274_n N_VGND_c_479_n 0.0181094f $X=3.57 $Y=1.465 $X2=0
+ $Y2=0
cc_238 N_A_431_368#_c_275_n N_VGND_c_479_n 0.00141269f $X=4.235 $Y=1.465 $X2=0
+ $Y2=0
cc_239 N_A_431_368#_M1007_g N_VGND_c_481_n 0.00364571f $X=4.235 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_431_368#_c_275_n N_VGND_c_481_n 8.29358e-19 $X=4.235 $Y=1.465 $X2=0
+ $Y2=0
cc_241 N_A_431_368#_c_270_n N_VGND_c_483_n 0.0146357f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_242 N_A_431_368#_M1001_g N_VGND_c_484_n 0.00434272f $X=3.805 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_431_368#_M1007_g N_VGND_c_484_n 0.00434272f $X=4.235 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_431_368#_M1001_g N_VGND_c_488_n 0.00825059f $X=3.805 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_431_368#_M1007_g N_VGND_c_488_n 0.00823934f $X=4.235 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_431_368#_c_270_n N_VGND_c_488_n 0.0121141f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_351_n N_X_c_402_n 0.0395285f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_248 N_VPWR_c_353_n N_X_c_402_n 0.00905805f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_249 N_VPWR_c_354_n N_X_c_402_n 0.0296638f $X=3.215 $Y=2.375 $X2=0 $Y2=0
cc_250 N_VPWR_c_347_n N_X_c_402_n 0.00749747f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_251 N_X_c_400_n N_VGND_c_479_n 0.018426f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_252 N_X_c_400_n N_VGND_c_481_n 0.0238012f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_253 N_X_c_400_n N_VGND_c_484_n 0.0144922f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_254 N_X_c_400_n N_VGND_c_488_n 0.0118826f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_255 N_A_27_74#_c_424_n N_VGND_M1011_d 0.00358162f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_256 N_A_27_74#_c_427_n N_VGND_M1003_d 0.00654166f $X=2.295 $Y=1.095 $X2=0
+ $Y2=0
cc_257 N_A_27_74#_c_423_n N_VGND_c_476_n 0.0191765f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_258 N_A_27_74#_c_424_n N_VGND_c_476_n 0.0248957f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_259 N_A_27_74#_c_426_n N_VGND_c_476_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_260 N_A_27_74#_c_426_n N_VGND_c_477_n 0.0144922f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_261 N_A_27_74#_c_426_n N_VGND_c_478_n 0.0182921f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_262 N_A_27_74#_c_427_n N_VGND_c_478_n 0.0345921f $X=2.295 $Y=1.095 $X2=0
+ $Y2=0
cc_263 N_A_27_74#_c_428_n N_VGND_c_478_n 0.0182921f $X=2.46 $Y=0.515 $X2=0 $Y2=0
cc_264 N_A_27_74#_c_423_n N_VGND_c_482_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_428_n N_VGND_c_483_n 0.014537f $X=2.46 $Y=0.515 $X2=0 $Y2=0
cc_266 N_A_27_74#_c_423_n N_VGND_c_488_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_267 N_A_27_74#_c_426_n N_VGND_c_488_n 0.0118826f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_268 N_A_27_74#_c_428_n N_VGND_c_488_n 0.011955f $X=2.46 $Y=0.515 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VPWR a_492_48# a_1200_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VPWR a_28_74# a_259_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 a_608_74# a_492_48# a_28_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 a_1598_400# CIN VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_28_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_2004_136# a_430_418# a_1857_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_1200_368# a_430_418# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_28_74# B a_608_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_1857_368# a_608_74# a_2004_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VPWR CIN a_1857_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_608_74# a_492_48# a_259_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VPWR a_2004_136# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_430_418# a_492_48# a_259_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X13 VGND a_28_74# a_259_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_430_418# a_492_48# a_28_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_28_74# B a_430_418# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X16 a_1967_384# a_1857_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_1200_368# a_608_74# COUT VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X18 VGND a_2004_136# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 COUT a_430_418# a_1598_400# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X20 VGND a_492_48# a_1200_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 a_1598_400# CIN VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 a_492_48# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 a_1967_384# a_608_74# a_2004_136# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X24 a_1967_384# a_1857_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X25 a_2004_136# a_430_418# a_1967_384# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 a_28_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_492_48# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 COUT a_608_74# a_1598_400# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 a_259_368# B a_608_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X30 a_259_368# B a_430_418# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 VGND CIN a_1857_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4_1 A B C D VGND VNB VPB VPWR X
X0 VPWR A a_96_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X1 a_335_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_96_74# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 VPWR C a_96_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X4 a_96_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 a_257_74# C a_335_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR a_96_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_179_74# B a_257_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_96_74# A a_179_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VGND a_96_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

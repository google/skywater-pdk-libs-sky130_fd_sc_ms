* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvn_1 A TE_B VGND VNB VPB VPWR Z
M1000 a_281_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=3.616e+11p ps=2.95e+06u
M1001 Z A a_281_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_281_100# a_22_46# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.564e+11p ps=2.36e+06u
M1003 Z A a_281_100# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 VPWR TE_B a_22_46# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1005 VGND TE_B a_22_46# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
.ends

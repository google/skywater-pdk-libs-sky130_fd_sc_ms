* File: sky130_fd_sc_ms__sdfxbp_2.pex.spice
* Created: Wed Sep  2 12:31:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_36_74# 1 2 9 13 15 17 20 23 24 25 29 37
+ 40 41
c92 40 0 2.15575e-19 $X=2.03 $Y=1.89
c93 37 0 1.99756e-19 $X=0.83 $Y=1.635
r94 41 49 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.89
+ $X2=2.03 $Y2=2.055
r95 40 43 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=1.89
+ $X2=2.03 $Y2=2.055
r96 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.89 $X2=2.03 $Y2=1.89
r97 35 37 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.75 $Y=1.635 $X2=0.83
+ $Y2=1.635
r98 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.635 $X2=0.75 $Y2=1.635
r99 26 29 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.17 $Y=0.54
+ $X2=0.325 $Y2=0.54
r100 24 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=2.055
+ $X2=2.03 $Y2=2.055
r101 24 25 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.865 $Y=2.055
+ $X2=0.915 $Y2=2.055
r102 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.83 $Y=1.97
+ $X2=0.915 $Y2=2.055
r103 22 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=1.8
+ $X2=0.83 $Y2=1.635
r104 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.83 $Y=1.8
+ $X2=0.83 $Y2=1.97
r105 18 35 15.6453 $w=3.28e-07 $l=4.48e-07 $layer=LI1_cond $X=0.302 $Y=1.635
+ $X2=0.75 $Y2=1.635
r106 18 31 4.60977 $w=3.28e-07 $l=1.32e-07 $layer=LI1_cond $X=0.302 $Y=1.635
+ $X2=0.17 $Y2=1.635
r107 18 20 16.1607 $w=4.33e-07 $l=6.1e-07 $layer=LI1_cond $X=0.302 $Y=1.8
+ $X2=0.302 $Y2=2.41
r108 17 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.47
+ $X2=0.17 $Y2=1.635
r109 16 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=0.54
r110 16 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=1.47
r111 15 36 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.635
+ $X2=0.75 $Y2=1.635
r112 13 49 206.016 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=2.04 $Y=2.585
+ $X2=2.04 $Y2=2.055
r113 7 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.04 $Y=1.47
+ $X2=0.965 $Y2=1.635
r114 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.04 $Y=1.47 $X2=1.04
+ $Y2=0.58
r115 2 20 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.21
+ $Y=2.265 $X2=0.355 $Y2=2.41
r116 1 29 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.37 $X2=0.325 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%SCE 2 3 4 5 7 8 10 11 13 15 16 18 19 20 24
+ 26 30 38
r76 32 34 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.27 $Y=1.065
+ $X2=0.54 $Y2=1.065
r77 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.065 $X2=1.91 $Y2=1.065
r78 26 30 6.311 $w=4.18e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=1.02 $X2=1.91
+ $Y2=1.02
r79 26 38 3.71646 $w=4.18e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.02
+ $X2=1.565 $Y2=1.02
r80 24 34 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.59 $Y=1.065 $X2=0.54
+ $Y2=1.065
r81 23 38 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=0.59 $Y=1.065
+ $X2=1.565 $Y2=1.065
r82 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.065 $X2=0.59 $Y2=1.065
r83 20 29 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.1 $Y=1.065
+ $X2=1.91 $Y2=1.065
r84 16 20 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.175 $Y=0.9
+ $X2=2.1 $Y2=1.065
r85 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.175 $Y=0.9
+ $X2=2.175 $Y2=0.58
r86 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.19
+ $X2=1.115 $Y2=2.585
r87 12 19 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.755 $Y=2.115
+ $X2=0.665 $Y2=2.115
r88 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.025 $Y=2.115
+ $X2=1.115 $Y2=2.19
r89 11 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.025 $Y=2.115
+ $X2=0.755 $Y2=2.115
r90 8 19 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=2.19
+ $X2=0.665 $Y2=2.115
r91 8 10 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.665 $Y=2.19
+ $X2=0.665 $Y2=2.585
r92 5 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.9 $X2=0.54
+ $Y2=1.065
r93 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.9 $X2=0.54
+ $Y2=0.58
r94 3 19 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.575 $Y=2.115
+ $X2=0.665 $Y2=2.115
r95 3 4 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.575 $Y=2.115
+ $X2=0.345 $Y2=2.115
r96 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.27 $Y=2.04
+ $X2=0.345 $Y2=2.115
r97 1 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.23
+ $X2=0.27 $Y2=1.065
r98 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.23 $X2=0.27
+ $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%D 3 7 9 12 13
c38 12 0 2.93225e-19 $X=1.49 $Y=1.635
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.635
+ $X2=1.49 $Y2=1.8
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.635
+ $X2=1.49 $Y2=1.47
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.635 $X2=1.49 $Y2=1.635
r42 9 13 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.635 $X2=1.49
+ $Y2=1.635
r43 7 15 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=1.535 $Y=2.585
+ $X2=1.535 $Y2=1.8
r44 3 14 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.43 $Y=0.58 $X2=1.43
+ $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%SCD 3 7 9 12 13
c40 12 0 6.78066e-20 $X=2.57 $Y=1.94
c41 7 0 1.30658e-19 $X=2.565 $Y=0.58
c42 3 0 1.22106e-19 $X=2.525 $Y=2.585
r43 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.94
+ $X2=2.57 $Y2=2.105
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.94
+ $X2=2.57 $Y2=1.775
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.94 $X2=2.57 $Y2=1.94
r46 9 13 3.12806 $w=3.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=2.035
+ $X2=2.58 $Y2=1.94
r47 7 14 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=2.565 $Y=0.58
+ $X2=2.565 $Y2=1.775
r48 3 15 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2.525 $Y=2.585
+ $X2=2.525 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%CLK 3 7 9 12
c38 9 0 1.30658e-19 $X=3.6 $Y=1.665
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.515 $X2=3.43 $Y2=1.515
r40 12 14 32.8636 $w=2.86e-07 $l=1.95e-07 $layer=POLY_cond $X=3.235 $Y=1.515
+ $X2=3.43 $Y2=1.515
r41 9 15 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.43
+ $Y2=1.565
r42 5 12 13.6159 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.68
+ $X2=3.235 $Y2=1.515
r43 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.235 $Y=1.68
+ $X2=3.235 $Y2=2.4
r44 1 12 26.965 $w=2.86e-07 $l=2.31571e-07 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.235 $Y2=1.515
r45 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.075 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_828_74# 1 2 9 13 15 17 20 24 25 28 30 31
+ 33 34 37 38 41 42 43 46 53 54 55 58 60 61 62 65 69
c194 65 0 1.41735e-19 $X=8.515 $Y=1.31
c195 61 0 8.50626e-20 $X=7.615 $Y=1.195
c196 53 0 5.59789e-20 $X=5.17 $Y=2.17
c197 33 0 1.21466e-19 $X=5.155 $Y=2.005
c198 13 0 1.1997e-19 $X=5.79 $Y=0.695
r199 69 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.515 $Y=1.39
+ $X2=8.515 $Y2=1.555
r200 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.515
+ $Y=1.39 $X2=8.515 $Y2=1.39
r201 65 68 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.515 $Y=1.31
+ $X2=8.515 $Y2=1.39
r202 61 76 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.615 $Y=1.195
+ $X2=7.48 $Y2=1.195
r203 60 63 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=7.65 $Y=1.195
+ $X2=7.65 $Y2=1.31
r204 60 62 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=1.195
+ $X2=7.65 $Y2=1.03
r205 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.615
+ $Y=1.195 $X2=7.615 $Y2=1.195
r206 58 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.21
+ $X2=5.84 $Y2=1.045
r207 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.21 $X2=5.84 $Y2=1.21
r208 55 57 16.8521 $w=2.57e-07 $l=3.55e-07 $layer=LI1_cond $X=5.915 $Y=0.855
+ $X2=5.915 $Y2=1.21
r209 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.17
+ $Y=2.17 $X2=5.17 $Y2=2.17
r210 47 63 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.78 $Y=1.31
+ $X2=7.65 $Y2=1.31
r211 46 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=1.31
+ $X2=8.515 $Y2=1.31
r212 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.35 $Y=1.31
+ $X2=7.78 $Y2=1.31
r213 44 62 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.605 $Y=0.425
+ $X2=7.605 $Y2=1.03
r214 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.52 $Y=0.34
+ $X2=7.605 $Y2=0.425
r215 42 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.52 $Y=0.34
+ $X2=7.01 $Y2=0.34
r216 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.925 $Y=0.425
+ $X2=7.01 $Y2=0.34
r217 40 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.925 $Y=0.425
+ $X2=6.925 $Y2=0.77
r218 39 55 3.1561 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0.855
+ $X2=5.915 $Y2=0.855
r219 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.84 $Y=0.855
+ $X2=6.925 $Y2=0.77
r220 38 39 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.84 $Y=0.855
+ $X2=6.08 $Y2=0.855
r221 37 55 5.43462 $w=2.57e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.995 $Y=0.77
+ $X2=5.915 $Y2=0.855
r222 36 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.995 $Y=0.425
+ $X2=5.995 $Y2=0.77
r223 35 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=0.34
+ $X2=5.155 $Y2=0.34
r224 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.91 $Y=0.34
+ $X2=5.995 $Y2=0.425
r225 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.91 $Y=0.34
+ $X2=5.24 $Y2=0.34
r226 33 52 0.582803 $w=3.14e-07 $l=1.5e-08 $layer=LI1_cond $X=5.155 $Y=2.072
+ $X2=5.17 $Y2=2.072
r227 33 49 18.0669 $w=3.14e-07 $l=4.65e-07 $layer=LI1_cond $X=5.155 $Y=2.072
+ $X2=4.69 $Y2=2.072
r228 32 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=0.34
r229 32 33 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=2.005
r230 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=5.155 $Y2=0.34
r231 30 31 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=4.445 $Y2=0.34
r232 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r233 26 28 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r234 24 25 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.395 $Y=1.99
+ $X2=8.395 $Y2=2.14
r235 24 82 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.425 $Y=1.99
+ $X2=8.425 $Y2=1.555
r236 20 25 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=8.38 $Y=2.75
+ $X2=8.38 $Y2=2.14
r237 15 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.48 $Y=1.03
+ $X2=7.48 $Y2=1.195
r238 15 17 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.48 $Y=1.03
+ $X2=7.48 $Y2=0.645
r239 13 74 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.79 $Y=0.695
+ $X2=5.79 $Y2=1.045
r240 7 53 57.4258 $w=2.56e-07 $l=3.78616e-07 $layer=POLY_cond $X=5.475 $Y=2.335
+ $X2=5.17 $Y2=2.17
r241 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.475 $Y=2.335
+ $X2=5.475 $Y2=2.705
r242 2 49 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=4.555
+ $Y=1.84 $X2=4.69 $Y2=2.01
r243 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_630_74# 1 2 9 11 13 15 16 20 22 28 32 35
+ 36 38 39 40 43 47 49 53 54 57 60 61 63 64 65 67 68 71 73 76 85 87
c200 73 0 5.59789e-20 $X=6.12 $Y=2.08
c201 43 0 3.61287e-20 $X=8.24 $Y=0.94
c202 40 0 1.21466e-19 $X=5.03 $Y=1.69
r203 77 87 20.917 $w=2.65e-07 $l=1.15e-07 $layer=POLY_cond $X=7.73 $Y=1.765
+ $X2=7.845 $Y2=1.765
r204 76 79 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=1.765
+ $X2=7.73 $Y2=1.93
r205 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.73
+ $Y=1.765 $X2=7.73 $Y2=1.765
r206 71 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.965 $Y=2.08
+ $X2=5.965 $Y2=2.245
r207 70 73 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.965 $Y=2.08
+ $X2=6.12 $Y2=2.08
r208 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.965
+ $Y=2.08 $X2=5.965 $Y2=2.08
r209 67 79 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=7.65 $Y=2.615
+ $X2=7.65 $Y2=1.93
r210 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.565 $Y=2.7
+ $X2=7.65 $Y2=2.615
r211 64 65 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.565 $Y=2.7
+ $X2=6.205 $Y2=2.7
r212 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.12 $Y=2.615
+ $X2=6.205 $Y2=2.7
r213 62 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.12 $Y=2.245
+ $X2=6.12 $Y2=2.08
r214 62 63 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.12 $Y=2.245
+ $X2=6.12 $Y2=2.615
r215 61 82 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.975 $Y=1.515
+ $X2=3.975 $Y2=1.69
r216 61 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.515
+ $X2=3.975 $Y2=1.35
r217 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.515 $X2=3.975 $Y2=1.515
r218 58 60 20.888 $w=2.38e-07 $l=4.35e-07 $layer=LI1_cond $X=3.975 $Y=1.95
+ $X2=3.975 $Y2=1.515
r219 57 68 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.975 $Y=1.47
+ $X2=3.975 $Y2=1.35
r220 57 60 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=3.975 $Y=1.47
+ $X2=3.975 $Y2=1.515
r221 55 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.94 $Y=1.18
+ $X2=3.94 $Y2=1.35
r222 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=1.095
+ $X2=3.94 $Y2=1.18
r223 53 54 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.855 $Y=1.095
+ $X2=3.455 $Y2=1.095
r224 49 58 6.82018 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=3.855 $Y=2.075
+ $X2=3.975 $Y2=1.95
r225 49 51 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=3.855 $Y=2.075
+ $X2=3.465 $Y2=2.075
r226 45 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.29 $Y=1.01
+ $X2=3.455 $Y2=1.095
r227 45 47 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.29 $Y=1.01
+ $X2=3.29 $Y2=0.515
r228 41 43 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=8.065 $Y=0.94
+ $X2=8.24 $Y2=0.94
r229 36 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.24 $Y=0.865
+ $X2=8.24 $Y2=0.94
r230 36 38 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.24 $Y=0.865
+ $X2=8.24 $Y2=0.58
r231 35 87 40.0151 $w=2.65e-07 $l=2.91033e-07 $layer=POLY_cond $X=8.065 $Y=1.6
+ $X2=7.845 $Y2=1.765
r232 34 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.065 $Y=1.015
+ $X2=8.065 $Y2=0.94
r233 34 35 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=8.065 $Y=1.015
+ $X2=8.065 $Y2=1.6
r234 30 87 11.8589 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.845 $Y=1.93
+ $X2=7.845 $Y2=1.765
r235 30 32 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=7.845 $Y=1.93
+ $X2=7.845 $Y2=2.54
r236 28 85 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=6.01 $Y=2.705
+ $X2=6.01 $Y2=2.245
r237 24 71 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.965 $Y=1.765
+ $X2=5.965 $Y2=2.08
r238 23 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.105 $Y=1.69
+ $X2=5.03 $Y2=1.69
r239 22 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.8 $Y=1.69
+ $X2=5.965 $Y2=1.765
r240 22 23 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.8 $Y=1.69
+ $X2=5.105 $Y2=1.69
r241 18 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.03 $Y=1.615
+ $X2=5.03 $Y2=1.69
r242 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=5.03 $Y=1.615
+ $X2=5.03 $Y2=0.695
r243 17 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.555 $Y=1.69
+ $X2=4.465 $Y2=1.69
r244 16 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.955 $Y=1.69
+ $X2=5.03 $Y2=1.69
r245 16 17 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.955 $Y=1.69
+ $X2=4.555 $Y2=1.69
r246 13 39 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.465 $Y=1.765
+ $X2=4.465 $Y2=1.69
r247 13 15 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=4.465 $Y=1.765
+ $X2=4.465 $Y2=2.4
r248 12 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.69
+ $X2=3.975 $Y2=1.69
r249 11 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.375 $Y=1.69
+ $X2=4.465 $Y2=1.69
r250 11 12 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=4.375 $Y=1.69
+ $X2=4.14 $Y2=1.69
r251 9 81 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.35
r252 2 51 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.84 $X2=3.465 $Y2=2.115
r253 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.37 $X2=3.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_1243_48# 1 2 9 13 15 18 22 27 28 30
c67 13 0 5.59221e-20 $X=6.43 $Y=2.705
c68 9 0 1.1651e-19 $X=6.29 $Y=0.58
r69 27 28 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=7.252 $Y=2.28
+ $X2=7.252 $Y2=2.115
r70 24 30 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.265 $Y=1.405
+ $X2=7.265 $Y2=1.257
r71 24 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.265 $Y=1.405
+ $X2=7.265 $Y2=2.115
r72 20 30 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.265 $Y=1.11
+ $X2=7.265 $Y2=1.257
r73 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.265 $Y=1.11
+ $X2=7.265 $Y2=0.765
r74 18 33 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.397 $Y=1.24
+ $X2=6.397 $Y2=1.405
r75 18 32 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.397 $Y=1.24
+ $X2=6.397 $Y2=1.075
r76 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.24 $X2=6.415 $Y2=1.24
r77 15 30 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=1.257
+ $X2=7.265 $Y2=1.257
r78 15 17 29.8854 $w=2.93e-07 $l=7.65e-07 $layer=LI1_cond $X=7.18 $Y=1.257
+ $X2=6.415 $Y2=1.257
r79 13 33 505.323 $w=1.8e-07 $l=1.3e-06 $layer=POLY_cond $X=6.43 $Y=2.705
+ $X2=6.43 $Y2=1.405
r80 9 32 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.29 $Y=0.58
+ $X2=6.29 $Y2=1.075
r81 2 27 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=2.12 $X2=7.29 $Y2=2.28
r82 1 22 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.37 $X2=7.265 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_1021_97# 1 2 9 13 16 19 22 25 27 28 30 34
c85 28 0 5.59221e-20 $X=5.685 $Y=2.475
c86 22 0 1.1651e-19 $X=5.575 $Y=0.695
r87 34 38 40.172 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=6.935 $Y=1.78
+ $X2=6.935 $Y2=1.945
r88 34 37 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=6.935 $Y=1.78
+ $X2=6.935 $Y2=1.615
r89 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.895
+ $Y=1.78 $X2=6.895 $Y2=1.78
r90 30 33 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=6.87 $Y=1.66
+ $X2=6.87 $Y2=1.78
r91 27 28 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.685 $Y=2.705
+ $X2=5.685 $Y2=2.475
r92 22 24 8.98601 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.575 $Y=0.695
+ $X2=5.575 $Y2=0.875
r93 20 25 1.34256 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.675 $Y=1.66
+ $X2=5.542 $Y2=1.66
r94 19 30 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.73 $Y=1.66 $X2=6.87
+ $Y2=1.66
r95 19 20 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=6.73 $Y=1.66
+ $X2=5.675 $Y2=1.66
r96 17 25 5.16603 $w=1.7e-07 $l=1.06325e-07 $layer=LI1_cond $X=5.59 $Y=1.745
+ $X2=5.542 $Y2=1.66
r97 17 28 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.59 $Y=1.745
+ $X2=5.59 $Y2=2.475
r98 16 25 5.16603 $w=1.7e-07 $l=1.05924e-07 $layer=LI1_cond $X=5.495 $Y=1.575
+ $X2=5.542 $Y2=1.66
r99 16 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.495 $Y=1.575
+ $X2=5.495 $Y2=0.875
r100 13 37 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.05 $Y=0.645
+ $X2=7.05 $Y2=1.615
r101 9 38 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=7.05 $Y=2.54
+ $X2=7.05 $Y2=1.945
r102 2 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.495 $X2=5.7 $Y2=2.705
r103 1 22 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.485 $X2=5.575 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_1711_48# 1 2 7 9 10 11 14 22 26 28 32 36
+ 38 42 46 48 49 50 53 57 60 62 65 66 69 73 74 76
c159 11 0 1.41735e-19 $X=8.705 $Y=0.94
r160 69 71 11.5626 $w=3.88e-07 $l=2.65e-07 $layer=LI1_cond $X=9.755 $Y=0.62
+ $X2=9.755 $Y2=0.885
r161 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.445
+ $Y=1.465 $X2=10.445 $Y2=1.465
r162 63 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.465
+ $X2=9.865 $Y2=1.465
r163 63 65 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.95 $Y=1.465
+ $X2=10.445 $Y2=1.465
r164 62 73 6.11814 $w=2.6e-07 $l=2.61151e-07 $layer=LI1_cond $X=9.865 $Y=1.94
+ $X2=9.775 $Y2=2.16
r165 61 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.63
+ $X2=9.865 $Y2=1.465
r166 61 62 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.865 $Y=1.63
+ $X2=9.865 $Y2=1.94
r167 60 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.3
+ $X2=9.865 $Y2=1.465
r168 60 71 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.865 $Y=1.3
+ $X2=9.865 $Y2=0.885
r169 55 73 6.11814 $w=2.6e-07 $l=2.2e-07 $layer=LI1_cond $X=9.775 $Y=2.38
+ $X2=9.775 $Y2=2.16
r170 55 57 14.3232 $w=3.48e-07 $l=4.35e-07 $layer=LI1_cond $X=9.775 $Y=2.38
+ $X2=9.775 $Y2=2.815
r171 53 77 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.875 $Y=2.215
+ $X2=8.875 $Y2=2.38
r172 53 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.875 $Y=2.215
+ $X2=8.875 $Y2=2.05
r173 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.875
+ $Y=2.215 $X2=8.875 $Y2=2.215
r174 50 73 0.606672 $w=3.2e-07 $l=2.02793e-07 $layer=LI1_cond $X=9.6 $Y=2.22
+ $X2=9.775 $Y2=2.16
r175 50 52 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=9.6 $Y=2.22
+ $X2=8.875 $Y2=2.22
r176 44 49 18.8402 $w=1.65e-07 $l=8.35165e-08 $layer=POLY_cond $X=11.99 $Y=1.3
+ $X2=11.972 $Y2=1.375
r177 44 46 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=11.99 $Y=1.3
+ $X2=11.99 $Y2=0.81
r178 40 49 18.8402 $w=1.65e-07 $l=7.59934e-08 $layer=POLY_cond $X=11.97 $Y=1.45
+ $X2=11.972 $Y2=1.375
r179 40 42 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=11.97 $Y=1.45
+ $X2=11.97 $Y2=2.34
r180 39 48 13.2179 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=11.075 $Y=1.375
+ $X2=10.982 $Y2=1.375
r181 38 49 6.66866 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=11.88 $Y=1.375
+ $X2=11.972 $Y2=1.375
r182 38 39 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=11.88 $Y=1.375
+ $X2=11.075 $Y2=1.375
r183 34 48 10.9219 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=11 $Y=1.3
+ $X2=10.982 $Y2=1.375
r184 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11 $Y=1.3 $X2=11
+ $Y2=0.74
r185 30 48 10.9219 $w=1.8e-07 $l=7.59934e-08 $layer=POLY_cond $X=10.98 $Y=1.45
+ $X2=10.982 $Y2=1.375
r186 30 32 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=10.98 $Y=1.45
+ $X2=10.98 $Y2=2.4
r187 29 66 7.86782 $w=1.5e-07 $l=1.40993e-07 $layer=POLY_cond $X=10.645 $Y=1.375
+ $X2=10.542 $Y2=1.465
r188 28 48 13.2179 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=10.89 $Y=1.375
+ $X2=10.982 $Y2=1.375
r189 28 29 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=10.89 $Y=1.375
+ $X2=10.645 $Y2=1.375
r190 24 66 16.8416 $w=1.5e-07 $l=1.78452e-07 $layer=POLY_cond $X=10.57 $Y=1.3
+ $X2=10.542 $Y2=1.465
r191 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.57 $Y=1.3
+ $X2=10.57 $Y2=0.74
r192 20 66 16.8416 $w=1.8e-07 $l=1.70895e-07 $layer=POLY_cond $X=10.53 $Y=1.63
+ $X2=10.542 $Y2=1.465
r193 20 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.53 $Y=1.63
+ $X2=10.53 $Y2=2.4
r194 16 76 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=8.965 $Y=1.015
+ $X2=8.965 $Y2=2.05
r195 14 77 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=8.8 $Y=2.75 $X2=8.8
+ $Y2=2.38
r196 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.89 $Y=0.94
+ $X2=8.965 $Y2=1.015
r197 10 11 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.89 $Y=0.94
+ $X2=8.705 $Y2=0.94
r198 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.63 $Y=0.865
+ $X2=8.705 $Y2=0.94
r199 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.63 $Y=0.865 $X2=8.63
+ $Y2=0.58
r200 2 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.96 $X2=9.765 $Y2=2.105
r201 2 57 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.96 $X2=9.765 $Y2=2.815
r202 1 69 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=9.585
+ $Y=0.37 $X2=9.725 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_1511_74# 1 2 9 12 16 18 22 24 25 27 28 31
+ 33 34 37 41 44
c105 34 0 3.61287e-20 $X=8.935 $Y=0.97
c106 31 0 8.50626e-20 $X=8.025 $Y=0.58
r107 41 45 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.385
+ $X2=9.455 $Y2=1.55
r108 41 44 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.385
+ $X2=9.455 $Y2=1.22
r109 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.445
+ $Y=1.385 $X2=9.445 $Y2=1.385
r110 37 40 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.445 $Y=1.14
+ $X2=9.445 $Y2=1.385
r111 34 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.935 $Y=0.97
+ $X2=8.935 $Y2=1.14
r112 31 32 17.365 $w=2.74e-07 $l=3.9e-07 $layer=LI1_cond $X=8.025 $Y=0.58
+ $X2=8.025 $Y2=0.97
r113 29 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=1.14
+ $X2=8.935 $Y2=1.14
r114 28 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.28 $Y=1.14
+ $X2=9.445 $Y2=1.14
r115 28 29 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.28 $Y=1.14
+ $X2=9.02 $Y2=1.14
r116 26 36 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=1.225
+ $X2=8.935 $Y2=1.14
r117 26 27 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.935 $Y=1.225
+ $X2=8.935 $Y2=1.72
r118 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.85 $Y=1.805
+ $X2=8.935 $Y2=1.72
r119 24 25 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=8.85 $Y=1.805
+ $X2=8.235 $Y2=1.805
r120 23 32 3.52985 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=0.97
+ $X2=8.025 $Y2=0.97
r121 22 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=0.97
+ $X2=8.935 $Y2=0.97
r122 22 23 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.85 $Y=0.97
+ $X2=8.19 $Y2=0.97
r123 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.15 $Y=1.89
+ $X2=8.235 $Y2=1.805
r124 20 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.15 $Y=1.89
+ $X2=8.15 $Y2=2.1
r125 16 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=2.265
+ $X2=8.07 $Y2=2.1
r126 16 18 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.07 $Y=2.265
+ $X2=8.07 $Y2=2.815
r127 12 45 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=9.54 $Y=2.46
+ $X2=9.54 $Y2=1.55
r128 9 44 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.51 $Y=0.74 $X2=9.51
+ $Y2=1.22
r129 2 18 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=7.935
+ $Y=2.12 $X2=8.07 $Y2=2.815
r130 2 16 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.935
+ $Y=2.12 $X2=8.07 $Y2=2.265
r131 1 31 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=7.555
+ $Y=0.37 $X2=8.025 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_2322_368# 1 2 9 13 17 21 25 29 35 38 43
c70 29 0 1.47924e-19 $X=11.745 $Y=1.985
r71 39 41 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=12.495 $Y=1.485
+ $X2=12.5 $Y2=1.485
r72 36 43 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=12.57 $Y=1.485
+ $X2=12.945 $Y2=1.485
r73 36 41 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=12.57 $Y=1.485
+ $X2=12.5 $Y2=1.485
r74 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.57
+ $Y=1.485 $X2=12.57 $Y2=1.485
r75 33 38 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=11.94 $Y=1.485
+ $X2=11.76 $Y2=1.485
r76 33 35 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=11.94 $Y=1.485
+ $X2=12.57 $Y2=1.485
r77 29 31 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.745 $Y=1.985
+ $X2=11.745 $Y2=2.695
r78 27 38 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=11.745 $Y=1.65
+ $X2=11.76 $Y2=1.485
r79 27 29 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.745 $Y=1.65
+ $X2=11.745 $Y2=1.985
r80 23 38 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=11.76 $Y=1.32
+ $X2=11.76 $Y2=1.485
r81 23 25 20.9681 $w=3.58e-07 $l=6.55e-07 $layer=LI1_cond $X=11.76 $Y=1.32
+ $X2=11.76 $Y2=0.665
r82 19 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.945 $Y=1.32
+ $X2=12.945 $Y2=1.485
r83 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.945 $Y=1.32
+ $X2=12.945 $Y2=0.76
r84 15 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.945 $Y=1.65
+ $X2=12.945 $Y2=1.485
r85 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=12.945 $Y=1.65
+ $X2=12.945 $Y2=2.4
r86 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.5 $Y=1.32
+ $X2=12.5 $Y2=1.485
r87 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.5 $Y=1.32
+ $X2=12.5 $Y2=0.76
r88 7 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.495 $Y=1.65
+ $X2=12.495 $Y2=1.485
r89 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=12.495 $Y=1.65
+ $X2=12.495 $Y2=2.4
r90 2 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=11.61
+ $Y=1.84 $X2=11.745 $Y2=2.695
r91 2 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.61
+ $Y=1.84 $X2=11.745 $Y2=1.985
r92 1 25 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=11.63
+ $Y=0.49 $X2=11.775 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 53
+ 56 60 64 66 69 70 72 73 75 78 82 83 85 97 108 116 120 125 131 134 137 140 144
r166 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r167 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r168 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r169 134 135 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r170 131 132 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r171 129 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r172 129 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r173 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r174 126 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.355 $Y=3.33
+ $X2=12.23 $Y2=3.33
r175 126 128 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.355 $Y=3.33
+ $X2=12.72 $Y2=3.33
r176 125 143 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=13.222 $Y2=3.33
r177 125 128 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=12.72 $Y2=3.33
r178 124 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r179 124 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r180 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r181 121 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.205 $Y2=3.33
r182 121 123 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.76 $Y2=3.33
r183 120 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.105 $Y=3.33
+ $X2=12.23 $Y2=3.33
r184 120 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=3.33
+ $X2=11.76 $Y2=3.33
r185 119 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r187 116 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=11.205 $Y2=3.33
r188 116 118 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=10.8 $Y2=3.33
r189 115 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r190 115 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r191 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r192 112 134 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.145 $Y2=3.33
r193 112 114 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.84 $Y2=3.33
r194 111 135 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r195 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r196 108 134 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=9.145 $Y2=3.33
r197 108 110 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r199 104 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r200 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r201 103 106 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r202 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 101 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.24 $Y2=3.33
r204 101 103 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 100 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r206 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r207 97 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=4.24 $Y2=3.33
r208 97 99 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=3.12 $Y2=3.33
r209 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r210 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r211 93 96 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 92 95 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r213 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r214 89 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r215 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r216 85 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 85 107 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r218 82 114 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=9.84 $Y2=3.33
r219 82 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.265 $Y2=3.33
r220 81 118 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.39 $Y=3.33
+ $X2=10.8 $Y2=3.33
r221 81 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.39 $Y=3.33
+ $X2=10.265 $Y2=3.33
r222 79 110 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.905 $Y=3.33
+ $X2=6.96 $Y2=3.33
r223 78 106 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.575 $Y=3.33
+ $X2=6.48 $Y2=3.33
r224 77 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=3.33
+ $X2=6.905 $Y2=3.33
r225 77 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=3.33
+ $X2=6.575 $Y2=3.33
r226 75 77 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6.74 $Y=3.04
+ $X2=6.74 $Y2=3.33
r227 72 95 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r228 72 73 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.88 $Y2=3.33
r229 71 99 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.09 $Y=3.33 $X2=3.12
+ $Y2=3.33
r230 71 73 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.09 $Y=3.33
+ $X2=2.88 $Y2=3.33
r231 69 88 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r233 68 92 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r234 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r235 64 143 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.222 $Y2=3.33
r236 64 66 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.405
r237 60 63 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.23 $Y=1.985
+ $X2=12.23 $Y2=2.815
r238 58 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.23 $Y=3.245
+ $X2=12.23 $Y2=3.33
r239 58 63 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.23 $Y=3.245
+ $X2=12.23 $Y2=2.815
r240 56 84 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=11.245 $Y=1.985
+ $X2=11.245 $Y2=2.14
r241 51 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=3.33
r242 51 53 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=2.4
r243 50 84 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.205 $Y=2.305
+ $X2=11.205 $Y2=2.14
r244 50 53 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=11.205 $Y=2.305
+ $X2=11.205 $Y2=2.4
r245 46 49 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.265 $Y=1.985
+ $X2=10.265 $Y2=2.815
r246 44 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=3.245
+ $X2=10.265 $Y2=3.33
r247 44 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.265 $Y=3.245
+ $X2=10.265 $Y2=2.815
r248 40 134 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=3.33
r249 40 42 9.02305 $w=5.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=2.815
r250 36 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=3.245
+ $X2=4.24 $Y2=3.33
r251 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.24 $Y=3.245
+ $X2=4.24 $Y2=2.805
r252 32 73 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=3.33
r253 32 34 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=2.875
r254 28 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r255 28 30 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.41
r256 9 66 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=13.035
+ $Y=1.84 $X2=13.17 $Y2=2.405
r257 8 63 600 $w=1.7e-07 $l=1.07488e-06 $layer=licon1_PDIFF $count=1 $X=12.06
+ $Y=1.84 $X2=12.27 $Y2=2.815
r258 8 60 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=12.06
+ $Y=1.84 $X2=12.27 $Y2=1.985
r259 7 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.07
+ $Y=1.84 $X2=11.205 $Y2=1.985
r260 7 53 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=11.07
+ $Y=1.84 $X2=11.205 $Y2=2.4
r261 6 49 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=2.815
r262 6 46 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=1.985
r263 5 42 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=8.89
+ $Y=2.54 $X2=9.145 $Y2=2.815
r264 4 75 600 $w=1.7e-07 $l=6.45697e-07 $layer=licon1_PDIFF $count=1 $X=6.52
+ $Y=2.495 $X2=6.74 $Y2=3.04
r265 3 38 600 $w=1.7e-07 $l=1.03496e-06 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=1.84 $X2=4.24 $Y2=2.805
r266 2 34 600 $w=1.7e-07 $l=7.30582e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=2.265 $X2=2.88 $Y2=2.875
r267 1 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.755
+ $Y=2.265 $X2=0.89 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%A_301_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 32 35 37 38 40 41 43
c122 24 0 6.78066e-20 $X=2.415 $Y=1.435
r123 43 46 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.21 $Y=2.58
+ $X2=5.21 $Y2=2.715
r124 38 42 23.0691 $w=2.14e-07 $l=4.25335e-07 $layer=LI1_cond $X=4.745 $Y=2.58
+ $X2=4.35 $Y2=2.517
r125 37 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.085 $Y=2.58
+ $X2=5.21 $Y2=2.58
r126 37 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.085 $Y=2.58
+ $X2=4.745 $Y2=2.58
r127 33 35 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.775 $Y=1.48
+ $X2=4.775 $Y2=0.76
r128 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.775 $Y2=1.48
r129 31 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.435 $Y2=1.565
r130 30 42 2.08775 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.35 $Y=2.37
+ $X2=4.35 $Y2=2.517
r131 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=1.65
+ $X2=4.435 $Y2=1.565
r132 29 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.35 $Y=1.65
+ $X2=4.35 $Y2=2.37
r133 28 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=2.455
+ $X2=3.01 $Y2=2.455
r134 27 42 5.39616 $w=2.14e-07 $l=1.11781e-07 $layer=LI1_cond $X=4.265 $Y=2.455
+ $X2=4.35 $Y2=2.517
r135 27 28 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.265 $Y=2.455
+ $X2=3.095 $Y2=2.455
r136 26 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=2.37
+ $X2=3.01 $Y2=2.455
r137 25 26 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=3.01 $Y=1.52
+ $X2=3.01 $Y2=2.37
r138 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.925 $Y=1.435
+ $X2=3.01 $Y2=1.52
r139 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.925 $Y=1.435
+ $X2=2.415 $Y2=1.435
r140 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=1.35
+ $X2=2.415 $Y2=1.435
r141 21 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.33 $Y=0.64
+ $X2=2.33 $Y2=1.35
r142 20 40 4.88517 $w=1.7e-07 $l=1.79374e-07 $layer=LI1_cond $X=1.98 $Y=2.455
+ $X2=1.815 $Y2=2.425
r143 19 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=2.455
+ $X2=3.01 $Y2=2.455
r144 19 20 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.925 $Y=2.455
+ $X2=1.98 $Y2=2.455
r145 13 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.245 $Y=0.515
+ $X2=2.33 $Y2=0.64
r146 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.245 $Y=0.515
+ $X2=1.8 $Y2=0.515
r147 4 46 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=2.495 $X2=5.25 $Y2=2.715
r148 3 40 300 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=2.265 $X2=1.815 $Y2=2.41
r149 2 35 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=4.68
+ $Y=0.485 $X2=4.815 $Y2=0.76
r150 1 15 182 $w=1.7e-07 $l=3.76298e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.8 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%Q 1 2 9 15 16 17 18 29
r39 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=10.785 $Y=0.965
+ $X2=10.785 $Y2=0.925
r40 18 31 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=10.785 $Y=0.987
+ $X2=10.785 $Y2=1.13
r41 18 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=10.785 $Y=0.987
+ $X2=10.785 $Y2=0.965
r42 18 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=10.785 $Y=0.902
+ $X2=10.785 $Y2=0.925
r43 17 18 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=10.785 $Y=0.515
+ $X2=10.785 $Y2=0.902
r44 15 16 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=10.77 $Y=1.8
+ $X2=10.77 $Y2=1.97
r45 15 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.865 $Y=1.8
+ $X2=10.865 $Y2=1.13
r46 9 11 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.715 $Y=1.985
+ $X2=10.715 $Y2=2.815
r47 9 16 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=10.715 $Y=1.985
+ $X2=10.715 $Y2=1.97
r48 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.755 $Y2=2.815
r49 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.755 $Y2=1.985
r50 1 17 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.645
+ $Y=0.37 $X2=10.785 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%Q_N 1 2 7 13 16 17 18
r28 30 31 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=13.195 $Y2=1.985
r29 27 30 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=12.695 $Y=1.985
+ $X2=12.72 $Y2=1.985
r30 22 31 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.82
+ $X2=13.195 $Y2=1.985
r31 18 31 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=13.2 $Y=1.985
+ $X2=13.195 $Y2=1.985
r32 17 22 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=13.195 $Y=1.665
+ $X2=13.195 $Y2=1.82
r33 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=13.195 $Y=1.295
+ $X2=13.195 $Y2=1.665
r34 15 16 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=13.195 $Y=1.15
+ $X2=13.195 $Y2=1.295
r35 11 27 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.695 $Y=2.15
+ $X2=12.695 $Y2=1.985
r36 11 13 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=12.695 $Y=2.15
+ $X2=12.695 $Y2=2.4
r37 7 15 6.82018 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=13.075 $Y=1.025
+ $X2=13.195 $Y2=1.15
r38 7 9 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=13.075 $Y=1.025
+ $X2=12.72 $Y2=1.025
r39 2 30 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.585
+ $Y=1.84 $X2=12.72 $Y2=1.985
r40 2 13 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=12.585
+ $Y=1.84 $X2=12.72 $Y2=2.4
r41 1 9 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=12.575
+ $Y=0.39 $X2=12.72 $Y2=0.985
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 32 36 42 46 50 54 59
+ 62 64 66 69 70 72 73 74 75 87 94 102 107 112 117 123 126 130 136 139 142 146
c159 46 0 1.1997e-19 $X=6.505 $Y=0.515
r160 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r161 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r162 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r163 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r164 130 133 9.0127 $w=7.08e-07 $l=5.35e-07 $layer=LI1_cond $X=9.035 $Y=0
+ $X2=9.035 $Y2=0.535
r165 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r166 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r167 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r168 121 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r169 121 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r170 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r171 118 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.45 $Y=0
+ $X2=12.285 $Y2=0
r172 118 120 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.45 $Y=0
+ $X2=12.72 $Y2=0
r173 117 145 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=13.217 $Y2=0
r174 117 120 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=12.72 $Y2=0
r175 116 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r176 116 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r177 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r178 113 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.38 $Y=0
+ $X2=11.255 $Y2=0
r179 113 115 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.38 $Y=0
+ $X2=11.76 $Y2=0
r180 112 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.12 $Y=0
+ $X2=12.285 $Y2=0
r181 112 115 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=12.12 $Y=0
+ $X2=11.76 $Y2=0
r182 111 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r183 111 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r184 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r185 108 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=0
+ $X2=10.285 $Y2=0
r186 108 110 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.45 $Y=0
+ $X2=10.8 $Y2=0
r187 107 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.13 $Y=0
+ $X2=11.255 $Y2=0
r188 107 110 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=11.13 $Y=0
+ $X2=10.8 $Y2=0
r189 106 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r190 106 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r191 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r192 103 130 9.41505 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=9.39 $Y=0
+ $X2=9.035 $Y2=0
r193 103 105 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.39 $Y=0
+ $X2=9.84 $Y2=0
r194 102 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.12 $Y=0
+ $X2=10.285 $Y2=0
r195 102 105 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.12 $Y=0
+ $X2=9.84 $Y2=0
r196 101 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r197 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r198 98 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.4 $Y2=0
r199 97 100 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r200 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r201 95 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=6.505 $Y2=0
r202 95 97 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.96
+ $Y2=0
r203 94 130 9.41505 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=8.68 $Y=0
+ $X2=9.035 $Y2=0
r204 94 100 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.68 $Y=0 $X2=8.4
+ $Y2=0
r205 93 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r206 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r207 90 93 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r208 89 92 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r209 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r210 87 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.505 $Y2=0
r211 87 92 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=6
+ $Y2=0
r212 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r213 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r214 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r215 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r216 80 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r217 80 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r218 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r219 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r220 77 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0
+ $X2=0.825 $Y2=0
r221 77 79 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r222 75 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.96 $Y2=0
r223 75 127 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r224 72 85 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r225 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.85
+ $Y2=0
r226 71 89 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.08
+ $Y2=0
r227 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.85
+ $Y2=0
r228 69 82 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.64
+ $Y2=0
r229 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.82
+ $Y2=0
r230 68 85 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r231 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.82
+ $Y2=0
r232 64 145 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=13.16 $Y=0.085
+ $X2=13.217 $Y2=0
r233 64 66 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=13.16 $Y=0.085
+ $X2=13.16 $Y2=0.55
r234 62 74 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=12.25 $Y=0.985
+ $X2=12.25 $Y2=0.73
r235 57 74 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.285 $Y=0.565
+ $X2=12.285 $Y2=0.73
r236 57 59 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.285 $Y=0.565
+ $X2=12.285 $Y2=0.55
r237 56 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.285 $Y=0.085
+ $X2=12.285 $Y2=0
r238 56 59 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=12.285 $Y=0.085
+ $X2=12.285 $Y2=0.55
r239 52 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=0.085
+ $X2=11.255 $Y2=0
r240 52 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.255 $Y=0.085
+ $X2=11.255 $Y2=0.515
r241 48 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0
r242 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.515
r243 44 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0.085
+ $X2=6.505 $Y2=0
r244 44 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.505 $Y=0.085
+ $X2=6.505 $Y2=0.515
r245 40 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0
r246 40 42 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0.595
r247 36 38 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.82 $Y=0.515
+ $X2=2.82 $Y2=0.965
r248 34 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0
r249 34 36 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0.515
r250 30 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r251 30 32 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.54
r252 9 66 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=13.02
+ $Y=0.39 $X2=13.16 $Y2=0.55
r253 8 62 182 $w=1.7e-07 $l=5.82301e-07 $layer=licon1_NDIFF $count=1 $X=12.065
+ $Y=0.49 $X2=12.255 $Y2=0.985
r254 8 59 182 $w=1.7e-07 $l=2.48193e-07 $layer=licon1_NDIFF $count=1 $X=12.065
+ $Y=0.49 $X2=12.285 $Y2=0.55
r255 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.075
+ $Y=0.37 $X2=11.215 $Y2=0.515
r256 6 50 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.14
+ $Y=0.37 $X2=10.285 $Y2=0.515
r257 5 133 91 $w=1.7e-07 $l=6.6742e-07 $layer=licon1_NDIFF $count=2 $X=8.705
+ $Y=0.37 $X2=9.295 $Y2=0.535
r258 4 46 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.365
+ $Y=0.37 $X2=6.505 $Y2=0.515
r259 3 42 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.85 $Y2=0.595
r260 2 38 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.86 $Y2=0.965
r261 2 36 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.86 $Y2=0.515
r262 1 32 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.37 $X2=0.825 $Y2=0.54
.ends


* File: sky130_fd_sc_ms__and4bb_4.pex.spice
* Created: Fri Aug 28 17:15:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4BB_4%B_N 1 3 6 8 9
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.615 $X2=0.405 $Y2=1.615
r29 9 14 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.405 $Y2=1.615
r30 8 14 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.405 $Y2=1.615
r31 4 13 38.5662 $w=2.97e-07 $l=2.00237e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.417 $Y2=1.615
r32 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.69
r33 1 13 48.8089 $w=2.97e-07 $l=2.95745e-07 $layer=POLY_cond $X=0.505 $Y=1.87
+ $X2=0.417 $Y2=1.615
r34 1 3 157.989 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=0.505 $Y=1.87
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_N 3 7 9 15
r33 13 15 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.055 $Y=1.615
+ $X2=1.17 $Y2=1.615
r34 11 13 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=0.925 $Y=1.615
+ $X2=1.055 $Y2=1.615
r35 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r36 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.78
+ $X2=1.055 $Y2=1.615
r37 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.055 $Y=1.78
+ $X2=1.055 $Y2=2.46
r38 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=0.925 $Y2=1.615
r39 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=0.925 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_200_74# 1 2 7 11 13 15 18 23 26 30 34 39
+ 40 49
c89 34 0 6.58453e-20 $X=1.525 $Y=0.42
c90 23 0 9.745e-20 $X=2.92 $Y=1.02
r91 48 49 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.905 $Y=1.6
+ $X2=2.92 $Y2=1.6
r92 47 48 66.5201 $w=3.6e-07 $l=4.15e-07 $layer=POLY_cond $X=2.49 $Y=1.6
+ $X2=2.905 $Y2=1.6
r93 46 47 32.8594 $w=3.6e-07 $l=2.05e-07 $layer=POLY_cond $X=2.285 $Y=1.6
+ $X2=2.49 $Y2=1.6
r94 35 40 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=0.42
+ $X2=1.525 $Y2=0.255
r95 34 37 9.44306 $w=5.62e-07 $l=4.35e-07 $layer=LI1_cond $X=1.367 $Y=0.42
+ $X2=1.367 $Y2=0.855
r96 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=0.42 $X2=1.525 $Y2=0.42
r97 31 46 30.455 $w=3.6e-07 $l=1.9e-07 $layer=POLY_cond $X=2.095 $Y=1.6
+ $X2=2.285 $Y2=1.6
r98 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.095
+ $Y=1.615 $X2=2.095 $Y2=1.615
r99 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.095 $Y=2.29
+ $X2=2.095 $Y2=1.615
r100 27 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.375
+ $X2=1.28 $Y2=2.375
r101 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.93 $Y=2.375
+ $X2=2.095 $Y2=2.29
r102 26 27 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.93 $Y=2.375
+ $X2=1.445 $Y2=2.375
r103 21 49 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.92 $Y=1.42
+ $X2=2.92 $Y2=1.6
r104 21 23 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.92 $Y=1.42 $X2=2.92
+ $Y2=1.02
r105 20 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.92 $Y=0.33
+ $X2=2.92 $Y2=1.02
r106 16 48 18.9685 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.905 $Y=1.78
+ $X2=2.905 $Y2=1.6
r107 16 18 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.905 $Y=1.78
+ $X2=2.905 $Y2=2.44
r108 13 47 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.49 $Y=1.42
+ $X2=2.49 $Y2=1.6
r109 13 15 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.49 $Y=1.42 $X2=2.49
+ $Y2=1.02
r110 9 46 18.9685 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.285 $Y=1.78
+ $X2=2.285 $Y2=1.6
r111 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.285 $Y=1.78
+ $X2=2.285 $Y2=2.44
r112 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.525 $Y2=0.255
r113 7 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.845 $Y=0.255
+ $X2=2.92 $Y2=0.33
r114 7 8 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=2.845 $Y=0.255
+ $X2=1.69 $Y2=0.255
r115 2 39 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=1.96 $X2=1.28 $Y2=2.455
r116 1 37 182 $w=1.7e-07 $l=5.80582e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_27_74# 1 2 10 13 18 21 24 26 29 31 33 35
+ 36 37 40 42 44 45 47 48 53 57
c132 42 0 2.63371e-20 $X=1.785 $Y=1.11
c133 24 0 3.95433e-21 $X=3.37 $Y=1.565
c134 13 0 1.77797e-19 $X=3.375 $Y=2.44
c135 10 0 2.67594e-19 $X=3.35 $Y=1.02
r136 55 57 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.785 $Y=0.84
+ $X2=1.945 $Y2=0.84
r137 52 53 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.59 $Y=1.195
+ $X2=1.785 $Y2=1.195
r138 48 59 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=3.44 $Y=0.42
+ $X2=3.35 $Y2=0.42
r139 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=0.42 $X2=3.44 $Y2=0.42
r140 45 47 49.2407 $w=3.28e-07 $l=1.41e-06 $layer=LI1_cond $X=2.03 $Y=0.42
+ $X2=3.44 $Y2=0.42
r141 44 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=0.755
+ $X2=1.945 $Y2=0.84
r142 43 45 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=0.585
+ $X2=2.03 $Y2=0.42
r143 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.945 $Y=0.585
+ $X2=1.945 $Y2=0.755
r144 42 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=1.11
+ $X2=1.785 $Y2=1.195
r145 41 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.925
+ $X2=1.785 $Y2=0.84
r146 41 42 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.785 $Y=0.925
+ $X2=1.785 $Y2=1.11
r147 39 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=1.28
+ $X2=1.59 $Y2=1.195
r148 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.59 $Y=1.28
+ $X2=1.59 $Y2=1.95
r149 38 51 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r150 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=2.035
+ $X2=1.59 $Y2=1.95
r151 37 38 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.505 $Y=2.035
+ $X2=0.445 $Y2=2.035
r152 35 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.195
+ $X2=1.59 $Y2=1.195
r153 35 36 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.505 $Y=1.195
+ $X2=0.365 $Y2=1.195
r154 31 51 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r155 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r156 27 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.365 $Y2=1.195
r157 27 29 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.24 $Y2=0.515
r158 25 26 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.825 $Y=1.415
+ $X2=3.825 $Y2=1.565
r159 23 24 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.37 $Y=1.415
+ $X2=3.37 $Y2=1.565
r160 21 26 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=3.855 $Y=2.44
+ $X2=3.855 $Y2=1.565
r161 18 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.78 $Y=1.02
+ $X2=3.78 $Y2=1.415
r162 15 48 65.0317 $w=2.52e-07 $l=4.14367e-07 $layer=POLY_cond $X=3.78 $Y=0.585
+ $X2=3.44 $Y2=0.42
r163 15 18 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.78 $Y=0.585
+ $X2=3.78 $Y2=1.02
r164 13 24 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=3.375 $Y=2.44
+ $X2=3.375 $Y2=1.565
r165 10 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.35 $Y=1.02
+ $X2=3.35 $Y2=1.415
r166 7 59 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=0.585
+ $X2=3.35 $Y2=0.42
r167 7 10 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.35 $Y=0.585
+ $X2=3.35 $Y2=1.02
r168 2 51 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r169 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r170 1 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%C 3 5 7 10 12 14 15 16 25
r53 23 25 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=5.27 $Y=1.615 $X2=5.47
+ $Y2=1.615
r54 22 23 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=4.855 $Y=1.615
+ $X2=5.27 $Y2=1.615
r55 21 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.84 $Y=1.615
+ $X2=4.855 $Y2=1.615
r56 19 21 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=4.405 $Y=1.615
+ $X2=4.84 $Y2=1.615
r57 15 16 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=5.47 $Y=1.615 $X2=6
+ $Y2=1.615
r58 15 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.47
+ $Y=1.615 $X2=5.47 $Y2=1.615
r59 12 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.27 $Y=1.45
+ $X2=5.27 $Y2=1.615
r60 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.27 $Y=1.45
+ $X2=5.27 $Y2=1.005
r61 8 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.78
+ $X2=4.855 $Y2=1.615
r62 8 10 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.855 $Y=1.78
+ $X2=4.855 $Y2=2.44
r63 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.45
+ $X2=4.84 $Y2=1.615
r64 5 7 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.84 $Y=1.45 $X2=4.84
+ $Y2=1.005
r65 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.78
+ $X2=4.405 $Y2=1.615
r66 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.405 $Y=1.78
+ $X2=4.405 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%D 3 7 11 15 17 25 26
c52 26 0 9.51185e-20 $X=6.73 $Y=1.515
c53 11 0 2.51603e-19 $X=6.69 $Y=0.79
r54 24 26 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.71 $Y=1.515 $X2=6.73
+ $Y2=1.515
r55 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.515 $X2=6.71 $Y2=1.515
r56 22 24 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.69 $Y=1.515 $X2=6.71
+ $Y2=1.515
r57 21 22 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.26 $Y=1.515
+ $X2=6.69 $Y2=1.515
r58 19 21 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.225 $Y=1.515
+ $X2=6.26 $Y2=1.515
r59 17 25 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.71 $Y2=1.565
r60 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.73 $Y=1.68
+ $X2=6.73 $Y2=1.515
r61 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.73 $Y=1.68
+ $X2=6.73 $Y2=2.34
r62 9 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.35
+ $X2=6.69 $Y2=1.515
r63 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.69 $Y=1.35 $X2=6.69
+ $Y2=0.79
r64 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.26 $Y=1.35
+ $X2=6.26 $Y2=1.515
r65 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.26 $Y=1.35 $X2=6.26
+ $Y2=0.79
r66 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.68
+ $X2=6.225 $Y2=1.515
r67 1 3 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=6.225 $Y=1.68
+ $X2=6.225 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_475_388# 1 2 3 4 5 18 22 26 30 34 38 40
+ 42 45 49 54 55 59 63 66 69 71 75 78 79 84 87 89 92 94 96 105
c172 89 0 1.54641e-19 $X=2.705 $Y=1.185
c173 78 0 1.51478e-19 $X=7.15 $Y=1.95
c174 54 0 2.58135e-19 $X=2.65 $Y=1.595
c175 49 0 5.89521e-20 $X=2.595 $Y=2.085
c176 22 0 1.60162e-19 $X=7.265 $Y=2.4
r177 105 106 0.728097 $w=3.31e-07 $l=5e-09 $layer=POLY_cond $X=8.615 $Y=1.53
+ $X2=8.62 $Y2=1.53
r178 89 91 7.39493 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.705 $Y=1.185
+ $X2=2.705 $Y2=1.36
r179 85 105 31.3082 $w=3.31e-07 $l=2.15e-07 $layer=POLY_cond $X=8.4 $Y=1.53
+ $X2=8.615 $Y2=1.53
r180 84 85 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.4
+ $Y=1.485 $X2=8.4 $Y2=1.485
r181 82 100 34.9486 $w=3.31e-07 $l=2.4e-07 $layer=POLY_cond $X=7.38 $Y=1.53
+ $X2=7.62 $Y2=1.53
r182 81 84 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=7.38 $Y=1.485
+ $X2=8.4 $Y2=1.485
r183 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.38
+ $Y=1.485 $X2=7.38 $Y2=1.485
r184 79 81 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.235 $Y=1.485
+ $X2=7.38 $Y2=1.485
r185 77 79 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.15 $Y=1.65
+ $X2=7.235 $Y2=1.485
r186 77 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.15 $Y=1.65 $X2=7.15
+ $Y2=1.95
r187 76 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=2.035
+ $X2=6.5 $Y2=2.035
r188 75 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.065 $Y=2.035
+ $X2=7.15 $Y2=1.95
r189 75 76 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.065 $Y=2.035
+ $X2=6.665 $Y2=2.035
r190 72 94 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.035
+ $X2=4.63 $Y2=2.035
r191 71 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=6.5 $Y2=2.035
r192 71 72 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=4.795 $Y2=2.035
r193 67 94 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=2.12
+ $X2=4.63 $Y2=2.035
r194 67 69 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.63 $Y=2.12
+ $X2=4.63 $Y2=2.795
r195 66 94 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=1.95
+ $X2=4.63 $Y2=2.035
r196 65 66 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.63 $Y=1.765
+ $X2=4.63 $Y2=1.95
r197 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=1.68
+ $X2=3.63 $Y2=1.68
r198 63 65 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.465 $Y=1.68
+ $X2=4.63 $Y2=1.765
r199 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.465 $Y=1.68
+ $X2=3.795 $Y2=1.68
r200 59 61 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.63 $Y=2.085
+ $X2=3.63 $Y2=2.795
r201 57 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=1.765
+ $X2=3.63 $Y2=1.68
r202 57 59 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.63 $Y=1.765
+ $X2=3.63 $Y2=2.085
r203 56 87 3.11956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=1.68
+ $X2=2.595 $Y2=1.68
r204 55 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=1.68
+ $X2=3.63 $Y2=1.68
r205 55 56 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.465 $Y=1.68
+ $X2=2.76 $Y2=1.68
r206 54 87 3.40559 $w=2.75e-07 $l=1.09087e-07 $layer=LI1_cond $X=2.65 $Y=1.595
+ $X2=2.595 $Y2=1.68
r207 54 91 12.3102 $w=2.18e-07 $l=2.35e-07 $layer=LI1_cond $X=2.65 $Y=1.595
+ $X2=2.65 $Y2=1.36
r208 49 51 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.595 $Y=2.085
+ $X2=2.595 $Y2=2.795
r209 47 87 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=1.68
r210 47 49 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=2.085
r211 43 106 21.295 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.62 $Y=1.32
+ $X2=8.62 $Y2=1.53
r212 43 45 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.62 $Y=1.32
+ $X2=8.62 $Y2=0.74
r213 40 105 17.0024 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.615 $Y=1.74
+ $X2=8.615 $Y2=1.53
r214 40 42 176.733 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=8.615 $Y=1.74
+ $X2=8.615 $Y2=2.4
r215 36 85 34.2205 $w=3.31e-07 $l=2.35e-07 $layer=POLY_cond $X=8.165 $Y=1.53
+ $X2=8.4 $Y2=1.53
r216 36 102 2.18429 $w=3.31e-07 $l=1.5e-08 $layer=POLY_cond $X=8.165 $Y=1.53
+ $X2=8.15 $Y2=1.53
r217 36 38 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.165 $Y=1.65
+ $X2=8.165 $Y2=2.4
r218 32 102 21.295 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.15 $Y=1.32
+ $X2=8.15 $Y2=1.53
r219 32 34 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.15 $Y=1.32
+ $X2=8.15 $Y2=0.74
r220 28 102 63.3444 $w=3.31e-07 $l=4.35e-07 $layer=POLY_cond $X=7.715 $Y=1.53
+ $X2=8.15 $Y2=1.53
r221 28 100 13.8338 $w=3.31e-07 $l=9.5e-08 $layer=POLY_cond $X=7.715 $Y=1.53
+ $X2=7.62 $Y2=1.53
r222 28 30 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.715 $Y=1.65
+ $X2=7.715 $Y2=2.4
r223 24 100 21.295 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.62 $Y=1.32
+ $X2=7.62 $Y2=1.53
r224 24 26 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.62 $Y=1.32
+ $X2=7.62 $Y2=0.74
r225 20 82 16.7462 $w=3.31e-07 $l=1.15e-07 $layer=POLY_cond $X=7.265 $Y=1.53
+ $X2=7.38 $Y2=1.53
r226 20 97 10.9215 $w=3.31e-07 $l=7.5e-08 $layer=POLY_cond $X=7.265 $Y=1.53
+ $X2=7.19 $Y2=1.53
r227 20 22 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.265 $Y=1.65
+ $X2=7.265 $Y2=2.4
r228 16 97 21.295 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.19 $Y=1.32
+ $X2=7.19 $Y2=1.53
r229 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.19 $Y=1.32
+ $X2=7.19 $Y2=0.74
r230 5 96 300 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=2 $X=6.315
+ $Y=1.94 $X2=6.5 $Y2=2.065
r231 4 94 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.94 $X2=4.63 $Y2=2.085
r232 4 69 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.94 $X2=4.63 $Y2=2.795
r233 3 61 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.94 $X2=3.63 $Y2=2.795
r234 3 59 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.94 $X2=3.63 $Y2=2.085
r235 2 51 400 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.94 $X2=2.595 $Y2=2.795
r236 2 49 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.94 $X2=2.595 $Y2=2.085
r237 1 89 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.7 $X2=2.705 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 41 49 55 57
+ 59 62 63 64 66 75 79 84 89 94 100 103 106 111 118 120 123 127
r120 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r121 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 115 118 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=2.852
+ $X2=6.165 $Y2=2.852
r124 115 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r125 113 115 9.43467 $w=1.123e-06 $l=8.7e-07 $layer=LI1_cond $X=5.13 $Y=2.852
+ $X2=6 $Y2=2.852
r126 110 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r127 109 113 0.976 $w=1.123e-06 $l=9e-08 $layer=LI1_cond $X=5.04 $Y=2.852
+ $X2=5.13 $Y2=2.852
r128 109 111 12.5495 $w=1.123e-06 $l=7.5e-08 $layer=LI1_cond $X=5.04 $Y=2.852
+ $X2=4.965 $Y2=2.852
r129 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r130 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r131 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r133 98 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r134 98 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r135 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r136 95 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=3.33
+ $X2=7.94 $Y2=3.33
r137 95 97 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.105 $Y=3.33
+ $X2=8.4 $Y2=3.33
r138 94 126 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.897 $Y2=3.33
r139 94 97 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.4 $Y2=3.33
r140 93 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r141 93 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r142 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r143 90 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.04 $Y2=3.33
r144 90 92 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 89 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.94 $Y2=3.33
r146 89 92 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r147 88 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r148 88 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r149 87 118 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=6.165 $Y2=3.33
r150 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r151 84 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=3.33
+ $X2=7.04 $Y2=3.33
r152 84 87 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.875 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 83 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r154 83 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r155 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r156 80 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.13 $Y2=3.33
r157 80 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.6 $Y2=3.33
r158 79 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.13 $Y2=3.33
r159 79 82 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 78 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r161 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 75 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.13 $Y2=3.33
r163 75 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r164 74 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r165 74 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r167 71 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r168 71 73 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r169 69 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r171 66 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r172 66 68 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r173 64 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r174 64 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 62 73 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=1.68 $Y2=3.33
r176 62 63 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=2.057 $Y2=3.33
r177 61 77 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.64 $Y2=3.33
r178 61 63 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.057 $Y2=3.33
r179 57 126 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.84 $Y=3.245
+ $X2=8.897 $Y2=3.33
r180 57 59 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.84 $Y=3.245
+ $X2=8.84 $Y2=2.405
r181 53 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=3.245
+ $X2=7.94 $Y2=3.33
r182 53 55 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=7.94 $Y=3.245
+ $X2=7.94 $Y2=2.405
r183 49 52 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=7.04 $Y=2.455
+ $X2=7.04 $Y2=2.815
r184 47 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=3.245
+ $X2=7.04 $Y2=3.33
r185 47 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.04 $Y=3.245
+ $X2=7.04 $Y2=2.815
r186 46 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.13 $Y2=3.33
r187 46 111 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.965 $Y2=3.33
r188 41 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.13 $Y=2.1
+ $X2=4.13 $Y2=2.795
r189 39 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=3.33
r190 39 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=2.795
r191 35 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.13 $Y=2.1
+ $X2=3.13 $Y2=2.795
r192 33 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r193 33 38 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.795
r194 29 63 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.057 $Y=3.245
+ $X2=2.057 $Y2=3.33
r195 29 31 17.0286 $w=3.33e-07 $l=4.95e-07 $layer=LI1_cond $X=2.057 $Y=3.245
+ $X2=2.057 $Y2=2.75
r196 25 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r197 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.455
r198 8 59 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.405
r199 7 55 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=7.805
+ $Y=1.84 $X2=7.94 $Y2=2.405
r200 6 52 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.84 $X2=7.04 $Y2=2.815
r201 6 49 600 $w=1.7e-07 $l=7.16607e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.84 $X2=7.04 $Y2=2.455
r202 5 115 200 $w=1.7e-07 $l=1.25377e-06 $layer=licon1_PDIFF $count=3 $X=4.945
+ $Y=1.94 $X2=6 $Y2=2.375
r203 5 113 200 $w=1.7e-07 $l=5.19326e-07 $layer=licon1_PDIFF $count=3 $X=4.945
+ $Y=1.94 $X2=5.13 $Y2=2.375
r204 4 44 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.94 $X2=4.13 $Y2=2.795
r205 4 41 400 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.94 $X2=4.13 $Y2=2.1
r206 3 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.995
+ $Y=1.94 $X2=3.13 $Y2=2.795
r207 3 35 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=2.995
+ $Y=1.94 $X2=3.13 $Y2=2.1
r208 2 31 600 $w=1.7e-07 $l=8.88679e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.94 $X2=2.055 $Y2=2.75
r209 1 27 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%X 1 2 3 4 15 17 19 22 23 27 28 33 34 35 36
+ 37 42 43
c63 27 0 1.28179e-19 $X=8.765 $Y=0.96
c64 22 0 1.0664e-19 $X=7.57 $Y=1.065
c65 17 0 1.60162e-19 $X=7.49 $Y=2.15
r66 37 43 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=1.82
r67 36 43 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.82
r68 35 36 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.665
r69 35 42 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.15
r70 34 42 4.58911 $w=2.3e-07 $l=1.9e-07 $layer=LI1_cond $X=8.88 $Y=0.96 $X2=8.88
+ $Y2=1.15
r71 32 33 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=0.96
+ $X2=8.24 $Y2=0.96
r72 28 32 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=8.43 $Y=0.96
+ $X2=8.405 $Y2=0.96
r73 27 34 2.77762 $w=3.8e-07 $l=1.15e-07 $layer=LI1_cond $X=8.765 $Y=0.96
+ $X2=8.88 $Y2=0.96
r74 27 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.765 $Y=0.96
+ $X2=8.43 $Y2=0.96
r75 24 30 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=1.985
+ $X2=7.49 $Y2=1.985
r76 24 26 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=7.575 $Y=1.985
+ $X2=8.39 $Y2=1.985
r77 23 37 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=8.765 $Y=1.985
+ $X2=8.88 $Y2=1.985
r78 23 26 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=8.765 $Y=1.985
+ $X2=8.39 $Y2=1.985
r79 22 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.57 $Y=1.065
+ $X2=8.24 $Y2=1.065
r80 17 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.49 $Y=2.15
+ $X2=7.49 $Y2=1.985
r81 17 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.49 $Y=2.15
+ $X2=7.49 $Y2=2.4
r82 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.405 $Y=0.98
+ $X2=7.57 $Y2=1.065
r83 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.405 $Y=0.98
+ $X2=7.405 $Y2=0.515
r84 4 26 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=1.985
r85 3 30 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.355
+ $Y=1.84 $X2=7.49 $Y2=1.985
r86 3 19 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=7.355
+ $Y=1.84 $X2=7.49 $Y2=2.4
r87 2 32 182 $w=1.7e-07 $l=6.63928e-07 $layer=licon1_NDIFF $count=1 $X=8.225
+ $Y=0.37 $X2=8.405 $Y2=0.95
r88 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.37 $X2=7.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43
+ 51 56 61 67 70 73 76 80
c97 5 0 1.28179e-19 $X=8.695 $Y=0.37
r98 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r99 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r100 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r101 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r102 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r104 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r105 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r106 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=7.905
+ $Y2=0
r107 62 64 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.4
+ $Y2=0
r108 61 79 4.77426 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.895
+ $Y2=0
r109 61 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.4
+ $Y2=0
r110 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r111 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r112 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r113 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.07 $Y=0 $X2=6.905
+ $Y2=0
r114 57 59 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.07 $Y=0 $X2=7.44
+ $Y2=0
r115 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.905
+ $Y2=0
r116 56 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.44
+ $Y2=0
r117 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r118 55 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r119 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r120 52 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.005
+ $Y2=0
r121 52 54 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.48
+ $Y2=0
r122 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=0 $X2=6.905
+ $Y2=0
r123 51 54 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.74 $Y=0 $X2=6.48
+ $Y2=0
r124 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r125 49 50 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r126 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r127 46 49 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.52
+ $Y2=0
r128 46 47 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r129 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r130 44 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r131 43 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.88 $Y=0 $X2=6.005
+ $Y2=0
r132 43 49 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.88 $Y=0 $X2=5.52
+ $Y2=0
r133 41 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r134 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r135 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r136 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r137 36 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r138 36 47 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r139 32 79 3.03431 $w=3.35e-07 $l=1.1025e-07 $layer=LI1_cond $X=8.837 $Y=0.085
+ $X2=8.895 $Y2=0
r140 32 34 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=8.837 $Y=0.085
+ $X2=8.837 $Y2=0.515
r141 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0
r142 28 30 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0.645
r143 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0
r144 24 26 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0.615
r145 20 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.085
+ $X2=6.005 $Y2=0
r146 20 22 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=6.005 $Y=0.085
+ $X2=6.005 $Y2=0.645
r147 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r148 16 18 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.495
r149 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.695
+ $Y=0.37 $X2=8.835 $Y2=0.515
r150 4 30 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.37 $X2=7.905 $Y2=0.645
r151 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.47 $X2=6.905 $Y2=0.615
r152 2 22 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=0.47 $X2=6.045 $Y2=0.645
r153 1 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_412_140# 1 2 3 11 12 13 18 19 26
c44 26 0 3.95433e-21 $X=3.995 $Y=1.185
c45 13 0 6.58453e-20 $X=2.37 $Y=0.84
r46 26 28 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.995 $Y=1.185
+ $X2=3.995 $Y2=1.34
r47 18 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.83 $Y=1.34
+ $X2=3.995 $Y2=1.34
r48 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.83 $Y=1.34
+ $X2=3.22 $Y2=1.34
r49 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.135 $Y=1.255
+ $X2=3.22 $Y2=1.34
r50 15 17 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.135 $Y=1.255
+ $X2=3.135 $Y2=1.055
r51 14 17 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.135 $Y=0.925
+ $X2=3.135 $Y2=1.055
r52 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.05 $Y=0.84
+ $X2=3.135 $Y2=0.925
r53 12 13 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.05 $Y=0.84
+ $X2=2.37 $Y2=0.84
r54 11 21 4.79607 $w=1.83e-07 $l=8e-08 $layer=LI1_cond $X=2.285 $Y=1.187
+ $X2=2.205 $Y2=1.187
r55 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.285 $Y=0.925
+ $X2=2.37 $Y2=0.84
r56 10 11 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=0.925
+ $X2=2.285 $Y2=1.095
r57 3 26 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.7 $X2=3.995 $Y2=1.185
r58 2 17 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.7 $X2=3.135 $Y2=1.055
r59 1 21 182 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.7 $X2=2.205 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_685_140# 1 2 11 14 15
c29 11 0 9.745e-20 $X=3.565 $Y=0.92
r30 14 15 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=0.802
+ $X2=4.89 $Y2=0.802
r31 8 11 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.65 $Y=0.84
+ $X2=3.525 $Y2=0.84
r32 8 15 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.65 $Y=0.84
+ $X2=4.89 $Y2=0.84
r33 2 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.685 $X2=5.055 $Y2=0.84
r34 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=3.425
+ $Y=0.7 $X2=3.565 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_4%A_882_137# 1 2 3 10 14 16 20 25 27
c44 20 0 1.44963e-19 $X=6.475 $Y=0.615
r45 23 25 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=1.22
+ $X2=4.72 $Y2=1.22
r46 18 20 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.435 $Y=1.01
+ $X2=6.435 $Y2=0.615
r47 17 27 7.02821 $w=1.7e-07 $l=1.47902e-07 $layer=LI1_cond $X=5.65 $Y=1.095
+ $X2=5.525 $Y2=1.145
r48 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.31 $Y=1.095
+ $X2=6.435 $Y2=1.01
r49 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.31 $Y=1.095
+ $X2=5.65 $Y2=1.095
r50 12 27 0.00168595 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=5.525 $Y=1.01
+ $X2=5.525 $Y2=1.145
r51 12 14 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=5.525 $Y=1.01
+ $X2=5.525 $Y2=0.83
r52 10 27 7.02821 $w=1.7e-07 $l=1.47902e-07 $layer=LI1_cond $X=5.4 $Y=1.195
+ $X2=5.525 $Y2=1.145
r53 10 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.4 $Y=1.195
+ $X2=4.72 $Y2=1.195
r54 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.335
+ $Y=0.47 $X2=6.475 $Y2=0.615
r55 2 27 182 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.685 $X2=5.485 $Y2=1.195
r56 2 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.685 $X2=5.485 $Y2=0.83
r57 1 23 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.685 $X2=4.555 $Y2=1.18
.ends


* File: sky130_fd_sc_ms__a32oi_1.pex.spice
* Created: Fri Aug 28 17:08:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A32OI_1%B2 3 5 7 8 15
r24 14 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.385
+ $X2=0.52 $Y2=1.385
r25 11 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.28 $Y=1.385
+ $X2=0.505 $Y2=1.385
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.385 $X2=0.28 $Y2=1.385
r27 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=1.295 $X2=0.28
+ $Y2=1.385
r28 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=1.385
r29 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.22 $X2=0.52
+ $Y2=0.74
r30 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.385
r31 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%B1 1 3 6 8 14
c32 8 0 1.62524e-19 $X=1.2 $Y=1.295
c33 6 0 1.68041e-19 $X=1.005 $Y=2.4
c34 1 0 1.47908e-19 $X=0.91 $Y=1.22
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.385 $X2=1.12 $Y2=1.385
r36 12 14 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.005 $Y=1.385
+ $X2=1.12 $Y2=1.385
r37 10 12 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.91 $Y=1.385
+ $X2=1.005 $Y2=1.385
r38 8 15 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.385
r39 4 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.55
+ $X2=1.005 $Y2=1.385
r40 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.005 $Y=1.55
+ $X2=1.005 $Y2=2.4
r41 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.22
+ $X2=0.91 $Y2=1.385
r42 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.91 $Y=1.22 $X2=0.91
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%A1 3 5 7 8 15
c33 8 0 1.47908e-19 $X=1.68 $Y=1.295
c34 5 0 1.62524e-19 $X=1.88 $Y=1.22
r35 13 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.88 $Y2=1.385
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.385 $X2=1.69 $Y2=1.385
r37 10 13 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.615 $Y=1.385
+ $X2=1.69 $Y2=1.385
r38 8 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.385
r39 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.22
+ $X2=1.88 $Y2=1.385
r40 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.88 $Y=1.22 $X2=1.88
+ $Y2=0.74
r41 1 10 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.55
+ $X2=1.615 $Y2=1.385
r42 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.615 $Y=1.55
+ $X2=1.615 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%A2 3 6 8 9 10 15 17
c40 17 0 3.79709e-20 $X=2.36 $Y=1.22
r41 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.385
+ $X2=2.36 $Y2=1.55
r42 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.385
+ $X2=2.36 $Y2=1.22
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.385 $X2=2.36 $Y2=1.385
r44 10 16 2.24265 $w=4.78e-07 $l=9e-08 $layer=LI1_cond $X=2.285 $Y=1.295
+ $X2=2.285 $Y2=1.385
r45 9 10 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.285 $Y=0.925
+ $X2=2.285 $Y2=1.295
r46 8 9 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.285 $Y=0.555
+ $X2=2.285 $Y2=0.925
r47 6 18 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.405 $Y=2.4
+ $X2=2.405 $Y2=1.55
r48 3 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.27 $Y=0.74 $X2=2.27
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%A3 3 6 8 11 13
c27 8 0 3.79709e-20 $X=3.12 $Y=1.295
r28 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.93 $Y=1.385
+ $X2=2.93 $Y2=1.55
r29 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.93 $Y=1.385
+ $X2=2.93 $Y2=1.22
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.385 $X2=2.93 $Y2=1.385
r31 8 12 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.93 $Y2=1.365
r32 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.855 $Y=2.4
+ $X2=2.855 $Y2=1.55
r33 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.84 $Y=0.74 $X2=2.84
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%A_27_368# 1 2 3 12 16 17 18 21 22 26 30 35
r50 33 34 6.99363 $w=3.14e-07 $l=1.8e-07 $layer=LI1_cond $X=1.28 $Y=2.225
+ $X2=1.28 $Y2=2.405
r51 28 35 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=2.655 $Y=2.49
+ $X2=2.63 $Y2=2.405
r52 28 30 13.3766 $w=2.78e-07 $l=3.25e-07 $layer=LI1_cond $X=2.655 $Y=2.49
+ $X2=2.655 $Y2=2.815
r53 24 35 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=2.32
+ $X2=2.63 $Y2=2.405
r54 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.63 $Y=2.32
+ $X2=2.63 $Y2=1.985
r55 23 34 4.32966 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.405
+ $X2=1.28 $Y2=2.405
r56 22 35 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=2.405
+ $X2=2.63 $Y2=2.405
r57 22 23 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.465 $Y=2.405
+ $X2=1.445 $Y2=2.405
r58 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.28 $Y=2.905 $X2=1.28
+ $Y2=2.815
r59 18 34 3.18267 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.49 $X2=1.28
+ $Y2=2.405
r60 18 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.28 $Y=2.49
+ $X2=1.28 $Y2=2.815
r61 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.905
r62 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r63 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r64 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r65 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r66 3 30 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.815
r67 3 26 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=1.985
r68 2 33 600 $w=1.7e-07 $l=4.68455e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.28 $Y2=2.225
r69 2 21 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.28 $Y2=2.815
r70 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r71 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%Y 1 2 8 11 13 15 19 20 23
c52 13 0 1.06273e-19 $X=0.785 $Y=0.68
c53 8 0 1.6439e-20 $X=0.7 $Y=1.72
r54 20 23 19.6393 $w=4.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.16 $Y=1.935
+ $X2=1.59 $Y2=1.935
r55 18 19 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.805
+ $X2=0.78 $Y2=1.805
r56 18 23 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.945 $Y=1.805
+ $X2=1.59 $Y2=1.805
r57 13 15 15.9477 $w=6.58e-07 $l=8.8e-07 $layer=LI1_cond $X=0.785 $Y=0.68
+ $X2=1.665 $Y2=0.68
r58 9 19 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.89 $X2=0.78
+ $Y2=1.805
r59 9 11 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.78 $Y=1.89 $X2=0.78
+ $Y2=1.985
r60 8 19 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.7 $Y=1.72
+ $X2=0.78 $Y2=1.805
r61 7 13 10.5067 $w=6.6e-07 $l=3.70068e-07 $layer=LI1_cond $X=0.7 $Y=1.01
+ $X2=0.785 $Y2=0.68
r62 7 8 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.7 $Y=1.01 $X2=0.7
+ $Y2=1.72
r63 2 11 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=1.985
r64 1 15 45.5 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_NDIFF $count=4 $X=0.985
+ $Y=0.37 $X2=1.665 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%VPWR 1 2 7 9 13 15 20 26 36
c39 26 0 1.68041e-19 $X=2.18 $Y=2.775
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 26 29 9.90781 $w=6.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.01 $Y=2.775
+ $X2=2.01 $Y2=3.33
r43 24 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 21 29 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.01 $Y2=3.33
r47 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 20 35 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r49 20 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 15 29 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=2.01 $Y2=3.33
r52 15 17 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 13 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 13 18 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 13 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=2.815
r57 7 35 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r58 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245 $X2=3.12
+ $Y2=2.815
r59 2 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.815
r60 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=1.985
r61 1 26 300 $w=1.7e-07 $l=1.14819e-06 $layer=licon1_PDIFF $count=2 $X=1.705
+ $Y=1.84 $X2=2.18 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_1%VGND 1 2 7 9 11 13 15 17 30
r31 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r32 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r34 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r36 20 23 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r37 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 18 26 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r39 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r40 17 29 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.125
+ $Y2=0
r41 17 23 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.64
+ $Y2=0
r42 15 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r43 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r44 11 29 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.125 $Y2=0
r45 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.515
r46 7 26 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r47 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r48 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.515
r49 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__sdfstp_4.pex.spice
* Created: Fri Aug 28 18:13:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%SCE 3 7 11 15 17 18 20 25 29 33
r77 25 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.645 $X2=0.69 $Y2=1.645
r78 21 33 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.88 $Y=1.415
+ $X2=2.01 $Y2=1.415
r79 20 23 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.88 $Y=1.415 $X2=1.88
+ $Y2=1.495
r80 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.415 $X2=1.88 $Y2=1.415
r81 18 25 9.23067 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.855 $Y=1.495
+ $X2=0.72 $Y2=1.58
r82 17 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.495
+ $X2=1.88 $Y2=1.495
r83 17 18 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.715 $Y=1.495
+ $X2=0.855 $Y2=1.495
r84 13 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.25
+ $X2=2.01 $Y2=1.415
r85 13 15 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.01 $Y=1.25
+ $X2=2.01 $Y2=0.58
r86 9 29 82.022 $w=3.03e-07 $l=6.07166e-07 $layer=POLY_cond $X=0.945 $Y=2.15
+ $X2=0.72 $Y2=1.645
r87 9 11 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=0.945 $Y=2.15
+ $X2=0.945 $Y2=2.64
r88 5 29 44.7447 $w=6.06e-07 $l=2.96226e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.72 $Y2=1.645
r89 5 7 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.495 $Y=1.48 $X2=0.495
+ $Y2=0.58
r90 1 29 82.022 $w=3.03e-07 $l=6.07166e-07 $layer=POLY_cond $X=0.495 $Y=2.15
+ $X2=0.72 $Y2=1.645
r91 1 3 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=2.15
+ $X2=0.495 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_27_74# 1 2 9 12 16 19 22 26 27 31 32 34
+ 36 38
c80 22 0 1.66495e-19 $X=1.785 $Y=2.405
r81 32 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.995
+ $X2=1.95 $Y2=2.16
r82 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.995 $X2=1.95 $Y2=1.995
r83 29 31 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=1.915 $Y=2.32
+ $X2=1.915 $Y2=1.995
r84 27 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.075
+ $X2=0.975 $Y2=0.91
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.075 $X2=0.975 $Y2=1.075
r86 24 34 0.94211 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=0.445 $Y=1.075
+ $X2=0.275 $Y2=1.075
r87 24 26 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.445 $Y=1.075
+ $X2=0.975 $Y2=1.075
r88 23 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.355 $Y=2.405
+ $X2=0.23 $Y2=2.405
r89 22 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.785 $Y=2.405
+ $X2=1.915 $Y2=2.32
r90 22 23 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.785 $Y=2.405
+ $X2=0.355 $Y2=2.405
r91 19 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.32 $X2=0.23
+ $Y2=2.405
r92 18 34 5.66538 $w=2.95e-07 $l=1.86145e-07 $layer=LI1_cond $X=0.23 $Y=1.24
+ $X2=0.275 $Y2=1.075
r93 18 19 49.7855 $w=2.48e-07 $l=1.08e-06 $layer=LI1_cond $X=0.23 $Y=1.24
+ $X2=0.23 $Y2=2.32
r94 14 34 5.66538 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=0.91
+ $X2=0.275 $Y2=1.075
r95 14 16 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=0.275 $Y=0.91
+ $X2=0.275 $Y2=0.58
r96 12 42 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=1.995 $Y=2.64
+ $X2=1.995 $Y2=2.16
r97 9 38 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.035 $Y=0.58
+ $X2=1.035 $Y2=0.91
r98 2 36 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.27 $Y2=2.465
r99 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%D 3 7 9 12 13
c41 12 0 4.43302e-20 $X=1.41 $Y=1.985
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.985
+ $X2=1.41 $Y2=2.15
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.985
+ $X2=1.41 $Y2=1.82
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.985 $X2=1.41 $Y2=1.985
r45 9 13 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.2 $Y=1.985 $X2=1.41
+ $Y2=1.985
r46 7 14 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.425 $Y=0.58
+ $X2=1.425 $Y2=1.82
r47 3 15 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=1.365 $Y=2.64
+ $X2=1.365 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%SCD 3 6 9 11 12 13 18 22
c45 11 0 1.07359e-19 $X=2.64 $Y=1.295
c46 9 0 1.66495e-19 $X=2.415 $Y=2.64
r47 22 24 41.7466 $w=5.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.592 $Y=1.945
+ $X2=2.592 $Y2=2.11
r48 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.945 $X2=2.695 $Y2=1.945
r49 18 20 47.5561 $w=5.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.592 $Y=1.265
+ $X2=2.592 $Y2=1.1
r50 13 23 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.695 $Y=2.035
+ $X2=2.695 $Y2=1.945
r51 12 23 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=2.695 $Y=1.665
+ $X2=2.695 $Y2=1.945
r52 11 12 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=2.695 $Y=1.265
+ $X2=2.695 $Y2=1.665
r53 11 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.265 $X2=2.695 $Y2=1.265
r54 9 24 206.016 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=2.415 $Y=2.64
+ $X2=2.415 $Y2=2.11
r55 6 22 10.2006 $w=5.35e-07 $l=1.02e-07 $layer=POLY_cond $X=2.592 $Y=1.843
+ $X2=2.592 $Y2=1.945
r56 5 18 10.2006 $w=5.35e-07 $l=1.02e-07 $layer=POLY_cond $X=2.592 $Y=1.367
+ $X2=2.592 $Y2=1.265
r57 5 6 47.6026 $w=5.35e-07 $l=4.76e-07 $layer=POLY_cond $X=2.592 $Y=1.367
+ $X2=2.592 $Y2=1.843
r58 3 20 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.4 $Y=0.58 $X2=2.4
+ $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%CLK 3 6 8 11 13
c38 6 0 1.07359e-19 $X=3.51 $Y=2.4
r39 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.385
+ $X2=3.49 $Y2=1.55
r40 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.385
+ $X2=3.49 $Y2=1.22
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.385 $X2=3.49 $Y2=1.385
r42 8 12 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.49
+ $Y2=1.365
r43 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.51 $Y=2.4 $X2=3.51
+ $Y2=1.55
r44 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.44 $Y=0.74 $X2=3.44
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_803_74# 1 2 9 11 15 19 20 21 23 24 26 28
+ 31 34 35 38 40 41 42 46 52 54 55 58 59 60 62 63 64 65 67 70 74 75 77 78 81 82
+ 87 88 93 97 104 106
c287 97 0 3.98141e-20 $X=10.6 $Y=1.97
c288 77 0 2.67659e-20 $X=5.665 $Y=1.94
c289 64 0 1.23112e-19 $X=7.545 $Y=2.035
c290 20 0 1.22616e-19 $X=9.375 $Y=1.16
r291 103 104 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.09 $Y=1.565
+ $X2=5.18 $Y2=1.565
r292 97 108 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=10.6 $Y=1.97
+ $X2=10.44 $Y2=1.97
r293 96 97 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.6
+ $Y=1.97 $X2=10.6 $Y2=1.97
r294 93 96 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=10.6 $Y=1.845
+ $X2=10.6 $Y2=1.97
r295 90 91 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=9.21 $Y=1.845
+ $X2=9.21 $Y2=1.865
r296 88 106 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=1.615
+ $X2=9.21 $Y2=1.45
r297 87 90 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=9.21 $Y=1.615
+ $X2=9.21 $Y2=1.845
r298 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.21
+ $Y=1.615 $X2=9.21 $Y2=1.615
r299 82 84 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.81 $Y=1.865
+ $X2=7.81 $Y2=2.035
r300 77 80 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=1.94
+ $X2=5.685 $Y2=2.105
r301 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.665
+ $Y=1.94 $X2=5.665 $Y2=1.94
r302 74 75 8.76268 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=4.945 $Y=1.095
+ $X2=4.945 $Y2=1.265
r303 70 72 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.235 $Y=2.78
+ $X2=4.235 $Y2=2.98
r304 68 90 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.375 $Y=1.845
+ $X2=9.21 $Y2=1.845
r305 67 93 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.435 $Y=1.845
+ $X2=10.6 $Y2=1.845
r306 67 68 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=10.435 $Y=1.845
+ $X2=9.375 $Y2=1.845
r307 66 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.895 $Y=1.865
+ $X2=7.81 $Y2=1.865
r308 65 91 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.865
+ $X2=9.21 $Y2=1.865
r309 65 66 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=9.045 $Y=1.865
+ $X2=7.895 $Y2=1.865
r310 63 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.81 $Y2=2.035
r311 63 64 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.545 $Y2=2.035
r312 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.46 $Y=2.12
+ $X2=7.545 $Y2=2.035
r313 61 62 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=7.46 $Y=2.12
+ $X2=7.46 $Y2=2.895
r314 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.375 $Y=2.98
+ $X2=7.46 $Y2=2.895
r315 59 60 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.375 $Y=2.98
+ $X2=6.865 $Y2=2.98
r316 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.78 $Y=2.895
+ $X2=6.865 $Y2=2.98
r317 57 58 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.78 $Y=2.46
+ $X2=6.78 $Y2=2.895
r318 56 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=2.375
+ $X2=5.745 $Y2=2.375
r319 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.695 $Y=2.375
+ $X2=6.78 $Y2=2.46
r320 55 56 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.695 $Y=2.375
+ $X2=5.83 $Y2=2.375
r321 53 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=2.46
+ $X2=5.745 $Y2=2.375
r322 53 54 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.745 $Y=2.46
+ $X2=5.745 $Y2=2.895
r323 52 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=2.29
+ $X2=5.745 $Y2=2.375
r324 52 80 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.745 $Y=2.29
+ $X2=5.745 $Y2=2.105
r325 49 74 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.055 $Y=0.425
+ $X2=5.055 $Y2=1.095
r326 47 103 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.9 $Y=1.565
+ $X2=5.09 $Y2=1.565
r327 46 75 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=4.89 $Y=1.565
+ $X2=4.89 $Y2=1.265
r328 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.565 $X2=4.9 $Y2=1.565
r329 43 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=2.98
+ $X2=4.235 $Y2=2.98
r330 42 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.66 $Y=2.98
+ $X2=5.745 $Y2=2.895
r331 42 43 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.66 $Y=2.98
+ $X2=4.4 $Y2=2.98
r332 40 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.97 $Y=0.34
+ $X2=5.055 $Y2=0.425
r333 40 41 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.97 $Y=0.34
+ $X2=4.24 $Y2=0.34
r334 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=0.425
+ $X2=4.24 $Y2=0.34
r335 36 38 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.155 $Y=0.425
+ $X2=4.155 $Y2=0.515
r336 33 78 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.665 $Y=1.73
+ $X2=5.665 $Y2=1.94
r337 33 34 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=5.665 $Y=1.73
+ $X2=5.665 $Y2=1.655
r338 29 108 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.44 $Y=2.135
+ $X2=10.44 $Y2=1.97
r339 29 31 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=10.44 $Y=2.135
+ $X2=10.44 $Y2=2.75
r340 26 28 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.16 $Y=1.085
+ $X2=10.16 $Y2=0.69
r341 25 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.805 $Y=1.16
+ $X2=9.73 $Y2=1.16
r342 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.085 $Y=1.16
+ $X2=10.16 $Y2=1.085
r343 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.085 $Y=1.16
+ $X2=9.805 $Y2=1.16
r344 21 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.73 $Y=1.085
+ $X2=9.73 $Y2=1.16
r345 21 23 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.73 $Y=1.085
+ $X2=9.73 $Y2=0.69
r346 19 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.655 $Y=1.16
+ $X2=9.73 $Y2=1.16
r347 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.655 $Y=1.16
+ $X2=9.375 $Y2=1.16
r348 17 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.3 $Y=1.235
+ $X2=9.375 $Y2=1.16
r349 17 106 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=9.3 $Y=1.235
+ $X2=9.3 $Y2=1.45
r350 13 34 13.5877 $w=2.4e-07 $l=8.66025e-08 $layer=POLY_cond $X=5.69 $Y=1.58
+ $X2=5.665 $Y2=1.655
r351 13 15 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=5.69 $Y=1.58
+ $X2=5.69 $Y2=0.615
r352 11 34 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.655
+ $X2=5.665 $Y2=1.655
r353 11 104 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.5 $Y=1.655
+ $X2=5.18 $Y2=1.655
r354 7 103 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.73
+ $X2=5.09 $Y2=1.565
r355 7 9 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=5.09 $Y=1.73
+ $X2=5.09 $Y2=2.495
r356 2 70 600 $w=1.7e-07 $l=1.02835e-06 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.84 $X2=4.235 $Y2=2.78
r357 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.015
+ $Y=0.37 $X2=4.155 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_1201_55# 1 2 9 12 16 18 22 26 28 32 35 36
+ 41 44
c88 44 0 2.67659e-20 $X=6.205 $Y=1.78
r89 42 44 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.26 $Y=1.265
+ $X2=6.26 $Y2=1.78
r90 36 45 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.945
+ $X2=6.205 $Y2=2.11
r91 36 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.945
+ $X2=6.205 $Y2=1.78
r92 35 38 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.205 $Y=1.945
+ $X2=6.205 $Y2=2.035
r93 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.205
+ $Y=1.945 $X2=6.205 $Y2=1.945
r94 32 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.1
+ $X2=6.17 $Y2=1.265
r95 32 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.1
+ $X2=6.17 $Y2=0.935
r96 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.17
+ $Y=1.1 $X2=6.17 $Y2=1.1
r97 28 31 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.17 $Y=0.855
+ $X2=6.17 $Y2=1.1
r98 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.12 $Y=2.12
+ $X2=7.12 $Y2=2.495
r99 20 22 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.935 $Y=0.77
+ $X2=6.935 $Y2=0.58
r100 19 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=2.035
+ $X2=6.205 $Y2=2.035
r101 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.035 $Y=2.035
+ $X2=7.12 $Y2=2.12
r102 18 19 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.035 $Y=2.035
+ $X2=6.37 $Y2=2.035
r103 17 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=0.855
+ $X2=6.17 $Y2=0.855
r104 16 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.77 $Y=0.855
+ $X2=6.935 $Y2=0.77
r105 16 17 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.77 $Y=0.855
+ $X2=6.335 $Y2=0.855
r106 12 45 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=6.13 $Y=2.495
+ $X2=6.13 $Y2=2.11
r107 9 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.08 $Y=0.615
+ $X2=6.08 $Y2=0.935
r108 2 26 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=6.955
+ $Y=2.285 $X2=7.12 $Y2=2.495
r109 1 22 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.79
+ $Y=0.37 $X2=6.935 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_1017_81# 1 2 9 11 13 16 18 20 23 25 27 31
+ 32 35 37 41 43 45 47 48 49 53 56 66
c164 23 0 7.59542e-20 $X=8.475 $Y=2.285
c165 9 0 1.23112e-19 $X=6.865 $Y=2.495
r166 65 66 27.3299 $w=2.91e-07 $l=1.65e-07 $layer=POLY_cond $X=8.31 $Y=1.267
+ $X2=8.475 $Y2=1.267
r167 60 65 34.7835 $w=2.91e-07 $l=2.1e-07 $layer=POLY_cond $X=8.1 $Y=1.267
+ $X2=8.31 $Y2=1.267
r168 60 63 12.4227 $w=2.91e-07 $l=7.5e-08 $layer=POLY_cond $X=8.1 $Y=1.267
+ $X2=8.025 $Y2=1.267
r169 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.1
+ $Y=1.285 $X2=8.1 $Y2=1.285
r170 56 59 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.1 $Y=1.195 $X2=8.1
+ $Y2=1.285
r171 52 54 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.79 $Y=1.275
+ $X2=6.79 $Y2=1.52
r172 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.79
+ $Y=1.275 $X2=6.79 $Y2=1.275
r173 49 52 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.79 $Y=1.195 $X2=6.79
+ $Y2=1.275
r174 46 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=1.195
+ $X2=6.79 $Y2=1.195
r175 45 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.935 $Y=1.195
+ $X2=8.1 $Y2=1.195
r176 45 46 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=7.935 $Y=1.195
+ $X2=6.955 $Y2=1.195
r177 44 47 2.76166 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=5.64 $Y=1.52
+ $X2=5.42 $Y2=1.52
r178 43 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=1.52
+ $X2=6.79 $Y2=1.52
r179 43 44 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=6.625 $Y=1.52
+ $X2=5.64 $Y2=1.52
r180 39 47 3.70735 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=5.475 $Y=1.435
+ $X2=5.42 $Y2=1.52
r181 39 41 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=5.475 $Y=1.435
+ $X2=5.475 $Y2=0.615
r182 35 48 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=5.34 $Y=2.415
+ $X2=5.34 $Y2=2.275
r183 35 37 3.49849 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=2.415
+ $X2=5.34 $Y2=2.5
r184 33 47 3.70735 $w=2.5e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.285 $Y=1.605
+ $X2=5.42 $Y2=1.52
r185 33 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.285 $Y=1.605
+ $X2=5.285 $Y2=2.275
r186 31 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.79 $Y=1.615
+ $X2=6.79 $Y2=1.275
r187 31 32 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.79 $Y=1.615
+ $X2=6.79 $Y2=1.78
r188 25 66 43.8935 $w=2.91e-07 $l=3.44173e-07 $layer=POLY_cond $X=8.74 $Y=1.085
+ $X2=8.475 $Y2=1.267
r189 25 27 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.74 $Y=1.085
+ $X2=8.74 $Y2=0.69
r190 21 66 14.0159 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=8.475 $Y=1.45
+ $X2=8.475 $Y2=1.267
r191 21 23 324.573 $w=1.8e-07 $l=8.35e-07 $layer=POLY_cond $X=8.475 $Y=1.45
+ $X2=8.475 $Y2=2.285
r192 18 65 18.2534 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=8.31 $Y=1.085
+ $X2=8.31 $Y2=1.267
r193 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.31 $Y=1.085
+ $X2=8.31 $Y2=0.69
r194 14 63 14.0159 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=8.025 $Y=1.45
+ $X2=8.025 $Y2=1.267
r195 14 16 324.573 $w=1.8e-07 $l=8.35e-07 $layer=POLY_cond $X=8.025 $Y=1.45
+ $X2=8.025 $Y2=2.285
r196 11 53 79.2329 $w=2.19e-07 $l=5.61872e-07 $layer=POLY_cond $X=7.15 $Y=0.865
+ $X2=6.79 $Y2=1.275
r197 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.15 $Y=0.865
+ $X2=7.15 $Y2=0.58
r198 9 32 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=6.865 $Y=2.495
+ $X2=6.865 $Y2=1.78
r199 2 37 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=5.18
+ $Y=2.285 $X2=5.315 $Y2=2.5
r200 1 41 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=5.085
+ $Y=0.405 $X2=5.475 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%SET_B 3 7 10 13 17 19 20 21 26 32 33 36 37
c132 26 0 1.12416e-19 $X=11.76 $Y=1.665
c133 20 0 6.13349e-20 $X=11.615 $Y=1.665
c134 10 0 7.95967e-20 $X=11.612 $Y=1.953
c135 3 0 1.49331e-19 $X=7.345 $Y=2.495
r136 36 38 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=11.612 $Y=1.635
+ $X2=11.612 $Y2=1.47
r137 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.635
+ $Y=1.635 $X2=11.635 $Y2=1.635
r138 31 33 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.36 $Y=1.615
+ $X2=7.54 $Y2=1.615
r139 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.36
+ $Y=1.615 $X2=7.36 $Y2=1.615
r140 28 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.345 $Y=1.615
+ $X2=7.36 $Y2=1.615
r141 26 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=1.665
+ $X2=11.76 $Y2=1.665
r142 23 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=1.665
r143 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.665
+ $X2=7.44 $Y2=1.665
r144 20 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=11.76 $Y2=1.665
r145 20 21 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=7.585 $Y2=1.665
r146 17 38 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=11.6 $Y=0.58
+ $X2=11.6 $Y2=1.47
r147 13 19 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=11.515 $Y=2.75
+ $X2=11.515 $Y2=2.14
r148 10 19 42.8297 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=11.612 $Y=1.953
+ $X2=11.612 $Y2=2.14
r149 9 36 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=11.612 $Y=1.657
+ $X2=11.612 $Y2=1.635
r150 9 10 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=11.612 $Y=1.657
+ $X2=11.612 $Y2=1.953
r151 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.54 $Y=1.45
+ $X2=7.54 $Y2=1.615
r152 5 7 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.54 $Y=1.45 $X2=7.54
+ $Y2=0.58
r153 1 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.78
+ $X2=7.345 $Y2=1.615
r154 1 3 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=7.345 $Y=1.78
+ $X2=7.345 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_616_74# 1 2 9 13 16 18 20 21 22 23 24 27
+ 31 33 35 37 38 43 44 45 48 52 54 55 58 61 62 63 68 71 76
c192 20 0 1.31023e-19 $X=4.53 $Y=3.075
r193 72 74 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.94 $Y=1.515
+ $X2=3.96 $Y2=1.515
r194 69 76 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=4.05 $Y=1.515
+ $X2=4.45 $Y2=1.515
r195 69 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.05 $Y=1.515
+ $X2=3.96 $Y2=1.515
r196 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r197 66 68 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.515
r198 63 65 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.175 $Y=1.945
+ $X2=3.285 $Y2=1.945
r199 62 66 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=4.05 $Y2=1.82
r200 62 65 27.6586 $w=2.48e-07 $l=6e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=3.285 $Y2=1.945
r201 61 63 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.09 $Y=1.82
+ $X2=3.175 $Y2=1.945
r202 61 71 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.09 $Y=1.82
+ $X2=3.09 $Y2=1.01
r203 56 71 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=3.197 $Y=0.818
+ $X2=3.197 $Y2=1.01
r204 56 58 9.06988 $w=3.83e-07 $l=3.03e-07 $layer=LI1_cond $X=3.197 $Y=0.818
+ $X2=3.197 $Y2=0.515
r205 50 52 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=4.45 $Y=2.045
+ $X2=4.53 $Y2=2.045
r206 46 48 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=10.67 $Y=1.445
+ $X2=10.67 $Y2=0.58
r207 44 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.595 $Y=1.52
+ $X2=10.67 $Y2=1.445
r208 44 45 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=10.595 $Y=1.52
+ $X2=10.025 $Y2=1.52
r209 41 43 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=9.935 $Y=3.075
+ $X2=9.935 $Y2=2.54
r210 40 45 22.7899 $w=1.97e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.935 $Y=1.685
+ $X2=10.025 $Y2=1.52
r211 40 43 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=9.935 $Y=1.685
+ $X2=9.935 $Y2=2.54
r212 39 55 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.575 $Y=3.15
+ $X2=9.485 $Y2=3.15
r213 38 41 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.845 $Y=3.15
+ $X2=9.935 $Y2=3.075
r214 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.845 $Y=3.15
+ $X2=9.575 $Y2=3.15
r215 35 55 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.485 $Y=3.075
+ $X2=9.485 $Y2=3.15
r216 35 37 143.261 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=9.485 $Y=3.075
+ $X2=9.485 $Y2=2.54
r217 34 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.715 $Y=3.15
+ $X2=5.625 $Y2=3.15
r218 33 55 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.395 $Y=3.15
+ $X2=9.485 $Y2=3.15
r219 33 34 1886.98 $w=1.5e-07 $l=3.68e-06 $layer=POLY_cond $X=9.395 $Y=3.15
+ $X2=5.715 $Y2=3.15
r220 29 54 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.625 $Y=3.075
+ $X2=5.625 $Y2=3.15
r221 29 31 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=5.625 $Y=3.075
+ $X2=5.625 $Y2=2.685
r222 25 27 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=5.01 $Y=1.04
+ $X2=5.01 $Y2=0.615
r223 23 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.535 $Y=3.15
+ $X2=5.625 $Y2=3.15
r224 23 24 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=5.535 $Y=3.15
+ $X2=4.605 $Y2=3.15
r225 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.935 $Y=1.115
+ $X2=5.01 $Y2=1.04
r226 21 22 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.935 $Y=1.115
+ $X2=4.525 $Y2=1.115
r227 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.53 $Y=3.075
+ $X2=4.605 $Y2=3.15
r228 19 52 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.53 $Y=2.12
+ $X2=4.53 $Y2=2.045
r229 19 20 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=4.53 $Y=2.12
+ $X2=4.53 $Y2=3.075
r230 18 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.45 $Y=1.97
+ $X2=4.45 $Y2=2.045
r231 17 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.45 $Y=1.68
+ $X2=4.45 $Y2=1.515
r232 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.45 $Y=1.68
+ $X2=4.45 $Y2=1.97
r233 16 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.45 $Y=1.35
+ $X2=4.45 $Y2=1.515
r234 15 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.45 $Y=1.19
+ $X2=4.525 $Y2=1.115
r235 15 16 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.45 $Y=1.19
+ $X2=4.45 $Y2=1.35
r236 11 74 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=1.68
+ $X2=3.96 $Y2=1.515
r237 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.96 $Y=1.68
+ $X2=3.96 $Y2=2.4
r238 7 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.35
+ $X2=3.94 $Y2=1.515
r239 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.94 $Y=1.35 $X2=3.94
+ $Y2=0.74
r240 2 65 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.84 $X2=3.285 $Y2=1.985
r241 1 58 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.08
+ $Y=0.37 $X2=3.225 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_2191_180# 1 2 9 13 14 18 21 23 24 28 33
+ 35 38 41
c96 33 0 1.14206e-19 $X=12.465 $Y=2.815
c97 28 0 1.71901e-19 $X=11.12 $Y=1.065
r98 36 38 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.465 $Y=2.265
+ $X2=12.625 $Y2=2.265
r99 31 33 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.3 $Y=2.815
+ $X2=12.465 $Y2=2.815
r100 28 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.12 $Y=1.065
+ $X2=11.12 $Y2=1.23
r101 28 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.12 $Y=1.065
+ $X2=11.12 $Y2=0.9
r102 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.12
+ $Y=1.065 $X2=11.12 $Y2=1.065
r103 24 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.12 $Y=0.985
+ $X2=11.12 $Y2=1.065
r104 23 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.625 $Y=2.18
+ $X2=12.625 $Y2=2.265
r105 22 35 3.351 $w=2.8e-07 $l=1.46458e-07 $layer=LI1_cond $X=12.625 $Y=1.07
+ $X2=12.515 $Y2=0.985
r106 22 23 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=12.625 $Y=1.07
+ $X2=12.625 $Y2=2.18
r107 21 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=2.65
+ $X2=12.465 $Y2=2.815
r108 20 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.465 $Y=2.35
+ $X2=12.465 $Y2=2.265
r109 20 21 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.465 $Y=2.35
+ $X2=12.465 $Y2=2.65
r110 16 35 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=12.515 $Y=0.9
+ $X2=12.515 $Y2=0.985
r111 16 18 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=12.515 $Y=0.9
+ $X2=12.515 $Y2=0.58
r112 15 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.285 $Y=0.985
+ $X2=11.12 $Y2=0.985
r113 14 35 3.18746 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.32 $Y=0.985
+ $X2=12.515 $Y2=0.985
r114 14 15 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=12.32 $Y=0.985
+ $X2=11.285 $Y2=0.985
r115 13 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.06 $Y=0.58
+ $X2=11.06 $Y2=0.9
r116 9 42 590.839 $w=1.8e-07 $l=1.52e-06 $layer=POLY_cond $X=11.065 $Y=2.75
+ $X2=11.065 $Y2=1.23
r117 2 31 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=12.155
+ $Y=2.54 $X2=12.3 $Y2=2.815
r118 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.345
+ $Y=0.37 $X2=12.485 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_1823_524# 1 2 3 4 5 18 22 24 26 28 31 33
+ 35 42 44 46 47 51 55 56 57 58 59 61 62 66 70 71 74 76 80 82 84
c198 58 0 2.62796e-19 $X=10.935 $Y=1.485
c199 33 0 2.05112e-20 $X=13.48 $Y=2.04
c200 26 0 1.14206e-19 $X=13.03 $Y=2.04
r201 87 88 34.5038 $w=5.75e-07 $l=7.5e-08 $layer=POLY_cond $X=12.327 $Y=1.965
+ $X2=12.327 $Y2=2.04
r202 76 78 7.28509 $w=2.78e-07 $l=1.77e-07 $layer=LI1_cond $X=9.235 $Y=2.79
+ $X2=9.235 $Y2=2.967
r203 74 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.125 $Y=2.31
+ $X2=12.125 $Y2=2.395
r204 74 84 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.125 $Y=2.31
+ $X2=12.125 $Y2=2.01
r205 71 87 42.8024 $w=5.75e-07 $l=4.6e-07 $layer=POLY_cond $X=12.327 $Y=1.505
+ $X2=12.327 $Y2=1.965
r206 71 86 48.7424 $w=5.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.327 $Y=1.505
+ $X2=12.327 $Y2=1.34
r207 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.205
+ $Y=1.505 $X2=12.205 $Y2=1.505
r208 68 84 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.205 $Y=1.845
+ $X2=12.205 $Y2=2.01
r209 68 70 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=12.205 $Y=1.845
+ $X2=12.205 $Y2=1.505
r210 64 82 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.74 $Y=2.395
+ $X2=12.125 $Y2=2.395
r211 64 66 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=11.74 $Y=2.48
+ $X2=11.74 $Y2=2.75
r212 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.105 $Y=2.395
+ $X2=11.02 $Y2=2.395
r213 62 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.575 $Y=2.395
+ $X2=11.74 $Y2=2.395
r214 62 63 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=11.575 $Y=2.395
+ $X2=11.105 $Y2=2.395
r215 61 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.02 $Y=2.31
+ $X2=11.02 $Y2=2.395
r216 60 61 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.02 $Y=1.57
+ $X2=11.02 $Y2=2.31
r217 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.935 $Y=1.485
+ $X2=11.02 $Y2=1.57
r218 58 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.935 $Y=1.485
+ $X2=10.54 $Y2=1.485
r219 56 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.935 $Y=2.395
+ $X2=11.02 $Y2=2.395
r220 56 57 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.935 $Y=2.395
+ $X2=10.375 $Y2=2.395
r221 53 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.375 $Y=1.4
+ $X2=10.54 $Y2=1.485
r222 53 55 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=10.375 $Y=1.4
+ $X2=10.375 $Y2=0.515
r223 52 55 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.375 $Y=0.425
+ $X2=10.375 $Y2=0.515
r224 49 51 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=10.21 $Y=2.86
+ $X2=10.21 $Y2=2.745
r225 48 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.21 $Y=2.48
+ $X2=10.375 $Y2=2.395
r226 48 51 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=10.21 $Y=2.48
+ $X2=10.21 $Y2=2.745
r227 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.21 $Y=0.34
+ $X2=10.375 $Y2=0.425
r228 46 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.21 $Y=0.34
+ $X2=9.68 $Y2=0.34
r229 45 78 2.30834 $w=2.15e-07 $l=1.4e-07 $layer=LI1_cond $X=9.375 $Y=2.967
+ $X2=9.235 $Y2=2.967
r230 44 49 7.21882 $w=2.15e-07 $l=2.11849e-07 $layer=LI1_cond $X=10.045 $Y=2.967
+ $X2=10.21 $Y2=2.86
r231 44 45 35.9133 $w=2.13e-07 $l=6.7e-07 $layer=LI1_cond $X=10.045 $Y=2.967
+ $X2=9.375 $Y2=2.967
r232 40 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.515 $Y=0.425
+ $X2=9.68 $Y2=0.34
r233 40 42 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.515 $Y=0.425
+ $X2=9.515 $Y2=0.515
r234 33 37 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=13.48 $Y=1.965
+ $X2=13.26 $Y2=1.965
r235 33 35 133.889 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=13.48 $Y=2.04
+ $X2=13.48 $Y2=2.54
r236 29 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.26 $Y=1.89
+ $X2=13.26 $Y2=1.965
r237 29 31 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=13.26 $Y=1.89
+ $X2=13.26 $Y2=0.74
r238 26 37 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=13.03 $Y=1.965
+ $X2=13.26 $Y2=1.965
r239 26 28 133.889 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=13.03 $Y=2.04
+ $X2=13.03 $Y2=2.54
r240 25 87 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=12.615 $Y=1.965
+ $X2=12.327 $Y2=1.965
r241 24 26 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.94 $Y=1.965
+ $X2=13.03 $Y2=1.965
r242 24 25 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=12.94 $Y=1.965
+ $X2=12.615 $Y2=1.965
r243 22 88 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=12.525 $Y=2.75
+ $X2=12.525 $Y2=2.04
r244 18 86 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=12.27 $Y=0.58
+ $X2=12.27 $Y2=1.34
r245 5 66 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.605
+ $Y=2.54 $X2=11.74 $Y2=2.75
r246 4 51 600 $w=1.7e-07 $l=7.11512e-07 $layer=licon1_PDIFF $count=1 $X=10.025
+ $Y=2.12 $X2=10.21 $Y2=2.745
r247 3 76 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=9.115
+ $Y=2.62 $X2=9.26 $Y2=2.79
r248 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.235
+ $Y=0.37 $X2=10.375 $Y2=0.515
r249 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.37
+ $Y=0.37 $X2=9.515 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_2580_74# 1 2 9 13 17 21 25 29 31 35 39 41
+ 44 48 55 58 68
c115 41 0 1.68497e-19 $X=15.312 $Y=1.395
c116 35 0 2.40437e-20 $X=15.275 $Y=0.74
c117 25 0 2.92295e-20 $X=14.845 $Y=0.74
r118 67 68 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=14.885 $Y=1.485
+ $X2=14.975 $Y2=1.485
r119 66 67 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=14.845 $Y=1.485
+ $X2=14.885 $Y2=1.485
r120 63 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=14.345 $Y=1.485
+ $X2=14.435 $Y2=1.485
r121 62 63 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=13.985 $Y=1.485
+ $X2=14.345 $Y2=1.485
r122 56 66 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=14.53 $Y=1.485
+ $X2=14.845 $Y2=1.485
r123 56 64 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=14.53 $Y=1.485
+ $X2=14.435 $Y2=1.485
r124 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14.53
+ $Y=1.485 $X2=14.53 $Y2=1.485
r125 53 62 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=13.85 $Y=1.485
+ $X2=13.985 $Y2=1.485
r126 53 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.85 $Y=1.485
+ $X2=13.76 $Y2=1.485
r127 52 55 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.85 $Y=1.485
+ $X2=14.53 $Y2=1.485
r128 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.85
+ $Y=1.485 $X2=13.85 $Y2=1.485
r129 50 58 0.364692 $w=3.3e-07 $l=5.3619e-07 $layer=LI1_cond $X=13.34 $Y=1.485
+ $X2=12.88 $Y2=1.32
r130 50 52 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=13.34 $Y=1.485
+ $X2=13.85 $Y2=1.485
r131 46 58 6.46576 $w=2.5e-07 $l=5.14174e-07 $layer=LI1_cond $X=13.255 $Y=1.65
+ $X2=12.88 $Y2=1.32
r132 46 48 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=13.255 $Y=1.65
+ $X2=13.255 $Y2=2.265
r133 42 58 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=13.045 $Y=1.32
+ $X2=12.88 $Y2=1.32
r134 42 44 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=13.045 $Y=1.32
+ $X2=13.045 $Y2=0.515
r135 37 41 18.8402 $w=1.65e-07 $l=8.57321e-08 $layer=POLY_cond $X=15.335 $Y=1.47
+ $X2=15.312 $Y2=1.395
r136 37 39 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=15.335 $Y=1.47
+ $X2=15.335 $Y2=2.4
r137 33 41 18.8402 $w=1.65e-07 $l=9.16515e-08 $layer=POLY_cond $X=15.275 $Y=1.32
+ $X2=15.312 $Y2=1.395
r138 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=15.275 $Y=1.32
+ $X2=15.275 $Y2=0.74
r139 31 41 6.66866 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=15.2 $Y=1.395
+ $X2=15.312 $Y2=1.395
r140 31 68 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=15.2 $Y=1.395
+ $X2=14.975 $Y2=1.395
r141 27 67 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.885 $Y=1.65
+ $X2=14.885 $Y2=1.485
r142 27 29 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=14.885 $Y=1.65
+ $X2=14.885 $Y2=2.4
r143 23 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.845 $Y=1.32
+ $X2=14.845 $Y2=1.485
r144 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=14.845 $Y=1.32
+ $X2=14.845 $Y2=0.74
r145 19 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.435 $Y=1.65
+ $X2=14.435 $Y2=1.485
r146 19 21 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=14.435 $Y=1.65
+ $X2=14.435 $Y2=2.4
r147 15 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.345 $Y=1.32
+ $X2=14.345 $Y2=1.485
r148 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=14.345 $Y=1.32
+ $X2=14.345 $Y2=0.74
r149 11 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.985 $Y=1.65
+ $X2=13.985 $Y2=1.485
r150 11 13 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=13.985 $Y=1.65
+ $X2=13.985 $Y2=2.4
r151 7 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.76 $Y=1.32
+ $X2=13.76 $Y2=1.485
r152 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=13.76 $Y=1.32
+ $X2=13.76 $Y2=0.74
r153 2 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=13.12
+ $Y=2.12 $X2=13.255 $Y2=2.265
r154 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.9
+ $Y=0.37 $X2=13.045 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 42 46 50
+ 54 58 62 66 70 74 76 78 83 84 86 87 88 90 95 100 115 122 127 132 137 143 146
+ 149 152 155 158 161 164 168
c209 46 0 1.31023e-19 $X=3.735 $Y=2.78
r210 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r211 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r212 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r213 158 159 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r214 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r215 152 153 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r216 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r217 147 150 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r218 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r219 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r220 141 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r221 141 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=14.64 $Y2=3.33
r222 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r223 138 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.825 $Y=3.33
+ $X2=14.66 $Y2=3.33
r224 138 140 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.825 $Y=3.33
+ $X2=15.12 $Y2=3.33
r225 137 167 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.395 $Y=3.33
+ $X2=15.617 $Y2=3.33
r226 137 140 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.395 $Y=3.33
+ $X2=15.12 $Y2=3.33
r227 136 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r228 136 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r229 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r230 133 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.87 $Y=3.33
+ $X2=13.705 $Y2=3.33
r231 133 135 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.87 $Y=3.33
+ $X2=14.16 $Y2=3.33
r232 132 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.66 $Y2=3.33
r233 132 135 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.16 $Y2=3.33
r234 131 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r235 131 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r236 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r237 128 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.97 $Y=3.33
+ $X2=12.845 $Y2=3.33
r238 128 130 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=12.97 $Y=3.33
+ $X2=13.2 $Y2=3.33
r239 127 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.705 $Y2=3.33
r240 127 130 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r241 126 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r242 126 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r243 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r244 123 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.25 $Y2=3.33
r245 123 125 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.76 $Y2=3.33
r246 122 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=12.845 $Y2=3.33
r247 122 125 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r248 121 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r249 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r250 118 121 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r251 117 120 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r252 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r253 115 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.125 $Y=3.33
+ $X2=11.25 $Y2=3.33
r254 115 120 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.125 $Y=3.33
+ $X2=10.8 $Y2=3.33
r255 114 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r256 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r257 111 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r258 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r259 108 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.525 $Y=3.33
+ $X2=6.4 $Y2=3.33
r260 108 110 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=6.525 $Y=3.33
+ $X2=7.44 $Y2=3.33
r261 107 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r262 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r263 104 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r264 104 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r265 103 106 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r266 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r267 101 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=3.33
+ $X2=3.735 $Y2=3.33
r268 101 103 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.9 $Y=3.33
+ $X2=4.08 $Y2=3.33
r269 100 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.4 $Y2=3.33
r270 100 106 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r271 99 147 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r272 99 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r273 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r274 96 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r275 96 98 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r276 95 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.725 $Y2=3.33
r277 95 98 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r278 93 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r279 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r280 90 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r281 90 92 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r282 88 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r283 88 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r284 86 113 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.4 $Y2=3.33
r285 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.7 $Y2=3.33
r286 85 117 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.865 $Y=3.33
+ $X2=8.88 $Y2=3.33
r287 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.865 $Y=3.33
+ $X2=8.7 $Y2=3.33
r288 83 110 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r289 83 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.8 $Y2=3.33
r290 82 113 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=8.4 $Y2=3.33
r291 82 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=7.8 $Y2=3.33
r292 78 81 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=15.56 $Y=2.115
+ $X2=15.56 $Y2=2.815
r293 76 167 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.56 $Y=3.245
+ $X2=15.617 $Y2=3.33
r294 76 81 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.56 $Y=3.245
+ $X2=15.56 $Y2=2.815
r295 72 164 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.66 $Y=3.245
+ $X2=14.66 $Y2=3.33
r296 72 74 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=14.66 $Y=3.245
+ $X2=14.66 $Y2=2.405
r297 68 161 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=3.33
r298 68 70 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=2.265
r299 64 158 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.845 $Y=3.245
+ $X2=12.845 $Y2=3.33
r300 64 66 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=12.845 $Y=3.245
+ $X2=12.845 $Y2=2.75
r301 60 155 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.25 $Y=3.245
+ $X2=11.25 $Y2=3.33
r302 60 62 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.25 $Y=3.245
+ $X2=11.25 $Y2=2.815
r303 56 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.7 $Y=3.245 $X2=8.7
+ $Y2=3.33
r304 56 58 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.7 $Y=3.245
+ $X2=8.7 $Y2=2.55
r305 52 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.8 $Y=3.245 $X2=7.8
+ $Y2=3.33
r306 52 54 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.8 $Y=3.245
+ $X2=7.8 $Y2=2.505
r307 48 152 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=3.245
+ $X2=6.4 $Y2=3.33
r308 48 50 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=6.4 $Y=3.245 $X2=6.4
+ $Y2=2.795
r309 44 149 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=3.245
+ $X2=3.735 $Y2=3.33
r310 44 46 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.735 $Y=3.245
+ $X2=3.735 $Y2=2.78
r311 43 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.725 $Y2=3.33
r312 42 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=3.33
+ $X2=3.735 $Y2=3.33
r313 42 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.57 $Y=3.33
+ $X2=2.89 $Y2=3.33
r314 38 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r315 38 40 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.995
r316 34 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r317 34 36 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.78
r318 11 81 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=15.425
+ $Y=1.84 $X2=15.56 $Y2=2.815
r319 11 78 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=15.425
+ $Y=1.84 $X2=15.56 $Y2=2.115
r320 10 74 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=14.525
+ $Y=1.84 $X2=14.66 $Y2=2.405
r321 9 70 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=13.57
+ $Y=2.12 $X2=13.705 $Y2=2.265
r322 8 66 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=12.615
+ $Y=2.54 $X2=12.805 $Y2=2.75
r323 7 62 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=11.155
+ $Y=2.54 $X2=11.29 $Y2=2.815
r324 6 58 600 $w=1.7e-07 $l=7.49466e-07 $layer=licon1_PDIFF $count=1 $X=8.565
+ $Y=1.865 $X2=8.7 $Y2=2.55
r325 5 54 600 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_PDIFF $count=1 $X=7.435
+ $Y=2.285 $X2=7.8 $Y2=2.505
r326 4 50 600 $w=1.7e-07 $l=6.10164e-07 $layer=licon1_PDIFF $count=1 $X=6.22
+ $Y=2.285 $X2=6.44 $Y2=2.795
r327 3 46 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=3.6
+ $Y=1.84 $X2=3.735 $Y2=2.78
r328 2 40 600 $w=1.7e-07 $l=7.77255e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=2.32 $X2=2.725 $Y2=2.995
r329 1 36 600 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.32 $X2=0.72 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_291_464# 1 2 3 4 13 18 19 20 22 23 25 28
+ 32 34 37 44 46
c126 22 0 4.43302e-20 $X=2.3 $Y=2.49
r127 46 48 4.07466 $w=5.09e-07 $l=1.7e-07 $layer=LI1_cond $X=4.72 $Y=2.325
+ $X2=4.72 $Y2=2.495
r128 41 44 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.495 $Y=0.76
+ $X2=4.715 $Y2=0.76
r129 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.09 $Y=2.325
+ $X2=3.09 $Y2=2.575
r130 30 32 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.715 $Y=0.575
+ $X2=1.875 $Y2=0.575
r131 28 46 15.9959 $w=5.09e-07 $l=5.25595e-07 $layer=LI1_cond $X=4.495 $Y=1.9
+ $X2=4.72 $Y2=2.325
r132 27 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.925
+ $X2=4.495 $Y2=0.76
r133 27 28 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=4.495 $Y=0.925
+ $X2=4.495 $Y2=1.9
r134 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.175 $Y=2.325
+ $X2=3.09 $Y2=2.325
r135 25 46 7.26882 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.41 $Y=2.325
+ $X2=4.72 $Y2=2.325
r136 25 26 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.41 $Y=2.325
+ $X2=3.175 $Y2=2.325
r137 24 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.575
+ $X2=2.3 $Y2=2.575
r138 23 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=2.575
+ $X2=3.09 $Y2=2.575
r139 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.005 $Y=2.575
+ $X2=2.385 $Y2=2.575
r140 22 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.575
r141 21 22 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.3 $Y=1.08
+ $X2=2.3 $Y2=2.49
r142 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=2.3 $Y2=1.08
r143 19 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=1.96 $Y2=0.995
r144 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.875 $Y=0.91
+ $X2=1.96 $Y2=0.995
r145 17 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.875 $Y2=0.575
r146 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.875 $Y2=0.91
r147 13 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.3 $Y=2.785
+ $X2=2.3 $Y2=2.575
r148 13 15 24.6623 $w=2.48e-07 $l=5.35e-07 $layer=LI1_cond $X=2.215 $Y=2.785
+ $X2=1.68 $Y2=2.785
r149 4 48 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=2.285 $X2=4.865 $Y2=2.495
r150 3 15 600 $w=1.7e-07 $l=5.25595e-07 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=2.32 $X2=1.68 $Y2=2.745
r151 2 44 182 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.405 $X2=4.715 $Y2=0.76
r152 1 30 182 $w=1.7e-07 $l=3.005e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.715 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_1623_373# 1 2 7 9 11 18
c33 9 0 7.59542e-20 $X=8.25 $Y=2.55
c34 7 0 1.49331e-19 $X=8.225 $Y=2.29
r35 12 16 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.365 $Y=2.205
+ $X2=8.225 $Y2=2.205
r36 11 18 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=9.545 $Y=2.205
+ $X2=9.71 $Y2=2.195
r37 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=9.545 $Y=2.205
+ $X2=8.365 $Y2=2.205
r38 7 16 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.225 $Y=2.29
+ $X2=8.225 $Y2=2.205
r39 7 9 10.7013 $w=2.78e-07 $l=2.6e-07 $layer=LI1_cond $X=8.225 $Y=2.29
+ $X2=8.225 $Y2=2.55
r40 2 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=2.12 $X2=9.71 $Y2=2.265
r41 1 16 600 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=1 $X=8.115
+ $Y=1.865 $X2=8.25 $Y2=2.205
r42 1 9 600 $w=1.7e-07 $l=7.49466e-07 $layer=licon1_PDIFF $count=1 $X=8.115
+ $Y=1.865 $X2=8.25 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 31 33 35 39
+ 43 45 48
c80 35 0 2.92295e-20 $X=15.485 $Y=1.355
c81 21 0 2.40437e-20 $X=14.895 $Y=1.065
c82 17 0 2.05112e-20 $X=14.185 $Y=2.15
r83 45 48 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.6 $Y=1.695 $X2=15.6
+ $Y2=1.61
r84 45 48 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=15.6 $Y=1.595
+ $X2=15.6 $Y2=1.61
r85 44 45 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=15.6 $Y=1.44
+ $X2=15.6 $Y2=1.595
r86 39 40 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=15.06 $Y=1.065
+ $X2=15.06 $Y2=1.355
r87 36 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.225 $Y=1.355
+ $X2=15.06 $Y2=1.355
r88 35 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=15.485 $Y=1.355
+ $X2=15.6 $Y2=1.44
r89 35 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=15.485 $Y=1.355
+ $X2=15.225 $Y2=1.355
r90 34 43 3.70735 $w=2.5e-07 $l=2.23495e-07 $layer=LI1_cond $X=15.195 $Y=1.695
+ $X2=15.11 $Y2=1.88
r91 33 45 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=15.485 $Y=1.695
+ $X2=15.6 $Y2=1.695
r92 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=15.485 $Y=1.695
+ $X2=15.195 $Y2=1.695
r93 29 43 2.76166 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=15.11 $Y=2.15
+ $X2=15.11 $Y2=1.88
r94 29 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=15.11 $Y=2.15
+ $X2=15.11 $Y2=2.4
r95 25 39 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=15.06 $Y=0.98
+ $X2=15.06 $Y2=1.065
r96 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=15.06 $Y=0.98
+ $X2=15.06 $Y2=0.515
r97 24 38 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=14.325 $Y=1.985
+ $X2=14.185 $Y2=1.985
r98 23 43 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=15.025 $Y=1.985
+ $X2=15.11 $Y2=1.88
r99 23 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=15.025 $Y=1.985
+ $X2=14.325 $Y2=1.985
r100 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.895 $Y=1.065
+ $X2=15.06 $Y2=1.065
r101 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.895 $Y=1.065
+ $X2=14.225 $Y2=1.065
r102 17 38 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.185 $Y=2.15
+ $X2=14.185 $Y2=1.985
r103 17 19 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=14.185 $Y=2.15
+ $X2=14.185 $Y2=2.4
r104 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.06 $Y=0.98
+ $X2=14.225 $Y2=1.065
r105 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=14.06 $Y=0.98
+ $X2=14.06 $Y2=0.515
r106 4 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.975
+ $Y=1.84 $X2=15.11 $Y2=1.985
r107 4 31 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=14.975
+ $Y=1.84 $X2=15.11 $Y2=2.4
r108 3 38 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.075
+ $Y=1.84 $X2=14.21 $Y2=1.985
r109 3 19 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=14.075
+ $Y=1.84 $X2=14.21 $Y2=2.4
r110 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.92
+ $Y=0.37 $X2=15.06 $Y2=0.515
r111 1 15 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=13.835
+ $Y=0.37 $X2=14.06 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%VGND 1 2 3 4 5 6 7 8 9 10 33 37 39 43 47 51
+ 57 61 65 69 71 73 76 77 78 80 85 93 101 106 111 126 130 136 139 142 145 148
+ 151 154 157 161
c176 73 0 1.68497e-19 $X=15.56 $Y=0.515
r177 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r178 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r179 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r180 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r181 145 146 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r182 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r183 140 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r184 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r185 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r186 134 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=15.6 $Y2=0
r187 134 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=14.64 $Y2=0
r188 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r189 131 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.725 $Y=0
+ $X2=14.56 $Y2=0
r190 131 133 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=14.725 $Y=0
+ $X2=15.12 $Y2=0
r191 130 160 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.395 $Y=0
+ $X2=15.617 $Y2=0
r192 130 133 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.395 $Y=0
+ $X2=15.12 $Y2=0
r193 129 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r194 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r195 126 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.395 $Y=0
+ $X2=14.56 $Y2=0
r196 126 128 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=14.395 $Y=0
+ $X2=14.16 $Y2=0
r197 125 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r198 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r199 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r200 122 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r201 121 124 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r202 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r203 119 154 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=12.15 $Y=0
+ $X2=11.9 $Y2=0
r204 119 121 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=12.15 $Y=0
+ $X2=12.24 $Y2=0
r205 118 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r206 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r207 115 118 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r208 115 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r209 114 117 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r210 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r211 112 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.12 $Y=0
+ $X2=8.955 $Y2=0
r212 112 114 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.12 $Y=0
+ $X2=9.36 $Y2=0
r213 111 154 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.9 $Y2=0
r214 111 117 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.28 $Y2=0
r215 110 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r216 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r217 107 148 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.26 $Y=0
+ $X2=7.925 $Y2=0
r218 107 109 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.26 $Y=0 $X2=8.4
+ $Y2=0
r219 106 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.79 $Y=0
+ $X2=8.955 $Y2=0
r220 106 109 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.79 $Y=0 $X2=8.4
+ $Y2=0
r221 105 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.48 $Y2=0
r222 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r223 102 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.54 $Y=0
+ $X2=6.375 $Y2=0
r224 102 104 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=6.54 $Y=0 $X2=7.44
+ $Y2=0
r225 101 148 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=7.925 $Y2=0
r226 101 104 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.59 $Y=0 $X2=7.44
+ $Y2=0
r227 100 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r228 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r229 97 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r230 97 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r231 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r232 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r233 94 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0
+ $X2=3.725 $Y2=0
r234 94 96 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.08
+ $Y2=0
r235 93 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=6.375 $Y2=0
r236 93 99 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.21 $Y=0 $X2=6
+ $Y2=0
r237 92 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r238 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r239 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r240 89 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r241 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r242 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r243 86 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.78 $Y2=0
r244 86 88 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r245 85 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0
+ $X2=2.615 $Y2=0
r246 85 91 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.16
+ $Y2=0
r247 83 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r248 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r249 80 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.78 $Y2=0
r250 80 82 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r251 78 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r252 78 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r253 78 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r254 76 124 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=13.38 $Y=0
+ $X2=13.2 $Y2=0
r255 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.38 $Y=0
+ $X2=13.545 $Y2=0
r256 75 128 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=13.71 $Y=0
+ $X2=14.16 $Y2=0
r257 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.71 $Y=0
+ $X2=13.545 $Y2=0
r258 71 160 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.56 $Y=0.085
+ $X2=15.617 $Y2=0
r259 71 73 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.56 $Y=0.085
+ $X2=15.56 $Y2=0.515
r260 67 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.56 $Y=0.085
+ $X2=14.56 $Y2=0
r261 67 69 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=14.56 $Y=0.085
+ $X2=14.56 $Y2=0.645
r262 63 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.545 $Y=0.085
+ $X2=13.545 $Y2=0
r263 63 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.545 $Y=0.085
+ $X2=13.545 $Y2=0.515
r264 59 154 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.9 $Y=0.085
+ $X2=11.9 $Y2=0
r265 59 61 10.2863 $w=4.98e-07 $l=4.3e-07 $layer=LI1_cond $X=11.9 $Y=0.085
+ $X2=11.9 $Y2=0.515
r266 55 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=0.085
+ $X2=8.955 $Y2=0
r267 55 57 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.955 $Y=0.085
+ $X2=8.955 $Y2=0.515
r268 51 53 6.06965 $w=6.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.925 $Y=0.495
+ $X2=7.925 $Y2=0.835
r269 49 148 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.925 $Y=0.085
+ $X2=7.925 $Y2=0
r270 49 51 7.31929 $w=6.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.925 $Y=0.085
+ $X2=7.925 $Y2=0.495
r271 45 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0
r272 45 47 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0.395
r273 41 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0
r274 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0.515
r275 40 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0
+ $X2=2.615 $Y2=0
r276 39 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=0
+ $X2=3.725 $Y2=0
r277 39 40 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=2.78
+ $Y2=0
r278 35 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0
r279 35 37 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.545
r280 31 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r281 31 33 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.545
r282 10 73 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=15.35
+ $Y=0.37 $X2=15.56 $Y2=0.515
r283 9 69 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=14.42
+ $Y=0.37 $X2=14.56 $Y2=0.645
r284 8 65 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=13.335
+ $Y=0.37 $X2=13.545 $Y2=0.515
r285 7 61 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=11.675
+ $Y=0.37 $X2=11.9 $Y2=0.515
r286 6 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.815
+ $Y=0.37 $X2=8.955 $Y2=0.515
r287 5 53 121.333 $w=1.7e-07 $l=6.73498e-07 $layer=licon1_NDIFF $count=1
+ $X=7.615 $Y=0.37 $X2=8.095 $Y2=0.835
r288 5 51 121.333 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=1
+ $X=7.615 $Y=0.37 $X2=8.095 $Y2=0.495
r289 4 47 182 $w=1.7e-07 $l=2.24944e-07 $layer=licon1_NDIFF $count=1 $X=6.155
+ $Y=0.405 $X2=6.375 $Y2=0.395
r290 3 43 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.515
+ $Y=0.37 $X2=3.725 $Y2=0.515
r291 2 37 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.37 $X2=2.615 $Y2=0.545
r292 1 33 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_4%A_1677_74# 1 2 9 11 12 15
c36 9 0 1.22616e-19 $X=8.525 $Y=0.515
r37 13 15 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.945 $Y=1.11
+ $X2=9.945 $Y2=0.81
r38 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.86 $Y=1.195
+ $X2=9.945 $Y2=1.11
r39 11 12 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=9.86 $Y=1.195
+ $X2=8.61 $Y2=1.195
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.525 $Y=1.11
+ $X2=8.61 $Y2=1.195
r41 7 9 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=8.525 $Y=1.11
+ $X2=8.525 $Y2=0.515
r42 2 15 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=9.805
+ $Y=0.37 $X2=9.945 $Y2=0.81
r43 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.385
+ $Y=0.37 $X2=8.525 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__a32o_4.pxi.spice
* Created: Wed Sep  2 11:55:53 2020
* 
x_PM_SKY130_FD_SC_MS__A32O_4%A_83_283# N_A_83_283#_M1001_d N_A_83_283#_M1025_d
+ N_A_83_283#_M1015_s N_A_83_283#_M1019_s N_A_83_283#_M1003_g
+ N_A_83_283#_c_149_n N_A_83_283#_M1007_g N_A_83_283#_c_150_n
+ N_A_83_283#_M1008_g N_A_83_283#_M1004_g N_A_83_283#_M1005_g
+ N_A_83_283#_M1014_g N_A_83_283#_M1006_g N_A_83_283#_M1023_g
+ N_A_83_283#_c_153_n N_A_83_283#_c_164_n N_A_83_283#_c_165_n
+ N_A_83_283#_c_230_p N_A_83_283#_c_166_n N_A_83_283#_c_154_n
+ N_A_83_283#_c_155_n N_A_83_283#_c_156_n N_A_83_283#_c_168_n
+ N_A_83_283#_c_169_n N_A_83_283#_c_157_n N_A_83_283#_c_158_n
+ PM_SKY130_FD_SC_MS__A32O_4%A_83_283#
x_PM_SKY130_FD_SC_MS__A32O_4%B2 N_B2_M1000_g N_B2_M1015_g N_B2_c_326_n
+ N_B2_M1022_g N_B2_c_340_n N_B2_M1020_g N_B2_c_327_n N_B2_c_328_n N_B2_c_329_n
+ N_B2_c_330_n N_B2_c_331_n N_B2_c_332_n N_B2_c_333_n N_B2_c_334_n B2
+ N_B2_c_336_n N_B2_c_337_n N_B2_c_338_n PM_SKY130_FD_SC_MS__A32O_4%B2
x_PM_SKY130_FD_SC_MS__A32O_4%B1 N_B1_M1001_g N_B1_c_436_n N_B1_M1018_g
+ N_B1_c_433_n N_B1_M1021_g N_B1_c_437_n N_B1_M1019_g B1 B1 N_B1_c_435_n
+ PM_SKY130_FD_SC_MS__A32O_4%B1
x_PM_SKY130_FD_SC_MS__A32O_4%A2 N_A2_M1010_g N_A2_M1009_g N_A2_M1024_g
+ N_A2_M1011_g N_A2_c_490_n N_A2_c_497_n N_A2_c_498_n N_A2_c_552_p N_A2_c_499_n
+ N_A2_c_491_n N_A2_c_492_n N_A2_c_493_n A2 N_A2_c_494_n
+ PM_SKY130_FD_SC_MS__A32O_4%A2
x_PM_SKY130_FD_SC_MS__A32O_4%A1 N_A1_M1016_g N_A1_M1025_g N_A1_M1026_g
+ N_A1_M1027_g A1 N_A1_c_599_n PM_SKY130_FD_SC_MS__A32O_4%A1
x_PM_SKY130_FD_SC_MS__A32O_4%A3 N_A3_M1002_g N_A3_M1013_g N_A3_M1017_g
+ N_A3_M1012_g A3 A3 N_A3_c_652_n PM_SKY130_FD_SC_MS__A32O_4%A3
x_PM_SKY130_FD_SC_MS__A32O_4%VPWR N_VPWR_M1003_s N_VPWR_M1004_s N_VPWR_M1006_s
+ N_VPWR_M1010_d N_VPWR_M1027_s N_VPWR_M1013_s N_VPWR_c_700_n N_VPWR_c_701_n
+ N_VPWR_c_702_n N_VPWR_c_703_n N_VPWR_c_704_n N_VPWR_c_705_n N_VPWR_c_706_n
+ VPWR N_VPWR_c_707_n N_VPWR_c_708_n N_VPWR_c_709_n N_VPWR_c_710_n
+ N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_699_n N_VPWR_c_714_n N_VPWR_c_715_n
+ N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_718_n PM_SKY130_FD_SC_MS__A32O_4%VPWR
x_PM_SKY130_FD_SC_MS__A32O_4%X N_X_M1007_d N_X_M1014_d N_X_M1003_d N_X_M1005_d
+ N_X_c_819_n N_X_c_810_n N_X_c_811_n N_X_c_812_n N_X_c_816_n N_X_c_817_n
+ N_X_c_813_n N_X_c_830_n N_X_c_834_n N_X_c_839_n N_X_c_818_n N_X_c_814_n
+ N_X_c_848_n N_X_c_849_n X PM_SKY130_FD_SC_MS__A32O_4%X
x_PM_SKY130_FD_SC_MS__A32O_4%A_509_392# N_A_509_392#_M1015_d
+ N_A_509_392#_M1018_d N_A_509_392#_M1020_d N_A_509_392#_M1016_d
+ N_A_509_392#_M1011_s N_A_509_392#_M1017_d N_A_509_392#_c_879_n
+ N_A_509_392#_c_880_n N_A_509_392#_c_881_n N_A_509_392#_c_897_n
+ N_A_509_392#_c_882_n N_A_509_392#_c_915_n N_A_509_392#_c_920_n
+ N_A_509_392#_c_883_n N_A_509_392#_c_928_n N_A_509_392#_c_884_n
+ N_A_509_392#_c_885_n N_A_509_392#_c_886_n N_A_509_392#_c_887_n
+ N_A_509_392#_c_888_n N_A_509_392#_c_889_n N_A_509_392#_c_933_n
+ N_A_509_392#_c_936_n PM_SKY130_FD_SC_MS__A32O_4%A_509_392#
x_PM_SKY130_FD_SC_MS__A32O_4%VGND N_VGND_M1007_s N_VGND_M1008_s N_VGND_M1023_s
+ N_VGND_M1022_s N_VGND_M1002_s N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n
+ N_VGND_c_989_n N_VGND_c_990_n N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n
+ VGND N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n
+ N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n
+ PM_SKY130_FD_SC_MS__A32O_4%VGND
x_PM_SKY130_FD_SC_MS__A32O_4%A_587_110# N_A_587_110#_M1000_d
+ N_A_587_110#_M1021_s N_A_587_110#_c_1079_n N_A_587_110#_c_1075_n
+ PM_SKY130_FD_SC_MS__A32O_4%A_587_110#
x_PM_SKY130_FD_SC_MS__A32O_4%A_992_122# N_A_992_122#_M1009_d
+ N_A_992_122#_M1024_d N_A_992_122#_M1012_d N_A_992_122#_c_1098_n
+ N_A_992_122#_c_1099_n N_A_992_122#_c_1100_n N_A_992_122#_c_1101_n
+ N_A_992_122#_c_1102_n N_A_992_122#_c_1103_n N_A_992_122#_c_1104_n
+ PM_SKY130_FD_SC_MS__A32O_4%A_992_122#
x_PM_SKY130_FD_SC_MS__A32O_4%A_1079_122# N_A_1079_122#_M1009_s
+ N_A_1079_122#_M1026_s N_A_1079_122#_c_1146_n N_A_1079_122#_c_1147_n
+ N_A_1079_122#_c_1148_n PM_SKY130_FD_SC_MS__A32O_4%A_1079_122#
cc_1 VNB N_A_83_283#_c_149_n 0.0162789f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.265
cc_2 VNB N_A_83_283#_c_150_n 0.0150928f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.265
cc_3 VNB N_A_83_283#_M1014_g 0.0202081f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.82
cc_4 VNB N_A_83_283#_M1023_g 0.0210256f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.82
cc_5 VNB N_A_83_283#_c_153_n 0.00571863f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.515
cc_6 VNB N_A_83_283#_c_154_n 0.00711934f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=1.95
cc_7 VNB N_A_83_283#_c_155_n 0.0111495f $X=-0.19 $Y=-0.245 $X2=5.8 $Y2=1.195
cc_8 VNB N_A_83_283#_c_156_n 0.00111139f $X=-0.19 $Y=-0.245 $X2=4.055 $Y2=1.195
cc_9 VNB N_A_83_283#_c_157_n 0.00227768f $X=-0.19 $Y=-0.245 $X2=5.965 $Y2=1.1
cc_10 VNB N_A_83_283#_c_158_n 0.0901281f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.472
cc_11 VNB N_B2_M1000_g 0.025871f $X=-0.19 $Y=-0.245 $X2=3.005 $Y2=1.96
cc_12 VNB N_B2_c_326_n 0.018238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B2_c_327_n 0.0291913f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_B2_c_328_n 0.0271649f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.82
cc_15 VNB N_B2_c_329_n 0.028259f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.265
cc_16 VNB N_B2_c_330_n 0.0150968f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_17 VNB N_B2_c_331_n 0.014764f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.68
cc_18 VNB N_B2_c_332_n 0.0237932f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.35
cc_19 VNB N_B2_c_333_n 0.0028535f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.82
cc_20 VNB N_B2_c_334_n 0.0031746f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.82
cc_21 VNB B2 0.00406528f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.35
cc_22 VNB N_B2_c_336_n 0.0291119f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.515
cc_23 VNB N_B2_c_337_n 0.0375518f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.68
cc_24 VNB N_B2_c_338_n 0.00800773f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=2.035
cc_25 VNB N_B1_M1001_g 0.0269902f $X=-0.19 $Y=-0.245 $X2=3.005 $Y2=1.96
cc_26 VNB N_B1_c_433_n 0.0173453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB B1 0.00445875f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB N_B1_c_435_n 0.0449866f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_29 VNB N_A2_M1009_g 0.0238027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_M1024_g 0.0213634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_490_n 6.33868e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.265
cc_32 VNB N_A2_c_491_n 0.0062281f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_33 VNB N_A2_c_492_n 0.00386552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_493_n 0.0183892f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.35
cc_35 VNB N_A2_c_494_n 0.0192509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A1_M1025_g 0.0204951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A1_M1026_g 0.0215724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB A1 0.00164534f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.265
cc_39 VNB N_A1_c_599_n 0.0250312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A3_M1002_g 0.0223605f $X=-0.19 $Y=-0.245 $X2=3.005 $Y2=1.96
cc_41 VNB N_A3_M1012_g 0.0313057f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_42 VNB A3 0.0123861f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.82
cc_43 VNB N_A3_c_652_n 0.0317816f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_44 VNB N_VPWR_c_699_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.472
cc_45 VNB N_X_c_810_n 0.0103681f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_46 VNB N_X_c_811_n 0.00236302f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_47 VNB N_X_c_812_n 0.00978528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_X_c_813_n 0.00265478f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_49 VNB N_X_c_814_n 0.00274556f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=2.4
cc_50 VNB X 0.0145337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_986_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_987_n 0.0263097f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.82
cc_53 VNB N_VGND_c_988_n 0.00908353f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.82
cc_54 VNB N_VGND_c_989_n 0.0133287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_990_n 0.0104913f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_56 VNB N_VGND_c_991_n 0.0211664f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.82
cc_57 VNB N_VGND_c_992_n 0.051306f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.82
cc_58 VNB N_VGND_c_993_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.82
cc_59 VNB N_VGND_c_994_n 0.0158697f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.515
cc_60 VNB N_VGND_c_995_n 0.0190672f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.515
cc_61 VNB N_VGND_c_996_n 0.0581589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_997_n 0.0201171f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=2.035
cc_63 VNB N_VGND_c_998_n 0.469086f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=2.115
cc_64 VNB N_VGND_c_999_n 0.00788625f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.472
cc_65 VNB N_VGND_c_1000_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.472
cc_66 VNB N_VGND_c_1001_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.472
cc_67 VNB N_A_587_110#_c_1075_n 0.00306396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_992_122#_c_1098_n 0.00828124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_992_122#_c_1099_n 0.0393952f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_70 VNB N_A_992_122#_c_1100_n 0.00467155f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_71 VNB N_A_992_122#_c_1101_n 0.00357252f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.82
cc_72 VNB N_A_992_122#_c_1102_n 0.0152974f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.265
cc_73 VNB N_A_992_122#_c_1103_n 0.00325088f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.82
cc_74 VNB N_A_992_122#_c_1104_n 0.0231985f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_75 VNB N_A_1079_122#_c_1146_n 0.00318029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1079_122#_c_1147_n 0.00185919f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.68
cc_77 VNB N_A_1079_122#_c_1148_n 0.00820929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VPB N_A_83_283#_M1003_g 0.02574f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_79 VPB N_A_83_283#_M1004_g 0.021252f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_80 VPB N_A_83_283#_M1005_g 0.0217904f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_81 VPB N_A_83_283#_M1006_g 0.0238741f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=2.4
cc_82 VPB N_A_83_283#_c_153_n 4.74324e-19 $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.515
cc_83 VPB N_A_83_283#_c_164_n 0.00314662f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.95
cc_84 VPB N_A_83_283#_c_165_n 0.0199466f $X=-0.19 $Y=1.66 $X2=3.025 $Y2=2.035
cc_85 VPB N_A_83_283#_c_166_n 0.00306854f $X=-0.19 $Y=1.66 $X2=3.885 $Y2=2.035
cc_86 VPB N_A_83_283#_c_154_n 0.00173705f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.95
cc_87 VPB N_A_83_283#_c_168_n 0.00252767f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=2.115
cc_88 VPB N_A_83_283#_c_169_n 0.00344672f $X=-0.19 $Y=1.66 $X2=4.19 $Y2=2.115
cc_89 VPB N_A_83_283#_c_158_n 0.0130754f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.472
cc_90 VPB N_B2_M1015_g 0.026911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_B2_c_340_n 0.0201591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_B2_c_330_n 0.0153061f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_93 VPB B2 0.00297837f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.35
cc_94 VPB N_B2_c_336_n 0.0205201f $X=-0.19 $Y=1.66 $X2=1.15 $Y2=1.515
cc_95 VPB N_B1_c_436_n 0.0184998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_B1_c_437_n 0.0179606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB B1 9.67622e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_98 VPB N_B1_c_435_n 0.0116253f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_99 VPB N_A2_M1010_g 0.0247876f $X=-0.19 $Y=1.66 $X2=3.005 $Y2=1.96
cc_100 VPB N_A2_M1011_g 0.0237945f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_101 VPB N_A2_c_497_n 0.00156767f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.82
cc_102 VPB N_A2_c_498_n 0.0116484f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.82
cc_103 VPB N_A2_c_499_n 0.00346252f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.82
cc_104 VPB N_A2_c_491_n 0.00273065f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_105 VPB N_A2_c_492_n 0.00176577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A2_c_493_n 0.0104366f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.35
cc_107 VPB N_A2_c_494_n 0.0151783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A1_M1016_g 0.0246227f $X=-0.19 $Y=1.66 $X2=3.005 $Y2=1.96
cc_109 VPB N_A1_M1027_g 0.023717f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_110 VPB A1 8.93752e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.265
cc_111 VPB N_A1_c_599_n 0.0143889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A3_M1013_g 0.0232436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A3_M1017_g 0.0318882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB A3 0.00792154f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.82
cc_115 VPB N_A3_c_652_n 0.0193992f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_116 VPB N_VPWR_c_700_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.82
cc_117 VPB N_VPWR_c_701_n 0.0563241f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.82
cc_118 VPB N_VPWR_c_702_n 0.00493781f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.68
cc_119 VPB N_VPWR_c_703_n 0.0118381f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.35
cc_120 VPB N_VPWR_c_704_n 0.00967519f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.68
cc_121 VPB N_VPWR_c_705_n 0.00543991f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.35
cc_122 VPB N_VPWR_c_706_n 0.00830039f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.515
cc_123 VPB N_VPWR_c_707_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_708_n 0.0172495f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.95
cc_125 VPB N_VPWR_c_709_n 0.0695125f $X=-0.19 $Y=1.66 $X2=3.885 $Y2=2.035
cc_126 VPB N_VPWR_c_710_n 0.0190672f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=2.035
cc_127 VPB N_VPWR_c_711_n 0.0172495f $X=-0.19 $Y=1.66 $X2=4.12 $Y2=2.035
cc_128 VPB N_VPWR_c_712_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.472
cc_129 VPB N_VPWR_c_699_n 0.0908165f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.472
cc_130 VPB N_VPWR_c_714_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.472
cc_131 VPB N_VPWR_c_715_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_716_n 0.00776418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_717_n 0.00670444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_718_n 0.00535984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_X_c_816_n 0.00151227f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.82
cc_136 VPB N_X_c_817_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.82
cc_137 VPB N_X_c_818_n 0.0023803f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.82
cc_138 VPB N_A_509_392#_c_879_n 0.00556001f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.82
cc_139 VPB N_A_509_392#_c_880_n 0.00241371f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_140 VPB N_A_509_392#_c_881_n 0.00413156f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_141 VPB N_A_509_392#_c_882_n 0.00715159f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_142 VPB N_A_509_392#_c_883_n 0.00612471f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.35
cc_143 VPB N_A_509_392#_c_884_n 0.0023803f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.515
cc_144 VPB N_A_509_392#_c_885_n 0.00249468f $X=-0.19 $Y=1.66 $X2=1.15 $Y2=1.515
cc_145 VPB N_A_509_392#_c_886_n 0.0097335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_509_392#_c_887_n 0.0352562f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.515
cc_147 VPB N_A_509_392#_c_888_n 0.0021839f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.68
cc_148 VPB N_A_509_392#_c_889_n 0.00245421f $X=-0.19 $Y=1.66 $X2=3.025 $Y2=2.035
cc_149 N_A_83_283#_c_164_n N_B2_M1015_g 0.003634f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_150 N_A_83_283#_c_165_n N_B2_M1015_g 0.0215484f $X=3.025 $Y=2.035 $X2=0 $Y2=0
cc_151 N_A_83_283#_c_154_n N_B2_c_326_n 0.00415276f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_152 N_A_83_283#_c_155_n N_B2_c_326_n 0.0133537f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_153 N_A_83_283#_c_169_n N_B2_c_326_n 0.00347275f $X=4.19 $Y=2.115 $X2=0 $Y2=0
cc_154 N_A_83_283#_c_169_n N_B2_c_340_n 0.0128864f $X=4.19 $Y=2.115 $X2=0 $Y2=0
cc_155 N_A_83_283#_c_154_n N_B2_c_328_n 0.00147539f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_83_283#_c_155_n N_B2_c_328_n 0.00430946f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_157 N_A_83_283#_c_154_n N_B2_c_330_n 0.00371436f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_158 N_A_83_283#_c_155_n N_B2_c_330_n 0.00394231f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_159 N_A_83_283#_c_155_n N_B2_c_331_n 0.0141855f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_160 N_A_83_283#_c_155_n N_B2_c_334_n 0.00422907f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_161 N_A_83_283#_c_153_n B2 0.0121195f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A_83_283#_c_164_n B2 0.00466494f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_163 N_A_83_283#_c_165_n B2 0.0254853f $X=3.025 $Y=2.035 $X2=0 $Y2=0
cc_164 N_A_83_283#_c_158_n B2 2.64894e-19 $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_165 N_A_83_283#_c_153_n N_B2_c_336_n 0.00221274f $X=2.015 $Y=1.515 $X2=0
+ $Y2=0
cc_166 N_A_83_283#_c_164_n N_B2_c_336_n 8.49292e-19 $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_83_283#_c_165_n N_B2_c_336_n 0.00224502f $X=3.025 $Y=2.035 $X2=0
+ $Y2=0
cc_168 N_A_83_283#_c_158_n N_B2_c_336_n 0.00615543f $X=1.905 $Y=1.472 $X2=0
+ $Y2=0
cc_169 N_A_83_283#_M1023_g N_B2_c_338_n 0.00475662f $X=1.95 $Y=0.82 $X2=0 $Y2=0
cc_170 N_A_83_283#_c_153_n N_B2_c_338_n 0.00476787f $X=2.015 $Y=1.515 $X2=0
+ $Y2=0
cc_171 N_A_83_283#_c_158_n N_B2_c_338_n 4.38111e-19 $X=1.905 $Y=1.472 $X2=0
+ $Y2=0
cc_172 N_A_83_283#_c_156_n N_B1_M1001_g 0.00296691f $X=4.055 $Y=1.195 $X2=0
+ $Y2=0
cc_173 N_A_83_283#_c_166_n N_B1_c_436_n 0.0132272f $X=3.885 $Y=2.035 $X2=0 $Y2=0
cc_174 N_A_83_283#_c_154_n N_B1_c_436_n 5.19647e-19 $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_175 N_A_83_283#_c_168_n N_B1_c_436_n 0.0111054f $X=3.19 $Y=2.115 $X2=0 $Y2=0
cc_176 N_A_83_283#_c_154_n N_B1_c_433_n 0.0106813f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_177 N_A_83_283#_c_156_n N_B1_c_433_n 0.0109713f $X=4.055 $Y=1.195 $X2=0 $Y2=0
cc_178 N_A_83_283#_c_166_n N_B1_c_437_n 0.00652003f $X=3.885 $Y=2.035 $X2=0
+ $Y2=0
cc_179 N_A_83_283#_c_154_n N_B1_c_437_n 0.00287293f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_180 N_A_83_283#_c_168_n N_B1_c_437_n 4.55692e-19 $X=3.19 $Y=2.115 $X2=0 $Y2=0
cc_181 N_A_83_283#_c_169_n N_B1_c_437_n 0.00814929f $X=4.19 $Y=2.115 $X2=0 $Y2=0
cc_182 N_A_83_283#_c_165_n B1 0.00154806f $X=3.025 $Y=2.035 $X2=0 $Y2=0
cc_183 N_A_83_283#_c_166_n B1 0.0264615f $X=3.885 $Y=2.035 $X2=0 $Y2=0
cc_184 N_A_83_283#_c_154_n B1 0.0260237f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_185 N_A_83_283#_c_156_n B1 0.020325f $X=4.055 $Y=1.195 $X2=0 $Y2=0
cc_186 N_A_83_283#_c_168_n B1 0.0289327f $X=3.19 $Y=2.115 $X2=0 $Y2=0
cc_187 N_A_83_283#_c_166_n N_B1_c_435_n 0.00401172f $X=3.885 $Y=2.035 $X2=0
+ $Y2=0
cc_188 N_A_83_283#_c_154_n N_B1_c_435_n 0.00947853f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_189 N_A_83_283#_c_156_n N_B1_c_435_n 0.00463794f $X=4.055 $Y=1.195 $X2=0
+ $Y2=0
cc_190 N_A_83_283#_c_168_n N_B1_c_435_n 5.65925e-19 $X=3.19 $Y=2.115 $X2=0 $Y2=0
cc_191 N_A_83_283#_c_155_n N_A2_M1009_g 0.015229f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_192 N_A_83_283#_c_157_n N_A2_M1009_g 8.67208e-19 $X=5.965 $Y=1.1 $X2=0 $Y2=0
cc_193 N_A_83_283#_c_155_n N_A2_c_490_n 0.0120417f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_194 N_A_83_283#_c_155_n N_A2_c_498_n 0.00804233f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_195 N_A_83_283#_c_157_n N_A2_c_498_n 3.19435e-19 $X=5.965 $Y=1.1 $X2=0 $Y2=0
cc_196 N_A_83_283#_c_154_n N_A2_c_491_n 0.0148327f $X=3.97 $Y=1.95 $X2=0 $Y2=0
cc_197 N_A_83_283#_c_155_n N_A2_c_491_n 0.0520648f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_198 N_A_83_283#_c_155_n N_A2_c_494_n 0.00460348f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_199 N_A_83_283#_c_155_n N_A1_M1025_g 0.00914156f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_200 N_A_83_283#_c_157_n N_A1_M1025_g 0.00505973f $X=5.965 $Y=1.1 $X2=0 $Y2=0
cc_201 N_A_83_283#_c_157_n N_A1_M1026_g 0.00492104f $X=5.965 $Y=1.1 $X2=0 $Y2=0
cc_202 N_A_83_283#_c_155_n A1 0.0119328f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_203 N_A_83_283#_c_157_n A1 0.0249237f $X=5.965 $Y=1.1 $X2=0 $Y2=0
cc_204 N_A_83_283#_c_155_n N_A1_c_599_n 0.00105442f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_205 N_A_83_283#_c_157_n N_A1_c_599_n 0.00228249f $X=5.965 $Y=1.1 $X2=0 $Y2=0
cc_206 N_A_83_283#_c_164_n N_VPWR_M1006_s 0.00255376f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_207 N_A_83_283#_c_165_n N_VPWR_M1006_s 0.00516953f $X=3.025 $Y=2.035 $X2=0
+ $Y2=0
cc_208 N_A_83_283#_c_230_p N_VPWR_M1006_s 0.00264469f $X=2.185 $Y=2.035 $X2=0
+ $Y2=0
cc_209 N_A_83_283#_M1003_g N_VPWR_c_701_n 0.00517389f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_210 N_A_83_283#_M1003_g N_VPWR_c_702_n 6.08595e-19 $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_83_283#_M1004_g N_VPWR_c_702_n 0.0155441f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_83_283#_M1005_g N_VPWR_c_702_n 0.0024353f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A_83_283#_M1005_g N_VPWR_c_703_n 4.96657e-19 $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_214 N_A_83_283#_M1006_g N_VPWR_c_703_n 0.014135f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_83_283#_c_153_n N_VPWR_c_703_n 0.00111188f $X=2.015 $Y=1.515 $X2=0
+ $Y2=0
cc_216 N_A_83_283#_c_165_n N_VPWR_c_703_n 0.00889054f $X=3.025 $Y=2.035 $X2=0
+ $Y2=0
cc_217 N_A_83_283#_c_230_p N_VPWR_c_703_n 0.0119464f $X=2.185 $Y=2.035 $X2=0
+ $Y2=0
cc_218 N_A_83_283#_M1003_g N_VPWR_c_707_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_83_283#_M1004_g N_VPWR_c_707_n 0.00460063f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_220 N_A_83_283#_M1005_g N_VPWR_c_708_n 0.00520371f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_221 N_A_83_283#_M1006_g N_VPWR_c_708_n 0.00460063f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_222 N_A_83_283#_M1003_g N_VPWR_c_699_n 0.00986008f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_223 N_A_83_283#_M1004_g N_VPWR_c_699_n 0.00908554f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_83_283#_M1005_g N_VPWR_c_699_n 0.00981712f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_225 N_A_83_283#_M1006_g N_VPWR_c_699_n 0.00908554f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_226 N_A_83_283#_c_149_n N_X_c_819_n 0.0166532f $X=0.495 $Y=1.265 $X2=0 $Y2=0
cc_227 N_A_83_283#_c_153_n N_X_c_811_n 0.0144067f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A_83_283#_c_158_n N_X_c_811_n 0.0252063f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_229 N_A_83_283#_M1003_g N_X_c_816_n 0.00770588f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A_83_283#_M1004_g N_X_c_816_n 0.00411725f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A_83_283#_c_153_n N_X_c_816_n 0.00223325f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_232 N_A_83_283#_c_158_n N_X_c_816_n 0.00445965f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_233 N_A_83_283#_M1003_g N_X_c_817_n 0.012903f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A_83_283#_M1004_g N_X_c_817_n 3.68116e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_83_283#_c_149_n N_X_c_813_n 7.4531e-19 $X=0.495 $Y=1.265 $X2=0 $Y2=0
cc_236 N_A_83_283#_c_150_n N_X_c_813_n 7.4531e-19 $X=0.94 $Y=1.265 $X2=0 $Y2=0
cc_237 N_A_83_283#_M1004_g N_X_c_830_n 0.0163066f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A_83_283#_M1005_g N_X_c_830_n 0.0132272f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_83_283#_c_153_n N_X_c_830_n 0.0344509f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A_83_283#_c_158_n N_X_c_830_n 0.00313888f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_241 N_A_83_283#_c_150_n N_X_c_834_n 0.0172454f $X=0.94 $Y=1.265 $X2=0 $Y2=0
cc_242 N_A_83_283#_M1014_g N_X_c_834_n 0.0151224f $X=1.52 $Y=0.82 $X2=0 $Y2=0
cc_243 N_A_83_283#_M1023_g N_X_c_834_n 0.00302177f $X=1.95 $Y=0.82 $X2=0 $Y2=0
cc_244 N_A_83_283#_c_153_n N_X_c_834_n 0.0615598f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_245 N_A_83_283#_c_158_n N_X_c_834_n 0.0086557f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_246 N_A_83_283#_M1005_g N_X_c_839_n 8.84614e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_83_283#_c_153_n N_X_c_839_n 0.0187792f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A_83_283#_c_158_n N_X_c_839_n 0.00229382f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_249 N_A_83_283#_M1004_g N_X_c_818_n 8.57327e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_83_283#_M1005_g N_X_c_818_n 0.0134225f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A_83_283#_M1006_g N_X_c_818_n 4.96772e-19 $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A_83_283#_c_150_n N_X_c_814_n 7.69011e-19 $X=0.94 $Y=1.265 $X2=0 $Y2=0
cc_253 N_A_83_283#_M1014_g N_X_c_814_n 0.00774615f $X=1.52 $Y=0.82 $X2=0 $Y2=0
cc_254 N_A_83_283#_M1023_g N_X_c_814_n 0.00618839f $X=1.95 $Y=0.82 $X2=0 $Y2=0
cc_255 N_A_83_283#_M1003_g N_X_c_848_n 0.00213632f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A_83_283#_c_158_n N_X_c_849_n 0.00346273f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_257 N_A_83_283#_c_149_n X 0.00966807f $X=0.495 $Y=1.265 $X2=0 $Y2=0
cc_258 N_A_83_283#_c_153_n X 0.00381558f $X=2.015 $Y=1.515 $X2=0 $Y2=0
cc_259 N_A_83_283#_c_158_n X 0.00234311f $X=1.905 $Y=1.472 $X2=0 $Y2=0
cc_260 N_A_83_283#_c_165_n N_A_509_392#_M1015_d 0.0032506f $X=3.025 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_261 N_A_83_283#_c_166_n N_A_509_392#_M1018_d 0.00218982f $X=3.885 $Y=2.035
+ $X2=0 $Y2=0
cc_262 N_A_83_283#_M1006_g N_A_509_392#_c_879_n 0.00111873f $X=1.905 $Y=2.4
+ $X2=0 $Y2=0
cc_263 N_A_83_283#_c_165_n N_A_509_392#_c_879_n 0.0219146f $X=3.025 $Y=2.035
+ $X2=0 $Y2=0
cc_264 N_A_83_283#_M1015_s N_A_509_392#_c_880_n 0.00218982f $X=3.005 $Y=1.96
+ $X2=0 $Y2=0
cc_265 N_A_83_283#_c_168_n N_A_509_392#_c_880_n 0.0177084f $X=3.19 $Y=2.115
+ $X2=0 $Y2=0
cc_266 N_A_83_283#_M1006_g N_A_509_392#_c_881_n 6.08298e-19 $X=1.905 $Y=2.4
+ $X2=0 $Y2=0
cc_267 N_A_83_283#_c_166_n N_A_509_392#_c_897_n 0.0189268f $X=3.885 $Y=2.035
+ $X2=0 $Y2=0
cc_268 N_A_83_283#_M1019_s N_A_509_392#_c_882_n 0.00218982f $X=4.005 $Y=1.96
+ $X2=0 $Y2=0
cc_269 N_A_83_283#_c_169_n N_A_509_392#_c_882_n 0.0177084f $X=4.19 $Y=2.115
+ $X2=0 $Y2=0
cc_270 N_A_83_283#_c_169_n N_A_509_392#_c_889_n 0.0466785f $X=4.19 $Y=2.115
+ $X2=0 $Y2=0
cc_271 N_A_83_283#_c_155_n N_VGND_M1022_s 0.00411123f $X=5.8 $Y=1.195 $X2=0
+ $Y2=0
cc_272 N_A_83_283#_c_149_n N_VGND_c_987_n 0.00861216f $X=0.495 $Y=1.265 $X2=0
+ $Y2=0
cc_273 N_A_83_283#_c_150_n N_VGND_c_987_n 3.63144e-19 $X=0.94 $Y=1.265 $X2=0
+ $Y2=0
cc_274 N_A_83_283#_c_149_n N_VGND_c_988_n 3.62248e-19 $X=0.495 $Y=1.265 $X2=0
+ $Y2=0
cc_275 N_A_83_283#_c_150_n N_VGND_c_988_n 0.0078948f $X=0.94 $Y=1.265 $X2=0
+ $Y2=0
cc_276 N_A_83_283#_M1014_g N_VGND_c_988_n 0.0040012f $X=1.52 $Y=0.82 $X2=0 $Y2=0
cc_277 N_A_83_283#_M1023_g N_VGND_c_989_n 0.0178705f $X=1.95 $Y=0.82 $X2=0 $Y2=0
cc_278 N_A_83_283#_c_153_n N_VGND_c_989_n 0.00998409f $X=2.015 $Y=1.515 $X2=0
+ $Y2=0
cc_279 N_A_83_283#_c_155_n N_VGND_c_990_n 0.0285408f $X=5.8 $Y=1.195 $X2=0 $Y2=0
cc_280 N_A_83_283#_c_149_n N_VGND_c_994_n 0.00432588f $X=0.495 $Y=1.265 $X2=0
+ $Y2=0
cc_281 N_A_83_283#_c_150_n N_VGND_c_994_n 0.00432588f $X=0.94 $Y=1.265 $X2=0
+ $Y2=0
cc_282 N_A_83_283#_M1014_g N_VGND_c_995_n 0.00497955f $X=1.52 $Y=0.82 $X2=0
+ $Y2=0
cc_283 N_A_83_283#_M1023_g N_VGND_c_995_n 0.00497955f $X=1.95 $Y=0.82 $X2=0
+ $Y2=0
cc_284 N_A_83_283#_c_149_n N_VGND_c_998_n 0.00437282f $X=0.495 $Y=1.265 $X2=0
+ $Y2=0
cc_285 N_A_83_283#_c_150_n N_VGND_c_998_n 0.00437282f $X=0.94 $Y=1.265 $X2=0
+ $Y2=0
cc_286 N_A_83_283#_M1014_g N_VGND_c_998_n 0.00520574f $X=1.52 $Y=0.82 $X2=0
+ $Y2=0
cc_287 N_A_83_283#_M1023_g N_VGND_c_998_n 0.00520574f $X=1.95 $Y=0.82 $X2=0
+ $Y2=0
cc_288 N_A_83_283#_c_154_n N_A_587_110#_M1021_s 6.02464e-19 $X=3.97 $Y=1.95
+ $X2=0 $Y2=0
cc_289 N_A_83_283#_c_155_n N_A_587_110#_M1021_s 0.0012905f $X=5.8 $Y=1.195 $X2=0
+ $Y2=0
cc_290 N_A_83_283#_c_156_n N_A_587_110#_M1021_s 0.00141439f $X=4.055 $Y=1.195
+ $X2=0 $Y2=0
cc_291 N_A_83_283#_M1001_d N_A_587_110#_c_1079_n 0.00586822f $X=3.365 $Y=0.55
+ $X2=0 $Y2=0
cc_292 N_A_83_283#_c_155_n N_A_587_110#_c_1079_n 0.0044508f $X=5.8 $Y=1.195
+ $X2=0 $Y2=0
cc_293 N_A_83_283#_c_156_n N_A_587_110#_c_1079_n 0.0370778f $X=4.055 $Y=1.195
+ $X2=0 $Y2=0
cc_294 N_A_83_283#_c_156_n N_A_587_110#_c_1075_n 0.00499071f $X=4.055 $Y=1.195
+ $X2=0 $Y2=0
cc_295 N_A_83_283#_c_155_n N_A_992_122#_M1009_d 0.00242368f $X=5.8 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_296 N_A_83_283#_c_155_n N_A_992_122#_c_1098_n 0.0201666f $X=5.8 $Y=1.195
+ $X2=0 $Y2=0
cc_297 N_A_83_283#_c_155_n N_A_1079_122#_M1009_s 0.00176461f $X=5.8 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_298 N_A_83_283#_M1025_d N_A_1079_122#_c_1146_n 0.00169276f $X=5.825 $Y=0.61
+ $X2=0 $Y2=0
cc_299 N_A_83_283#_c_155_n N_A_1079_122#_c_1146_n 0.00478439f $X=5.8 $Y=1.195
+ $X2=0 $Y2=0
cc_300 N_A_83_283#_c_157_n N_A_1079_122#_c_1146_n 0.0161743f $X=5.965 $Y=1.1
+ $X2=0 $Y2=0
cc_301 N_A_83_283#_c_155_n N_A_1079_122#_c_1147_n 0.0144832f $X=5.8 $Y=1.195
+ $X2=0 $Y2=0
cc_302 N_A_83_283#_c_157_n N_A_1079_122#_c_1148_n 0.0127348f $X=5.965 $Y=1.1
+ $X2=0 $Y2=0
cc_303 N_B2_M1000_g N_B1_M1001_g 0.0176613f $X=2.86 $Y=0.87 $X2=0 $Y2=0
cc_304 N_B2_c_332_n N_B1_M1001_g 0.00548812f $X=4.085 $Y=0.34 $X2=0 $Y2=0
cc_305 N_B2_c_337_n N_B1_M1001_g 0.00339207f $X=4.415 $Y=0.42 $X2=0 $Y2=0
cc_306 N_B2_M1015_g N_B1_c_436_n 0.0149287f $X=2.915 $Y=2.46 $X2=0 $Y2=0
cc_307 N_B2_c_326_n N_B1_c_433_n 0.0234859f $X=4.23 $Y=0.585 $X2=0 $Y2=0
cc_308 N_B2_c_332_n N_B1_c_433_n 0.00437843f $X=4.085 $Y=0.34 $X2=0 $Y2=0
cc_309 N_B2_c_337_n N_B1_c_433_n 0.00137701f $X=4.415 $Y=0.42 $X2=0 $Y2=0
cc_310 N_B2_c_340_n N_B1_c_437_n 0.0118685f $X=4.415 $Y=1.855 $X2=0 $Y2=0
cc_311 B2 B1 0.0262736f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_312 N_B2_c_336_n B1 0.00339157f $X=2.915 $Y=1.615 $X2=0 $Y2=0
cc_313 N_B2_c_330_n N_B1_c_435_n 0.0118685f $X=4.705 $Y=1.78 $X2=0 $Y2=0
cc_314 B2 N_B1_c_435_n 2.10201e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_315 N_B2_c_336_n N_B1_c_435_n 0.0247329f $X=2.915 $Y=1.615 $X2=0 $Y2=0
cc_316 N_B2_c_340_n N_A2_M1010_g 0.0195499f $X=4.415 $Y=1.855 $X2=0 $Y2=0
cc_317 N_B2_c_330_n N_A2_M1010_g 0.0107041f $X=4.705 $Y=1.78 $X2=0 $Y2=0
cc_318 N_B2_c_327_n N_A2_M1009_g 0.0178376f $X=4.735 $Y=0.51 $X2=0 $Y2=0
cc_319 N_B2_c_328_n N_A2_M1009_g 0.00715928f $X=4.705 $Y=1.705 $X2=0 $Y2=0
cc_320 N_B2_c_340_n N_A2_c_497_n 3.97731e-19 $X=4.415 $Y=1.855 $X2=0 $Y2=0
cc_321 N_B2_c_330_n N_A2_c_497_n 3.34079e-19 $X=4.705 $Y=1.78 $X2=0 $Y2=0
cc_322 N_B2_c_328_n N_A2_c_491_n 0.0121365f $X=4.705 $Y=1.705 $X2=0 $Y2=0
cc_323 N_B2_c_330_n N_A2_c_491_n 0.0162275f $X=4.705 $Y=1.78 $X2=0 $Y2=0
cc_324 N_B2_c_331_n N_A2_c_491_n 6.63248e-19 $X=4.81 $Y=1.155 $X2=0 $Y2=0
cc_325 N_B2_c_328_n N_A2_c_494_n 0.0107041f $X=4.705 $Y=1.705 $X2=0 $Y2=0
cc_326 N_B2_M1015_g N_VPWR_c_703_n 0.00200483f $X=2.915 $Y=2.46 $X2=0 $Y2=0
cc_327 N_B2_M1015_g N_VPWR_c_709_n 0.00333896f $X=2.915 $Y=2.46 $X2=0 $Y2=0
cc_328 N_B2_c_340_n N_VPWR_c_709_n 0.00333926f $X=4.415 $Y=1.855 $X2=0 $Y2=0
cc_329 N_B2_M1015_g N_VPWR_c_699_n 0.00428385f $X=2.915 $Y=2.46 $X2=0 $Y2=0
cc_330 N_B2_c_340_n N_VPWR_c_699_n 0.0042525f $X=4.415 $Y=1.855 $X2=0 $Y2=0
cc_331 N_B2_M1015_g N_A_509_392#_c_879_n 0.00935952f $X=2.915 $Y=2.46 $X2=0
+ $Y2=0
cc_332 N_B2_M1015_g N_A_509_392#_c_880_n 0.0118818f $X=2.915 $Y=2.46 $X2=0 $Y2=0
cc_333 N_B2_M1015_g N_A_509_392#_c_881_n 0.00291744f $X=2.915 $Y=2.46 $X2=0
+ $Y2=0
cc_334 N_B2_c_340_n N_A_509_392#_c_897_n 7.8508e-19 $X=4.415 $Y=1.855 $X2=0
+ $Y2=0
cc_335 N_B2_c_340_n N_A_509_392#_c_882_n 0.0157614f $X=4.415 $Y=1.855 $X2=0
+ $Y2=0
cc_336 N_B2_c_340_n N_A_509_392#_c_889_n 0.0133598f $X=4.415 $Y=1.855 $X2=0
+ $Y2=0
cc_337 N_B2_c_330_n N_A_509_392#_c_889_n 0.00515135f $X=4.705 $Y=1.78 $X2=0
+ $Y2=0
cc_338 N_B2_c_338_n N_VGND_M1023_s 0.0114021f $X=2.67 $Y=1.45 $X2=0 $Y2=0
cc_339 N_B2_M1000_g N_VGND_c_989_n 0.00129931f $X=2.86 $Y=0.87 $X2=0 $Y2=0
cc_340 N_B2_c_333_n N_VGND_c_989_n 0.0150384f $X=2.74 $Y=0.34 $X2=0 $Y2=0
cc_341 N_B2_c_338_n N_VGND_c_989_n 0.0580184f $X=2.67 $Y=1.45 $X2=0 $Y2=0
cc_342 N_B2_c_326_n N_VGND_c_990_n 0.0032883f $X=4.23 $Y=0.585 $X2=0 $Y2=0
cc_343 N_B2_c_327_n N_VGND_c_990_n 0.0107093f $X=4.735 $Y=0.51 $X2=0 $Y2=0
cc_344 N_B2_c_329_n N_VGND_c_990_n 0.00846666f $X=4.81 $Y=1.08 $X2=0 $Y2=0
cc_345 N_B2_c_331_n N_VGND_c_990_n 0.00262004f $X=4.81 $Y=1.155 $X2=0 $Y2=0
cc_346 N_B2_c_334_n N_VGND_c_990_n 0.028447f $X=4.25 $Y=0.34 $X2=0 $Y2=0
cc_347 N_B2_c_337_n N_VGND_c_990_n 0.00832206f $X=4.415 $Y=0.42 $X2=0 $Y2=0
cc_348 N_B2_M1000_g N_VGND_c_992_n 6.29586e-19 $X=2.86 $Y=0.87 $X2=0 $Y2=0
cc_349 N_B2_c_327_n N_VGND_c_992_n 0.00296597f $X=4.735 $Y=0.51 $X2=0 $Y2=0
cc_350 N_B2_c_332_n N_VGND_c_992_n 0.0866135f $X=4.085 $Y=0.34 $X2=0 $Y2=0
cc_351 N_B2_c_333_n N_VGND_c_992_n 0.0121867f $X=2.74 $Y=0.34 $X2=0 $Y2=0
cc_352 N_B2_c_334_n N_VGND_c_992_n 0.0212434f $X=4.25 $Y=0.34 $X2=0 $Y2=0
cc_353 N_B2_c_337_n N_VGND_c_992_n 0.00213713f $X=4.415 $Y=0.42 $X2=0 $Y2=0
cc_354 N_B2_c_327_n N_VGND_c_996_n 0.00387605f $X=4.735 $Y=0.51 $X2=0 $Y2=0
cc_355 N_B2_c_327_n N_VGND_c_998_n 0.00865339f $X=4.735 $Y=0.51 $X2=0 $Y2=0
cc_356 N_B2_c_332_n N_VGND_c_998_n 0.0505651f $X=4.085 $Y=0.34 $X2=0 $Y2=0
cc_357 N_B2_c_333_n N_VGND_c_998_n 0.00660921f $X=2.74 $Y=0.34 $X2=0 $Y2=0
cc_358 N_B2_c_334_n N_VGND_c_998_n 0.0123341f $X=4.25 $Y=0.34 $X2=0 $Y2=0
cc_359 N_B2_c_326_n N_A_587_110#_c_1079_n 0.00240721f $X=4.23 $Y=0.585 $X2=0
+ $Y2=0
cc_360 N_B2_c_332_n N_A_587_110#_c_1079_n 0.0303947f $X=4.085 $Y=0.34 $X2=0
+ $Y2=0
cc_361 N_B2_c_334_n N_A_587_110#_c_1079_n 0.00471774f $X=4.25 $Y=0.34 $X2=0
+ $Y2=0
cc_362 N_B2_c_337_n N_A_587_110#_c_1079_n 3.62043e-19 $X=4.415 $Y=0.42 $X2=0
+ $Y2=0
cc_363 N_B2_M1000_g N_A_587_110#_c_1075_n 0.00833353f $X=2.86 $Y=0.87 $X2=0
+ $Y2=0
cc_364 N_B2_c_332_n N_A_587_110#_c_1075_n 0.0203882f $X=4.085 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_B2_c_336_n N_A_587_110#_c_1075_n 0.00308615f $X=2.915 $Y=1.615 $X2=0
+ $Y2=0
cc_366 N_B2_c_338_n N_A_587_110#_c_1075_n 0.0237911f $X=2.67 $Y=1.45 $X2=0 $Y2=0
cc_367 N_B2_c_327_n N_A_992_122#_c_1098_n 0.00556037f $X=4.735 $Y=0.51 $X2=0
+ $Y2=0
cc_368 N_B1_c_436_n N_VPWR_c_709_n 0.00333926f $X=3.415 $Y=1.855 $X2=0 $Y2=0
cc_369 N_B1_c_437_n N_VPWR_c_709_n 0.00333896f $X=3.915 $Y=1.855 $X2=0 $Y2=0
cc_370 N_B1_c_436_n N_VPWR_c_699_n 0.00423742f $X=3.415 $Y=1.855 $X2=0 $Y2=0
cc_371 N_B1_c_437_n N_VPWR_c_699_n 0.0042374f $X=3.915 $Y=1.855 $X2=0 $Y2=0
cc_372 N_B1_c_436_n N_A_509_392#_c_879_n 5.24303e-19 $X=3.415 $Y=1.855 $X2=0
+ $Y2=0
cc_373 N_B1_c_436_n N_A_509_392#_c_880_n 0.0144686f $X=3.415 $Y=1.855 $X2=0
+ $Y2=0
cc_374 N_B1_c_437_n N_A_509_392#_c_897_n 0.00899947f $X=3.915 $Y=1.855 $X2=0
+ $Y2=0
cc_375 N_B1_c_437_n N_A_509_392#_c_882_n 0.0118818f $X=3.915 $Y=1.855 $X2=0
+ $Y2=0
cc_376 N_B1_c_437_n N_A_509_392#_c_888_n 0.00214324f $X=3.915 $Y=1.855 $X2=0
+ $Y2=0
cc_377 N_B1_M1001_g N_VGND_c_992_n 6.29586e-19 $X=3.29 $Y=0.87 $X2=0 $Y2=0
cc_378 N_B1_M1001_g N_A_587_110#_c_1079_n 0.0105309f $X=3.29 $Y=0.87 $X2=0 $Y2=0
cc_379 N_B1_c_433_n N_A_587_110#_c_1079_n 0.00899967f $X=3.8 $Y=1.45 $X2=0 $Y2=0
cc_380 B1 N_A_587_110#_c_1079_n 0.00436875f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_381 N_B1_M1001_g N_A_587_110#_c_1075_n 0.00950294f $X=3.29 $Y=0.87 $X2=0
+ $Y2=0
cc_382 N_B1_c_433_n N_A_587_110#_c_1075_n 0.00137982f $X=3.8 $Y=1.45 $X2=0 $Y2=0
cc_383 B1 N_A_587_110#_c_1075_n 0.015912f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A2_M1010_g N_A1_M1016_g 0.0274307f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_385 N_A2_c_497_n N_A1_M1016_g 0.00295955f $X=5.265 $Y=1.95 $X2=0 $Y2=0
cc_386 N_A2_c_498_n N_A1_M1016_g 0.0125511f $X=6.425 $Y=2.035 $X2=0 $Y2=0
cc_387 N_A2_c_494_n N_A1_M1016_g 0.00945217f $X=5.32 $Y=1.635 $X2=0 $Y2=0
cc_388 N_A2_M1009_g N_A1_M1025_g 0.0291177f $X=5.32 $Y=0.93 $X2=0 $Y2=0
cc_389 N_A2_M1024_g N_A1_M1026_g 0.0194846f $X=6.69 $Y=0.93 $X2=0 $Y2=0
cc_390 N_A2_c_492_n N_A1_M1026_g 2.1371e-19 $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_391 N_A2_c_493_n N_A1_M1026_g 4.8841e-19 $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_392 N_A2_c_498_n N_A1_M1027_g 0.0167078f $X=6.425 $Y=2.035 $X2=0 $Y2=0
cc_393 N_A2_M1009_g A1 0.00131772f $X=5.32 $Y=0.93 $X2=0 $Y2=0
cc_394 N_A2_c_490_n A1 0.0167955f $X=5.265 $Y=1.79 $X2=0 $Y2=0
cc_395 N_A2_c_498_n A1 0.0353667f $X=6.425 $Y=2.035 $X2=0 $Y2=0
cc_396 N_A2_c_499_n A1 4.45324e-19 $X=6.51 $Y=1.95 $X2=0 $Y2=0
cc_397 N_A2_c_492_n A1 0.0168753f $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_398 N_A2_c_493_n A1 2.81631e-19 $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_399 N_A2_M1009_g N_A1_c_599_n 0.00945217f $X=5.32 $Y=0.93 $X2=0 $Y2=0
cc_400 N_A2_M1011_g N_A1_c_599_n 0.0327743f $X=6.705 $Y=2.46 $X2=0 $Y2=0
cc_401 N_A2_c_490_n N_A1_c_599_n 4.25448e-19 $X=5.265 $Y=1.79 $X2=0 $Y2=0
cc_402 N_A2_c_498_n N_A1_c_599_n 0.00250566f $X=6.425 $Y=2.035 $X2=0 $Y2=0
cc_403 N_A2_c_499_n N_A1_c_599_n 0.00385971f $X=6.51 $Y=1.95 $X2=0 $Y2=0
cc_404 N_A2_c_492_n N_A1_c_599_n 0.00278666f $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_405 N_A2_c_493_n N_A1_c_599_n 0.0209592f $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_406 N_A2_M1024_g N_A3_M1002_g 0.0136615f $X=6.69 $Y=0.93 $X2=0 $Y2=0
cc_407 N_A2_c_493_n N_A3_M1002_g 0.0181723f $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_408 N_A2_c_499_n A3 3.31897e-19 $X=6.51 $Y=1.95 $X2=0 $Y2=0
cc_409 N_A2_c_492_n A3 0.0195876f $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_410 N_A2_c_493_n A3 4.03387e-19 $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_411 N_A2_M1011_g N_A3_c_652_n 0.0150137f $X=6.705 $Y=2.46 $X2=0 $Y2=0
cc_412 N_A2_c_492_n N_A3_c_652_n 4.02409e-19 $X=6.66 $Y=1.605 $X2=0 $Y2=0
cc_413 N_A2_c_498_n N_VPWR_M1010_d 0.00299596f $X=6.425 $Y=2.035 $X2=0 $Y2=0
cc_414 N_A2_c_552_p N_VPWR_M1010_d 0.00103027f $X=5.35 $Y=2.035 $X2=0 $Y2=0
cc_415 N_A2_c_498_n N_VPWR_M1027_s 0.00308605f $X=6.425 $Y=2.035 $X2=0 $Y2=0
cc_416 N_A2_M1010_g N_VPWR_c_704_n 0.00200073f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_417 N_A2_M1011_g N_VPWR_c_705_n 0.00846267f $X=6.705 $Y=2.46 $X2=0 $Y2=0
cc_418 N_A2_M1010_g N_VPWR_c_709_n 0.00553757f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_419 N_A2_M1011_g N_VPWR_c_711_n 0.00460063f $X=6.705 $Y=2.46 $X2=0 $Y2=0
cc_420 N_A2_M1010_g N_VPWR_c_699_n 0.0109123f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_421 N_A2_M1011_g N_VPWR_c_699_n 0.00908665f $X=6.705 $Y=2.46 $X2=0 $Y2=0
cc_422 N_A2_c_498_n N_A_509_392#_M1016_d 0.00187091f $X=6.425 $Y=2.035 $X2=0
+ $Y2=0
cc_423 N_A2_M1010_g N_A_509_392#_c_882_n 0.00211513f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_424 N_A2_M1010_g N_A_509_392#_c_915_n 0.0192057f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_425 N_A2_c_498_n N_A_509_392#_c_915_n 0.0266572f $X=6.425 $Y=2.035 $X2=0
+ $Y2=0
cc_426 N_A2_c_552_p N_A_509_392#_c_915_n 0.00901441f $X=5.35 $Y=2.035 $X2=0
+ $Y2=0
cc_427 N_A2_c_491_n N_A_509_392#_c_915_n 0.00720107f $X=5.18 $Y=1.63 $X2=0 $Y2=0
cc_428 N_A2_c_494_n N_A_509_392#_c_915_n 5.25024e-19 $X=5.32 $Y=1.635 $X2=0
+ $Y2=0
cc_429 N_A2_M1011_g N_A_509_392#_c_920_n 0.0138845f $X=6.705 $Y=2.46 $X2=0 $Y2=0
cc_430 N_A2_c_498_n N_A_509_392#_c_920_n 0.0277459f $X=6.425 $Y=2.035 $X2=0
+ $Y2=0
cc_431 N_A2_c_492_n N_A_509_392#_c_920_n 0.00461576f $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_432 N_A2_c_493_n N_A_509_392#_c_920_n 2.90147e-19 $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_433 N_A2_M1011_g N_A_509_392#_c_883_n 0.00245062f $X=6.705 $Y=2.46 $X2=0
+ $Y2=0
cc_434 N_A2_c_498_n N_A_509_392#_c_883_n 0.00761666f $X=6.425 $Y=2.035 $X2=0
+ $Y2=0
cc_435 N_A2_c_492_n N_A_509_392#_c_883_n 0.00462064f $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_436 N_A2_c_493_n N_A_509_392#_c_883_n 6.90659e-19 $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_437 N_A2_M1011_g N_A_509_392#_c_928_n 0.00335669f $X=6.705 $Y=2.46 $X2=0
+ $Y2=0
cc_438 N_A2_M1011_g N_A_509_392#_c_884_n 3.13895e-19 $X=6.705 $Y=2.46 $X2=0
+ $Y2=0
cc_439 N_A2_M1010_g N_A_509_392#_c_889_n 0.0151205f $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_440 N_A2_c_552_p N_A_509_392#_c_889_n 0.00963908f $X=5.35 $Y=2.035 $X2=0
+ $Y2=0
cc_441 N_A2_c_491_n N_A_509_392#_c_889_n 0.0276176f $X=5.18 $Y=1.63 $X2=0 $Y2=0
cc_442 N_A2_M1010_g N_A_509_392#_c_933_n 6.29986e-19 $X=5.11 $Y=2.46 $X2=0 $Y2=0
cc_443 N_A2_M1011_g N_A_509_392#_c_933_n 6.96091e-19 $X=6.705 $Y=2.46 $X2=0
+ $Y2=0
cc_444 N_A2_c_498_n N_A_509_392#_c_933_n 0.0171308f $X=6.425 $Y=2.035 $X2=0
+ $Y2=0
cc_445 N_A2_M1011_g N_A_509_392#_c_936_n 0.00186115f $X=6.705 $Y=2.46 $X2=0
+ $Y2=0
cc_446 N_A2_M1024_g N_VGND_c_996_n 2.28603e-19 $X=6.69 $Y=0.93 $X2=0 $Y2=0
cc_447 N_A2_M1009_g N_A_992_122#_c_1098_n 0.00319542f $X=5.32 $Y=0.93 $X2=0
+ $Y2=0
cc_448 N_A2_M1009_g N_A_992_122#_c_1099_n 0.00665247f $X=5.32 $Y=0.93 $X2=0
+ $Y2=0
cc_449 N_A2_M1024_g N_A_992_122#_c_1099_n 0.00586193f $X=6.69 $Y=0.93 $X2=0
+ $Y2=0
cc_450 N_A2_M1024_g N_A_992_122#_c_1101_n 0.00912122f $X=6.69 $Y=0.93 $X2=0
+ $Y2=0
cc_451 N_A2_M1024_g N_A_992_122#_c_1103_n 0.00237179f $X=6.69 $Y=0.93 $X2=0
+ $Y2=0
cc_452 N_A2_c_492_n N_A_992_122#_c_1103_n 0.00701349f $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_453 N_A2_c_493_n N_A_992_122#_c_1103_n 0.00151606f $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_454 N_A2_M1009_g N_A_1079_122#_c_1147_n 0.0042312f $X=5.32 $Y=0.93 $X2=0
+ $Y2=0
cc_455 N_A2_M1024_g N_A_1079_122#_c_1148_n 0.00365046f $X=6.69 $Y=0.93 $X2=0
+ $Y2=0
cc_456 N_A2_c_492_n N_A_1079_122#_c_1148_n 0.0115827f $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_457 N_A2_c_493_n N_A_1079_122#_c_1148_n 0.00148807f $X=6.66 $Y=1.605 $X2=0
+ $Y2=0
cc_458 N_A1_M1016_g N_VPWR_c_704_n 0.00462216f $X=5.725 $Y=2.46 $X2=0 $Y2=0
cc_459 N_A1_M1027_g N_VPWR_c_705_n 0.00222098f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_460 N_A1_M1016_g N_VPWR_c_710_n 0.00522932f $X=5.725 $Y=2.46 $X2=0 $Y2=0
cc_461 N_A1_M1027_g N_VPWR_c_710_n 0.0054279f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_462 N_A1_M1016_g N_VPWR_c_699_n 0.00985386f $X=5.725 $Y=2.46 $X2=0 $Y2=0
cc_463 N_A1_M1027_g N_VPWR_c_699_n 0.0105603f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_464 N_A1_M1016_g N_A_509_392#_c_915_n 0.0134752f $X=5.725 $Y=2.46 $X2=0 $Y2=0
cc_465 N_A1_M1027_g N_A_509_392#_c_920_n 0.0144393f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_466 N_A1_M1027_g N_A_509_392#_c_928_n 7.87188e-19 $X=6.195 $Y=2.46 $X2=0
+ $Y2=0
cc_467 N_A1_M1016_g N_A_509_392#_c_933_n 0.00860098f $X=5.725 $Y=2.46 $X2=0
+ $Y2=0
cc_468 N_A1_M1027_g N_A_509_392#_c_933_n 0.00678294f $X=6.195 $Y=2.46 $X2=0
+ $Y2=0
cc_469 N_A1_M1025_g N_A_992_122#_c_1099_n 0.00452619f $X=5.75 $Y=0.93 $X2=0
+ $Y2=0
cc_470 N_A1_M1026_g N_A_992_122#_c_1099_n 0.00452619f $X=6.18 $Y=0.93 $X2=0
+ $Y2=0
cc_471 N_A1_M1026_g N_A_992_122#_c_1101_n 5.92696e-19 $X=6.18 $Y=0.93 $X2=0
+ $Y2=0
cc_472 N_A1_M1025_g N_A_1079_122#_c_1146_n 0.008467f $X=5.75 $Y=0.93 $X2=0 $Y2=0
cc_473 N_A1_M1026_g N_A_1079_122#_c_1146_n 0.011549f $X=6.18 $Y=0.93 $X2=0 $Y2=0
cc_474 N_A3_M1013_g N_VPWR_c_705_n 3.87154e-19 $X=7.155 $Y=2.46 $X2=0 $Y2=0
cc_475 N_A3_M1013_g N_VPWR_c_706_n 0.00170765f $X=7.155 $Y=2.46 $X2=0 $Y2=0
cc_476 N_A3_M1017_g N_VPWR_c_706_n 0.00325025f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_477 N_A3_M1013_g N_VPWR_c_711_n 0.00520371f $X=7.155 $Y=2.46 $X2=0 $Y2=0
cc_478 N_A3_M1017_g N_VPWR_c_712_n 0.005209f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_479 N_A3_M1013_g N_VPWR_c_699_n 0.00981823f $X=7.155 $Y=2.46 $X2=0 $Y2=0
cc_480 N_A3_M1017_g N_VPWR_c_699_n 0.00985824f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_481 N_A3_M1013_g N_A_509_392#_c_883_n 0.00100213f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_482 A3 N_A_509_392#_c_883_n 0.00239474f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_483 N_A3_M1013_g N_A_509_392#_c_928_n 0.0033929f $X=7.155 $Y=2.46 $X2=0 $Y2=0
cc_484 N_A3_M1017_g N_A_509_392#_c_928_n 4.45329e-19 $X=7.655 $Y=2.46 $X2=0
+ $Y2=0
cc_485 N_A3_M1013_g N_A_509_392#_c_884_n 0.00669715f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_486 N_A3_M1013_g N_A_509_392#_c_885_n 0.0132272f $X=7.155 $Y=2.46 $X2=0 $Y2=0
cc_487 N_A3_M1017_g N_A_509_392#_c_885_n 0.0132272f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_488 A3 N_A_509_392#_c_885_n 0.045409f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_489 N_A3_c_652_n N_A_509_392#_c_885_n 0.00313888f $X=7.665 $Y=1.615 $X2=0
+ $Y2=0
cc_490 N_A3_M1017_g N_A_509_392#_c_886_n 0.00108119f $X=7.655 $Y=2.46 $X2=0
+ $Y2=0
cc_491 A3 N_A_509_392#_c_886_n 0.0277596f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_492 N_A3_c_652_n N_A_509_392#_c_886_n 0.0016307f $X=7.665 $Y=1.615 $X2=0
+ $Y2=0
cc_493 N_A3_M1013_g N_A_509_392#_c_887_n 6.10838e-19 $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_494 N_A3_M1017_g N_A_509_392#_c_887_n 0.0118584f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_495 N_A3_M1013_g N_A_509_392#_c_936_n 0.00192359f $X=7.155 $Y=2.46 $X2=0
+ $Y2=0
cc_496 N_A3_M1002_g N_VGND_c_991_n 0.00733698f $X=7.14 $Y=0.93 $X2=0 $Y2=0
cc_497 N_A3_M1012_g N_VGND_c_991_n 0.00508523f $X=7.665 $Y=0.93 $X2=0 $Y2=0
cc_498 N_A3_M1002_g N_VGND_c_996_n 0.00351846f $X=7.14 $Y=0.93 $X2=0 $Y2=0
cc_499 N_A3_M1012_g N_VGND_c_997_n 0.00407419f $X=7.665 $Y=0.93 $X2=0 $Y2=0
cc_500 N_A3_M1002_g N_VGND_c_998_n 0.00397821f $X=7.14 $Y=0.93 $X2=0 $Y2=0
cc_501 N_A3_M1012_g N_VGND_c_998_n 0.00473597f $X=7.665 $Y=0.93 $X2=0 $Y2=0
cc_502 N_A3_M1002_g N_A_992_122#_c_1101_n 0.00580529f $X=7.14 $Y=0.93 $X2=0
+ $Y2=0
cc_503 N_A3_M1002_g N_A_992_122#_c_1102_n 0.0128803f $X=7.14 $Y=0.93 $X2=0 $Y2=0
cc_504 N_A3_M1012_g N_A_992_122#_c_1102_n 0.0126425f $X=7.665 $Y=0.93 $X2=0
+ $Y2=0
cc_505 A3 N_A_992_122#_c_1102_n 0.0723776f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_506 N_A3_c_652_n N_A_992_122#_c_1102_n 0.00631331f $X=7.665 $Y=1.615 $X2=0
+ $Y2=0
cc_507 N_A3_M1002_g N_A_992_122#_c_1104_n 8.48859e-19 $X=7.14 $Y=0.93 $X2=0
+ $Y2=0
cc_508 N_A3_M1012_g N_A_992_122#_c_1104_n 0.0076648f $X=7.665 $Y=0.93 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_701_n N_X_c_811_n 7.22336e-19 $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_510 N_VPWR_c_701_n N_X_c_812_n 0.0216434f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_511 N_VPWR_c_701_n N_X_c_816_n 0.00159165f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_512 N_VPWR_c_701_n N_X_c_817_n 0.0309546f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_513 N_VPWR_c_702_n N_X_c_817_n 0.0267028f $X=1.18 $Y=2.295 $X2=0 $Y2=0
cc_514 N_VPWR_c_707_n N_X_c_817_n 0.0109793f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_515 N_VPWR_c_699_n N_X_c_817_n 0.00901959f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_M1004_s N_X_c_830_n 0.0040648f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_517 N_VPWR_c_702_n N_X_c_830_n 0.0189268f $X=1.18 $Y=2.295 $X2=0 $Y2=0
cc_518 N_VPWR_c_702_n N_X_c_818_n 0.0312603f $X=1.18 $Y=2.295 $X2=0 $Y2=0
cc_519 N_VPWR_c_703_n N_X_c_818_n 0.0282236f $X=2.13 $Y=2.405 $X2=0 $Y2=0
cc_520 N_VPWR_c_708_n N_X_c_818_n 0.0133949f $X=1.965 $Y=3.33 $X2=0 $Y2=0
cc_521 N_VPWR_c_699_n N_X_c_818_n 0.0102507f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_522 N_VPWR_c_703_n N_A_509_392#_c_879_n 0.0414286f $X=2.13 $Y=2.405 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_709_n N_A_509_392#_c_880_n 0.0421443f $X=5.21 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_699_n N_A_509_392#_c_880_n 0.0236813f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_703_n N_A_509_392#_c_881_n 0.0121616f $X=2.13 $Y=2.405 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_709_n N_A_509_392#_c_881_n 0.0235512f $X=5.21 $Y=3.33 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_699_n N_A_509_392#_c_881_n 0.0126924f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_704_n N_A_509_392#_c_882_n 0.00883727f $X=5.39 $Y=2.755 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_709_n N_A_509_392#_c_882_n 0.0703102f $X=5.21 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_699_n N_A_509_392#_c_882_n 0.0391428f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_M1010_d N_A_509_392#_c_915_n 0.00735111f $X=5.2 $Y=1.96 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_704_n N_A_509_392#_c_915_n 0.0261161f $X=5.39 $Y=2.755 $X2=0
+ $Y2=0
cc_533 N_VPWR_M1027_s N_A_509_392#_c_920_n 0.00452367f $X=6.285 $Y=1.96 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_705_n N_A_509_392#_c_920_n 0.0197404f $X=6.465 $Y=2.795 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_705_n N_A_509_392#_c_884_n 0.0156521f $X=6.465 $Y=2.795 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_706_n N_A_509_392#_c_884_n 0.0213046f $X=7.38 $Y=2.455 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_711_n N_A_509_392#_c_884_n 0.0133949f $X=7.265 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_699_n N_A_509_392#_c_884_n 0.0102507f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_M1013_s N_A_509_392#_c_885_n 0.00218982f $X=7.245 $Y=1.96 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_706_n N_A_509_392#_c_885_n 0.0167599f $X=7.38 $Y=2.455 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_706_n N_A_509_392#_c_887_n 0.0266615f $X=7.38 $Y=2.455 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_712_n N_A_509_392#_c_887_n 0.014549f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_c_699_n N_A_509_392#_c_887_n 0.0119743f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_709_n N_A_509_392#_c_888_n 0.0235512f $X=5.21 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_699_n N_A_509_392#_c_888_n 0.0126924f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_705_n N_A_509_392#_c_933_n 0.0215129f $X=6.465 $Y=2.795 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_710_n N_A_509_392#_c_933_n 0.00883515f $X=6.285 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_699_n N_A_509_392#_c_933_n 0.0112505f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_X_c_810_n N_VGND_M1007_s 0.00389177f $X=0.355 $Y=1.055 $X2=-0.19
+ $Y2=-0.245
cc_550 N_X_c_834_n N_VGND_M1008_s 0.0071582f $X=1.57 $Y=1.055 $X2=0 $Y2=0
cc_551 N_X_c_819_n N_VGND_c_987_n 0.00246556f $X=0.615 $Y=1.055 $X2=0 $Y2=0
cc_552 N_X_c_810_n N_VGND_c_987_n 0.020861f $X=0.355 $Y=1.055 $X2=0 $Y2=0
cc_553 N_X_c_813_n N_VGND_c_987_n 0.0146425f $X=0.715 $Y=0.575 $X2=0 $Y2=0
cc_554 N_X_c_813_n N_VGND_c_988_n 0.015086f $X=0.715 $Y=0.575 $X2=0 $Y2=0
cc_555 N_X_c_834_n N_VGND_c_988_n 0.0282307f $X=1.57 $Y=1.055 $X2=0 $Y2=0
cc_556 N_X_c_814_n N_VGND_c_988_n 0.0131993f $X=1.735 $Y=0.595 $X2=0 $Y2=0
cc_557 N_X_c_814_n N_VGND_c_989_n 0.0195142f $X=1.735 $Y=0.595 $X2=0 $Y2=0
cc_558 N_X_c_813_n N_VGND_c_994_n 0.00729225f $X=0.715 $Y=0.575 $X2=0 $Y2=0
cc_559 N_X_c_814_n N_VGND_c_995_n 0.0109286f $X=1.735 $Y=0.595 $X2=0 $Y2=0
cc_560 N_X_c_813_n N_VGND_c_998_n 0.00722011f $X=0.715 $Y=0.575 $X2=0 $Y2=0
cc_561 N_X_c_814_n N_VGND_c_998_n 0.011467f $X=1.735 $Y=0.595 $X2=0 $Y2=0
cc_562 N_A_509_392#_c_886_n N_A_992_122#_c_1102_n 3.53329e-19 $X=7.88 $Y=2.12
+ $X2=0 $Y2=0
cc_563 N_A_509_392#_c_883_n N_A_992_122#_c_1103_n 0.00582992f $X=6.93 $Y=2.12
+ $X2=0 $Y2=0
cc_564 N_VGND_c_998_n N_A_587_110#_c_1079_n 0.0025026f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_565 N_VGND_c_990_n N_A_992_122#_c_1098_n 0.0363805f $X=4.67 $Y=0.755 $X2=0
+ $Y2=0
cc_566 N_VGND_c_991_n N_A_992_122#_c_1099_n 0.0134785f $X=7.365 $Y=0.755 $X2=0
+ $Y2=0
cc_567 N_VGND_c_996_n N_A_992_122#_c_1099_n 0.117712f $X=7.19 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_998_n N_A_992_122#_c_1099_n 0.067988f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_569 N_VGND_c_990_n N_A_992_122#_c_1100_n 0.0135234f $X=4.67 $Y=0.755 $X2=0
+ $Y2=0
cc_570 N_VGND_c_996_n N_A_992_122#_c_1100_n 0.0179316f $X=7.19 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_998_n N_A_992_122#_c_1100_n 0.00972129f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_991_n N_A_992_122#_c_1101_n 0.0338465f $X=7.365 $Y=0.755 $X2=0
+ $Y2=0
cc_573 N_VGND_M1002_s N_A_992_122#_c_1102_n 0.00296556f $X=7.215 $Y=0.61 $X2=0
+ $Y2=0
cc_574 N_VGND_c_991_n N_A_992_122#_c_1102_n 0.0220515f $X=7.365 $Y=0.755 $X2=0
+ $Y2=0
cc_575 N_VGND_c_991_n N_A_992_122#_c_1104_n 0.0131817f $X=7.365 $Y=0.755 $X2=0
+ $Y2=0
cc_576 N_VGND_c_997_n N_A_992_122#_c_1104_n 0.00725695f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_c_998_n N_A_992_122#_c_1104_n 0.0102594f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_578 N_A_992_122#_c_1099_n N_A_1079_122#_c_1146_n 0.0478568f $X=6.74 $Y=0.34
+ $X2=0 $Y2=0
cc_579 N_A_992_122#_c_1098_n N_A_1079_122#_c_1147_n 0.0123866f $X=5.105 $Y=0.765
+ $X2=0 $Y2=0
cc_580 N_A_992_122#_c_1099_n N_A_1079_122#_c_1147_n 0.0185146f $X=6.74 $Y=0.34
+ $X2=0 $Y2=0
cc_581 N_A_992_122#_c_1099_n N_A_1079_122#_c_1148_n 0.0197406f $X=6.74 $Y=0.34
+ $X2=0 $Y2=0
cc_582 N_A_992_122#_c_1101_n N_A_1079_122#_c_1148_n 0.00649205f $X=6.905
+ $Y=0.755 $X2=0 $Y2=0
cc_583 N_A_992_122#_c_1103_n N_A_1079_122#_c_1148_n 0.00756924f $X=6.99 $Y=1.185
+ $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__a221oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_297_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2432e+12p pd=1.118e+07u as=8.848e+11p ps=8.3e+06u
M1001 VGND B2 a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=7.696e+11p pd=6.52e+06u as=4.44e+11p ps=4.16e+06u
M1002 VPWR A2 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_293_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.362e+11p ps=8.18e+06u
M1004 a_675_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=7.03e+11p pd=4.86e+06u as=0p ps=0u
M1005 a_297_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A1 a_675_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_675_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_293_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_29_368# B2 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1872e+12p pd=1.108e+07u as=0p ps=0u
M1011 a_297_368# B2 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_29_368# B1 a_297_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_675_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1017 a_29_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_297_368# B1 a_29_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__o22ai_1.pex.spice
* Created: Fri Aug 28 17:58:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O22AI_1%B1 1 3 6 8 13
r28 11 13 36.4894 $w=2.84e-07 $l=2.15e-07 $layer=POLY_cond $X=0.28 $Y=1.385
+ $X2=0.495 $Y2=1.385
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.385 $X2=0.28 $Y2=1.385
r30 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=1.295 $X2=0.28
+ $Y2=1.385
r31 4 13 23.7606 $w=2.84e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.635 $Y=1.55
+ $X2=0.495 $Y2=1.385
r32 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.635 $Y=1.55
+ $X2=0.635 $Y2=2.4
r33 1 13 17.6835 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r34 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%B2 3 7 9 12 13
c31 3 0 9.97888e-20 $X=1.055 $Y=2.4
r32 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.13 $Y2=1.68
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.13 $Y2=1.35
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.515 $X2=1.13 $Y2=1.515
r35 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.515
r36 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.22 $Y=0.74 $X2=1.22
+ $Y2=1.35
r37 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.055 $Y=2.4
+ $X2=1.055 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%A2 3 7 9 12 13
c39 13 0 9.97888e-20 $X=1.7 $Y=1.515
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.515
+ $X2=1.7 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.515
+ $X2=1.7 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.515 $X2=1.7 $Y2=1.515
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.7
+ $Y2=1.515
r44 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.72 $Y=0.74 $X2=1.72
+ $Y2=1.35
r45 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.625 $Y=2.4
+ $X2=1.625 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%A1 3 7 10 11 12 16
r32 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.61
+ $Y=1.465 $X2=2.61 $Y2=1.465
r33 12 17 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.54 $X2=2.61
+ $Y2=1.54
r34 11 17 11.2132 $w=4.78e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=1.54
+ $X2=2.61 $Y2=1.54
r35 9 16 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.365 $Y=1.465
+ $X2=2.61 $Y2=1.465
r36 9 10 3.90195 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.365 $Y=1.465
+ $X2=2.235 $Y2=1.465
r37 5 10 34.7346 $w=1.65e-07 $l=1.90526e-07 $layer=POLY_cond $X=2.29 $Y=1.3
+ $X2=2.235 $Y2=1.465
r38 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.29 $Y=1.3 $X2=2.29
+ $Y2=0.74
r39 1 10 34.7346 $w=1.65e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.195 $Y=1.63
+ $X2=2.235 $Y2=1.465
r40 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.195 $Y=1.63
+ $X2=2.195 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%VPWR 1 2 7 9 15 19 20 21 22 33
r26 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r29 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 27 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 24 35 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r34 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 22 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 22 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 20 29 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.42 $Y2=3.33
r39 19 32 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=2.42 $Y2=3.33
r41 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.42 $Y=2.115 $X2=2.42
+ $Y2=2.815
r42 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=3.245
+ $X2=2.42 $Y2=3.33
r43 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.42 $Y=3.245
+ $X2=2.42 $Y2=2.815
r44 9 12 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.29 $Y=1.985
+ $X2=0.29 $Y2=2.815
r45 7 35 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.227 $Y2=3.33
r46 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.815
r47 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.84 $X2=2.42 $Y2=2.815
r48 2 15 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.84 $X2=2.42 $Y2=2.115
r49 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r50 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%Y 1 2 10 13 14 18 19
r31 18 19 12.4206 $w=9.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.087 $Y=2.115
+ $X2=1.087 $Y2=1.95
r32 14 25 0.527568 $w=9.23e-07 $l=4e-08 $layer=LI1_cond $X=1.087 $Y=2.775
+ $X2=1.087 $Y2=2.815
r33 13 14 4.88 $w=9.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.087 $Y=2.405
+ $X2=1.087 $Y2=2.775
r34 13 18 3.82486 $w=9.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.087 $Y=2.405
+ $X2=1.087 $Y2=2.115
r35 12 19 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r36 10 12 12.5466 $w=4.48e-07 $l=2.9e-07 $layer=LI1_cond $X=0.84 $Y=0.84
+ $X2=0.84 $Y2=1.13
r37 2 25 400 $w=1.7e-07 $l=1.06577e-06 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.335 $Y2=2.815
r38 2 18 400 $w=1.7e-07 $l=3.57596e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.335 $Y2=2.115
r39 1 10 182 $w=1.7e-07 $l=5.95693e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.855 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%A_27_74# 1 2 3 12 14 15 19 20 21 24
r41 22 24 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.505 $Y=0.96
+ $X2=2.505 $Y2=0.515
r42 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.34 $Y=1.045
+ $X2=2.505 $Y2=0.96
r43 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.34 $Y=1.045
+ $X2=1.67 $Y2=1.045
r44 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.505 $Y=0.96
+ $X2=1.67 $Y2=1.045
r45 17 19 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.505 $Y=0.96
+ $X2=1.505 $Y2=0.515
r46 16 19 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.505 $Y=0.485
+ $X2=1.505 $Y2=0.515
r47 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.34 $Y=0.4
+ $X2=1.505 $Y2=0.485
r48 14 15 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.34 $Y=0.4
+ $X2=0.445 $Y2=0.4
r49 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.485
+ $X2=0.445 $Y2=0.4
r50 10 12 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.28 $Y=0.485 $X2=0.28
+ $Y2=0.515
r51 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.37 $X2=2.505 $Y2=0.515
r52 2 19 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.295
+ $Y=0.37 $X2=1.505 $Y2=0.515
r53 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O22AI_1%VGND 1 6 9 10 11 21 22
r25 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r26 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r27 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r28 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r29 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r31 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.24
+ $Y2=0
r32 9 18 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=1.68
+ $Y2=0
r33 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=0 $X2=2.005
+ $Y2=0
r34 8 21 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.64
+ $Y2=0
r35 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.005
+ $Y2=0
r36 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0
r37 4 6 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0.625
r38 1 6 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=1.795
+ $Y=0.37 $X2=2.005 $Y2=0.625
.ends


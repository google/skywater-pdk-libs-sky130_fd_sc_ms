* File: sky130_fd_sc_ms__a2111oi_4.pxi.spice
* Created: Wed Sep  2 11:49:52 2020
* 
x_PM_SKY130_FD_SC_MS__A2111OI_4%D1 N_D1_M1021_g N_D1_M1022_g N_D1_M1026_g
+ N_D1_c_142_n N_D1_M1017_g N_D1_c_143_n N_D1_M1029_g N_D1_M1031_g D1 D1 D1
+ N_D1_c_145_n N_D1_c_146_n PM_SKY130_FD_SC_MS__A2111OI_4%D1
x_PM_SKY130_FD_SC_MS__A2111OI_4%C1 N_C1_M1016_g N_C1_c_212_n N_C1_M1000_g
+ N_C1_M1025_g N_C1_M1002_g N_C1_M1004_g N_C1_M1006_g C1 C1 N_C1_c_210_n
+ N_C1_c_211_n PM_SKY130_FD_SC_MS__A2111OI_4%C1
x_PM_SKY130_FD_SC_MS__A2111OI_4%B1 N_B1_M1013_g N_B1_M1019_g N_B1_M1012_g
+ N_B1_M1014_g N_B1_M1020_g N_B1_M1024_g B1 B1 B1 N_B1_c_287_n N_B1_c_288_n
+ PM_SKY130_FD_SC_MS__A2111OI_4%B1
x_PM_SKY130_FD_SC_MS__A2111OI_4%A1 N_A1_M1001_g N_A1_M1009_g N_A1_M1003_g
+ N_A1_M1011_g N_A1_M1028_g N_A1_M1030_g N_A1_M1032_g N_A1_M1033_g A1 A1 A1
+ N_A1_c_360_n PM_SKY130_FD_SC_MS__A2111OI_4%A1
x_PM_SKY130_FD_SC_MS__A2111OI_4%A2 N_A2_M1007_g N_A2_M1005_g N_A2_M1018_g
+ N_A2_M1008_g N_A2_M1023_g N_A2_M1010_g N_A2_M1027_g N_A2_M1015_g A2 A2 A2
+ N_A2_c_445_n N_A2_c_440_n PM_SKY130_FD_SC_MS__A2111OI_4%A2
x_PM_SKY130_FD_SC_MS__A2111OI_4%A_29_368# N_A_29_368#_M1021_s
+ N_A_29_368#_M1022_s N_A_29_368#_M1031_s N_A_29_368#_M1002_s
+ N_A_29_368#_M1006_s N_A_29_368#_c_511_n N_A_29_368#_c_512_n
+ N_A_29_368#_c_513_n N_A_29_368#_c_546_p N_A_29_368#_c_514_n
+ N_A_29_368#_c_521_n N_A_29_368#_c_522_n N_A_29_368#_c_528_n
+ N_A_29_368#_c_555_p N_A_29_368#_c_532_n N_A_29_368#_c_515_n
+ N_A_29_368#_c_536_n N_A_29_368#_c_516_n
+ PM_SKY130_FD_SC_MS__A2111OI_4%A_29_368#
x_PM_SKY130_FD_SC_MS__A2111OI_4%Y N_Y_M1017_d N_Y_M1016_d N_Y_M1013_d
+ N_Y_M1009_s N_Y_M1030_s N_Y_M1021_d N_Y_M1026_d N_Y_c_570_n N_Y_c_571_n
+ N_Y_c_583_n N_Y_c_592_n N_Y_c_584_n N_Y_c_600_n N_Y_c_572_n N_Y_c_604_n
+ N_Y_c_573_n N_Y_c_574_n N_Y_c_575_n N_Y_c_576_n N_Y_c_585_n N_Y_c_610_n
+ N_Y_c_577_n N_Y_c_578_n N_Y_c_579_n N_Y_c_580_n N_Y_c_581_n Y Y N_Y_c_587_n Y
+ PM_SKY130_FD_SC_MS__A2111OI_4%Y
x_PM_SKY130_FD_SC_MS__A2111OI_4%A_477_368# N_A_477_368#_M1000_d
+ N_A_477_368#_M1004_d N_A_477_368#_M1012_d N_A_477_368#_M1020_d
+ N_A_477_368#_c_701_n N_A_477_368#_c_695_n N_A_477_368#_c_696_n
+ N_A_477_368#_c_707_n N_A_477_368#_c_697_n N_A_477_368#_c_714_n
+ N_A_477_368#_c_698_n N_A_477_368#_c_720_n N_A_477_368#_c_699_n
+ N_A_477_368#_c_700_n PM_SKY130_FD_SC_MS__A2111OI_4%A_477_368#
x_PM_SKY130_FD_SC_MS__A2111OI_4%A_853_368# N_A_853_368#_M1012_s
+ N_A_853_368#_M1014_s N_A_853_368#_M1024_s N_A_853_368#_M1003_s
+ N_A_853_368#_M1032_s N_A_853_368#_M1008_s N_A_853_368#_M1015_s
+ N_A_853_368#_c_757_n N_A_853_368#_c_758_n N_A_853_368#_c_767_n
+ N_A_853_368#_c_813_n N_A_853_368#_c_771_n N_A_853_368#_c_759_n
+ N_A_853_368#_c_777_n N_A_853_368#_c_760_n N_A_853_368#_c_781_n
+ N_A_853_368#_c_761_n N_A_853_368#_c_788_n N_A_853_368#_c_762_n
+ N_A_853_368#_c_796_n N_A_853_368#_c_763_n N_A_853_368#_c_764_n
+ N_A_853_368#_c_775_n N_A_853_368#_c_785_n N_A_853_368#_c_787_n
+ N_A_853_368#_c_802_n PM_SKY130_FD_SC_MS__A2111OI_4%A_853_368#
x_PM_SKY130_FD_SC_MS__A2111OI_4%VPWR N_VPWR_M1001_d N_VPWR_M1028_d
+ N_VPWR_M1005_d N_VPWR_M1010_d N_VPWR_c_845_n N_VPWR_c_846_n N_VPWR_c_847_n
+ N_VPWR_c_848_n N_VPWR_c_849_n N_VPWR_c_850_n N_VPWR_c_851_n VPWR
+ N_VPWR_c_852_n N_VPWR_c_853_n N_VPWR_c_854_n N_VPWR_c_844_n N_VPWR_c_856_n
+ N_VPWR_c_857_n N_VPWR_c_858_n PM_SKY130_FD_SC_MS__A2111OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A2111OI_4%VGND N_VGND_M1017_s N_VGND_M1029_s
+ N_VGND_M1025_s N_VGND_M1019_s N_VGND_M1007_s N_VGND_M1023_s N_VGND_c_959_n
+ N_VGND_c_960_n N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n N_VGND_c_964_n
+ N_VGND_c_965_n N_VGND_c_966_n VGND N_VGND_c_967_n N_VGND_c_968_n
+ N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n
+ N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n
+ PM_SKY130_FD_SC_MS__A2111OI_4%VGND
x_PM_SKY130_FD_SC_MS__A2111OI_4%A_1228_74# N_A_1228_74#_M1009_d
+ N_A_1228_74#_M1011_d N_A_1228_74#_M1033_d N_A_1228_74#_M1018_d
+ N_A_1228_74#_M1027_d N_A_1228_74#_c_1062_n N_A_1228_74#_c_1063_n
+ N_A_1228_74#_c_1064_n N_A_1228_74#_c_1065_n N_A_1228_74#_c_1066_n
+ N_A_1228_74#_c_1067_n N_A_1228_74#_c_1068_n N_A_1228_74#_c_1069_n
+ N_A_1228_74#_c_1070_n N_A_1228_74#_c_1071_n N_A_1228_74#_c_1072_n
+ PM_SKY130_FD_SC_MS__A2111OI_4%A_1228_74#
cc_1 VNB N_D1_M1021_g 0.00630099f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_D1_M1022_g 0.00579577f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_3 VNB N_D1_M1026_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_4 VNB N_D1_c_142_n 0.0208421f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.22
cc_5 VNB N_D1_c_143_n 0.0162859f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.22
cc_6 VNB N_D1_M1031_g 0.00610499f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_7 VNB N_D1_c_145_n 0.0126583f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_8 VNB N_D1_c_146_n 0.102905f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.385
cc_9 VNB N_C1_M1016_g 0.0218891f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_C1_M1025_g 0.0273339f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_11 VNB N_C1_c_210_n 0.0953563f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.385
cc_12 VNB N_C1_c_211_n 0.00205555f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_13 VNB N_B1_M1013_g 0.0288572f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_14 VNB N_B1_M1019_g 0.0305521f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_15 VNB N_B1_c_287_n 0.124966f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_16 VNB N_B1_c_288_n 0.00264168f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.385
cc_17 VNB N_A1_M1009_g 0.0326041f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_18 VNB N_A1_M1011_g 0.0232165f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_19 VNB N_A1_M1030_g 0.0233981f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A1_M1033_g 0.0240711f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_21 VNB A1 0.00465397f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.385
cc_22 VNB N_A1_c_360_n 0.0706289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1007_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_24 VNB N_A2_M1018_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_25 VNB N_A2_M1023_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.55
cc_26 VNB N_A2_M1027_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_c_440_n 0.0833513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_570_n 0.0224339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_571_n 0.0130653f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_30 VNB N_Y_c_572_n 0.00210053f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_31 VNB N_Y_c_573_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_574_n 0.0118592f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.365
cc_33 VNB N_Y_c_575_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_576_n 0.00249052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_577_n 0.00242779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_578_n 0.00507892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_579_n 0.0762531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_580_n 0.00228886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_581_n 0.00250929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB Y 0.0375295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_844_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_959_n 0.0211662f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_43 VNB N_VGND_c_960_n 0.00259973f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_44 VNB N_VGND_c_961_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_962_n 0.0264859f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_46 VNB N_VGND_c_963_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.385
cc_47 VNB N_VGND_c_964_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_48 VNB N_VGND_c_965_n 0.0151212f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.385
cc_49 VNB N_VGND_c_966_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_50 VNB N_VGND_c_967_n 0.0346017f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.365
cc_51 VNB N_VGND_c_968_n 0.0938841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_969_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_970_n 0.0197776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_971_n 0.573484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_972_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_973_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_974_n 0.037009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_975_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_976_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_977_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1228_74#_c_1062_n 0.00310413f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=0.74
cc_62 VNB N_A_1228_74#_c_1063_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_63 VNB N_A_1228_74#_c_1064_n 0.00460553f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.21
cc_64 VNB N_A_1228_74#_c_1065_n 0.00406794f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.21
cc_65 VNB N_A_1228_74#_c_1066_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1228_74#_c_1067_n 0.0158169f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_67 VNB N_A_1228_74#_c_1068_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.395
+ $Y2=1.385
cc_68 VNB N_A_1228_74#_c_1069_n 0.0157537f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_69 VNB N_A_1228_74#_c_1070_n 0.00301978f $X=-0.19 $Y=-0.245 $X2=1.845
+ $Y2=1.385
cc_70 VNB N_A_1228_74#_c_1071_n 0.0017805f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_71 VNB N_A_1228_74#_c_1072_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.365
cc_72 VPB N_D1_M1021_g 0.0248758f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_73 VPB N_D1_M1022_g 0.0205287f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_74 VPB N_D1_M1026_g 0.0205309f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_75 VPB N_D1_M1031_g 0.0219013f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_76 VPB N_C1_c_212_n 0.0162581f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.55
cc_77 VPB N_C1_M1002_g 0.0196343f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_78 VPB N_C1_M1004_g 0.0182882f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_79 VPB N_C1_M1006_g 0.0233819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_C1_c_210_n 0.0200303f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.385
cc_81 VPB N_C1_c_211_n 0.00813053f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_82 VPB N_B1_M1012_g 0.0249106f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_83 VPB N_B1_M1014_g 0.0196343f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_84 VPB N_B1_M1020_g 0.0196343f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.55
cc_85 VPB N_B1_M1024_g 0.0204768f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_86 VPB N_B1_c_287_n 0.0305745f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_87 VPB N_B1_c_288_n 0.0126405f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.385
cc_88 VPB N_A1_M1001_g 0.0208086f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_89 VPB N_A1_M1003_g 0.0198928f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_90 VPB N_A1_M1028_g 0.0198928f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.55
cc_91 VPB N_A1_M1032_g 0.0202413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB A1 0.00976217f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.385
cc_93 VPB N_A1_c_360_n 0.0116093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A2_M1005_g 0.0207949f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_95 VPB N_A2_M1008_g 0.020498f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_96 VPB N_A2_M1010_g 0.0204973f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_97 VPB N_A2_M1015_g 0.0281481f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.385
cc_98 VPB N_A2_c_445_n 0.00755622f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.365
cc_99 VPB N_A2_c_440_n 0.0124528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_29_368#_c_511_n 0.0325715f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_101 VPB N_A_29_368#_c_512_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_102 VPB N_A_29_368#_c_513_n 0.00932809f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_103 VPB N_A_29_368#_c_514_n 0.00423682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_29_368#_c_515_n 0.00123754f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.385
cc_105 VPB N_A_29_368#_c_516_n 0.01417f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.365
cc_106 VPB N_Y_c_583_n 0.00168332f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_107 VPB N_Y_c_584_n 0.00530403f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.385
cc_108 VPB N_Y_c_585_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB Y 0.00287511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_Y_c_587_n 0.00758256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_477_368#_c_695_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_112 VPB N_A_477_368#_c_696_n 0.00247907f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_113 VPB N_A_477_368#_c_697_n 0.0160187f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_114 VPB N_A_477_368#_c_698_n 0.00388794f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_115 VPB N_A_477_368#_c_699_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.385
cc_116 VPB N_A_477_368#_c_700_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.385
cc_117 VPB N_A_853_368#_c_757_n 0.00170943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_853_368#_c_758_n 0.00536257f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_119 VPB N_A_853_368#_c_759_n 0.00179576f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.385
cc_120 VPB N_A_853_368#_c_760_n 0.00179594f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.385
cc_121 VPB N_A_853_368#_c_761_n 0.00179594f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.365
cc_122 VPB N_A_853_368#_c_762_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_853_368#_c_763_n 0.0185501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_853_368#_c_764_n 0.0345796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_845_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_126 VPB N_VPWR_c_846_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_127 VPB N_VPWR_c_847_n 0.00261791f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_128 VPB N_VPWR_c_848_n 0.0048755f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_129 VPB N_VPWR_c_849_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_130 VPB N_VPWR_c_850_n 0.152843f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.385
cc_131 VPB N_VPWR_c_851_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.385
cc_132 VPB N_VPWR_c_852_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.385
cc_133 VPB N_VPWR_c_853_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_854_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_844_n 0.100814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_856_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_857_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_858_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 N_D1_c_143_n N_C1_M1016_g 0.0174718f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_140 N_D1_c_145_n N_C1_M1016_g 0.00131191f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_141 N_D1_M1031_g N_C1_c_210_n 0.0155982f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_142 N_D1_c_145_n N_C1_c_210_n 3.91262e-19 $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_143 N_D1_c_146_n N_C1_c_210_n 0.0299006f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_144 N_D1_M1031_g N_C1_c_211_n 4.54361e-19 $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_145 N_D1_c_145_n N_C1_c_211_n 0.00980746f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_146 N_D1_c_146_n N_C1_c_211_n 0.00152517f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_147 N_D1_M1021_g N_A_29_368#_c_512_n 0.0149445f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_148 N_D1_M1022_g N_A_29_368#_c_512_n 0.0140221f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_149 N_D1_M1026_g N_A_29_368#_c_514_n 0.0140221f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_150 N_D1_M1031_g N_A_29_368#_c_514_n 0.0135505f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_151 N_D1_M1031_g N_A_29_368#_c_521_n 0.0034531f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_152 N_D1_M1026_g N_A_29_368#_c_522_n 7.23726e-19 $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_153 N_D1_M1031_g N_A_29_368#_c_522_n 0.011184f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_154 N_D1_c_142_n N_Y_c_570_n 0.0116578f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_155 N_D1_c_145_n N_Y_c_570_n 0.0722866f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_156 N_D1_c_146_n N_Y_c_570_n 0.0106615f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_157 N_D1_M1021_g N_Y_c_583_n 0.0184993f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_158 N_D1_M1021_g N_Y_c_592_n 0.0185855f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_159 N_D1_M1022_g N_Y_c_592_n 0.0139272f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_160 N_D1_M1026_g N_Y_c_592_n 6.45773e-19 $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_161 N_D1_M1022_g N_Y_c_584_n 0.0128923f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_162 N_D1_M1026_g N_Y_c_584_n 0.014881f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_163 N_D1_M1031_g N_Y_c_584_n 0.00278382f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_164 N_D1_c_145_n N_Y_c_584_n 0.0631462f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_165 N_D1_c_146_n N_Y_c_584_n 0.00411446f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_166 N_D1_M1022_g N_Y_c_600_n 6.48223e-19 $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_167 N_D1_M1026_g N_Y_c_600_n 0.0133704f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_168 N_D1_c_142_n N_Y_c_572_n 4.50863e-19 $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_169 N_D1_c_143_n N_Y_c_572_n 4.50863e-19 $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_170 N_D1_c_143_n N_Y_c_604_n 0.00957073f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_171 N_D1_c_145_n N_Y_c_604_n 0.0131073f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_172 N_D1_M1021_g N_Y_c_585_n 0.00228751f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_173 N_D1_M1022_g N_Y_c_585_n 0.00228751f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_174 N_D1_c_145_n N_Y_c_585_n 0.0277828f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_175 N_D1_c_146_n N_Y_c_585_n 0.00209661f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_176 N_D1_c_145_n N_Y_c_610_n 0.0146818f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_177 N_D1_c_146_n N_Y_c_610_n 7.07126e-19 $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_178 N_D1_c_145_n Y 0.0267576f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_179 N_D1_c_146_n Y 0.0172295f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_180 N_D1_M1021_g N_VPWR_c_850_n 0.00333926f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_181 N_D1_M1022_g N_VPWR_c_850_n 0.00333926f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_182 N_D1_M1026_g N_VPWR_c_850_n 0.00333926f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_183 N_D1_M1031_g N_VPWR_c_850_n 0.00333896f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_184 N_D1_M1021_g N_VPWR_c_844_n 0.00426394f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_185 N_D1_M1022_g N_VPWR_c_844_n 0.00422687f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_186 N_D1_M1026_g N_VPWR_c_844_n 0.00422687f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_187 N_D1_M1031_g N_VPWR_c_844_n 0.00422796f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_188 N_D1_c_142_n N_VGND_c_959_n 0.00850375f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_189 N_D1_c_143_n N_VGND_c_959_n 3.67997e-19 $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_190 N_D1_c_142_n N_VGND_c_960_n 3.67997e-19 $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_191 N_D1_c_143_n N_VGND_c_960_n 0.0074045f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_192 N_D1_c_142_n N_VGND_c_965_n 0.00383152f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_193 N_D1_c_143_n N_VGND_c_965_n 0.00383152f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_194 N_D1_c_142_n N_VGND_c_971_n 0.00383967f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_195 N_D1_c_143_n N_VGND_c_971_n 0.00383967f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_196 N_C1_c_210_n N_B1_M1013_g 0.01353f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_197 N_C1_c_210_n N_B1_c_287_n 0.00780189f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_198 N_C1_c_211_n N_B1_c_287_n 0.00157841f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_199 N_C1_c_210_n N_B1_c_288_n 0.00440879f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_200 N_C1_c_212_n N_A_29_368#_c_514_n 0.00347444f $X=2.295 $Y=1.77 $X2=0 $Y2=0
cc_201 N_C1_c_212_n N_A_29_368#_c_521_n 0.00102889f $X=2.295 $Y=1.77 $X2=0 $Y2=0
cc_202 N_C1_c_212_n N_A_29_368#_c_522_n 0.0111124f $X=2.295 $Y=1.77 $X2=0 $Y2=0
cc_203 N_C1_M1002_g N_A_29_368#_c_522_n 4.41999e-19 $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_204 N_C1_c_212_n N_A_29_368#_c_528_n 0.012931f $X=2.295 $Y=1.77 $X2=0 $Y2=0
cc_205 N_C1_M1002_g N_A_29_368#_c_528_n 0.0142562f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_206 N_C1_c_210_n N_A_29_368#_c_528_n 4.87549e-19 $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_207 N_C1_c_211_n N_A_29_368#_c_528_n 0.0422425f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_208 N_C1_M1004_g N_A_29_368#_c_532_n 0.0142562f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_209 N_C1_M1006_g N_A_29_368#_c_532_n 0.0163597f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_210 N_C1_c_210_n N_A_29_368#_c_532_n 5.25345e-19 $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_211 N_C1_c_211_n N_A_29_368#_c_532_n 0.0293818f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_212 N_C1_c_210_n N_A_29_368#_c_536_n 5.54061e-19 $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_213 N_C1_c_211_n N_A_29_368#_c_536_n 0.0170101f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_214 N_C1_M1004_g N_A_29_368#_c_516_n 6.1989e-19 $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_215 N_C1_M1006_g N_A_29_368#_c_516_n 0.00579521f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_216 N_C1_c_211_n N_Y_c_584_n 0.00219619f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_217 N_C1_M1016_g N_Y_c_604_n 0.0108637f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_218 N_C1_c_211_n N_Y_c_604_n 0.00539983f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_219 N_C1_M1016_g N_Y_c_573_n 3.97481e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_220 N_C1_M1025_g N_Y_c_573_n 0.00615586f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_221 N_C1_M1025_g N_Y_c_574_n 0.0142398f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_222 N_C1_c_210_n N_Y_c_574_n 0.0290405f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_223 N_C1_c_211_n N_Y_c_574_n 0.0662651f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_224 N_C1_M1016_g N_Y_c_577_n 0.00177693f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_225 N_C1_M1025_g N_Y_c_577_n 0.00906122f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_226 N_C1_c_210_n N_Y_c_577_n 0.00264009f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_227 N_C1_c_211_n N_Y_c_577_n 0.0211949f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_228 N_C1_M1002_g N_A_477_368#_c_701_n 0.00861945f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_229 N_C1_M1004_g N_A_477_368#_c_701_n 5.55068e-19 $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_230 N_C1_M1002_g N_A_477_368#_c_695_n 0.0116345f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_231 N_C1_M1004_g N_A_477_368#_c_695_n 0.0115958f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_232 N_C1_c_212_n N_A_477_368#_c_696_n 0.00100838f $X=2.295 $Y=1.77 $X2=0
+ $Y2=0
cc_233 N_C1_M1002_g N_A_477_368#_c_696_n 0.001619f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_234 N_C1_M1002_g N_A_477_368#_c_707_n 5.53268e-19 $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_235 N_C1_M1004_g N_A_477_368#_c_707_n 0.00891111f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_236 N_C1_M1006_g N_A_477_368#_c_707_n 0.0133813f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_237 N_C1_M1006_g N_A_477_368#_c_697_n 0.0137576f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_238 N_C1_M1004_g N_A_477_368#_c_699_n 0.00194226f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_239 N_C1_M1006_g N_A_477_368#_c_699_n 0.00194226f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_240 N_C1_c_212_n N_VPWR_c_850_n 0.00517089f $X=2.295 $Y=1.77 $X2=0 $Y2=0
cc_241 N_C1_M1002_g N_VPWR_c_850_n 0.00333896f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_242 N_C1_M1004_g N_VPWR_c_850_n 0.00333896f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_243 N_C1_M1006_g N_VPWR_c_850_n 0.00333896f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_244 N_C1_c_212_n N_VPWR_c_844_n 0.00978686f $X=2.295 $Y=1.77 $X2=0 $Y2=0
cc_245 N_C1_M1002_g N_VPWR_c_844_n 0.00422685f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_246 N_C1_M1004_g N_VPWR_c_844_n 0.00422685f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_247 N_C1_M1006_g N_VPWR_c_844_n 0.00427818f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_248 N_C1_M1016_g N_VGND_c_960_n 0.00766594f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_249 N_C1_M1025_g N_VGND_c_960_n 4.39708e-19 $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_250 N_C1_M1016_g N_VGND_c_971_n 0.00383967f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_251 N_C1_M1025_g N_VGND_c_971_n 0.00825037f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_252 N_C1_M1016_g N_VGND_c_973_n 0.00383152f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_253 N_C1_M1025_g N_VGND_c_973_n 0.00434272f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_254 N_C1_M1025_g N_VGND_c_974_n 0.00597094f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B1_M1024_g N_A1_M1001_g 0.0148524f $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B1_c_287_n A1 4.61559e-19 $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_257 N_B1_c_288_n A1 0.0190385f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_258 N_B1_c_287_n N_A1_c_360_n 0.0148524f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_259 N_B1_c_288_n N_A1_c_360_n 0.00189297f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_260 N_B1_M1012_g N_A_29_368#_c_516_n 0.00209241f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B1_c_287_n N_A_29_368#_c_516_n 0.00251593f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_262 N_B1_M1013_g N_Y_c_574_n 0.0149534f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_263 N_B1_M1013_g N_Y_c_575_n 0.0118293f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_264 N_B1_M1019_g N_Y_c_575_n 3.97481e-19 $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_265 N_B1_M1013_g N_Y_c_578_n 0.0040828f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B1_c_287_n N_Y_c_578_n 0.00423267f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_267 N_B1_c_288_n N_Y_c_578_n 0.00386581f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_268 N_B1_M1019_g N_Y_c_579_n 0.0166073f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B1_c_287_n N_Y_c_579_n 0.0398662f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_270 N_B1_c_288_n N_Y_c_579_n 0.135914f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_271 N_B1_M1012_g N_A_477_368#_c_697_n 0.0137576f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_272 N_B1_M1012_g N_A_477_368#_c_714_n 0.0135563f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_273 N_B1_M1014_g N_A_477_368#_c_714_n 0.00908611f $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_274 N_B1_M1020_g N_A_477_368#_c_714_n 5.53268e-19 $X=5.535 $Y=2.4 $X2=0 $Y2=0
cc_275 N_B1_M1014_g N_A_477_368#_c_698_n 0.0116345f $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_276 N_B1_M1020_g N_A_477_368#_c_698_n 0.0135768f $X=5.535 $Y=2.4 $X2=0 $Y2=0
cc_277 N_B1_M1024_g N_A_477_368#_c_698_n 0.0041969f $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_278 N_B1_M1014_g N_A_477_368#_c_720_n 5.53268e-19 $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_279 N_B1_M1020_g N_A_477_368#_c_720_n 0.00908611f $X=5.535 $Y=2.4 $X2=0 $Y2=0
cc_280 N_B1_M1024_g N_A_477_368#_c_720_n 0.00816355f $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_281 N_B1_M1012_g N_A_477_368#_c_700_n 0.00194226f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_282 N_B1_M1014_g N_A_477_368#_c_700_n 0.00194226f $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_283 N_B1_c_287_n N_A_853_368#_c_757_n 0.00262904f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_284 N_B1_c_288_n N_A_853_368#_c_757_n 0.0204386f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_285 N_B1_M1012_g N_A_853_368#_c_767_n 0.0142562f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_286 N_B1_M1014_g N_A_853_368#_c_767_n 0.0142562f $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_287 N_B1_c_287_n N_A_853_368#_c_767_n 4.90767e-19 $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_288 N_B1_c_288_n N_A_853_368#_c_767_n 0.045298f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_289 N_B1_M1020_g N_A_853_368#_c_771_n 0.0142562f $X=5.535 $Y=2.4 $X2=0 $Y2=0
cc_290 N_B1_M1024_g N_A_853_368#_c_771_n 0.0142562f $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_291 N_B1_c_287_n N_A_853_368#_c_771_n 4.90767e-19 $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_292 N_B1_c_288_n N_A_853_368#_c_771_n 0.0444314f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_293 N_B1_c_287_n N_A_853_368#_c_775_n 5.54777e-19 $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_294 N_B1_c_288_n N_A_853_368#_c_775_n 0.0170101f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_295 N_B1_M1024_g N_VPWR_c_845_n 5.80674e-19 $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_296 N_B1_M1012_g N_VPWR_c_850_n 0.00333896f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_297 N_B1_M1014_g N_VPWR_c_850_n 0.00333896f $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_298 N_B1_M1020_g N_VPWR_c_850_n 0.00333896f $X=5.535 $Y=2.4 $X2=0 $Y2=0
cc_299 N_B1_M1024_g N_VPWR_c_850_n 0.00517089f $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_300 N_B1_M1012_g N_VPWR_c_844_n 0.00427818f $X=4.635 $Y=2.4 $X2=0 $Y2=0
cc_301 N_B1_M1014_g N_VPWR_c_844_n 0.00422685f $X=5.085 $Y=2.4 $X2=0 $Y2=0
cc_302 N_B1_M1020_g N_VPWR_c_844_n 0.00422685f $X=5.535 $Y=2.4 $X2=0 $Y2=0
cc_303 N_B1_M1024_g N_VPWR_c_844_n 0.00978686f $X=5.985 $Y=2.4 $X2=0 $Y2=0
cc_304 N_B1_M1013_g N_VGND_c_961_n 0.00434272f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_305 N_B1_M1019_g N_VGND_c_961_n 0.00383152f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_306 N_B1_M1013_g N_VGND_c_962_n 5.07239e-19 $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_307 N_B1_M1019_g N_VGND_c_962_n 0.0117017f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_308 N_B1_M1013_g N_VGND_c_971_n 0.00825037f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_309 N_B1_M1019_g N_VGND_c_971_n 0.0075754f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B1_M1013_g N_VGND_c_974_n 0.00597094f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A1_M1033_g N_A2_M1007_g 0.019323f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A1_M1032_g N_A2_M1005_g 0.0145057f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_313 A1 N_A2_c_445_n 0.0381127f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_314 N_A1_c_360_n N_A2_c_445_n 3.70592e-19 $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_315 A1 N_A2_c_440_n 0.00355468f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_316 N_A1_c_360_n N_A2_c_440_n 0.0145057f $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_317 N_A1_M1011_g N_Y_c_576_n 0.00939349f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A1_M1030_g N_Y_c_576_n 0.0106855f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_319 A1 N_Y_c_576_n 0.0330906f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A1_c_360_n N_Y_c_576_n 0.00233206f $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_321 N_A1_M1009_g N_Y_c_579_n 0.0123964f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_322 A1 N_Y_c_579_n 0.0342389f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_323 N_A1_c_360_n N_Y_c_579_n 0.00338169f $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_324 N_A1_M1009_g N_Y_c_580_n 0.0110564f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A1_M1011_g N_Y_c_580_n 0.00548858f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A1_M1030_g N_Y_c_580_n 6.61345e-19 $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A1_c_360_n N_Y_c_580_n 0.00252767f $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_328 N_A1_M1011_g N_Y_c_581_n 5.30577e-19 $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_M1030_g N_Y_c_581_n 0.0045607f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1033_g N_Y_c_581_n 0.00463734f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_331 A1 N_Y_c_581_n 0.0218587f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A1_c_360_n N_Y_c_581_n 0.00229269f $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_333 N_A1_M1001_g N_A_477_368#_c_698_n 2.99783e-19 $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_334 N_A1_M1001_g N_A_853_368#_c_777_n 0.0172931f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A1_M1003_g N_A_853_368#_c_777_n 0.0142562f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_336 A1 N_A_853_368#_c_777_n 0.0381041f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_337 N_A1_c_360_n N_A_853_368#_c_777_n 4.8724e-19 $X=7.79 $Y=1.515 $X2=0 $Y2=0
cc_338 N_A1_M1028_g N_A_853_368#_c_781_n 0.0142562f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_339 N_A1_M1032_g N_A_853_368#_c_781_n 0.0142562f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_340 A1 N_A_853_368#_c_781_n 0.0478981f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_341 N_A1_c_360_n N_A_853_368#_c_781_n 4.90062e-19 $X=7.79 $Y=1.515 $X2=0
+ $Y2=0
cc_342 A1 N_A_853_368#_c_785_n 0.0143992f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_343 N_A1_c_360_n N_A_853_368#_c_785_n 5.52655e-19 $X=7.79 $Y=1.515 $X2=0
+ $Y2=0
cc_344 A1 N_A_853_368#_c_787_n 0.00940956f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_345 N_A1_M1001_g N_VPWR_c_845_n 0.0134031f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_346 N_A1_M1003_g N_VPWR_c_845_n 0.0133668f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_347 N_A1_M1028_g N_VPWR_c_845_n 5.41206e-19 $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A1_M1003_g N_VPWR_c_846_n 0.00460063f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_349 N_A1_M1028_g N_VPWR_c_846_n 0.00460063f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_350 N_A1_M1003_g N_VPWR_c_847_n 5.41206e-19 $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A1_M1028_g N_VPWR_c_847_n 0.0133668f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A1_M1032_g N_VPWR_c_847_n 0.0133668f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_353 N_A1_M1032_g N_VPWR_c_848_n 5.43099e-19 $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_354 N_A1_M1001_g N_VPWR_c_850_n 0.00460063f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_355 N_A1_M1032_g N_VPWR_c_852_n 0.00460063f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_356 N_A1_M1001_g N_VPWR_c_844_n 0.00908665f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A1_M1003_g N_VPWR_c_844_n 0.00908554f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_358 N_A1_M1028_g N_VPWR_c_844_n 0.00908554f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A1_M1032_g N_VPWR_c_844_n 0.00908665f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A1_M1033_g N_VGND_c_963_n 6.35276e-19 $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_361 N_A1_M1009_g N_VGND_c_968_n 0.00291649f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A1_M1011_g N_VGND_c_968_n 0.00291649f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A1_M1030_g N_VGND_c_968_n 0.00291649f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A1_M1033_g N_VGND_c_968_n 0.00291649f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_365 N_A1_M1009_g N_VGND_c_971_n 0.0036412f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A1_M1011_g N_VGND_c_971_n 0.00359121f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A1_M1030_g N_VGND_c_971_n 0.00359121f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A1_M1033_g N_VGND_c_971_n 0.00359219f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A1_M1030_g N_A_1228_74#_c_1062_n 0.010822f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A1_M1033_g N_A_1228_74#_c_1062_n 0.0142063f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A1_M1033_g N_A_1228_74#_c_1065_n 0.00174382f $X=7.79 $Y=0.74 $X2=0
+ $Y2=0
cc_372 A1 N_A_1228_74#_c_1065_n 0.0103694f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_373 N_A1_M1009_g N_A_1228_74#_c_1070_n 0.0113038f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A1_M1011_g N_A_1228_74#_c_1070_n 0.0109057f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A2_M1005_g N_A_853_368#_c_788_n 0.0160581f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_376 N_A2_M1008_g N_A_853_368#_c_788_n 0.012931f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_377 N_A2_c_445_n N_A_853_368#_c_788_n 0.0370319f $X=9.39 $Y=1.515 $X2=0 $Y2=0
cc_378 N_A2_c_440_n N_A_853_368#_c_788_n 4.89356e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_379 N_A2_M1005_g N_A_853_368#_c_762_n 6.74232e-19 $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_380 N_A2_M1008_g N_A_853_368#_c_762_n 0.0121949f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_381 N_A2_M1010_g N_A_853_368#_c_762_n 0.0121949f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_382 N_A2_M1015_g N_A_853_368#_c_762_n 6.74232e-19 $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_383 N_A2_M1010_g N_A_853_368#_c_796_n 0.012931f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_384 N_A2_M1015_g N_A_853_368#_c_796_n 0.0177335f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_385 N_A2_c_445_n N_A_853_368#_c_796_n 0.0326541f $X=9.39 $Y=1.515 $X2=0 $Y2=0
cc_386 N_A2_c_440_n N_A_853_368#_c_796_n 4.86535e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_387 N_A2_M1015_g N_A_853_368#_c_763_n 8.13654e-19 $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_388 N_A2_M1015_g N_A_853_368#_c_764_n 0.00147311f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_389 N_A2_M1008_g N_A_853_368#_c_802_n 8.84614e-19 $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_390 N_A2_M1010_g N_A_853_368#_c_802_n 8.84614e-19 $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_391 N_A2_c_445_n N_A_853_368#_c_802_n 0.0235495f $X=9.39 $Y=1.515 $X2=0 $Y2=0
cc_392 N_A2_c_440_n N_A_853_368#_c_802_n 5.51948e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_393 N_A2_M1005_g N_VPWR_c_847_n 5.41206e-19 $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_394 N_A2_M1005_g N_VPWR_c_848_n 0.0124151f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_395 N_A2_M1008_g N_VPWR_c_848_n 0.002979f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_396 N_A2_M1010_g N_VPWR_c_849_n 0.002979f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A2_M1015_g N_VPWR_c_849_n 0.0153844f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A2_M1005_g N_VPWR_c_852_n 0.00460063f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_399 N_A2_M1008_g N_VPWR_c_853_n 0.005209f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_400 N_A2_M1010_g N_VPWR_c_853_n 0.005209f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_401 N_A2_M1015_g N_VPWR_c_854_n 0.00460063f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_402 N_A2_M1005_g N_VPWR_c_844_n 0.00908665f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_403 N_A2_M1008_g N_VPWR_c_844_n 0.00982266f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_404 N_A2_M1010_g N_VPWR_c_844_n 0.00982266f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_405 N_A2_M1015_g N_VPWR_c_844_n 0.00912261f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A2_M1007_g N_VGND_c_963_n 0.010782f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A2_M1018_g N_VGND_c_963_n 0.0106755f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_408 N_A2_M1023_g N_VGND_c_963_n 4.71636e-19 $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A2_M1018_g N_VGND_c_964_n 4.71636e-19 $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_410 N_A2_M1023_g N_VGND_c_964_n 0.0106755f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_411 N_A2_M1027_g N_VGND_c_964_n 0.0137191f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_412 N_A2_M1007_g N_VGND_c_968_n 0.00383152f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_413 N_A2_M1018_g N_VGND_c_969_n 0.00383152f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_414 N_A2_M1023_g N_VGND_c_969_n 0.00383152f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A2_M1027_g N_VGND_c_970_n 0.00383152f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A2_M1007_g N_VGND_c_971_n 0.00757637f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_417 N_A2_M1018_g N_VGND_c_971_n 0.0075754f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_418 N_A2_M1023_g N_VGND_c_971_n 0.0075754f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_419 N_A2_M1027_g N_VGND_c_971_n 0.00761428f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_420 N_A2_M1007_g N_A_1228_74#_c_1064_n 0.0147292f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_421 N_A2_M1018_g N_A_1228_74#_c_1064_n 0.0130453f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_422 N_A2_c_445_n N_A_1228_74#_c_1064_n 0.0431743f $X=9.39 $Y=1.515 $X2=0
+ $Y2=0
cc_423 N_A2_c_440_n N_A_1228_74#_c_1064_n 0.00236025f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_424 N_A2_M1018_g N_A_1228_74#_c_1066_n 3.92313e-19 $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_425 N_A2_M1023_g N_A_1228_74#_c_1066_n 3.92313e-19 $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_426 N_A2_M1023_g N_A_1228_74#_c_1067_n 0.0130918f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A2_M1027_g N_A_1228_74#_c_1067_n 0.0145697f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A2_c_445_n N_A_1228_74#_c_1067_n 0.0453632f $X=9.39 $Y=1.515 $X2=0
+ $Y2=0
cc_429 N_A2_c_440_n N_A_1228_74#_c_1067_n 0.00647684f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_430 N_A2_M1027_g N_A_1228_74#_c_1068_n 0.00159319f $X=9.51 $Y=0.74 $X2=0
+ $Y2=0
cc_431 N_A2_c_445_n N_A_1228_74#_c_1072_n 0.0146029f $X=9.39 $Y=1.515 $X2=0
+ $Y2=0
cc_432 N_A2_c_440_n N_A_1228_74#_c_1072_n 0.00252677f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_433 N_A_29_368#_c_512_n N_Y_M1021_d 0.00165831f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_434 N_A_29_368#_c_514_n N_Y_M1026_d 0.00165831f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_435 N_A_29_368#_c_512_n N_Y_c_592_n 0.0159318f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_436 N_A_29_368#_M1022_s N_Y_c_584_n 0.00165831f $X=1.035 $Y=1.84 $X2=0 $Y2=0
cc_437 N_A_29_368#_c_546_p N_Y_c_584_n 0.0126919f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_438 N_A_29_368#_c_514_n N_Y_c_600_n 0.0139027f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_439 N_A_29_368#_c_516_n N_Y_c_574_n 0.0104493f $X=3.87 $Y=2.05 $X2=0 $Y2=0
cc_440 N_A_29_368#_M1021_s N_Y_c_587_n 0.00246785f $X=0.145 $Y=1.84 $X2=0 $Y2=0
cc_441 N_A_29_368#_c_511_n N_Y_c_587_n 0.0201299f $X=0.27 $Y=2.225 $X2=0 $Y2=0
cc_442 N_A_29_368#_c_528_n N_A_477_368#_M1000_d 0.00314376f $X=2.855 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_443 N_A_29_368#_c_532_n N_A_477_368#_M1004_d 0.0031345f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_444 N_A_29_368#_c_528_n N_A_477_368#_c_701_n 0.0148589f $X=2.855 $Y=2.035
+ $X2=0 $Y2=0
cc_445 N_A_29_368#_M1002_s N_A_477_368#_c_695_n 0.00165831f $X=2.835 $Y=1.84
+ $X2=0 $Y2=0
cc_446 N_A_29_368#_c_555_p N_A_477_368#_c_695_n 0.0118736f $X=2.97 $Y=2.57 $X2=0
+ $Y2=0
cc_447 N_A_29_368#_c_514_n N_A_477_368#_c_696_n 0.0110621f $X=1.905 $Y=2.99
+ $X2=0 $Y2=0
cc_448 N_A_29_368#_c_532_n N_A_477_368#_c_707_n 0.0170259f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_449 N_A_29_368#_M1006_s N_A_477_368#_c_697_n 0.00239704f $X=3.735 $Y=1.84
+ $X2=0 $Y2=0
cc_450 N_A_29_368#_c_516_n N_A_477_368#_c_697_n 0.0185322f $X=3.87 $Y=2.05 $X2=0
+ $Y2=0
cc_451 N_A_29_368#_c_516_n N_A_853_368#_c_757_n 0.0137126f $X=3.87 $Y=2.05 $X2=0
+ $Y2=0
cc_452 N_A_29_368#_c_516_n N_A_853_368#_c_758_n 0.0430072f $X=3.87 $Y=2.05 $X2=0
+ $Y2=0
cc_453 N_A_29_368#_c_512_n N_VPWR_c_850_n 0.0459191f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_454 N_A_29_368#_c_513_n N_VPWR_c_850_n 0.0178855f $X=0.355 $Y=2.99 $X2=0
+ $Y2=0
cc_455 N_A_29_368#_c_514_n N_VPWR_c_850_n 0.0643017f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_456 N_A_29_368#_c_515_n N_VPWR_c_850_n 0.0121867f $X=1.17 $Y=2.99 $X2=0 $Y2=0
cc_457 N_A_29_368#_c_512_n N_VPWR_c_844_n 0.0258001f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_458 N_A_29_368#_c_513_n N_VPWR_c_844_n 0.00971414f $X=0.355 $Y=2.99 $X2=0
+ $Y2=0
cc_459 N_A_29_368#_c_514_n N_VPWR_c_844_n 0.0354845f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_460 N_A_29_368#_c_515_n N_VPWR_c_844_n 0.00660921f $X=1.17 $Y=2.99 $X2=0
+ $Y2=0
cc_461 N_Y_c_570_n N_VGND_M1017_s 0.00473729f $X=1.53 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_462 N_Y_c_604_n N_VGND_M1029_s 0.00807452f $X=2.39 $Y=0.925 $X2=0 $Y2=0
cc_463 N_Y_c_574_n N_VGND_M1025_s 0.0158527f $X=4.07 $Y=1.095 $X2=0 $Y2=0
cc_464 N_Y_c_579_n N_VGND_M1019_s 0.00285432f $X=6.55 $Y=0.975 $X2=0 $Y2=0
cc_465 N_Y_c_570_n N_VGND_c_959_n 0.0215198f $X=1.53 $Y=0.925 $X2=0 $Y2=0
cc_466 N_Y_c_572_n N_VGND_c_959_n 0.0135953f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_467 N_Y_c_572_n N_VGND_c_960_n 0.0135953f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_468 N_Y_c_604_n N_VGND_c_960_n 0.0167019f $X=2.39 $Y=0.925 $X2=0 $Y2=0
cc_469 N_Y_c_573_n N_VGND_c_960_n 0.0121972f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_470 N_Y_c_575_n N_VGND_c_961_n 0.0109942f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_471 N_Y_c_575_n N_VGND_c_962_n 0.0170358f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_472 N_Y_c_579_n N_VGND_c_962_n 0.022285f $X=6.55 $Y=0.975 $X2=0 $Y2=0
cc_473 N_Y_c_572_n N_VGND_c_965_n 0.00814895f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_474 N_Y_c_570_n N_VGND_c_971_n 0.0293519f $X=1.53 $Y=0.925 $X2=0 $Y2=0
cc_475 N_Y_c_571_n N_VGND_c_971_n 0.00906892f $X=0.355 $Y=0.925 $X2=0 $Y2=0
cc_476 N_Y_c_572_n N_VGND_c_971_n 0.00627841f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_477 N_Y_c_604_n N_VGND_c_971_n 0.0116543f $X=2.39 $Y=0.925 $X2=0 $Y2=0
cc_478 N_Y_c_573_n N_VGND_c_971_n 0.00904371f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_479 N_Y_c_575_n N_VGND_c_971_n 0.00904371f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_480 N_Y_c_573_n N_VGND_c_973_n 0.0109942f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_481 N_Y_c_573_n N_VGND_c_974_n 0.0185534f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_482 N_Y_c_574_n N_VGND_c_974_n 0.0863478f $X=4.07 $Y=1.095 $X2=0 $Y2=0
cc_483 N_Y_c_575_n N_VGND_c_974_n 0.0185534f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_484 N_Y_c_579_n N_A_1228_74#_M1009_d 0.00392596f $X=6.55 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_485 N_Y_c_576_n N_A_1228_74#_M1011_d 0.00205565f $X=7.41 $Y=1.022 $X2=0 $Y2=0
cc_486 N_Y_M1030_s N_A_1228_74#_c_1062_n 0.00178571f $X=7.435 $Y=0.37 $X2=0
+ $Y2=0
cc_487 N_Y_c_576_n N_A_1228_74#_c_1062_n 0.00540301f $X=7.41 $Y=1.022 $X2=0
+ $Y2=0
cc_488 N_Y_c_581_n N_A_1228_74#_c_1062_n 0.0161432f $X=7.575 $Y=0.95 $X2=0 $Y2=0
cc_489 N_Y_c_581_n N_A_1228_74#_c_1065_n 0.00517071f $X=7.575 $Y=0.95 $X2=0
+ $Y2=0
cc_490 N_Y_c_579_n N_A_1228_74#_c_1069_n 0.0128721f $X=6.55 $Y=0.975 $X2=0 $Y2=0
cc_491 N_Y_M1009_s N_A_1228_74#_c_1070_n 0.00179007f $X=6.575 $Y=0.37 $X2=0
+ $Y2=0
cc_492 N_Y_c_576_n N_A_1228_74#_c_1070_n 0.00538156f $X=7.41 $Y=1.022 $X2=0
+ $Y2=0
cc_493 N_Y_c_579_n N_A_1228_74#_c_1070_n 0.00465091f $X=6.55 $Y=0.975 $X2=0
+ $Y2=0
cc_494 N_Y_c_580_n N_A_1228_74#_c_1070_n 0.0163588f $X=6.88 $Y=0.975 $X2=0 $Y2=0
cc_495 N_Y_c_576_n N_A_1228_74#_c_1071_n 0.0101598f $X=7.41 $Y=1.022 $X2=0 $Y2=0
cc_496 N_A_477_368#_c_697_n N_A_853_368#_M1012_s 0.00266942f $X=4.695 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_497 N_A_477_368#_c_698_n N_A_853_368#_M1014_s 0.00165831f $X=5.595 $Y=2.99
+ $X2=0 $Y2=0
cc_498 N_A_477_368#_c_697_n N_A_853_368#_c_758_n 0.0184743f $X=4.695 $Y=2.99
+ $X2=0 $Y2=0
cc_499 N_A_477_368#_M1012_d N_A_853_368#_c_767_n 0.00314376f $X=4.725 $Y=1.84
+ $X2=0 $Y2=0
cc_500 N_A_477_368#_c_714_n N_A_853_368#_c_767_n 0.0170259f $X=4.86 $Y=2.405
+ $X2=0 $Y2=0
cc_501 N_A_477_368#_c_698_n N_A_853_368#_c_813_n 0.0118736f $X=5.595 $Y=2.99
+ $X2=0 $Y2=0
cc_502 N_A_477_368#_M1020_d N_A_853_368#_c_771_n 0.00314376f $X=5.625 $Y=1.84
+ $X2=0 $Y2=0
cc_503 N_A_477_368#_c_720_n N_A_853_368#_c_771_n 0.0170259f $X=5.76 $Y=2.405
+ $X2=0 $Y2=0
cc_504 N_A_477_368#_c_698_n N_A_853_368#_c_759_n 0.00341172f $X=5.595 $Y=2.99
+ $X2=0 $Y2=0
cc_505 N_A_477_368#_c_698_n N_VPWR_c_845_n 0.00279016f $X=5.595 $Y=2.99 $X2=0
+ $Y2=0
cc_506 N_A_477_368#_c_695_n N_VPWR_c_850_n 0.0357927f $X=3.255 $Y=2.99 $X2=0
+ $Y2=0
cc_507 N_A_477_368#_c_696_n N_VPWR_c_850_n 0.0178163f $X=2.685 $Y=2.99 $X2=0
+ $Y2=0
cc_508 N_A_477_368#_c_697_n N_VPWR_c_850_n 0.0705786f $X=4.695 $Y=2.99 $X2=0
+ $Y2=0
cc_509 N_A_477_368#_c_698_n N_VPWR_c_850_n 0.0592384f $X=5.595 $Y=2.99 $X2=0
+ $Y2=0
cc_510 N_A_477_368#_c_699_n N_VPWR_c_850_n 0.0234458f $X=3.42 $Y=2.99 $X2=0
+ $Y2=0
cc_511 N_A_477_368#_c_700_n N_VPWR_c_850_n 0.0234458f $X=4.86 $Y=2.99 $X2=0
+ $Y2=0
cc_512 N_A_477_368#_c_695_n N_VPWR_c_844_n 0.0200586f $X=3.255 $Y=2.99 $X2=0
+ $Y2=0
cc_513 N_A_477_368#_c_696_n N_VPWR_c_844_n 0.00958215f $X=2.685 $Y=2.99 $X2=0
+ $Y2=0
cc_514 N_A_477_368#_c_697_n N_VPWR_c_844_n 0.0403615f $X=4.695 $Y=2.99 $X2=0
+ $Y2=0
cc_515 N_A_477_368#_c_698_n N_VPWR_c_844_n 0.0326137f $X=5.595 $Y=2.99 $X2=0
+ $Y2=0
cc_516 N_A_477_368#_c_699_n N_VPWR_c_844_n 0.0125551f $X=3.42 $Y=2.99 $X2=0
+ $Y2=0
cc_517 N_A_477_368#_c_700_n N_VPWR_c_844_n 0.0125551f $X=4.86 $Y=2.99 $X2=0
+ $Y2=0
cc_518 N_A_853_368#_c_777_n N_VPWR_M1001_d 0.00314376f $X=7.025 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_519 N_A_853_368#_c_781_n N_VPWR_M1028_d 0.00314376f $X=7.925 $Y=2.035 $X2=0
+ $Y2=0
cc_520 N_A_853_368#_c_788_n N_VPWR_M1005_d 0.00314376f $X=8.745 $Y=2.035 $X2=0
+ $Y2=0
cc_521 N_A_853_368#_c_796_n N_VPWR_M1010_d 0.00314376f $X=9.725 $Y=2.035 $X2=0
+ $Y2=0
cc_522 N_A_853_368#_c_759_n N_VPWR_c_845_n 0.0233699f $X=6.21 $Y=2.43 $X2=0
+ $Y2=0
cc_523 N_A_853_368#_c_777_n N_VPWR_c_845_n 0.0170259f $X=7.025 $Y=2.035 $X2=0
+ $Y2=0
cc_524 N_A_853_368#_c_760_n N_VPWR_c_845_n 0.0233699f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_525 N_A_853_368#_c_760_n N_VPWR_c_846_n 0.00749631f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_526 N_A_853_368#_c_760_n N_VPWR_c_847_n 0.0233699f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_527 N_A_853_368#_c_781_n N_VPWR_c_847_n 0.0170259f $X=7.925 $Y=2.035 $X2=0
+ $Y2=0
cc_528 N_A_853_368#_c_761_n N_VPWR_c_847_n 0.0233699f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_529 N_A_853_368#_c_761_n N_VPWR_c_848_n 0.022423f $X=8.01 $Y=2.43 $X2=0 $Y2=0
cc_530 N_A_853_368#_c_788_n N_VPWR_c_848_n 0.0148589f $X=8.745 $Y=2.035 $X2=0
+ $Y2=0
cc_531 N_A_853_368#_c_762_n N_VPWR_c_848_n 0.0234083f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_532 N_A_853_368#_c_762_n N_VPWR_c_849_n 0.0234083f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_533 N_A_853_368#_c_796_n N_VPWR_c_849_n 0.0148589f $X=9.725 $Y=2.035 $X2=0
+ $Y2=0
cc_534 N_A_853_368#_c_764_n N_VPWR_c_849_n 0.0224614f $X=9.81 $Y=2.4 $X2=0 $Y2=0
cc_535 N_A_853_368#_c_759_n N_VPWR_c_850_n 0.00749631f $X=6.21 $Y=2.43 $X2=0
+ $Y2=0
cc_536 N_A_853_368#_c_761_n N_VPWR_c_852_n 0.00749631f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_537 N_A_853_368#_c_762_n N_VPWR_c_853_n 0.0144623f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_538 N_A_853_368#_c_764_n N_VPWR_c_854_n 0.011066f $X=9.81 $Y=2.4 $X2=0 $Y2=0
cc_539 N_A_853_368#_c_759_n N_VPWR_c_844_n 0.0062048f $X=6.21 $Y=2.43 $X2=0
+ $Y2=0
cc_540 N_A_853_368#_c_760_n N_VPWR_c_844_n 0.0062048f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_541 N_A_853_368#_c_761_n N_VPWR_c_844_n 0.0062048f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_542 N_A_853_368#_c_762_n N_VPWR_c_844_n 0.0118344f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_543 N_A_853_368#_c_764_n N_VPWR_c_844_n 0.00915947f $X=9.81 $Y=2.4 $X2=0
+ $Y2=0
cc_544 N_A_853_368#_c_763_n N_A_1228_74#_c_1067_n 0.00609927f $X=9.85 $Y=2.12
+ $X2=0 $Y2=0
cc_545 N_VGND_c_963_n N_A_1228_74#_c_1063_n 0.00985092f $X=8.435 $Y=0.675 $X2=0
+ $Y2=0
cc_546 N_VGND_c_968_n N_A_1228_74#_c_1063_n 0.00758556f $X=8.27 $Y=0 $X2=0 $Y2=0
cc_547 N_VGND_c_971_n N_A_1228_74#_c_1063_n 0.00627867f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_548 N_VGND_M1007_s N_A_1228_74#_c_1064_n 0.00176461f $X=8.295 $Y=0.37 $X2=0
+ $Y2=0
cc_549 N_VGND_c_963_n N_A_1228_74#_c_1064_n 0.0170777f $X=8.435 $Y=0.675 $X2=0
+ $Y2=0
cc_550 N_VGND_c_963_n N_A_1228_74#_c_1066_n 0.0182488f $X=8.435 $Y=0.675 $X2=0
+ $Y2=0
cc_551 N_VGND_c_964_n N_A_1228_74#_c_1066_n 0.0182488f $X=9.295 $Y=0.675 $X2=0
+ $Y2=0
cc_552 N_VGND_c_969_n N_A_1228_74#_c_1066_n 0.00749631f $X=9.13 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_971_n N_A_1228_74#_c_1066_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_554 N_VGND_M1023_s N_A_1228_74#_c_1067_n 0.00176461f $X=9.155 $Y=0.37 $X2=0
+ $Y2=0
cc_555 N_VGND_c_964_n N_A_1228_74#_c_1067_n 0.0170777f $X=9.295 $Y=0.675 $X2=0
+ $Y2=0
cc_556 N_VGND_c_964_n N_A_1228_74#_c_1068_n 0.0182902f $X=9.295 $Y=0.675 $X2=0
+ $Y2=0
cc_557 N_VGND_c_970_n N_A_1228_74#_c_1068_n 0.011066f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_c_971_n N_A_1228_74#_c_1068_n 0.00915947f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_968_n N_A_1228_74#_c_1069_n 0.0732673f $X=8.27 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_c_971_n N_A_1228_74#_c_1069_n 0.0615998f $X=9.84 $Y=0 $X2=0 $Y2=0

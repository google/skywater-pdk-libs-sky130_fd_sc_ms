* File: sky130_fd_sc_ms__sdfbbn_1.spice
* Created: Fri Aug 28 18:10:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfbbn_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfbbn_1  VNB VPB SCD D SCE CLK_N SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK_N	CLK_N
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1006 A_119_119# N_SCD_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1034 N_A_197_119#_M1034_d N_SCE_M1034_g A_119_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_305_119# N_D_M1002_g N_A_197_119#_M1034_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=31.428 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_353_93#_M1035_g A_305_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1449 AS=0.0504 PD=1.11 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_A_353_93#_M1021_d N_SCE_M1021_g N_VGND_M1035_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1449 PD=1.41 PS=1.11 NRD=0 NRS=117.132 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_CLK_N_M1018_g N_A_662_82#_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.2109 PD=1.41 PS=2.05 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1019 N_A_867_82#_M1019_d N_A_662_82#_M1019_g N_VGND_M1018_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.3219 AS=0.19615 PD=2.35 PS=1.41 NRD=12.156 NRS=34.056 M=1
+ R=4.93333 SA=75000.8 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1025 A_1151_119# N_A_977_243#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1020 N_A_1162_497#_M1020_d N_A_662_82#_M1020_g A_1151_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_197_119#_M1003_d N_A_867_82#_M1003_g N_A_1162_497#_M1020_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=21.42 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_977_243#_M1005_d N_A_1162_497#_M1005_g N_A_1434_78#_M1005_s VNB
+ NLOWVT L=0.15 W=0.55 AD=0.1045 AS=0.2602 PD=0.93 PS=2.24 NRD=4.908 NRS=91.212
+ M=1 R=3.66667 SA=75000.3 SB=75004.9 A=0.0825 P=1.4 MULT=1
MM1045 N_A_1434_78#_M1045_d N_A_1579_258#_M1045_g N_A_977_243#_M1005_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.125125 AS=0.1045 PD=1.005 PS=0.93 NRD=15.264 NRS=0
+ M=1 R=3.66667 SA=75000.8 SB=75004.4 A=0.0825 P=1.4 MULT=1
MM1026 N_VGND_M1026_d N_SET_B_M1026_g N_A_1434_78#_M1045_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.11275 AS=0.125125 PD=0.96 PS=1.005 NRD=0 NRS=22.908 M=1 R=3.66667
+ SA=75001.4 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1042 A_1876_119# N_A_977_243#_M1042_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.066 AS=0.11275 PD=0.79 PS=0.96 NRD=14.172 NRS=28.356 M=1 R=3.66667
+ SA=75002 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1027 N_A_1954_119#_M1027_d N_A_662_82#_M1027_g A_1876_119# VNB NLOWVT L=0.15
+ W=0.55 AD=0.272562 AS=0.066 PD=1.64433 PS=0.79 NRD=0 NRS=14.172 M=1 R=3.66667
+ SA=75002.4 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1040 A_2164_119# N_A_867_82#_M1040_g N_A_1954_119#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0819 AS=0.208138 PD=0.81 PS=1.25567 NRD=39.996 NRS=32.856 M=1
+ R=2.8 SA=75003.4 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_2133_410#_M1010_g A_2164_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.128218 AS=0.0819 PD=0.99931 PS=0.81 NRD=71.508 NRS=39.996 M=1 R=2.8
+ SA=75004 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_2392_74#_M1009_d N_SET_B_M1009_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.225907 PD=1.02 PS=1.76069 NRD=0 NRS=40.584 M=1 R=4.93333
+ SA=75002.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1039 N_A_2133_410#_M1039_d N_A_1579_258#_M1039_g N_A_2392_74#_M1009_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1406 AS=0.1036 PD=1.12 PS=1.02 NRD=16.212 NRS=0 M=1
+ R=4.93333 SA=75003.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1032 N_A_2392_74#_M1032_d N_A_1954_119#_M1032_g N_A_2133_410#_M1039_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.2875 AS=0.1406 PD=2.33 PS=1.12 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75003.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_RESET_B_M1004_g N_A_1579_258#_M1004_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.132372 AS=0.1197 PD=0.970345 PS=1.41 NRD=74.328 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1007 N_Q_N_M1007_d N_A_2133_410#_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.233228 PD=2.05 PS=1.70966 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_2133_410#_M1024_g N_A_3078_384#_M1024_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=17.988 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1038 N_Q_M1038_d N_A_3078_384#_M1038_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.144644 PD=2.05 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_SCD_M1008_g N_A_27_464#_M1008_s VPB PSHORT L=0.18 W=0.64
+ AD=0.096 AS=0.1792 PD=0.94 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1036 A_215_464# N_SCE_M1036_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.096 PD=0.88 PS=0.94 NRD=19.9955 NRS=7.683 M=1 R=3.55556
+ SA=90000.7 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1011 N_A_197_119#_M1011_d N_D_M1011_g A_215_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.1
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1013 N_A_27_464#_M1013_d N_A_353_93#_M1013_g N_A_197_119#_M1011_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.176 AS=0.0864 PD=1.83 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90001.5 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1000 N_A_353_93#_M1000_d N_SCE_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.1792 PD=1.84 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1029 N_VPWR_M1029_d N_CLK_N_M1029_g N_A_662_82#_M1029_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1033 N_A_867_82#_M1033_d N_A_662_82#_M1033_g N_VPWR_M1029_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1031 A_1084_497# N_A_977_243#_M1031_g N_VPWR_M1031_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=23.443 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1014 N_A_1162_497#_M1014_d N_A_867_82#_M1014_g A_1084_497# VPB PSHORT L=0.18
+ W=0.42 AD=0.0834849 AS=0.0441 PD=0.788491 PS=0.63 NRD=39.8531 NRS=23.443 M=1
+ R=2.33333 SA=90000.6 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1017 N_A_197_119#_M1017_d N_A_662_82#_M1017_g N_A_1162_497#_M1014_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.2112 AS=0.127215 PD=1.94 PS=1.20151 NRD=13.8491 NRS=0 M=1
+ R=3.55556 SA=90000.8 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1037 A_1531_424# N_A_1162_497#_M1037_g N_A_977_243#_M1037_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1008 AS=0.378 PD=1.08 PS=2.58 NRD=15.2281 NRS=0 M=1 R=4.66667
+ SA=90000.4 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1041 N_VPWR_M1041_d N_A_1579_258#_M1041_g A_1531_424# VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1008 PD=1.11 PS=1.08 NRD=0 NRS=15.2281 M=1 R=4.66667 SA=90000.8
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1044 N_A_977_243#_M1044_d N_SET_B_M1044_g N_VPWR_M1041_d VPB PSHORT L=0.18
+ W=0.84 AD=0.231 AS=0.1134 PD=2.23 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667 SA=90001.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1001 A_1906_424# N_A_977_243#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.0882 AS=0.2352 PD=1.05 PS=2.24 NRD=11.7215 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1015 N_A_1954_119#_M1015_d N_A_867_82#_M1015_g A_1906_424# VPB PSHORT L=0.18
+ W=0.84 AD=0.1778 AS=0.0882 PD=1.59333 PS=1.05 NRD=0 NRS=11.7215 M=1 R=4.66667
+ SA=90000.6 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1030 A_2091_508# N_A_662_82#_M1030_g N_A_1954_119#_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0889 PD=0.63 PS=0.796667 NRD=23.443 NRS=37.5088 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1012 N_VPWR_M1012_d N_A_2133_410#_M1012_g A_2091_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.22145 AS=0.0441 PD=2.04 PS=0.63 NRD=221.507 NRS=23.443 M=1 R=2.33333
+ SA=90001.5 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1028 N_VPWR_M1028_d N_SET_B_M1028_g N_A_2133_410#_M1028_s VPB PSHORT L=0.18
+ W=1 AD=0.254075 AS=0.28 PD=1.675 PS=2.56 NRD=39.203 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1023 A_2512_392# N_A_1579_258#_M1023_g N_VPWR_M1028_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.254075 PD=1.24 PS=1.675 NRD=12.7853 NRS=39.203 M=1 R=5.55556
+ SA=90000.8 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1046 N_A_2133_410#_M1046_d N_A_1954_119#_M1046_g A_2512_392# VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90001.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1047 N_VPWR_M1047_d N_RESET_B_M1047_g N_A_1579_258#_M1047_s VPB PSHORT L=0.18
+ W=0.64 AD=0.190255 AS=0.3529 PD=1.27273 PS=3.68 NRD=0 NRS=152.793 M=1
+ R=3.55556 SA=90000.2 SB=90001 A=0.1152 P=1.64 MULT=1
MM1043 N_Q_N_M1043_d N_A_2133_410#_M1043_g N_VPWR_M1047_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.332945 PD=2.8 PS=2.22727 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_A_2133_410#_M1016_g N_A_3078_384#_M1016_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1614 AS=0.2352 PD=1.26429 PS=2.24 NRD=19.1484 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1022 N_Q_M1022_d N_A_3078_384#_M1022_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2152 PD=2.8 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX48_noxref VNB VPB NWDIODE A=32.1616 P=38.3
c_197 VNB 0 1.86341e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sdfbbn_1.pxi.spice"
*
.ends
*
*

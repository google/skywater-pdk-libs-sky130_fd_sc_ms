* File: sky130_fd_sc_ms__dfbbn_1.pex.spice
* Created: Fri Aug 28 17:21:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFBBN_1%CLK_N 3 7 9 13 15
c34 3 0 1.52998e-19 $X=0.495 $Y=2.4
r35 12 15 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.33 $Y=1.465
+ $X2=0.495 $Y2=1.465
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.465 $X2=0.33 $Y2=1.465
r37 9 13 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=0.31 $Y=1.665 $X2=0.31
+ $Y2=1.465
r38 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r39 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r40 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=1.465
r41 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%D 3 7 9 10 17
r41 15 17 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.01 $Y=1.345 $X2=2.09
+ $Y2=1.345
r42 13 15 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=2.01 $Y2=1.345
r43 9 10 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.09 $Y=1.345
+ $X2=2.64 $Y2=1.345
r44 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.345 $X2=2.09 $Y2=1.345
r45 5 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.51
+ $X2=2.01 $Y2=1.345
r46 5 7 472.282 $w=1.8e-07 $l=1.215e-06 $layer=POLY_cond $X=2.01 $Y=1.51
+ $X2=2.01 $Y2=2.725
r47 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.915 $Y2=1.345
r48 1 3 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.915 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_474_405# 1 2 3 12 16 20 24 27 28 29 31 32
+ 33 34 38 40 44 49 51 57 62 69
c179 69 0 3.07191e-20 $X=6.41 $Y=1.795
c180 16 0 1.47675e-19 $X=2.61 $Y=2.725
r181 49 65 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.535 $Y=2.19
+ $X2=2.535 $Y2=2.355
r182 49 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.535 $Y=2.19
+ $X2=2.535 $Y2=2.025
r183 48 51 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.535 $Y=2.19
+ $X2=2.72 $Y2=2.19
r184 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=2.19 $X2=2.535 $Y2=2.19
r185 45 69 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.285 $Y=1.795
+ $X2=6.41 $Y2=1.795
r186 45 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.285 $Y=1.795
+ $X2=6.195 $Y2=1.795
r187 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.285
+ $Y=1.795 $X2=6.285 $Y2=1.795
r188 42 44 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.285 $Y=2.32
+ $X2=6.285 $Y2=1.795
r189 41 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.82 $Y=2.405
+ $X2=5.695 $Y2=2.405
r190 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.12 $Y=2.405
+ $X2=6.285 $Y2=2.32
r191 40 41 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.12 $Y=2.405
+ $X2=5.82 $Y2=2.405
r192 36 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.49
+ $X2=5.695 $Y2=2.405
r193 36 38 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=5.695 $Y=2.49
+ $X2=5.695 $Y2=2.815
r194 34 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.57 $Y=2.405
+ $X2=5.695 $Y2=2.405
r195 34 57 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.57 $Y=2.405
+ $X2=4.815 $Y2=2.405
r196 33 57 5.18835 $w=1.83e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=2.397
+ $X2=4.815 $Y2=2.397
r197 33 54 21.8821 $w=1.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.73 $Y=2.397
+ $X2=4.365 $Y2=2.397
r198 32 60 8.61582 $w=3.54e-07 $l=3.44601e-07 $layer=LI1_cond $X=4.73 $Y=1.165
+ $X2=4.98 $Y2=0.94
r199 32 33 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=4.73 $Y=1.165
+ $X2=4.73 $Y2=2.305
r200 31 54 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.365 $Y=2.905
+ $X2=4.365 $Y2=2.49
r201 28 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.2 $Y=2.99
+ $X2=4.365 $Y2=2.905
r202 28 29 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=4.2 $Y=2.99
+ $X2=2.805 $Y2=2.99
r203 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=2.905
+ $X2=2.805 $Y2=2.99
r204 26 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=2.355
+ $X2=2.72 $Y2=2.19
r205 26 27 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.72 $Y=2.355
+ $X2=2.72 $Y2=2.905
r206 22 69 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.41 $Y=1.96
+ $X2=6.41 $Y2=1.795
r207 22 24 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.41 $Y=1.96
+ $X2=6.41 $Y2=2.54
r208 18 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=1.795
r209 18 20 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=0.87
r210 16 65 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.61 $Y=2.725
+ $X2=2.61 $Y2=2.355
r211 12 64 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.54 $Y=0.805
+ $X2=2.54 $Y2=2.025
r212 3 62 600 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=1 $X=5.52
+ $Y=2.12 $X2=5.655 $Y2=2.405
r213 3 38 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=5.52
+ $Y=2.12 $X2=5.655 $Y2=2.815
r214 2 54 300 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_PDIFF $count=2 $X=4.235
+ $Y=2.12 $X2=4.365 $Y2=2.39
r215 1 60 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.595 $X2=4.98 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_200_74# 1 2 9 13 16 18 20 24 27 31 32 34
+ 35 36 38 41 42 44 46 47 51 55 56 57 58 59 60 66 73 74 75 82
c228 82 0 1.02788e-19 $X=7.98 $Y=1.395
c229 74 0 5.14108e-20 $X=3.35 $Y=1.29
c230 60 0 7.83046e-20 $X=3.265 $Y=1.295
c231 59 0 7.98666e-20 $X=6.815 $Y=1.295
c232 58 0 1.63798e-20 $X=3.107 $Y=1.77
c233 55 0 1.52998e-19 $X=1.17 $Y=1.985
c234 47 0 8.92848e-20 $X=6.875 $Y=1.765
c235 38 0 9.67413e-20 $X=3.107 $Y=1.685
c236 36 0 1.55193e-19 $X=2.125 $Y=1.77
c237 18 0 1.47104e-19 $X=7.98 $Y=1.23
r238 73 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.29
+ $X2=3.35 $Y2=1.125
r239 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.29 $X2=3.35 $Y2=1.29
r240 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.295
+ $X2=6.96 $Y2=1.295
r241 63 74 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=1.29
+ $X2=3.35 $Y2=1.29
r242 63 84 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=3.12 $Y=1.29
+ $X2=3.107 $Y2=1.29
r243 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r244 60 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.295
+ $X2=3.12 $Y2=1.295
r245 59 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=6.96 $Y2=1.295
r246 59 60 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=3.265 $Y2=1.295
r247 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.33 $Y=1.82
+ $X2=1.33 $Y2=1.13
r248 55 56 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=1.985
+ $X2=1.21 $Y2=1.82
r249 52 82 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=7.775 $Y=1.395
+ $X2=7.98 $Y2=1.395
r250 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.775
+ $Y=1.395 $X2=7.775 $Y2=1.395
r251 49 67 3.34605 $w=3.8e-07 $l=1.83e-07 $layer=LI1_cond $X=7.075 $Y=1.37
+ $X2=6.892 $Y2=1.37
r252 49 51 21.2292 $w=3.78e-07 $l=7e-07 $layer=LI1_cond $X=7.075 $Y=1.37
+ $X2=7.775 $Y2=1.37
r253 47 79 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.875 $Y=1.765
+ $X2=6.875 $Y2=1.93
r254 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.875
+ $Y=1.765 $X2=6.875 $Y2=1.765
r255 44 67 3.47404 $w=3.65e-07 $l=1.9e-07 $layer=LI1_cond $X=6.892 $Y=1.56
+ $X2=6.892 $Y2=1.37
r256 44 46 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=6.892 $Y=1.56
+ $X2=6.892 $Y2=1.765
r257 42 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=2.19
+ $X2=3.075 $Y2=2.355
r258 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.075
+ $Y=2.19 $X2=3.075 $Y2=2.19
r259 39 58 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.855
+ $X2=3.107 $Y2=1.77
r260 39 41 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=3.107 $Y=1.855
+ $X2=3.107 $Y2=2.19
r261 38 58 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.685
+ $X2=3.107 $Y2=1.77
r262 37 84 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=3.107 $Y=1.455
+ $X2=3.107 $Y2=1.29
r263 37 38 10.0023 $w=2.63e-07 $l=2.3e-07 $layer=LI1_cond $X=3.107 $Y=1.455
+ $X2=3.107 $Y2=1.685
r264 35 58 2.98021 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=3.107 $Y2=1.77
r265 35 36 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=2.125 $Y2=1.77
r266 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.04 $Y=1.855
+ $X2=2.125 $Y2=1.77
r267 33 34 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=2.04 $Y=1.855
+ $X2=2.04 $Y2=2.905
r268 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=2.04 $Y2=2.905
r269 31 32 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=1.415 $Y2=2.99
r270 25 57 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.235 $Y=0.95
+ $X2=1.235 $Y2=1.13
r271 25 27 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=1.235 $Y=0.95
+ $X2=1.235 $Y2=0.515
r272 22 32 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=1.21 $Y=2.905
+ $X2=1.415 $Y2=2.99
r273 22 24 2.52975 $w=4.08e-07 $l=9e-08 $layer=LI1_cond $X=1.21 $Y=2.905
+ $X2=1.21 $Y2=2.815
r274 21 55 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=1.21 $Y=2.025
+ $X2=1.21 $Y2=1.985
r275 21 24 22.2056 $w=4.08e-07 $l=7.9e-07 $layer=LI1_cond $X=1.21 $Y=2.025
+ $X2=1.21 $Y2=2.815
r276 18 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.98 $Y=1.23
+ $X2=7.98 $Y2=1.395
r277 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.98 $Y=1.23
+ $X2=7.98 $Y2=0.91
r278 16 79 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.8 $Y=2.54 $X2=6.8
+ $Y2=1.93
r279 13 75 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.33 $Y=0.805
+ $X2=3.33 $Y2=1.125
r280 9 71 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.03 $Y=2.725
+ $X2=3.03 $Y2=2.355
r281 2 55 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=1.985
r282 2 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=2.815
r283 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_595_119# 1 2 7 11 15 17 18 22 25 27 29 34
+ 38
c106 38 0 6.77906e-20 $X=3.975 $Y=1.47
c107 34 0 7.83046e-20 $X=3.72 $Y=1.595
c108 29 0 7.98666e-20 $X=3.115 $Y=0.775
c109 18 0 1.47675e-19 $X=3.41 $Y=2.65
c110 11 0 1.21772e-19 $X=4.59 $Y=2.54
r111 37 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.975 $Y=1.56
+ $X2=3.975 $Y2=1.47
r112 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.56 $X2=3.975 $Y2=1.56
r113 34 36 9.48476 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.72 $Y=1.595
+ $X2=3.975 $Y2=1.595
r114 29 31 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.115 $Y=0.775
+ $X2=3.115 $Y2=0.87
r115 27 34 4.5877 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.72 $Y=1.395 $X2=3.72
+ $Y2=1.595
r116 26 27 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.72 $Y=0.955
+ $X2=3.72 $Y2=1.395
r117 24 34 8.3689 $w=3.28e-07 $l=3.09233e-07 $layer=LI1_cond $X=3.495 $Y=1.795
+ $X2=3.72 $Y2=1.595
r118 24 25 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.495 $Y=1.795
+ $X2=3.495 $Y2=2.565
r119 23 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=0.87
+ $X2=3.115 $Y2=0.87
r120 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.635 $Y=0.87
+ $X2=3.72 $Y2=0.955
r121 22 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.635 $Y=0.87
+ $X2=3.28 $Y2=0.87
r122 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=2.65
+ $X2=3.495 $Y2=2.565
r123 18 20 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.41 $Y=2.65
+ $X2=3.285 $Y2=2.65
r124 13 17 18.8402 $w=1.65e-07 $l=1.00623e-07 $layer=POLY_cond $X=4.695 $Y=1.395
+ $X2=4.635 $Y2=1.47
r125 13 15 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.695 $Y=1.395
+ $X2=4.695 $Y2=0.87
r126 9 17 18.8402 $w=1.65e-07 $l=9.48683e-08 $layer=POLY_cond $X=4.59 $Y=1.545
+ $X2=4.635 $Y2=1.47
r127 9 11 386.766 $w=1.8e-07 $l=9.95e-07 $layer=POLY_cond $X=4.59 $Y=1.545
+ $X2=4.59 $Y2=2.54
r128 8 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.47
+ $X2=3.975 $Y2=1.47
r129 7 17 6.66866 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.5 $Y=1.47
+ $X2=4.635 $Y2=1.47
r130 7 8 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.5 $Y=1.47 $X2=4.14
+ $Y2=1.47
r131 2 20 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=2.515 $X2=3.285 $Y2=2.65
r132 1 29 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.595 $X2=3.115 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_978_357# 1 2 7 9 13 17 20 22 25 26 27 29
+ 30 31 34 35 37 40 43 45 47 49 55 56 59
c180 55 0 1.32454e-19 $X=9.465 $Y=1.02
c181 49 0 1.21772e-19 $X=5.125 $Y=1.42
c182 47 0 1.48333e-19 $X=10.685 $Y=2.035
c183 35 0 5.09967e-20 $X=9.465 $Y=1.395
c184 34 0 3.62021e-19 $X=9.465 $Y=1.395
c185 31 0 1.47104e-19 $X=8.545 $Y=1.02
c186 22 0 7.44062e-20 $X=6.315 $Y=1.42
c187 7 0 7.90569e-20 $X=4.98 $Y=1.935
r188 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=1.5 $X2=5.145 $Y2=1.5
r189 49 52 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=5.125 $Y=1.42
+ $X2=5.125 $Y2=1.5
r190 45 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.515 $Y=2.035
+ $X2=10.685 $Y2=2.035
r191 41 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.515 $Y=1.02
+ $X2=10.43 $Y2=1.02
r192 41 43 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=10.515 $Y=1.02
+ $X2=10.725 $Y2=1.02
r193 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.43 $Y=1.95
+ $X2=10.515 $Y2=2.035
r194 39 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.43 $Y=1.105
+ $X2=10.43 $Y2=1.02
r195 39 40 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=10.43 $Y=1.105
+ $X2=10.43 $Y2=1.95
r196 38 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=1.02
+ $X2=9.465 $Y2=1.02
r197 37 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=1.02
+ $X2=10.43 $Y2=1.02
r198 37 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=10.345 $Y=1.02
+ $X2=9.63 $Y2=1.02
r199 35 60 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.465 $Y=1.395
+ $X2=9.465 $Y2=1.56
r200 35 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.465 $Y=1.395
+ $X2=9.465 $Y2=1.23
r201 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.465
+ $Y=1.395 $X2=9.465 $Y2=1.395
r202 32 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.465 $Y=1.105
+ $X2=9.465 $Y2=1.02
r203 32 34 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.465 $Y=1.105
+ $X2=9.465 $Y2=1.395
r204 30 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.3 $Y=1.02
+ $X2=9.465 $Y2=1.02
r205 30 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.3 $Y=1.02
+ $X2=8.545 $Y2=1.02
r206 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.46 $Y=0.935
+ $X2=8.545 $Y2=1.02
r207 28 29 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.46 $Y=0.51
+ $X2=8.46 $Y2=0.935
r208 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.375 $Y=0.425
+ $X2=8.46 $Y2=0.51
r209 26 27 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=8.375 $Y=0.425
+ $X2=6.485 $Y2=0.425
r210 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.4 $Y=0.51
+ $X2=6.485 $Y2=0.425
r211 24 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=6.4 $Y=0.51
+ $X2=6.4 $Y2=1.335
r212 23 49 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.265 $Y=1.42
+ $X2=5.125 $Y2=1.42
r213 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.315 $Y=1.42
+ $X2=6.4 $Y2=1.335
r214 22 23 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=6.315 $Y=1.42
+ $X2=5.265 $Y2=1.42
r215 20 60 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=9.51 $Y=2.46 $X2=9.51
+ $Y2=1.56
r216 17 59 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.445 $Y=0.75
+ $X2=9.445 $Y2=1.23
r217 11 53 38.8824 $w=2.71e-07 $l=2.07123e-07 $layer=POLY_cond $X=5.195 $Y=1.335
+ $X2=5.1 $Y2=1.5
r218 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.195 $Y=1.335
+ $X2=5.195 $Y2=0.87
r219 7 53 82.8133 $w=2.71e-07 $l=4.9135e-07 $layer=POLY_cond $X=4.98 $Y=1.935
+ $X2=5.1 $Y2=1.5
r220 7 9 235.169 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=4.98 $Y=1.935
+ $X2=4.98 $Y2=2.54
r221 2 47 600 $w=1.7e-07 $l=2.51744e-07 $layer=licon1_PDIFF $count=1 $X=10.555
+ $Y=1.84 $X2=10.685 $Y2=2.035
r222 1 43 182 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_NDIFF $count=1 $X=10.595
+ $Y=0.745 $X2=10.725 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%SET_B 1 3 6 8 10 14 16 17 22 26 27 31
c132 17 0 2.35896e-19 $X=5.665 $Y=2.035
c133 16 0 4.10562e-20 $X=8.735 $Y=2.035
c134 14 0 5.31324e-20 $X=9.015 $Y=0.75
r135 31 35 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=8.895 $Y=1.415
+ $X2=8.895 $Y2=2.035
r136 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.895
+ $Y=1.415 $X2=8.895 $Y2=1.415
r137 26 28 1.56494 $w=3.08e-07 $l=1e-08 $layer=POLY_cond $X=5.685 $Y=1.827
+ $X2=5.695 $Y2=1.827
r138 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.685
+ $Y=1.795 $X2=5.685 $Y2=1.795
r139 22 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r140 20 27 8.8997 $w=3.29e-07 $l=2.94754e-07 $layer=LI1_cond $X=5.52 $Y=2.035
+ $X2=5.642 $Y2=1.795
r141 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r142 17 19 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r143 16 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r144 16 17 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.665 $Y2=2.035
r145 12 30 38.7084 $w=3.43e-07 $l=2.11069e-07 $layer=POLY_cond $X=9.015 $Y=1.25
+ $X2=8.91 $Y2=1.415
r146 12 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.015 $Y=1.25
+ $X2=9.015 $Y2=0.75
r147 8 30 34.0194 $w=3.43e-07 $l=1.74714e-07 $layer=POLY_cond $X=8.89 $Y=1.58
+ $X2=8.91 $Y2=1.415
r148 8 10 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=8.89 $Y=1.58
+ $X2=8.89 $Y2=2.46
r149 4 28 19.5884 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=5.695 $Y=1.63
+ $X2=5.695 $Y2=1.827
r150 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.695 $Y=1.63
+ $X2=5.695 $Y2=0.87
r151 1 26 39.9058 $w=3.08e-07 $l=3.39875e-07 $layer=POLY_cond $X=5.43 $Y=2.025
+ $X2=5.685 $Y2=1.827
r152 1 3 137.906 $w=1.8e-07 $l=5.15e-07 $layer=POLY_cond $X=5.43 $Y=2.025
+ $X2=5.43 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_27_74# 1 2 10 13 15 16 20 21 23 24 27 29
+ 34 35 36 39 41 43 44 45 46 48 52 54 55 56 59 61 67 68
c184 68 0 1.96015e-20 $X=0.96 $Y=1.465
c185 41 0 1.51042e-19 $X=7.34 $Y=2.75
c186 36 0 7.44062e-20 $X=6.745 $Y=1.27
c187 35 0 1.71071e-19 $X=7.25 $Y=1.27
c188 20 0 6.36774e-20 $X=2.9 $Y=0.805
r189 68 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.465
+ $X2=0.96 $Y2=1.63
r190 68 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.465
+ $X2=0.96 $Y2=1.3
r191 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.465 $X2=0.96 $Y2=1.465
r192 64 67 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.75 $Y=1.465
+ $X2=0.96 $Y2=1.465
r193 60 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.63
+ $X2=0.75 $Y2=1.465
r194 60 61 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.75 $Y=1.63
+ $X2=0.75 $Y2=1.95
r195 59 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.3
+ $X2=0.75 $Y2=1.465
r196 58 59 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.75 $Y=1.13
+ $X2=0.75 $Y2=1.3
r197 57 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.035
+ $X2=0.27 $Y2=2.035
r198 56 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.75 $Y2=1.95
r199 56 57 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.435 $Y2=2.035
r200 54 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=1.045
+ $X2=0.75 $Y2=1.13
r201 54 55 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.665 $Y=1.045
+ $X2=0.365 $Y2=1.045
r202 50 55 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r203 50 52 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r204 46 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.12 $X2=0.27
+ $Y2=2.035
r205 46 48 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.27 $Y=2.12
+ $X2=0.27 $Y2=2.815
r206 39 45 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.34 $Y=1.89 $X2=7.34
+ $Y2=1.8
r207 39 41 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=7.34 $Y=1.89
+ $X2=7.34 $Y2=2.75
r208 37 45 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.325 $Y=1.345
+ $X2=7.325 $Y2=1.8
r209 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.25 $Y=1.27
+ $X2=7.325 $Y2=1.345
r210 35 36 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.25 $Y=1.27
+ $X2=6.745 $Y2=1.27
r211 32 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.67 $Y=1.195
+ $X2=6.745 $Y2=1.27
r212 32 34 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.67 $Y=1.195
+ $X2=6.67 $Y2=0.845
r213 31 34 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.67 $Y=0.255
+ $X2=6.67 $Y2=0.845
r214 27 44 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.54 $Y=2.055
+ $X2=3.54 $Y2=1.965
r215 27 29 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=3.54 $Y=2.055
+ $X2=3.54 $Y2=2.725
r216 25 44 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.525 $Y=1.815
+ $X2=3.525 $Y2=1.965
r217 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.45 $Y=1.74
+ $X2=3.525 $Y2=1.815
r218 23 24 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3.45 $Y=1.74
+ $X2=2.975 $Y2=1.74
r219 22 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.975 $Y=0.18
+ $X2=2.9 $Y2=0.18
r220 21 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.595 $Y=0.18
+ $X2=6.67 $Y2=0.255
r221 21 22 1856.21 $w=1.5e-07 $l=3.62e-06 $layer=POLY_cond $X=6.595 $Y=0.18
+ $X2=2.975 $Y2=0.18
r222 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.9 $Y=1.665
+ $X2=2.975 $Y2=1.74
r223 18 20 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.9 $Y=1.665
+ $X2=2.9 $Y2=0.805
r224 17 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.9 $Y=0.255
+ $X2=2.9 $Y2=0.18
r225 17 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.9 $Y=0.255
+ $X2=2.9 $Y2=0.805
r226 15 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.825 $Y=0.18
+ $X2=2.9 $Y2=0.18
r227 15 16 935.798 $w=1.5e-07 $l=1.825e-06 $layer=POLY_cond $X=2.825 $Y=0.18
+ $X2=1 $Y2=0.18
r228 13 72 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.945 $Y=2.4
+ $X2=0.945 $Y2=1.63
r229 10 71 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=0.74
+ $X2=0.925 $Y2=1.3
r230 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=1 $Y2=0.18
r231 7 10 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=0.925 $Y2=0.74
r232 2 63 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.115
r233 2 48 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r234 1 52 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_1534_446# 1 2 3 12 16 20 24 26 29 31 32 34
+ 35 37 40 42 49 50 53 54 56 60 61 62 67 70 71 75 76 77
c203 76 0 1.9889e-19 $X=11.42 $Y=1.485
c204 67 0 5.76555e-20 $X=11.3 $Y=2.29
c205 56 0 5.31324e-20 $X=11.215 $Y=0.68
c206 49 0 1.02788e-19 $X=8.055 $Y=2.215
c207 20 0 1.48333e-19 $X=11.435 $Y=2.4
c208 1 0 1.81011e-19 $X=9.52 $Y=0.38
r209 75 78 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.4 $Y=1.485
+ $X2=11.4 $Y2=1.65
r210 75 77 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.4 $Y=1.485
+ $X2=11.4 $Y2=1.32
r211 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.42
+ $Y=1.485 $X2=11.42 $Y2=1.485
r212 69 71 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=2.805
+ $X2=8.83 $Y2=2.805
r213 69 70 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=2.805
+ $X2=8.5 $Y2=2.805
r214 67 78 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=11.3 $Y=2.29
+ $X2=11.3 $Y2=1.65
r215 64 77 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=11.3 $Y=0.765
+ $X2=11.3 $Y2=1.32
r216 63 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.32 $Y=2.375
+ $X2=10.155 $Y2=2.375
r217 62 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.215 $Y=2.375
+ $X2=11.3 $Y2=2.29
r218 62 63 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=11.215 $Y=2.375
+ $X2=10.32 $Y2=2.375
r219 60 73 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.155 $Y=2.46
+ $X2=10.155 $Y2=2.375
r220 60 61 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=10.155 $Y=2.46
+ $X2=10.155 $Y2=2.63
r221 56 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.215 $Y=0.68
+ $X2=11.3 $Y2=0.765
r222 56 58 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=11.215 $Y=0.68
+ $X2=9.68 $Y2=0.68
r223 54 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.99 $Y=2.715
+ $X2=10.155 $Y2=2.63
r224 54 71 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=9.99 $Y=2.715
+ $X2=8.83 $Y2=2.715
r225 53 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.22 $Y=2.715
+ $X2=8.5 $Y2=2.715
r226 50 81 54.6151 $w=2.78e-07 $l=3.15e-07 $layer=POLY_cond $X=8.055 $Y=2.215
+ $X2=8.37 $Y2=2.215
r227 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=2.215 $X2=8.055 $Y2=2.215
r228 47 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.055 $Y=2.63
+ $X2=8.22 $Y2=2.715
r229 47 49 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.055 $Y=2.63
+ $X2=8.055 $Y2=2.215
r230 38 40 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=12.19 $Y=0.94
+ $X2=12.465 $Y2=0.94
r231 35 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.465 $Y=0.865
+ $X2=12.465 $Y2=0.94
r232 35 37 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.465 $Y=0.865
+ $X2=12.465 $Y2=0.58
r233 32 43 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=12.42 $Y=1.9
+ $X2=12.19 $Y2=1.9
r234 32 34 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=12.42 $Y=1.975
+ $X2=12.42 $Y2=2.47
r235 31 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=1.825
+ $X2=12.19 $Y2=1.9
r236 30 42 35.9208 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=12.19 $Y=1.635
+ $X2=12.19 $Y2=1.477
r237 30 31 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.19 $Y=1.635
+ $X2=12.19 $Y2=1.825
r238 29 42 35.9208 $w=1.5e-07 $l=1.57e-07 $layer=POLY_cond $X=12.19 $Y=1.32
+ $X2=12.19 $Y2=1.477
r239 28 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=1.015
+ $X2=12.19 $Y2=0.94
r240 28 29 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=12.19 $Y=1.015
+ $X2=12.19 $Y2=1.32
r241 27 76 3.33671 $w=3.15e-07 $l=1.68953e-07 $layer=POLY_cond $X=11.585
+ $Y=1.477 $X2=11.42 $Y2=1.485
r242 26 42 4.4846 $w=3.15e-07 $l=7.5e-08 $layer=POLY_cond $X=12.115 $Y=1.477
+ $X2=12.19 $Y2=1.477
r243 26 27 97.0896 $w=3.15e-07 $l=5.3e-07 $layer=POLY_cond $X=12.115 $Y=1.477
+ $X2=11.585 $Y2=1.477
r244 22 76 33.6231 $w=1.65e-07 $l=2.03101e-07 $layer=POLY_cond $X=11.505 $Y=1.32
+ $X2=11.42 $Y2=1.485
r245 22 24 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=11.505 $Y=1.32
+ $X2=11.505 $Y2=0.795
r246 18 76 33.6231 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=11.435 $Y=1.65
+ $X2=11.42 $Y2=1.485
r247 18 20 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=11.435 $Y=1.65
+ $X2=11.435 $Y2=2.4
r248 14 81 17.1848 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.37 $Y=2.05
+ $X2=8.37 $Y2=2.215
r249 14 16 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=8.37 $Y=2.05
+ $X2=8.37 $Y2=0.91
r250 10 50 51.1475 $w=2.78e-07 $l=3.68375e-07 $layer=POLY_cond $X=7.76 $Y=2.38
+ $X2=8.055 $Y2=2.215
r251 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.76 $Y=2.38
+ $X2=7.76 $Y2=2.75
r252 3 73 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=10.02
+ $Y=1.96 $X2=10.155 $Y2=2.455
r253 2 69 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=1.96 $X2=8.665 $Y2=2.805
r254 1 58 182 $w=1.7e-07 $l=3.71484e-07 $layer=licon1_NDIFF $count=1 $X=9.52
+ $Y=0.38 $X2=9.68 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_1349_114# 1 2 9 13 15 23 27 28 30 31 34 35
+ 36 38 39 40 43 44 47 48 49
c153 48 0 7.86413e-20 $X=7.137 $Y=2.1
c154 30 0 1.39048e-19 $X=8.12 $Y=1.73
c155 28 0 1.72728e-19 $X=7.415 $Y=1.815
c156 15 0 1.06435e-20 $X=8.035 $Y=0.845
r157 47 48 9.86413 $w=5.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.137 $Y=2.265
+ $X2=7.137 $Y2=2.1
r158 44 52 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.005 $Y=1.585
+ $X2=10.005 $Y2=1.75
r159 44 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.005 $Y=1.585
+ $X2=10.005 $Y2=1.42
r160 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.005
+ $Y=1.585 $X2=10.005 $Y2=1.585
r161 41 43 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=10.005 $Y=1.95
+ $X2=10.005 $Y2=1.585
r162 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.84 $Y=2.035
+ $X2=10.005 $Y2=1.95
r163 39 40 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=9.84 $Y=2.035
+ $X2=9.4 $Y2=2.035
r164 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=2.12
+ $X2=9.4 $Y2=2.035
r165 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.315 $Y=2.12
+ $X2=9.315 $Y2=2.29
r166 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.23 $Y=2.375
+ $X2=9.315 $Y2=2.29
r167 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.23 $Y=2.375
+ $X2=8.56 $Y2=2.375
r168 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=2.29
+ $X2=8.56 $Y2=2.375
r169 33 34 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.475 $Y=1.9
+ $X2=8.475 $Y2=2.29
r170 32 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.205 $Y=1.815
+ $X2=8.12 $Y2=1.815
r171 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.39 $Y=1.815
+ $X2=8.475 $Y2=1.9
r172 31 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.39 $Y=1.815
+ $X2=8.205 $Y2=1.815
r173 30 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=1.73
+ $X2=8.12 $Y2=1.815
r174 29 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.12 $Y=1.01
+ $X2=8.12 $Y2=1.73
r175 27 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.035 $Y=1.815
+ $X2=8.12 $Y2=1.815
r176 27 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.035 $Y=1.815
+ $X2=7.415 $Y2=1.815
r177 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.33 $Y=1.9
+ $X2=7.415 $Y2=1.815
r178 25 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.33 $Y=1.9 $X2=7.33
+ $Y2=2.1
r179 21 47 2.41371 $w=5.53e-07 $l=1.12e-07 $layer=LI1_cond $X=7.137 $Y=2.377
+ $X2=7.137 $Y2=2.265
r180 21 23 9.43932 $w=5.53e-07 $l=4.38e-07 $layer=LI1_cond $X=7.137 $Y=2.377
+ $X2=7.137 $Y2=2.815
r181 17 20 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=6.885 $Y=0.845
+ $X2=7.685 $Y2=0.845
r182 15 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.035 $Y=0.845
+ $X2=8.12 $Y2=1.01
r183 15 20 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.035 $Y=0.845
+ $X2=7.685 $Y2=0.845
r184 13 52 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=9.93 $Y=2.46
+ $X2=9.93 $Y2=1.75
r185 9 51 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=9.915 $Y=0.75
+ $X2=9.915 $Y2=1.42
r186 2 47 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=2.12 $X2=7.025 $Y2=2.265
r187 2 23 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=2.12 $X2=7.025 $Y2=2.815
r188 1 20 121.333 $w=1.7e-07 $l=1.06869e-06 $layer=licon1_NDIFF $count=1
+ $X=6.745 $Y=0.57 $X2=7.685 $Y2=0.845
r189 1 17 121.333 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1
+ $X=6.745 $Y=0.57 $X2=6.885 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%RESET_B 3 7 9 12 13
c37 7 0 1.78363e-19 $X=10.94 $Y=0.955
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.85 $Y=1.515
+ $X2=10.85 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.85 $Y=1.515
+ $X2=10.85 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.85
+ $Y=1.515 $X2=10.85 $Y2=1.515
r41 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=10.85 $Y=1.665
+ $X2=10.85 $Y2=1.515
r42 7 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.94 $Y=0.955
+ $X2=10.94 $Y2=1.35
r43 3 15 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=10.91 $Y=2.16
+ $X2=10.91 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_2412_410# 1 2 9 13 15 16 19 23 27 30
c56 15 0 1.18517e-19 $X=12.855 $Y=1.42
r57 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.67
+ $Y=1.42 $X2=12.67 $Y2=1.42
r58 25 30 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.36 $Y=1.42
+ $X2=12.235 $Y2=1.42
r59 25 27 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=12.36 $Y=1.42
+ $X2=12.67 $Y2=1.42
r60 21 30 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=12.235 $Y=1.585
+ $X2=12.235 $Y2=1.42
r61 21 23 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=12.235 $Y=1.585
+ $X2=12.235 $Y2=2.195
r62 17 30 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=12.235 $Y=1.255
+ $X2=12.235 $Y2=1.42
r63 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=12.235 $Y=1.255
+ $X2=12.235 $Y2=0.58
r64 15 28 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=12.855 $Y=1.42
+ $X2=12.67 $Y2=1.42
r65 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.855 $Y=1.42
+ $X2=12.945 $Y2=1.42
r66 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.96 $Y=1.255
+ $X2=12.945 $Y2=1.42
r67 11 13 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.96 $Y=1.255
+ $X2=12.96 $Y2=0.74
r68 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=12.945 $Y=1.585
+ $X2=12.945 $Y2=1.42
r69 7 9 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=12.945 $Y=1.585
+ $X2=12.945 $Y2=2.4
r70 2 23 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.06
+ $Y=2.05 $X2=12.195 $Y2=2.195
r71 1 19 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=12.12
+ $Y=0.37 $X2=12.25 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 52 53
+ 55 56 57 59 71 79 83 88 93 100 101 104 107 110 117 124 127
c157 27 0 1.96015e-20 $X=0.72 $Y=2.455
r158 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r159 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r160 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 117 120 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.2 $Y=3.055
+ $X2=9.2 $Y2=3.33
r162 107 108 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r163 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 101 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r165 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r166 98 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.805 $Y=3.33
+ $X2=12.68 $Y2=3.33
r167 98 100 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.805 $Y=3.33
+ $X2=13.2 $Y2=3.33
r168 97 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r169 97 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r170 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r171 94 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.21 $Y2=3.33
r172 94 96 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=12.24 $Y2=3.33
r173 93 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.555 $Y=3.33
+ $X2=12.68 $Y2=3.33
r174 93 96 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.555 $Y=3.33
+ $X2=12.24 $Y2=3.33
r175 92 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r176 92 121 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.36 $Y2=3.33
r177 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r178 89 120 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.365 $Y=3.33
+ $X2=9.2 $Y2=3.33
r179 89 91 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=9.365 $Y=3.33
+ $X2=10.8 $Y2=3.33
r180 88 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=3.33
+ $X2=11.21 $Y2=3.33
r181 88 91 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.045 $Y=3.33
+ $X2=10.8 $Y2=3.33
r182 87 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r183 87 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=7.92 $Y2=3.33
r184 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r185 84 86 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.27 $Y=3.33
+ $X2=8.88 $Y2=3.33
r186 83 120 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.035 $Y=3.33
+ $X2=9.2 $Y2=3.33
r187 83 86 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=9.035 $Y=3.33
+ $X2=8.88 $Y2=3.33
r188 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r189 79 84 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=8.087 $Y=3.33
+ $X2=8.27 $Y2=3.33
r190 79 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r191 79 110 8.68279 $w=3.63e-07 $l=2.75e-07 $layer=LI1_cond $X=8.087 $Y=3.33
+ $X2=8.087 $Y2=3.055
r192 79 81 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=6.48 $Y2=3.33
r193 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r194 78 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r195 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r196 75 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.205 $Y2=3.33
r197 75 77 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.37 $Y=3.33 $X2=6
+ $Y2=3.33
r198 74 108 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r199 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r200 71 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=5.205 $Y2=3.33
r201 71 73 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r203 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r204 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r205 67 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r207 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r208 64 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.72 $Y2=3.33
r209 64 66 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r210 62 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r211 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r212 59 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.72 $Y2=3.33
r213 59 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r214 57 114 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=7.92 $Y2=3.33
r215 57 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r216 55 77 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.02 $Y=3.33 $X2=6
+ $Y2=3.33
r217 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.02 $Y=3.33
+ $X2=6.185 $Y2=3.33
r218 54 81 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.48 $Y2=3.33
r219 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.185 $Y2=3.33
r220 52 69 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r221 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.38 $Y2=3.33
r222 51 73 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.64 $Y2=3.33
r223 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.38 $Y2=3.33
r224 47 50 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=12.68 $Y=1.985
+ $X2=12.68 $Y2=2.4
r225 45 127 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.68 $Y=3.245
+ $X2=12.68 $Y2=3.33
r226 45 50 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=12.68 $Y=3.245
+ $X2=12.68 $Y2=2.4
r227 41 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=3.245
+ $X2=11.21 $Y2=3.33
r228 41 43 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=11.21 $Y=3.245
+ $X2=11.21 $Y2=2.805
r229 37 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.185 $Y=3.245
+ $X2=6.185 $Y2=3.33
r230 37 39 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.185 $Y=3.245
+ $X2=6.185 $Y2=2.78
r231 33 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=3.245
+ $X2=5.205 $Y2=3.33
r232 33 35 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.205 $Y=3.245
+ $X2=5.205 $Y2=2.78
r233 29 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r234 29 31 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.74
r235 25 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r236 25 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.455
r237 8 50 300 $w=1.7e-07 $l=4.42719e-07 $layer=licon1_PDIFF $count=2 $X=12.51
+ $Y=2.05 $X2=12.72 $Y2=2.4
r238 8 47 600 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=1 $X=12.51
+ $Y=2.05 $X2=12.72 $Y2=1.985
r239 7 43 600 $w=1.7e-07 $l=1.06484e-06 $layer=licon1_PDIFF $count=1 $X=11
+ $Y=1.84 $X2=11.21 $Y2=2.805
r240 6 117 600 $w=1.7e-07 $l=1.19997e-06 $layer=licon1_PDIFF $count=1 $X=8.98
+ $Y=1.96 $X2=9.2 $Y2=3.055
r241 5 110 600 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=1 $X=7.85
+ $Y=2.54 $X2=8.085 $Y2=3.055
r242 4 39 600 $w=1.7e-07 $l=7.2208e-07 $layer=licon1_PDIFF $count=1 $X=6.055
+ $Y=2.12 $X2=6.185 $Y2=2.78
r243 3 35 600 $w=1.7e-07 $l=7.24362e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=2.12 $X2=5.205 $Y2=2.78
r244 2 31 600 $w=1.7e-07 $l=3.76032e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=2.515 $X2=2.38 $Y2=2.74
r245 1 27 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_311_119# 1 2 3 4 15 18 20 21 22 27 30 31
+ 32 34 36 41 42 44 47
r121 45 47 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.06 $Y=1.08
+ $X2=4.39 $Y2=1.08
r122 41 42 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.57
+ $X2=1.685 $Y2=2.405
r123 39 42 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=1.67 $Y=1.01
+ $X2=1.67 $Y2=2.405
r124 38 39 5.26419 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.925
+ $X2=1.725 $Y2=1.01
r125 36 38 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=1.725 $Y=0.79
+ $X2=1.725 $Y2=0.925
r126 33 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.39 $Y=1.165
+ $X2=4.39 $Y2=1.08
r127 33 34 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.39 $Y=1.165
+ $X2=4.39 $Y2=1.965
r128 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.305 $Y=2.05
+ $X2=4.39 $Y2=1.965
r129 31 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.305 $Y=2.05
+ $X2=4 $Y2=2.05
r130 30 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=0.995
+ $X2=4.06 $Y2=1.08
r131 29 30 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.06 $Y=0.615
+ $X2=4.06 $Y2=0.995
r132 25 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.875 $Y=2.135
+ $X2=4 $Y2=2.05
r133 25 27 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=3.875 $Y=2.135
+ $X2=3.875 $Y2=2.57
r134 22 44 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=3.64 $Y=0.435
+ $X2=3.46 $Y2=0.435
r135 22 24 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=0.435
+ $X2=3.77 $Y2=0.435
r136 21 29 8.02311 $w=3.6e-07 $l=2.18403e-07 $layer=LI1_cond $X=3.975 $Y=0.435
+ $X2=4.06 $Y2=0.615
r137 21 24 6.56252 $w=3.58e-07 $l=2.05e-07 $layer=LI1_cond $X=3.975 $Y=0.435
+ $X2=3.77 $Y2=0.435
r138 20 44 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.75 $Y=0.34
+ $X2=3.46 $Y2=0.34
r139 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.665 $Y=0.425
+ $X2=2.75 $Y2=0.34
r140 17 18 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.665 $Y=0.425
+ $X2=2.665 $Y2=0.84
r141 16 38 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.865 $Y=0.925
+ $X2=1.725 $Y2=0.925
r142 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.58 $Y=0.925
+ $X2=2.665 $Y2=0.84
r143 15 16 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.58 $Y=0.925
+ $X2=1.865 $Y2=0.925
r144 4 27 600 $w=1.7e-07 $l=2.30868e-07 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=2.515 $X2=3.835 $Y2=2.57
r145 3 41 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=2.425 $X2=1.7 $Y2=2.57
r146 2 24 182 $w=1.7e-07 $l=3.96169e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.595 $X2=3.77 $Y2=0.53
r147 1 36 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.595 $X2=1.7 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%Q_N 1 2 9 13 14 15 16 23 33
c35 33 0 2.54845e-19 $X=11.75 $Y=1.82
c36 14 0 6.25621e-20 $X=11.675 $Y=1.95
c37 9 0 1.78363e-19 $X=11.72 $Y=0.57
r38 21 35 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=11.75 $Y=1.995
+ $X2=11.75 $Y2=1.985
r39 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=11.75 $Y=1.995
+ $X2=11.75 $Y2=2.035
r40 16 30 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=11.75 $Y=2.775
+ $X2=11.75 $Y2=2.815
r41 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.75 $Y=2.405
+ $X2=11.75 $Y2=2.775
r42 14 35 0.42805 $w=3.48e-07 $l=1.3e-08 $layer=LI1_cond $X=11.75 $Y=1.972
+ $X2=11.75 $Y2=1.985
r43 14 33 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=11.75 $Y=1.972
+ $X2=11.75 $Y2=1.82
r44 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=11.75 $Y=2.057
+ $X2=11.75 $Y2=2.405
r45 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=11.75 $Y=2.057
+ $X2=11.75 $Y2=2.035
r46 13 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.84 $Y=1.15
+ $X2=11.84 $Y2=1.82
r47 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.74 $Y=0.965
+ $X2=11.74 $Y2=1.15
r48 7 9 12.3031 $w=3.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.74 $Y=0.965
+ $X2=11.74 $Y2=0.57
r49 2 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.525
+ $Y=1.84 $X2=11.66 $Y2=1.985
r50 2 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.525
+ $Y=1.84 $X2=11.66 $Y2=2.815
r51 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.58
+ $Y=0.425 $X2=11.72 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%Q 1 2 7 8 9 10 11 12 13
r15 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.172 $Y=2.405
+ $X2=13.172 $Y2=2.775
r16 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=13.172 $Y=1.985
+ $X2=13.172 $Y2=2.405
r17 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=13.172 $Y=1.665
+ $X2=13.172 $Y2=1.985
r18 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.172 $Y=1.295
+ $X2=13.172 $Y2=1.665
r19 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.172 $Y=0.925
+ $X2=13.172 $Y2=1.295
r20 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=13.172 $Y=0.515
+ $X2=13.172 $Y2=0.925
r21 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.035
+ $Y=1.84 $X2=13.17 $Y2=2.815
r22 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.035
+ $Y=1.84 $X2=13.17 $Y2=1.985
r23 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.035
+ $Y=0.37 $X2=13.175 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 43 45 50
+ 55 63 71 76 83 84 87 90 93 96 99 102
r130 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r131 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r132 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r133 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r134 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r135 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r136 84 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r137 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r138 81 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.83 $Y=0
+ $X2=12.705 $Y2=0
r139 81 83 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.83 $Y=0 $X2=13.2
+ $Y2=0
r140 80 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r141 80 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.28 $Y2=0
r142 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r143 77 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=11.22 $Y2=0
r144 77 79 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=12.24 $Y2=0
r145 76 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.58 $Y=0
+ $X2=12.705 $Y2=0
r146 76 79 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.58 $Y=0
+ $X2=12.24 $Y2=0
r147 75 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r148 75 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=8.88 $Y2=0
r149 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r150 72 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=0 $X2=8.8
+ $Y2=0
r151 72 74 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=8.885 $Y=0
+ $X2=10.8 $Y2=0
r152 71 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.22 $Y2=0
r153 71 74 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.8 $Y2=0
r154 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r155 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r156 67 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r157 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r158 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r159 64 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=5.98
+ $Y2=0
r160 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=6.48 $Y2=0
r161 63 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=0 $X2=8.8
+ $Y2=0
r162 63 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.715 $Y=0 $X2=8.4
+ $Y2=0
r163 62 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r164 61 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r165 59 62 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.52 $Y2=0
r166 59 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r167 58 61 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r168 58 59 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r169 56 90 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.227
+ $Y2=0
r170 56 58 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.64
+ $Y2=0
r171 55 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.98
+ $Y2=0
r172 55 61 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.52
+ $Y2=0
r173 54 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r174 54 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r175 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r176 51 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r177 51 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=1.68 $Y2=0
r178 50 90 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.227 $Y2=0
r179 50 53 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r180 48 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r181 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r182 45 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r183 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r184 43 70 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r185 43 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r186 39 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.705 $Y=0.085
+ $X2=12.705 $Y2=0
r187 39 41 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=12.705 $Y=0.085
+ $X2=12.705 $Y2=0.58
r188 35 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0
r189 35 37 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0.34
r190 31 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.8 $Y=0.085 $X2=8.8
+ $Y2=0
r191 31 33 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=8.8 $Y=0.085
+ $X2=8.8 $Y2=0.56
r192 27 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=0.085
+ $X2=5.98 $Y2=0
r193 27 29 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=5.98 $Y=0.085
+ $X2=5.98 $Y2=0.87
r194 23 90 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.227 $Y=0.085
+ $X2=2.227 $Y2=0
r195 23 25 13.261 $w=3.63e-07 $l=4.2e-07 $layer=LI1_cond $X=2.227 $Y=0.085
+ $X2=2.227 $Y2=0.505
r196 19 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r197 19 21 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.625
r198 6 41 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.37 $X2=12.745 $Y2=0.58
r199 5 37 182 $w=1.7e-07 $l=4.97041e-07 $layer=licon1_NDIFF $count=1 $X=11.015
+ $Y=0.745 $X2=11.22 $Y2=0.34
r200 4 33 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=8.445
+ $Y=0.7 $X2=8.8 $Y2=0.56
r201 3 29 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=5.77
+ $Y=0.595 $X2=5.98 $Y2=0.87
r202 2 25 182 $w=1.7e-07 $l=2.7636e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.595 $X2=2.225 $Y2=0.505
r203 1 21 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_867_119# 1 2 9 11 12 15
r29 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.48 $Y=0.425
+ $X2=5.48 $Y2=0.87
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.315 $Y=0.34
+ $X2=5.48 $Y2=0.425
r31 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.315 $Y=0.34
+ $X2=4.645 $Y2=0.34
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.48 $Y=0.425
+ $X2=4.645 $Y2=0.34
r33 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.48 $Y=0.425
+ $X2=4.48 $Y2=0.74
r34 2 15 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=5.27
+ $Y=0.595 $X2=5.48 $Y2=0.87
r35 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.595 $X2=4.48 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBN_1%A_1818_76# 1 2 9 11 13
c20 9 0 5.09967e-20 $X=9.23 $Y=0.56
c21 1 0 3.13464e-19 $X=9.09 $Y=0.38
r22 11 13 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.315 $Y=0.34
+ $X2=10.195 $Y2=0.34
r23 7 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.19 $Y=0.425
+ $X2=9.315 $Y2=0.34
r24 7 9 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=9.19 $Y=0.425
+ $X2=9.19 $Y2=0.56
r25 2 13 182 $w=1.7e-07 $l=2.24109e-07 $layer=licon1_NDIFF $count=1 $X=9.99
+ $Y=0.38 $X2=10.195 $Y2=0.34
r26 1 9 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.09 $Y=0.38
+ $X2=9.23 $Y2=0.56
.ends


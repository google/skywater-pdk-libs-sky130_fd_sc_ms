* NGSPICE file created from sky130_fd_sc_ms__or3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__or3b_2 A B C_N VGND VNB VPB VPWR X
M1000 a_190_260# a_27_368# VGND VNB nlowvt w=640000u l=150000u
+  ad=4.064e+11p pd=3.83e+06u as=9.1395e+11p ps=6.95e+06u
M1001 a_461_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=9.8195e+11p ps=6.3e+06u
M1002 VPWR C_N a_27_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1003 a_545_368# B a_461_368# VPB pshort w=1e+06u l=180000u
+  ad=3.6e+11p pd=2.72e+06u as=0p ps=0u
M1004 X a_190_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1005 VGND C_N a_27_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 VGND B a_190_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_190_260# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_190_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_190_260# a_27_368# a_545_368# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1010 X a_190_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VPWR a_190_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a22oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__a22oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.430000 0.880000 1.780000 ;
        RECT 0.710000 1.780000 0.880000 1.950000 ;
        RECT 0.710000 1.950000 2.210000 2.120000 ;
        RECT 1.880000 1.430000 2.210000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.430000 1.420000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.090000 4.075000 1.260000 ;
        RECT 2.720000 1.260000 3.235000 1.550000 ;
        RECT 3.905000 1.260000 4.075000 1.300000 ;
        RECT 3.905000 1.300000 4.370000 1.630000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.430000 3.735000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.430200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.285000 0.350000 0.535000 1.090000 ;
        RECT 0.285000 1.090000 2.550000 1.260000 ;
        RECT 2.040000 0.810000 2.550000 1.090000 ;
        RECT 2.145000 0.350000 2.550000 0.810000 ;
        RECT 2.380000 1.260000 2.550000 1.720000 ;
        RECT 2.380000 1.720000 3.130000 1.890000 ;
        RECT 2.930000 1.890000 3.130000 1.950000 ;
        RECT 2.930000 1.950000 4.710000 2.120000 ;
        RECT 2.930000 2.120000 3.130000 2.735000 ;
        RECT 3.860000 2.120000 4.030000 2.735000 ;
        RECT 4.245000 0.350000 4.710000 1.130000 ;
        RECT 4.540000 1.130000 4.710000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.800000 0.085000 ;
        RECT 1.145000  0.085000 1.475000 0.580000 ;
        RECT 3.305000  0.085000 3.635000 0.580000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.800000 3.415000 ;
        RECT 0.740000 2.630000 0.990000 3.245000 ;
        RECT 1.690000 2.630000 2.230000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.290000 1.950000 0.540000 2.290000 ;
      RECT 0.290000 2.290000 2.730000 2.460000 ;
      RECT 0.290000 2.460000 0.540000 2.980000 ;
      RECT 0.715000 0.330000 0.965000 0.750000 ;
      RECT 0.715000 0.750000 1.815000 0.920000 ;
      RECT 1.190000 2.460000 1.520000 2.980000 ;
      RECT 1.645000 0.350000 1.975000 0.640000 ;
      RECT 1.645000 0.640000 1.815000 0.750000 ;
      RECT 2.400000 2.060000 2.730000 2.290000 ;
      RECT 2.400000 2.460000 2.730000 2.905000 ;
      RECT 2.400000 2.905000 4.560000 3.075000 ;
      RECT 2.835000 0.330000 3.135000 0.750000 ;
      RECT 2.835000 0.750000 4.065000 0.920000 ;
      RECT 3.330000 2.290000 3.660000 2.905000 ;
      RECT 3.815000 0.330000 4.065000 0.750000 ;
      RECT 4.230000 2.290000 4.560000 2.905000 ;
  END
END sky130_fd_sc_ms__a22oi_2

* NGSPICE file created from sky130_fd_sc_ms__dlxbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_887_270# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.3791e+12p pd=1.953e+07u as=3.024e+11p ps=2.78e+06u
M1001 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.0325e+12p ps=1.669e+07u
M1002 Q a_887_270# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 Q_N a_1442_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1004 VGND a_232_98# a_343_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.817e+11p ps=2.29e+06u
M1005 VPWR a_1442_94# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_817_392# a_232_98# a_647_79# VPB pshort w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=4.159e+11p ps=3.29e+06u
M1007 Q_N a_1442_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 VGND a_887_270# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_887_270# a_647_79# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1010 a_1442_94# a_887_270# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1011 a_568_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1012 a_569_79# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1013 a_647_79# a_232_98# a_569_79# VNB nlowvt w=640000u l=150000u
+  ad=3.952e+11p pd=2.9e+06u as=0p ps=0u
M1014 VGND a_1442_94# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_887_270# a_647_79# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 a_1442_94# a_887_270# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1017 a_647_79# a_343_74# a_568_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1019 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1020 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=3.066e+11p ps=2.41e+06u
M1021 VPWR a_887_270# a_817_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_887_270# a_839_123# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1023 VPWR a_232_98# a_343_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1024 Q a_887_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_839_123# a_343_74# a_647_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__dfxbp_2.spice
* Created: Fri Aug 28 17:24:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfxbp_2.pex.spice"
.subckt sky130_fd_sc_ms__dfxbp_2  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_CLK_M1031_g N_A_27_74#_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.20385 AS=0.2109 PD=1.355 PS=2.05 NRD=17.832 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1013 N_A_209_368#_M1013_d N_A_27_74#_M1013_g N_VGND_M1031_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.3252 AS=0.20385 PD=2.59 PS=1.355 NRD=62.34 NRS=4.86 M=1 R=4.93333
+ SA=75000.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1030 N_A_454_503#_M1030_d N_D_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.35635 PD=0.7 PS=2.6 NRD=0 NRS=226.692 M=1 R=2.8 SA=75000.5
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1032 N_A_561_445#_M1032_d N_A_27_74#_M1032_g N_A_454_503#_M1030_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0830375 AS=0.0588 PD=0.865 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1020 A_717_102# N_A_209_368#_M1020_g N_A_561_445#_M1032_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0830375 PD=0.66 PS=0.865 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75001.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_753_284#_M1002_g A_717_102# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0850825 AS=0.0504 PD=0.801031 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1005 N_A_753_284#_M1005_d N_A_561_445#_M1005_g N_VGND_M1002_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.1935 AS=0.111418 PD=1.49 PS=1.04897 NRD=64.752 NRS=2.172
+ M=1 R=3.66667 SA=75001.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1018 N_A_1003_424#_M1018_d N_A_209_368#_M1018_g N_A_753_284#_M1005_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.222296 AS=0.1935 PD=1.90515 PS=1.49 NRD=157.08
+ NRS=64.752 M=1 R=3.66667 SA=75002.3 SB=75001 A=0.0825 P=1.4 MULT=1
MM1000 A_1248_128# N_A_27_74#_M1000_g N_A_1003_424#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.169754 PD=0.63 PS=1.45485 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_1290_102#_M1009_g A_1248_128# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1533 AS=0.0441 PD=1.57 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_1003_424#_M1028_g N_A_1290_102#_M1028_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.12025 AS=0.2109 PD=1.065 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_Q_M1001_d N_A_1290_102#_M1001_g N_VGND_M1028_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12025 PD=1.02 PS=1.065 NRD=0 NRS=7.296 M=1 R=4.93333 SA=75000.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1019 N_Q_M1001_d N_A_1290_102#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_1290_102#_M1021_g N_A_1835_368#_M1021_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.118058 AS=0.15675 PD=0.976357 PS=1.67 NRD=27.816 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1003 N_Q_N_M1003_d N_A_1835_368#_M1003_g N_VGND_M1021_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.158842 PD=1.02 PS=1.31364 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_Q_N_M1003_d N_A_1835_368#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_27_74#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_A_209_368#_M1011_d N_A_27_74#_M1011_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1004 N_A_454_503#_M1004_d N_D_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=0.42
+ AD=0.099925 AS=0.3171 PD=1.065 PS=2.35 NRD=85.7935 NRS=328.32 M=1 R=2.33333
+ SA=90000.4 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1024 N_A_561_445#_M1024_d N_A_209_368#_M1024_g N_A_454_503#_M1004_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1134 AS=0.099925 PD=0.96 PS=1.065 NRD=65.6601 NRS=0 M=1
+ R=2.33333 SA=90000.4 SB=90004.5 A=0.0756 P=1.2 MULT=1
MM1012 A_705_445# N_A_27_74#_M1012_g N_A_561_445#_M1024_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.1134 PD=0.66 PS=0.96 NRD=30.4759 NRS=56.2829 M=1
+ R=2.33333 SA=90001.1 SB=90003.8 A=0.0756 P=1.2 MULT=1
MM1029 N_VPWR_M1029_d N_A_753_284#_M1029_g A_705_445# VPB PSHORT L=0.18 W=0.42
+ AD=0.131392 AS=0.0504 PD=1.01 PS=0.66 NRD=120.919 NRS=30.4759 M=1 R=2.33333
+ SA=90001.6 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1014 N_A_753_284#_M1014_d N_A_561_445#_M1014_g N_VPWR_M1029_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.262783 PD=1.11 PS=2.02 NRD=0 NRS=60.4593 M=1
+ R=4.66667 SA=90001.2 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1015 N_A_1003_424#_M1015_d N_A_27_74#_M1015_g N_A_753_284#_M1014_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.3108 AS=0.1134 PD=2.26667 PS=1.11 NRD=90.2851 NRS=0 M=1
+ R=4.66667 SA=90001.7 SB=90002 A=0.1512 P=2.04 MULT=1
MM1025 A_1211_479# N_A_209_368#_M1025_g N_A_1003_424#_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.08295 AS=0.1554 PD=0.815 PS=1.13333 NRD=66.8224 NRS=91.4474 M=1
+ R=2.33333 SA=90003 SB=90002.8 A=0.0756 P=1.2 MULT=1
MM1026 N_VPWR_M1026_d N_A_1290_102#_M1026_g A_1211_479# VPB PSHORT L=0.18 W=0.42
+ AD=0.0882 AS=0.08295 PD=0.813333 PS=0.815 NRD=0 NRS=66.8224 M=1 R=2.33333
+ SA=90003.6 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1008 N_A_1290_102#_M1008_d N_A_1003_424#_M1008_g N_VPWR_M1026_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.1764 PD=1.11 PS=1.62667 NRD=0 NRS=24.625 M=1
+ R=4.66667 SA=90002.1 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1017 N_A_1290_102#_M1008_d N_A_1003_424#_M1017_g N_VPWR_M1017_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.1578 PD=1.11 PS=1.26429 NRD=0 NRS=18.7544 M=1
+ R=4.66667 SA=90002.6 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1022 N_Q_M1022_d N_A_1290_102#_M1022_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2104 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1023 N_Q_M1022_d N_A_1290_102#_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_A_1290_102#_M1016_g N_A_1835_368#_M1016_s VPB PSHORT
+ L=0.18 W=1 AD=0.183302 AS=0.28 PD=1.39151 PS=2.56 NRD=16.0752 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1016_d N_A_1835_368#_M1007_g N_Q_N_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.205298 AS=0.1512 PD=1.55849 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1027 N_VPWR_M1027_d N_A_1835_368#_M1027_g N_Q_N_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3192 AS=0.1512 PD=2.81 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX33_noxref VNB VPB NWDIODE A=20.8198 P=27.12
c_135 VNB 0 8.25183e-20 $X=0 $Y=0
c_222 VPB 0 6.95252e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dfxbp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__or3b_1.spice
* Created: Fri Aug 28 18:07:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or3b_1.pex.spice"
.subckt sky130_fd_sc_ms__or3b_1  VNB VPB C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1007 N_A_127_74#_M1007_d N_C_N_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.1595 AS=0.1925 PD=1.68 PS=1.8 NRD=1.08 NRS=14.172 M=1 R=3.66667
+ SA=75000.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_A_127_74#_M1004_g N_A_239_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.1155 AS=0.15675 PD=0.97 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002 A=0.0825 P=1.4 MULT=1
MM1000 N_A_239_74#_M1000_d N_B_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.086625 AS=0.1155 PD=0.865 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.8 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_239_74#_M1000_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.162122 AS=0.086625 PD=1.1469 PS=0.865 NRD=31.632 NRS=7.632 M=1 R=3.66667
+ SA=75001.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1006 N_X_M1006_d N_A_239_74#_M1006_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.218128 PD=2.05 PS=1.5431 NRD=0 NRS=29.184 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_127_74#_M1008_d N_C_N_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2436 AS=0.2688 PD=2.26 PS=2.32 NRD=1.1623 NRS=8.1952 M=1 R=4.66667
+ SA=90000.2 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1009 A_371_391# N_A_127_74#_M1009_g N_A_239_74#_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1001 A_455_391# N_B_M1001_g A_371_391# VPB PSHORT L=0.18 W=1 AD=0.12 AS=0.12
+ PD=1.24 PS=1.24 NRD=12.7853 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90001.2
+ A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_455_391# VPB PSHORT L=0.18 W=1 AD=0.209717
+ AS=0.12 PD=1.43868 PS=1.24 NRD=15.7403 NRS=12.7853 M=1 R=5.55556 SA=90001
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_239_74#_M1003_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.234883 PD=2.8 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__or3b_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__bufinv_8.pxi.spice
* Created: Fri Aug 28 17:16:44 2020
* 
x_PM_SKY130_FD_SC_MS__BUFINV_8%A N_A_M1007_g N_A_M1023_g A N_A_c_117_n
+ N_A_c_118_n PM_SKY130_FD_SC_MS__BUFINV_8%A
x_PM_SKY130_FD_SC_MS__BUFINV_8%A_183_48# N_A_183_48#_M1010_d N_A_183_48#_M1019_d
+ N_A_183_48#_M1000_d N_A_183_48#_M1005_d N_A_183_48#_M1006_g
+ N_A_183_48#_M1001_g N_A_183_48#_M1009_g N_A_183_48#_M1002_g
+ N_A_183_48#_M1003_g N_A_183_48#_M1013_g N_A_183_48#_M1008_g
+ N_A_183_48#_M1014_g N_A_183_48#_M1011_g N_A_183_48#_M1018_g
+ N_A_183_48#_M1012_g N_A_183_48#_M1020_g N_A_183_48#_M1016_g
+ N_A_183_48#_M1021_g N_A_183_48#_M1017_g N_A_183_48#_M1022_g
+ N_A_183_48#_c_164_n N_A_183_48#_c_165_n N_A_183_48#_c_166_n
+ N_A_183_48#_c_167_n N_A_183_48#_c_168_n N_A_183_48#_c_194_p
+ N_A_183_48#_c_169_n N_A_183_48#_c_170_n N_A_183_48#_c_182_n
+ N_A_183_48#_c_183_n N_A_183_48#_c_171_n N_A_183_48#_c_184_n
+ N_A_183_48#_c_172_n PM_SKY130_FD_SC_MS__BUFINV_8%A_183_48#
x_PM_SKY130_FD_SC_MS__BUFINV_8%A_27_368# N_A_27_368#_M1023_s N_A_27_368#_M1007_s
+ N_A_27_368#_c_393_n N_A_27_368#_M1000_g N_A_27_368#_M1010_g
+ N_A_27_368#_M1004_g N_A_27_368#_M1015_g N_A_27_368#_c_385_n
+ N_A_27_368#_M1005_g N_A_27_368#_M1019_g N_A_27_368#_c_397_n
+ N_A_27_368#_c_388_n N_A_27_368#_c_389_n N_A_27_368#_c_390_n
+ N_A_27_368#_c_410_n N_A_27_368#_c_391_n N_A_27_368#_c_451_n
+ N_A_27_368#_c_462_n N_A_27_368#_c_399_n N_A_27_368#_c_400_n
+ N_A_27_368#_c_401_n N_A_27_368#_c_480_p N_A_27_368#_c_392_n
+ PM_SKY130_FD_SC_MS__BUFINV_8%A_27_368#
x_PM_SKY130_FD_SC_MS__BUFINV_8%VPWR N_VPWR_M1007_d N_VPWR_M1002_d N_VPWR_M1008_d
+ N_VPWR_M1012_d N_VPWR_M1017_d N_VPWR_M1004_s N_VPWR_c_538_n N_VPWR_c_539_n
+ N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n
+ N_VPWR_c_545_n VPWR N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n
+ N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_537_n N_VPWR_c_553_n
+ N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ PM_SKY130_FD_SC_MS__BUFINV_8%VPWR
x_PM_SKY130_FD_SC_MS__BUFINV_8%Y N_Y_M1006_d N_Y_M1013_d N_Y_M1018_d N_Y_M1021_d
+ N_Y_M1001_s N_Y_M1003_s N_Y_M1011_s N_Y_M1016_s N_Y_c_636_n N_Y_c_645_n
+ N_Y_c_637_n N_Y_c_638_n N_Y_c_639_n N_Y_c_640_n N_Y_c_641_n N_Y_c_680_n
+ N_Y_c_642_n N_Y_c_643_n Y Y Y Y PM_SKY130_FD_SC_MS__BUFINV_8%Y
x_PM_SKY130_FD_SC_MS__BUFINV_8%VGND N_VGND_M1023_d N_VGND_M1009_s N_VGND_M1014_s
+ N_VGND_M1020_s N_VGND_M1022_s N_VGND_M1015_s N_VGND_c_739_n N_VGND_c_740_n
+ N_VGND_c_741_n N_VGND_c_742_n N_VGND_c_743_n N_VGND_c_744_n VGND
+ N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n
+ N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n N_VGND_c_754_n
+ N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ PM_SKY130_FD_SC_MS__BUFINV_8%VGND
cc_1 VNB N_A_M1023_g 0.0327781f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_2 VNB N_A_c_117_n 0.0340561f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_3 VNB N_A_c_118_n 0.0147537f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_183_48#_M1006_g 0.0215966f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.68
cc_5 VNB N_A_183_48#_M1001_g 0.00151588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_183_48#_M1009_g 0.0213269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_183_48#_M1002_g 0.00142151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_183_48#_M1003_g 0.00154131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_183_48#_M1013_g 0.0211937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_183_48#_M1008_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_183_48#_M1014_g 0.0212282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_183_48#_M1011_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_183_48#_M1018_g 0.0217898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_183_48#_M1012_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_183_48#_M1020_g 0.0217898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_183_48#_M1016_g 0.00168816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_183_48#_M1021_g 0.022104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_183_48#_M1017_g 0.00181543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_183_48#_M1022_g 0.0231611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_183_48#_c_164_n 0.00862531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_183_48#_c_165_n 0.00197374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_183_48#_c_166_n 0.00209186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_183_48#_c_167_n 0.00496443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_183_48#_c_168_n 0.00313284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_183_48#_c_169_n 0.0227723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_183_48#_c_170_n 0.0220728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_183_48#_c_171_n 0.0104445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_183_48#_c_172_n 0.177993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_368#_M1010_g 0.0216729f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_30 VNB N_A_27_368#_M1004_g 4.21584e-19 $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_31 VNB N_A_27_368#_M1015_g 0.022431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_368#_c_385_n 0.0691761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_368#_M1005_g 5.97508e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_368#_M1019_g 0.0287448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_368#_c_388_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_368#_c_389_n 0.00538315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_368#_c_390_n 0.00909915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_368#_c_391_n 0.00862727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_368#_c_392_n 0.00269557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_537_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_636_n 0.00381057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_637_n 0.00195975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_638_n 0.00309972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_639_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_640_n 0.0053906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_641_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_642_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_643_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB Y 0.00257348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_739_n 0.00571296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_740_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_741_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_742_n 0.00516528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_743_n 0.00500818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_744_n 0.00570743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_745_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_746_n 0.0186748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_747_n 0.0150174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_748_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_749_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_750_n 0.0153775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_751_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_752_n 0.345062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_753_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_754_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_755_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_756_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_757_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_758_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VPB N_A_M1007_g 0.0289575f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_71 VPB N_A_c_117_n 0.00735861f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_72 VPB N_A_c_118_n 0.00730023f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_73 VPB N_A_183_48#_M1001_g 0.0219028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_183_48#_M1002_g 0.0208608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_183_48#_M1003_g 0.0214391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_183_48#_M1008_g 0.0214644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_183_48#_M1011_g 0.0214644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_183_48#_M1012_g 0.0214644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_183_48#_M1016_g 0.0229973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_183_48#_M1017_g 0.0241007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_183_48#_c_170_n 0.018854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_183_48#_c_182_n 0.0275857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_183_48#_c_183_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_183_48#_c_184_n 0.00704942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_27_368#_c_393_n 0.0184948f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_86 VPB N_A_27_368#_M1004_g 0.0214904f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.515
cc_87 VPB N_A_27_368#_c_385_n 0.00453292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_27_368#_M1005_g 0.0278853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_368#_c_397_n 0.0242446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_368#_c_391_n 0.00330443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_368#_c_399_n 0.00301616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_368#_c_400_n 0.00194157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_368#_c_401_n 0.0179584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_368#_c_392_n 0.00273704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_538_n 0.00568435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_539_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_540_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_541_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_542_n 0.00565985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_543_n 0.00565985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_544_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_545_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_546_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_547_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_548_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_549_n 0.0218958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_550_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_551_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_537_n 0.104262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_553_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_554_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_555_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_556_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_557_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_Y_c_645_n 0.0147266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 N_A_M1023_g N_A_183_48#_M1006_g 0.0228206f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_M1007_g N_A_183_48#_M1001_g 0.0226736f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_c_117_n N_A_183_48#_c_172_n 0.0226736f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A_M1007_g N_A_27_368#_c_397_n 0.00852848f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_M1023_g N_A_27_368#_c_388_n 0.00159319f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_M1023_g N_A_27_368#_c_389_n 0.0146911f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_c_117_n N_A_27_368#_c_389_n 7.98718e-19 $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_c_118_n N_A_27_368#_c_389_n 0.012562f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_c_117_n N_A_27_368#_c_390_n 0.00126636f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_c_118_n N_A_27_368#_c_390_n 0.0219605f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_M1007_g N_A_27_368#_c_410_n 0.0162204f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_c_118_n N_A_27_368#_c_410_n 0.00339179f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_M1023_g N_A_27_368#_c_391_n 0.00374261f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_c_117_n N_A_27_368#_c_391_n 0.00926348f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_c_118_n N_A_27_368#_c_391_n 0.0329132f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_M1007_g N_A_27_368#_c_401_n 0.00533924f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_c_117_n N_A_27_368#_c_401_n 0.00105714f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_118_n N_A_27_368#_c_401_n 0.0254422f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_M1007_g N_VPWR_c_538_n 0.00345319f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_M1007_g N_VPWR_c_546_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_M1007_g N_VPWR_c_537_n 0.00985902f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_M1023_g Y 3.41373e-19 $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_M1023_g Y 6.75874e-19 $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_M1023_g N_VGND_c_739_n 0.0132976f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_M1023_g N_VGND_c_745_n 0.00383152f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_M1023_g N_VGND_c_752_n 0.00761248f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_183_48#_c_183_n N_A_27_368#_c_393_n 0.0139051f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_143 N_A_183_48#_M1022_g N_A_27_368#_M1010_g 0.0189902f $X=4.3 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_183_48#_c_164_n N_A_27_368#_M1010_g 7.44057e-19 $X=4.65 $Y=1.465
+ $X2=0 $Y2=0
cc_145 N_A_183_48#_c_165_n N_A_27_368#_M1010_g 0.00529113f $X=4.735 $Y=1.3 $X2=0
+ $Y2=0
cc_146 N_A_183_48#_c_166_n N_A_27_368#_M1010_g 4.16154e-19 $X=5.02 $Y=0.515
+ $X2=0 $Y2=0
cc_147 N_A_183_48#_c_168_n N_A_27_368#_M1010_g 0.0132602f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_148 N_A_183_48#_c_194_p N_A_27_368#_M1004_g 0.013221f $X=5.795 $Y=2.225 $X2=0
+ $Y2=0
cc_149 N_A_183_48#_c_170_n N_A_27_368#_M1004_g 0.00101477f $X=5.96 $Y=1.985
+ $X2=0 $Y2=0
cc_150 N_A_183_48#_c_183_n N_A_27_368#_M1004_g 0.0119601f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_151 N_A_183_48#_c_165_n N_A_27_368#_M1015_g 9.46656e-19 $X=4.735 $Y=1.3 $X2=0
+ $Y2=0
cc_152 N_A_183_48#_c_166_n N_A_27_368#_M1015_g 4.16154e-19 $X=5.02 $Y=0.515
+ $X2=0 $Y2=0
cc_153 N_A_183_48#_c_167_n N_A_27_368#_M1015_g 0.0153525f $X=5.795 $Y=1.005
+ $X2=0 $Y2=0
cc_154 N_A_183_48#_c_169_n N_A_27_368#_M1015_g 5.56882e-19 $X=5.96 $Y=0.515
+ $X2=0 $Y2=0
cc_155 N_A_183_48#_c_170_n N_A_27_368#_M1015_g 8.9077e-19 $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A_183_48#_M1017_g N_A_27_368#_c_385_n 0.036748f $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_157 N_A_183_48#_c_164_n N_A_27_368#_c_385_n 0.0140069f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_158 N_A_183_48#_c_167_n N_A_27_368#_c_385_n 0.00120405f $X=5.795 $Y=1.005
+ $X2=0 $Y2=0
cc_159 N_A_183_48#_c_168_n N_A_27_368#_c_385_n 0.00135031f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_160 N_A_183_48#_c_194_p N_A_27_368#_c_385_n 4.93656e-19 $X=5.795 $Y=2.225
+ $X2=0 $Y2=0
cc_161 N_A_183_48#_c_170_n N_A_27_368#_c_385_n 0.0125303f $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_183_48#_c_183_n N_A_27_368#_c_385_n 3.12521e-19 $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_163 N_A_183_48#_c_172_n N_A_27_368#_c_385_n 0.0189902f $X=4.3 $Y=1.465 $X2=0
+ $Y2=0
cc_164 N_A_183_48#_c_194_p N_A_27_368#_M1005_g 0.0168909f $X=5.795 $Y=2.225
+ $X2=0 $Y2=0
cc_165 N_A_183_48#_c_170_n N_A_27_368#_M1005_g 0.0108941f $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_183_48#_c_182_n N_A_27_368#_M1005_g 9.97796e-19 $X=5.96 $Y=2.4 $X2=0
+ $Y2=0
cc_167 N_A_183_48#_c_183_n N_A_27_368#_M1005_g 6.3423e-19 $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_168 N_A_183_48#_c_184_n N_A_27_368#_M1005_g 0.00242337f $X=5.96 $Y=2.225
+ $X2=0 $Y2=0
cc_169 N_A_183_48#_c_167_n N_A_27_368#_M1019_g 0.0176987f $X=5.795 $Y=1.005
+ $X2=0 $Y2=0
cc_170 N_A_183_48#_c_169_n N_A_27_368#_M1019_g 0.00889319f $X=5.96 $Y=0.515
+ $X2=0 $Y2=0
cc_171 N_A_183_48#_c_170_n N_A_27_368#_M1019_g 0.00744164f $X=5.96 $Y=1.985
+ $X2=0 $Y2=0
cc_172 N_A_183_48#_c_171_n N_A_27_368#_M1019_g 9.50735e-19 $X=5.96 $Y=1.005
+ $X2=0 $Y2=0
cc_173 N_A_183_48#_M1006_g N_A_27_368#_c_389_n 0.00116372f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_183_48#_M1006_g N_A_27_368#_c_391_n 0.00814278f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_183_48#_M1001_g N_A_27_368#_c_451_n 0.0209348f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_176 N_A_183_48#_M1002_g N_A_27_368#_c_451_n 0.0162594f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_177 N_A_183_48#_M1003_g N_A_27_368#_c_451_n 0.0162741f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_178 N_A_183_48#_M1008_g N_A_27_368#_c_451_n 0.0162741f $X=2.355 $Y=2.4 $X2=0
+ $Y2=0
cc_179 N_A_183_48#_M1011_g N_A_27_368#_c_451_n 0.0162741f $X=2.805 $Y=2.4 $X2=0
+ $Y2=0
cc_180 N_A_183_48#_M1012_g N_A_27_368#_c_451_n 0.0162741f $X=3.255 $Y=2.4 $X2=0
+ $Y2=0
cc_181 N_A_183_48#_M1016_g N_A_27_368#_c_451_n 0.0169687f $X=3.705 $Y=2.4 $X2=0
+ $Y2=0
cc_182 N_A_183_48#_M1017_g N_A_27_368#_c_451_n 0.0186541f $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_183 N_A_183_48#_c_164_n N_A_27_368#_c_451_n 0.00405996f $X=4.65 $Y=1.465
+ $X2=0 $Y2=0
cc_184 N_A_183_48#_c_183_n N_A_27_368#_c_451_n 0.00976092f $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_185 N_A_183_48#_c_172_n N_A_27_368#_c_451_n 2.59519e-19 $X=4.3 $Y=1.465 $X2=0
+ $Y2=0
cc_186 N_A_183_48#_c_183_n N_A_27_368#_c_462_n 0.00531798f $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_187 N_A_183_48#_M1000_d N_A_27_368#_c_399_n 9.26908e-19 $X=4.875 $Y=1.84
+ $X2=0 $Y2=0
cc_188 N_A_183_48#_c_164_n N_A_27_368#_c_399_n 0.0197805f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_189 N_A_183_48#_c_168_n N_A_27_368#_c_399_n 0.0046576f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_190 N_A_183_48#_c_183_n N_A_27_368#_c_399_n 0.00696193f $X=5.01 $Y=2.305
+ $X2=0 $Y2=0
cc_191 N_A_183_48#_M1017_g N_A_27_368#_c_400_n 0.00108206f $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_192 N_A_183_48#_c_164_n N_A_27_368#_c_400_n 0.01491f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_193 N_A_183_48#_M1001_g N_A_27_368#_c_401_n 9.14596e-19 $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_194 N_A_183_48#_M1000_d N_A_27_368#_c_392_n 0.00137918f $X=4.875 $Y=1.84
+ $X2=0 $Y2=0
cc_195 N_A_183_48#_M1017_g N_A_27_368#_c_392_n 2.82703e-19 $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_196 N_A_183_48#_c_164_n N_A_27_368#_c_392_n 0.0259125f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_197 N_A_183_48#_c_168_n N_A_27_368#_c_392_n 0.0455162f $X=5.125 $Y=1.005
+ $X2=0 $Y2=0
cc_198 N_A_183_48#_c_194_p N_A_27_368#_c_392_n 0.0280472f $X=5.795 $Y=2.225
+ $X2=0 $Y2=0
cc_199 N_A_183_48#_c_170_n N_A_27_368#_c_392_n 0.0427206f $X=5.96 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_183_48#_c_183_n N_A_27_368#_c_392_n 0.011205f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_201 N_A_183_48#_c_172_n N_A_27_368#_c_392_n 2.27533e-19 $X=4.3 $Y=1.465 $X2=0
+ $Y2=0
cc_202 N_A_183_48#_c_194_p N_VPWR_M1004_s 0.00421004f $X=5.795 $Y=2.225 $X2=0
+ $Y2=0
cc_203 N_A_183_48#_M1001_g N_VPWR_c_538_n 0.0124551f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_183_48#_M1002_g N_VPWR_c_538_n 0.00149196f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_205 N_A_183_48#_M1001_g N_VPWR_c_539_n 0.00149196f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_206 N_A_183_48#_M1002_g N_VPWR_c_539_n 0.0124969f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_183_48#_M1003_g N_VPWR_c_539_n 0.0124969f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_183_48#_M1008_g N_VPWR_c_539_n 0.00149196f $X=2.355 $Y=2.4 $X2=0
+ $Y2=0
cc_209 N_A_183_48#_M1003_g N_VPWR_c_540_n 0.00149196f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_210 N_A_183_48#_M1008_g N_VPWR_c_540_n 0.0124969f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A_183_48#_M1011_g N_VPWR_c_540_n 0.0124969f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_183_48#_M1012_g N_VPWR_c_540_n 0.00149196f $X=3.255 $Y=2.4 $X2=0
+ $Y2=0
cc_213 N_A_183_48#_M1011_g N_VPWR_c_541_n 0.00149196f $X=2.805 $Y=2.4 $X2=0
+ $Y2=0
cc_214 N_A_183_48#_M1012_g N_VPWR_c_541_n 0.0124969f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_183_48#_M1016_g N_VPWR_c_541_n 0.0134899f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A_183_48#_M1017_g N_VPWR_c_541_n 0.00231482f $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_217 N_A_183_48#_M1016_g N_VPWR_c_542_n 0.00231482f $X=3.705 $Y=2.4 $X2=0
+ $Y2=0
cc_218 N_A_183_48#_M1017_g N_VPWR_c_542_n 0.0134481f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_183_48#_c_183_n N_VPWR_c_542_n 0.0157994f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_220 N_A_183_48#_c_194_p N_VPWR_c_543_n 0.0189268f $X=5.795 $Y=2.225 $X2=0
+ $Y2=0
cc_221 N_A_183_48#_c_182_n N_VPWR_c_543_n 0.0195323f $X=5.96 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_183_48#_c_183_n N_VPWR_c_543_n 0.0195517f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_223 N_A_183_48#_M1011_g N_VPWR_c_544_n 0.00460063f $X=2.805 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_183_48#_M1012_g N_VPWR_c_544_n 0.00460063f $X=3.255 $Y=2.4 $X2=0
+ $Y2=0
cc_225 N_A_183_48#_M1001_g N_VPWR_c_547_n 0.00460063f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_226 N_A_183_48#_M1002_g N_VPWR_c_547_n 0.00460063f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_227 N_A_183_48#_M1003_g N_VPWR_c_548_n 0.00460063f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_228 N_A_183_48#_M1008_g N_VPWR_c_548_n 0.00460063f $X=2.355 $Y=2.4 $X2=0
+ $Y2=0
cc_229 N_A_183_48#_M1016_g N_VPWR_c_549_n 0.00460063f $X=3.705 $Y=2.4 $X2=0
+ $Y2=0
cc_230 N_A_183_48#_M1017_g N_VPWR_c_549_n 0.00460063f $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_231 N_A_183_48#_c_183_n N_VPWR_c_550_n 0.0144623f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_232 N_A_183_48#_c_182_n N_VPWR_c_551_n 0.0124046f $X=5.96 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_183_48#_M1001_g N_VPWR_c_537_n 0.00908554f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_234 N_A_183_48#_M1002_g N_VPWR_c_537_n 0.00908554f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_235 N_A_183_48#_M1003_g N_VPWR_c_537_n 0.00908554f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_236 N_A_183_48#_M1008_g N_VPWR_c_537_n 0.00908554f $X=2.355 $Y=2.4 $X2=0
+ $Y2=0
cc_237 N_A_183_48#_M1011_g N_VPWR_c_537_n 0.00908554f $X=2.805 $Y=2.4 $X2=0
+ $Y2=0
cc_238 N_A_183_48#_M1012_g N_VPWR_c_537_n 0.00908554f $X=3.255 $Y=2.4 $X2=0
+ $Y2=0
cc_239 N_A_183_48#_M1016_g N_VPWR_c_537_n 0.00909733f $X=3.705 $Y=2.4 $X2=0
+ $Y2=0
cc_240 N_A_183_48#_M1017_g N_VPWR_c_537_n 0.00909733f $X=4.285 $Y=2.4 $X2=0
+ $Y2=0
cc_241 N_A_183_48#_c_182_n N_VPWR_c_537_n 0.0102675f $X=5.96 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A_183_48#_c_183_n N_VPWR_c_537_n 0.0118344f $X=5.01 $Y=2.305 $X2=0
+ $Y2=0
cc_243 N_A_183_48#_M1009_g N_Y_c_636_n 0.0154892f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_183_48#_M1013_g N_Y_c_636_n 0.0152302f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_183_48#_c_164_n N_Y_c_636_n 0.0299541f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_246 N_A_183_48#_c_172_n N_Y_c_636_n 0.00448425f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_247 N_A_183_48#_M1002_g N_Y_c_645_n 0.0135168f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_183_48#_M1003_g N_Y_c_645_n 0.0130762f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_183_48#_M1008_g N_Y_c_645_n 0.0130762f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_183_48#_M1011_g N_Y_c_645_n 0.0130762f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A_183_48#_M1012_g N_Y_c_645_n 0.0130762f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A_183_48#_M1016_g N_Y_c_645_n 0.0168814f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A_183_48#_M1017_g N_Y_c_645_n 0.00809268f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_183_48#_c_164_n N_Y_c_645_n 0.19572f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_255 N_A_183_48#_c_172_n N_Y_c_645_n 0.0160605f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_256 N_A_183_48#_M1013_g N_Y_c_637_n 3.99083e-19 $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_183_48#_M1014_g N_Y_c_637_n 3.99083e-19 $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_183_48#_M1014_g N_Y_c_638_n 0.0152302f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_183_48#_M1018_g N_Y_c_638_n 0.01369f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_183_48#_c_164_n N_Y_c_638_n 0.0507189f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_261 N_A_183_48#_c_172_n N_Y_c_638_n 0.00416134f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_262 N_A_183_48#_M1014_g N_Y_c_639_n 5.56882e-19 $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_183_48#_M1018_g N_Y_c_639_n 0.0082419f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_183_48#_M1020_g N_Y_c_639_n 0.00746139f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_183_48#_M1021_g N_Y_c_639_n 3.52398e-19 $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_183_48#_M1020_g N_Y_c_640_n 0.0115433f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_183_48#_M1021_g N_Y_c_640_n 0.0151263f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_183_48#_M1022_g N_Y_c_640_n 0.00323816f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_183_48#_c_164_n N_Y_c_640_n 0.0769774f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_270 N_A_183_48#_c_168_n N_Y_c_640_n 0.00764154f $X=5.125 $Y=1.005 $X2=0 $Y2=0
cc_271 N_A_183_48#_c_172_n N_Y_c_640_n 0.00832347f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_272 N_A_183_48#_M1021_g N_Y_c_641_n 0.00324276f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_183_48#_M1022_g N_Y_c_641_n 0.00946516f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_183_48#_c_168_n N_Y_c_641_n 0.00335458f $X=5.125 $Y=1.005 $X2=0 $Y2=0
cc_275 N_A_183_48#_M1001_g N_Y_c_680_n 0.00408251f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A_183_48#_M1002_g N_Y_c_680_n 0.00139868f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A_183_48#_c_164_n N_Y_c_642_n 0.0160251f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_278 N_A_183_48#_c_172_n N_Y_c_642_n 0.00244789f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_279 N_A_183_48#_M1018_g N_Y_c_643_n 0.00115621f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_183_48#_M1020_g N_Y_c_643_n 0.00257766f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_183_48#_M1021_g N_Y_c_643_n 2.50354e-19 $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_183_48#_c_164_n N_Y_c_643_n 0.0276081f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_283 N_A_183_48#_c_172_n N_Y_c_643_n 0.00256622f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_284 N_A_183_48#_M1006_g Y 0.00600697f $X=0.99 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_183_48#_M1009_g Y 0.00829833f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_183_48#_M1013_g Y 5.00623e-19 $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_183_48#_M1006_g Y 0.00377972f $X=0.99 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_183_48#_M1009_g Y 8.07377e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A_183_48#_M1006_g Y 0.00361253f $X=0.99 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_183_48#_M1001_g Y 0.00391162f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A_183_48#_M1009_g Y 0.00538497f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A_183_48#_M1002_g Y 0.00510363f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A_183_48#_M1003_g Y 7.94469e-19 $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A_183_48#_M1013_g Y 7.96256e-19 $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A_183_48#_c_164_n Y 0.0177955f $X=4.65 $Y=1.465 $X2=0 $Y2=0
cc_296 N_A_183_48#_c_172_n Y 0.0239221f $X=4.3 $Y=1.465 $X2=0 $Y2=0
cc_297 N_A_183_48#_c_168_n N_VGND_M1022_s 0.00318074f $X=5.125 $Y=1.005 $X2=0
+ $Y2=0
cc_298 N_A_183_48#_c_167_n N_VGND_M1015_s 0.00253871f $X=5.795 $Y=1.005 $X2=0
+ $Y2=0
cc_299 N_A_183_48#_M1006_g N_VGND_c_739_n 0.00233397f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_183_48#_M1009_g N_VGND_c_740_n 0.00365073f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_301 N_A_183_48#_M1013_g N_VGND_c_740_n 0.00799341f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_302 N_A_183_48#_M1014_g N_VGND_c_740_n 4.27258e-19 $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_183_48#_M1013_g N_VGND_c_741_n 4.27258e-19 $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_183_48#_M1014_g N_VGND_c_741_n 0.00792092f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_183_48#_M1018_g N_VGND_c_741_n 0.00365073f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_183_48#_M1020_g N_VGND_c_742_n 0.00406778f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_183_48#_M1021_g N_VGND_c_742_n 0.00979254f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A_183_48#_M1022_g N_VGND_c_742_n 4.87331e-19 $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A_183_48#_M1022_g N_VGND_c_743_n 0.00365073f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_183_48#_c_164_n N_VGND_c_743_n 0.00785549f $X=4.65 $Y=1.465 $X2=0
+ $Y2=0
cc_311 N_A_183_48#_c_166_n N_VGND_c_743_n 0.0142435f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_312 N_A_183_48#_c_168_n N_VGND_c_743_n 0.00333948f $X=5.125 $Y=1.005 $X2=0
+ $Y2=0
cc_313 N_A_183_48#_c_166_n N_VGND_c_744_n 0.0142435f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_314 N_A_183_48#_c_167_n N_VGND_c_744_n 0.0215485f $X=5.795 $Y=1.005 $X2=0
+ $Y2=0
cc_315 N_A_183_48#_c_169_n N_VGND_c_744_n 0.0142986f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_316 N_A_183_48#_M1006_g N_VGND_c_746_n 0.00456932f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_317 N_A_183_48#_M1009_g N_VGND_c_746_n 0.00434272f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_318 N_A_183_48#_M1013_g N_VGND_c_747_n 0.00383152f $X=1.94 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_183_48#_M1014_g N_VGND_c_747_n 0.00383152f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_320 N_A_183_48#_M1018_g N_VGND_c_748_n 0.00434272f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_321 N_A_183_48#_M1020_g N_VGND_c_748_n 0.00434272f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_183_48#_M1021_g N_VGND_c_749_n 0.00383152f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A_183_48#_M1022_g N_VGND_c_749_n 0.00434272f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A_183_48#_c_166_n N_VGND_c_750_n 0.00889602f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_325 N_A_183_48#_c_169_n N_VGND_c_751_n 0.0145639f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_326 N_A_183_48#_M1006_g N_VGND_c_752_n 0.00889942f $X=0.99 $Y=0.74 $X2=0
+ $Y2=0
cc_327 N_A_183_48#_M1009_g N_VGND_c_752_n 0.00820916f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_328 N_A_183_48#_M1013_g N_VGND_c_752_n 0.0075754f $X=1.94 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A_183_48#_M1014_g N_VGND_c_752_n 0.0075754f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A_183_48#_M1018_g N_VGND_c_752_n 0.00820718f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_331 N_A_183_48#_M1020_g N_VGND_c_752_n 0.00820718f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_183_48#_M1021_g N_VGND_c_752_n 0.00758198f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A_183_48#_M1022_g N_VGND_c_752_n 0.0082143f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A_183_48#_c_166_n N_VGND_c_752_n 0.00743504f $X=5.02 $Y=0.515 $X2=0
+ $Y2=0
cc_335 N_A_183_48#_c_169_n N_VGND_c_752_n 0.0119984f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_336 N_A_27_368#_c_410_n N_VPWR_M1007_d 0.00326865f $X=0.72 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_337 N_A_27_368#_c_391_n N_VPWR_M1007_d 0.00532598f $X=0.805 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_338 N_A_27_368#_c_480_p N_VPWR_M1007_d 0.00151608f $X=0.805 $Y=2.325
+ $X2=-0.19 $Y2=-0.245
cc_339 N_A_27_368#_c_451_n N_VPWR_M1002_d 0.00324075f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_340 N_A_27_368#_c_451_n N_VPWR_M1008_d 0.00324075f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_341 N_A_27_368#_c_451_n N_VPWR_M1012_d 0.00324075f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_342 N_A_27_368#_c_451_n N_VPWR_M1017_d 0.00335161f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_c_462_n N_VPWR_M1017_d 0.00337014f $X=4.48 $Y=2.24 $X2=0
+ $Y2=0
cc_344 N_A_27_368#_c_399_n N_VPWR_M1017_d 0.00144475f $X=4.99 $Y=1.885 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_400_n N_VPWR_M1017_d 5.9723e-19 $X=4.565 $Y=1.885 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_392_n N_VPWR_M1004_s 0.00283799f $X=5.475 $Y=1.485 $X2=0
+ $Y2=0
cc_347 N_A_27_368#_c_397_n N_VPWR_c_538_n 0.0157994f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_348 N_A_27_368#_c_410_n N_VPWR_c_538_n 0.00549591f $X=0.72 $Y=2.325 $X2=0
+ $Y2=0
cc_349 N_A_27_368#_c_451_n N_VPWR_c_538_n 0.00216696f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_350 N_A_27_368#_c_480_p N_VPWR_c_538_n 0.0123972f $X=0.805 $Y=2.325 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_451_n N_VPWR_c_539_n 0.0170259f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_451_n N_VPWR_c_540_n 0.0170259f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_451_n N_VPWR_c_541_n 0.0170259f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_393_n N_VPWR_c_542_n 0.00205601f $X=4.785 $Y=1.74 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_451_n N_VPWR_c_542_n 0.0140626f $X=4.395 $Y=2.325 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_399_n N_VPWR_c_542_n 0.0022621f $X=4.99 $Y=1.885 $X2=0
+ $Y2=0
cc_357 N_A_27_368#_M1004_g N_VPWR_c_543_n 0.00258607f $X=5.235 $Y=2.4 $X2=0
+ $Y2=0
cc_358 N_A_27_368#_M1005_g N_VPWR_c_543_n 0.0144643f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A_27_368#_c_397_n N_VPWR_c_546_n 0.014549f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_360 N_A_27_368#_c_393_n N_VPWR_c_550_n 0.005209f $X=4.785 $Y=1.74 $X2=0 $Y2=0
cc_361 N_A_27_368#_M1004_g N_VPWR_c_550_n 0.005209f $X=5.235 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A_27_368#_M1005_g N_VPWR_c_551_n 0.00460063f $X=5.735 $Y=2.4 $X2=0
+ $Y2=0
cc_363 N_A_27_368#_c_393_n N_VPWR_c_537_n 0.0098216f $X=4.785 $Y=1.74 $X2=0
+ $Y2=0
cc_364 N_A_27_368#_M1004_g N_VPWR_c_537_n 0.00982082f $X=5.235 $Y=2.4 $X2=0
+ $Y2=0
cc_365 N_A_27_368#_M1005_g N_VPWR_c_537_n 0.00912296f $X=5.735 $Y=2.4 $X2=0
+ $Y2=0
cc_366 N_A_27_368#_c_397_n N_VPWR_c_537_n 0.0119743f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_367 N_A_27_368#_c_451_n N_Y_M1001_s 0.00753096f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_368 N_A_27_368#_c_451_n N_Y_M1003_s 0.0075347f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_369 N_A_27_368#_c_451_n N_Y_M1011_s 0.0075347f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_370 N_A_27_368#_c_451_n N_Y_M1016_s 0.0141367f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_371 N_A_27_368#_c_451_n N_Y_c_645_n 0.156272f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_372 N_A_27_368#_c_400_n N_Y_c_645_n 0.00889661f $X=4.565 $Y=1.885 $X2=0 $Y2=0
cc_373 N_A_27_368#_M1010_g N_Y_c_641_n 6.39165e-19 $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A_27_368#_c_391_n N_Y_c_680_n 0.012847f $X=0.805 $Y=2.24 $X2=0 $Y2=0
cc_375 N_A_27_368#_c_451_n N_Y_c_680_n 0.017094f $X=4.395 $Y=2.325 $X2=0 $Y2=0
cc_376 N_A_27_368#_c_389_n Y 0.00596854f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_377 N_A_27_368#_c_389_n Y 0.00417827f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_378 N_A_27_368#_c_391_n Y 0.0464398f $X=0.805 $Y=2.24 $X2=0 $Y2=0
cc_379 N_A_27_368#_c_389_n N_VGND_M1023_d 0.00286042f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_368#_c_388_n N_VGND_c_739_n 0.0182902f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_381 N_A_27_368#_c_389_n N_VGND_c_739_n 0.02058f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_382 N_A_27_368#_M1010_g N_VGND_c_743_n 0.00796521f $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_383 N_A_27_368#_M1015_g N_VGND_c_743_n 4.26797e-19 $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_27_368#_M1010_g N_VGND_c_744_n 4.26797e-19 $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A_27_368#_M1015_g N_VGND_c_744_n 0.00796521f $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_386 N_A_27_368#_M1019_g N_VGND_c_744_n 0.00503266f $X=5.745 $Y=0.74 $X2=0
+ $Y2=0
cc_387 N_A_27_368#_c_388_n N_VGND_c_745_n 0.011066f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_388 N_A_27_368#_M1010_g N_VGND_c_750_n 0.00383152f $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_389 N_A_27_368#_M1015_g N_VGND_c_750_n 0.00383152f $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_390 N_A_27_368#_M1019_g N_VGND_c_751_n 0.00434272f $X=5.745 $Y=0.74 $X2=0
+ $Y2=0
cc_391 N_A_27_368#_M1010_g N_VGND_c_752_n 0.00757689f $X=4.8 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A_27_368#_M1015_g N_VGND_c_752_n 0.00757689f $X=5.245 $Y=0.74 $X2=0
+ $Y2=0
cc_393 N_A_27_368#_M1019_g N_VGND_c_752_n 0.00824376f $X=5.745 $Y=0.74 $X2=0
+ $Y2=0
cc_394 N_A_27_368#_c_388_n N_VGND_c_752_n 0.00915947f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_395 N_VPWR_M1002_d N_Y_c_645_n 0.00168622f $X=1.545 $Y=1.84 $X2=0 $Y2=0
cc_396 N_VPWR_M1008_d N_Y_c_645_n 0.00168622f $X=2.445 $Y=1.84 $X2=0 $Y2=0
cc_397 N_VPWR_M1012_d N_Y_c_645_n 0.00168622f $X=3.345 $Y=1.84 $X2=0 $Y2=0
cc_398 N_Y_c_636_n N_VGND_M1009_s 0.00253871f $X=2.06 $Y=1.005 $X2=0 $Y2=0
cc_399 N_Y_c_638_n N_VGND_M1014_s 0.00253871f $X=2.92 $Y=1.005 $X2=0 $Y2=0
cc_400 N_Y_c_640_n N_VGND_M1020_s 0.00250873f $X=3.92 $Y=1.045 $X2=0 $Y2=0
cc_401 Y N_VGND_c_739_n 0.0191764f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_402 N_Y_c_636_n N_VGND_c_740_n 0.0215485f $X=2.06 $Y=1.005 $X2=0 $Y2=0
cc_403 N_Y_c_637_n N_VGND_c_740_n 0.0142351f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_404 Y N_VGND_c_740_n 0.0142986f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_405 N_Y_c_637_n N_VGND_c_741_n 0.0142351f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_406 N_Y_c_638_n N_VGND_c_741_n 0.0215485f $X=2.92 $Y=1.005 $X2=0 $Y2=0
cc_407 N_Y_c_639_n N_VGND_c_741_n 0.0142986f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_408 N_Y_c_639_n N_VGND_c_742_n 0.0173003f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_409 N_Y_c_640_n N_VGND_c_742_n 0.0209867f $X=3.92 $Y=1.045 $X2=0 $Y2=0
cc_410 N_Y_c_641_n N_VGND_c_742_n 0.0173003f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_411 N_Y_c_641_n N_VGND_c_743_n 0.0142986f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_412 Y N_VGND_c_746_n 0.014552f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_413 N_Y_c_637_n N_VGND_c_747_n 0.00838873f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_414 N_Y_c_639_n N_VGND_c_748_n 0.0144922f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_415 N_Y_c_641_n N_VGND_c_749_n 0.0145639f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_416 N_Y_c_637_n N_VGND_c_752_n 0.00694347f $X=2.155 $Y=0.515 $X2=0 $Y2=0
cc_417 N_Y_c_639_n N_VGND_c_752_n 0.0118826f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_418 N_Y_c_641_n N_VGND_c_752_n 0.0119984f $X=4.085 $Y=0.515 $X2=0 $Y2=0
cc_419 Y N_VGND_c_752_n 0.0119791f $X=1.115 $Y=0.47 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1555_410# a_1335_112# a_1934_392# VPB pshort w=1e+06u l=180000u
+  ad=5.45e+11p pd=5.09e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR a_1555_410# a_2516_368# VPB pshort w=1e+06u l=180000u
+  ad=3.0275e+12p pd=2.579e+07u as=2.65e+11p ps=2.53e+06u
M1002 a_1507_508# a_27_74# a_1335_112# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.688e+11p ps=2.4e+06u
M1003 a_1240_125# a_473_405# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.90125e+11p pd=1.88e+06u as=2.06398e+12p ps=1.857e+07u
M1004 a_1640_138# a_200_74# a_1335_112# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=6.1e+11p ps=3.85e+06u
M1005 VGND SET_B a_867_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.4925e+11p ps=3.47e+06u
M1006 a_933_424# a_601_119# a_473_405# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=4.452e+11p ps=4.42e+06u
M1007 a_867_125# a_975_322# a_473_405# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.54e+11p ps=1.66e+06u
M1008 Q a_2516_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1009 a_1832_74# a_1335_112# a_1555_410# VNB nlowvt w=740000u l=150000u
+  ad=4.979e+11p pd=4.43e+06u as=2.368e+11p ps=2.12e+06u
M1010 a_1832_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_311_119# a_27_74# a_601_119# VPB pshort w=420000u l=180000u
+  ad=3.3075e+11p pd=3.39e+06u as=1.386e+11p ps=1.5e+06u
M1012 VPWR RESET_B a_975_322# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1013 VPWR a_1555_410# a_1507_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_473_405# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q_N a_1555_410# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1016 Q a_2516_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1017 VGND D a_311_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=5.0085e+11p ps=3.93e+06u
M1018 a_539_503# a_473_405# VPWR VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1019 VPWR a_1555_410# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_2516_368# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1934_392# a_975_322# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1335_112# a_200_74# a_1315_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.016e+11p ps=2.16e+06u
M1023 VGND a_1555_410# a_1640_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1555_410# a_975_322# a_1832_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR D a_311_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND RESET_B a_975_322# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1027 VPWR SET_B a_1555_410# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_311_119# a_200_74# a_601_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1029 VPWR a_975_322# a_933_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_601_119# a_200_74# a_539_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_1555_410# a_2516_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1032 VGND a_2516_368# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR CLK_N a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1034 a_200_74# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1035 VGND a_1555_410# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1036 a_529_119# a_473_405# VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1037 VGND CLK_N a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1038 a_200_74# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1039 a_1335_112# a_27_74# a_1240_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_473_405# a_601_119# a_867_125# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1315_424# a_473_405# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_601_119# a_27_74# a_529_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Q_N a_1555_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__ebufn_1.spice
* Created: Fri Aug 28 17:31:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__ebufn_1.pex.spice"
.subckt sky130_fd_sc_ms__ebufn_1  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_TE_B_M1007_g N_A_27_404#_M1007_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.0825 AS=0.15675 PD=0.85 PS=1.67 NRD=2.172 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_A_229_74#_M1002_d N_A_M1002_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.0825 PD=1.63 PS=0.85 NRD=0 NRS=2.172 M=1 R=3.66667 SA=75000.7
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 A_569_74# N_A_27_404#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_Z_M1006_d N_A_229_74#_M1006_g A_569_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_TE_B_M1000_g N_A_27_404#_M1000_s VPB PSHORT L=0.18
+ W=0.84 AD=0.21525 AS=0.2352 PD=1.49 PS=2.24 NRD=47.1815 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1003 N_A_229_74#_M1003_d N_A_M1003_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=0.84
+ AD=0.2436 AS=0.21525 PD=2.26 PS=1.49 NRD=0 NRS=47.1815 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1001 A_569_368# N_TE_B_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1344 AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1004 N_Z_M1004_d N_A_229_74#_M1004_g A_569_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1344 PD=2.8 PS=1.36 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__ebufn_1.pxi.spice"
*
.ends
*
*

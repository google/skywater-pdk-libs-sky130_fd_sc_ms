* File: sky130_fd_sc_ms__sdlclkp_1.spice
* Created: Wed Sep  2 12:32:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdlclkp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdlclkp_1  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1013 N_A_114_112#_M1013_d N_SCE_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.15675 PD=0.83 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1012 N_VGND_M1012_d N_GATE_M1012_g N_A_114_112#_M1013_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.161184 AS=0.077 PD=1.20233 PS=0.83 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_A_318_74#_M1003_d N_A_288_48#_M1003_g N_VGND_M1012_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_566_74#_M1017_d N_A_288_48#_M1017_g N_A_114_112#_M1017_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.10467 AS=0.29425 PD=1.02629 PS=2.17 NRD=0 NRS=54.54 M=1
+ R=3.66667 SA=75000.5 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1015 A_667_80# N_A_318_74#_M1015_g N_A_566_74#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0799299 PD=0.63 PS=0.783711 NRD=14.28 NRS=22.848 M=1
+ R=2.8 SA=75001 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_709_54#_M1016_g A_667_80# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109562 AS=0.0441 PD=0.919655 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1010 N_A_709_54#_M1010_d N_A_566_74#_M1010_g N_VGND_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.193038 PD=2.04 PS=1.62034 NRD=0 NRS=40.536 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_CLK_M1005_g N_A_288_48#_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.2072 PD=1.14217 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1006 A_1166_94# N_CLK_M1006_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.108058 PD=0.85 PS=0.987826 NRD=9.372 NRS=8.436 M=1 R=4.26667
+ SA=75000.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_1238_94#_M1007_d N_A_709_54#_M1007_g A_1166_94# VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75001 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 N_GCLK_M1019_d N_A_1238_94#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.2664 PD=2.04 PS=2.2 NRD=0 NRS=12.156 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 A_119_424# N_SCE_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.0882 AS=0.2352 PD=1.05 PS=2.24 NRD=11.7215 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1000 N_A_114_112#_M1000_d N_GATE_M1000_g A_119_424# VPB PSHORT L=0.18 W=0.84
+ AD=0.2352 AS=0.0882 PD=2.24 PS=1.05 NRD=0 NRS=11.7215 M=1 R=4.66667 SA=90000.6
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1021 N_A_318_74#_M1021_d N_A_288_48#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.3907 PD=2.24 PS=2.99 NRD=0 NRS=96.1754 M=1 R=4.66667
+ SA=90000.3 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1011 N_A_566_74#_M1011_d N_A_318_74#_M1011_g N_A_114_112#_M1011_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.194717 AS=0.2352 PD=1.78667 PS=2.24 NRD=0 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1002 A_725_492# N_A_288_48#_M1002_g N_A_566_74#_M1011_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0973583 PD=0.63 PS=0.893333 NRD=23.443 NRS=37.5088 M=1
+ R=2.33333 SA=90000.5 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1018 N_VPWR_M1018_d N_A_709_54#_M1018_g A_725_492# VPB PSHORT L=0.18 W=0.42
+ AD=0.0849545 AS=0.0441 PD=0.788182 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333
+ SA=90000.9 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1001 N_A_709_54#_M1001_d N_A_566_74#_M1001_g N_VPWR_M1018_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.226545 PD=2.8 PS=2.10182 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1020_d N_CLK_M1020_g N_A_288_48#_M1020_s VPB PSHORT L=0.18 W=0.84
+ AD=0.269225 AS=0.2352 PD=1.645 PS=2.24 NRD=62.252 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1004 N_A_1238_94#_M1004_d N_CLK_M1004_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.269225 PD=1.11 PS=1.645 NRD=0 NRS=62.252 M=1 R=4.66667
+ SA=90000.9 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1009 N_VPWR_M1009_d N_A_709_54#_M1009_g N_A_1238_94#_M1004_d VPB PSHORT L=0.18
+ W=0.84 AD=0.147 AS=0.1134 PD=1.23857 PS=1.11 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90001.3 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1014 N_GCLK_M1014_d N_A_1238_94#_M1014_g N_VPWR_M1009_d VPB PSHORT L=0.18
+ W=1.12 AD=0.4088 AS=0.196 PD=2.97 PS=1.65143 NRD=14.0658 NRS=0 M=1 R=6.22222
+ SA=90001.4 SB=90000.3 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.0772 P=20
*
.include "sky130_fd_sc_ms__sdlclkp_1.pxi.spice"
*
.ends
*
*

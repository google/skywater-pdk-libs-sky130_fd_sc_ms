* File: sky130_fd_sc_ms__dlygate4sd2_1.pxi.spice
* Created: Fri Aug 28 17:30:39 2020
* 
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A N_A_M1003_g N_A_M1001_g A A N_A_c_67_n
+ PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_28_74# N_A_28_74#_M1003_s
+ N_A_28_74#_M1001_s N_A_28_74#_M1007_g N_A_28_74#_M1002_g N_A_28_74#_c_98_n
+ N_A_28_74#_c_104_n N_A_28_74#_c_105_n N_A_28_74#_c_106_n N_A_28_74#_c_99_n
+ N_A_28_74#_c_100_n N_A_28_74#_c_101_n N_A_28_74#_c_102_n
+ PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_28_74#
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_288_74# N_A_288_74#_M1002_d
+ N_A_288_74#_M1007_d N_A_288_74#_M1006_g N_A_288_74#_M1004_g
+ N_A_288_74#_c_159_n N_A_288_74#_c_160_n N_A_288_74#_c_161_n
+ N_A_288_74#_c_162_n N_A_288_74#_c_166_n N_A_288_74#_c_163_n
+ N_A_288_74#_c_164_n PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_288_74#
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_405_138# N_A_405_138#_M1004_s
+ N_A_405_138#_M1006_s N_A_405_138#_M1000_g N_A_405_138#_M1005_g
+ N_A_405_138#_c_216_n N_A_405_138#_c_222_n N_A_405_138#_c_217_n
+ N_A_405_138#_c_218_n N_A_405_138#_c_219_n N_A_405_138#_c_224_n
+ N_A_405_138#_c_220_n PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_405_138#
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%VPWR N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n VPWR
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_274_n N_VPWR_c_282_n
+ PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%VPWR
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%X N_X_M1005_d N_X_M1000_d X X X X X X X
+ N_X_c_310_n X X N_X_c_314_n PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%X
x_PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%VGND N_VGND_M1003_d N_VGND_M1004_d
+ N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n N_VGND_c_334_n VGND
+ N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n
+ PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%VGND
cc_1 VNB N_A_M1003_g 0.0470899f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_M1001_g 0.00890285f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_3 VNB A 0.0265853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_67_n 0.0358668f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_M1002_g 0.0395543f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_6 VNB N_A_28_74#_c_98_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.52
cc_7 VNB N_A_28_74#_c_99_n 0.0206633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_28_74#_c_100_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_74#_c_101_n 0.00140945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_74#_c_102_n 0.0616725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_288_74#_M1006_g 0.00282418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_288_74#_M1004_g 0.0313942f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_13 VNB N_A_288_74#_c_159_n 0.014798f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.52
cc_14 VNB N_A_288_74#_c_160_n 0.0208388f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_15 VNB N_A_288_74#_c_161_n 0.0219379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_288_74#_c_162_n 0.0631267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_288_74#_c_163_n 0.0020102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_288_74#_c_164_n 0.00336402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_405_138#_M1000_g 0.00188052f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_A_405_138#_M1005_g 0.0275176f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_21 VNB N_A_405_138#_c_216_n 0.00382325f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_22 VNB N_A_405_138#_c_217_n 0.00323188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_405_138#_c_218_n 2.9305e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_405_138#_c_219_n 0.00926587f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.665
cc_25 VNB N_A_405_138#_c_220_n 0.0339153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_274_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0286532f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_X_c_310_n 0.029118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.0145768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_331_n 0.00984339f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_VGND_c_332_n 0.0187989f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_32 VNB N_VGND_c_333_n 0.0567418f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_33 VNB N_VGND_c_334_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.52
cc_34 VNB N_VGND_c_335_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_336_n 0.0205885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_337_n 0.253672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_338_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_M1001_g 0.0678332f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_39 VPB A 0.0146632f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_40 VPB N_A_28_74#_M1007_g 0.0329704f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_41 VPB N_A_28_74#_c_104_n 0.0222074f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_42 VPB N_A_28_74#_c_105_n 0.00180999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_28_74#_c_106_n 0.0109668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_28_74#_c_101_n 0.0017204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_28_74#_c_102_n 0.02099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_288_74#_M1006_g 0.0367294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_288_74#_c_166_n 0.0125296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_288_74#_c_163_n 0.0217942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_405_138#_M1000_g 0.02702f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_50 VPB N_A_405_138#_c_222_n 0.00303941f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.52
cc_51 VPB N_A_405_138#_c_218_n 0.00160201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_405_138#_c_224_n 0.00800757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_275_n 0.0156916f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_54 VPB N_VPWR_c_276_n 0.0110042f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_55 VPB N_VPWR_c_277_n 0.0596029f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_56 VPB N_VPWR_c_278_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_279_n 0.0190092f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.665
cc_58 VPB N_VPWR_c_280_n 0.0200102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_274_n 0.109013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_282_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB X 0.00819691f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_62 VPB X 0.0507672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_X_c_314_n 0.014629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_A_28_74#_M1007_g 0.0136756f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_A_28_74#_M1002_g 0.00808739f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_A_28_74#_c_98_n 0.0127782f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_A_28_74#_c_104_n 0.00641825f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_68 N_A_M1001_g N_A_28_74#_c_105_n 0.0199916f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_69 A N_A_28_74#_c_105_n 0.0262324f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_c_67_n N_A_28_74#_c_105_n 6.49888e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_71 A N_A_28_74#_c_106_n 0.0280303f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_A_28_74#_c_99_n 0.0120856f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_73 A N_A_28_74#_c_99_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_c_67_n N_A_28_74#_c_99_n 0.00146766f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_A_28_74#_c_100_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_76 A N_A_28_74#_c_100_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_A_28_74#_c_101_n 0.0025292f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_A_28_74#_c_101_n 0.0039553f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_79 A N_A_28_74#_c_101_n 0.0413255f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_c_67_n N_A_28_74#_c_101_n 0.00110303f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_81 N_A_M1003_g N_A_28_74#_c_102_n 0.0021171f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_82 N_A_M1001_g N_A_28_74#_c_102_n 0.00881686f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_83 A N_A_28_74#_c_102_n 0.00372609f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A_c_67_n N_A_28_74#_c_102_n 0.0208886f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_85 N_A_M1001_g N_VPWR_c_275_n 0.0130994f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_VPWR_c_279_n 0.00500714f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_VPWR_c_274_n 0.00551156f $X=0.495 $Y=2.545 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VGND_c_331_n 0.00293875f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VGND_c_335_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_90 N_A_M1003_g N_VGND_c_337_n 0.00456437f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_91 N_A_28_74#_M1002_g N_A_288_74#_c_159_n 0.00938998f $X=1.35 $Y=0.58 $X2=0
+ $Y2=0
cc_92 N_A_28_74#_M1002_g N_A_288_74#_c_160_n 0.00883481f $X=1.35 $Y=0.58 $X2=0
+ $Y2=0
cc_93 N_A_28_74#_c_99_n N_A_288_74#_c_160_n 0.0164122f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_94 N_A_28_74#_c_101_n N_A_288_74#_c_160_n 0.0277104f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_95 N_A_28_74#_c_102_n N_A_288_74#_c_160_n 0.00609936f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_96 N_A_28_74#_c_102_n N_A_288_74#_c_162_n 0.00416224f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_97 N_A_28_74#_M1007_g N_A_288_74#_c_166_n 0.00903431f $X=1.32 $Y=2.46 $X2=0
+ $Y2=0
cc_98 N_A_28_74#_c_101_n N_A_288_74#_c_163_n 0.0295243f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_99 N_A_28_74#_c_102_n N_A_288_74#_c_163_n 0.0182179f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_100 N_A_28_74#_c_101_n N_A_288_74#_c_164_n 0.0193935f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_101 N_A_28_74#_c_102_n N_A_288_74#_c_164_n 0.00352926f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_102 N_A_28_74#_c_105_n N_VPWR_M1001_d 0.0234374f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_28_74#_c_101_n N_VPWR_M1001_d 0.00114873f $X=1.14 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_28_74#_M1007_g N_VPWR_c_275_n 0.0146599f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_105 N_A_28_74#_c_105_n N_VPWR_c_275_n 0.0237211f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_106 N_A_28_74#_M1007_g N_VPWR_c_277_n 0.00742301f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_107 N_A_28_74#_c_104_n N_VPWR_c_279_n 0.00578326f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_108 N_A_28_74#_M1007_g N_VPWR_c_274_n 0.0142438f $X=1.32 $Y=2.46 $X2=0 $Y2=0
cc_109 N_A_28_74#_c_104_n N_VPWR_c_274_n 0.00940928f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_110 N_A_28_74#_M1002_g N_VGND_c_331_n 0.00497305f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_111 N_A_28_74#_c_98_n N_VGND_c_331_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_112 N_A_28_74#_c_99_n N_VGND_c_331_n 0.0255952f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_113 N_A_28_74#_M1002_g N_VGND_c_333_n 0.00524396f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_114 N_A_28_74#_c_98_n N_VGND_c_335_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_115 N_A_28_74#_M1002_g N_VGND_c_337_n 0.0087053f $X=1.35 $Y=0.58 $X2=0 $Y2=0
cc_116 N_A_28_74#_c_98_n N_VGND_c_337_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_117 N_A_28_74#_c_99_n N_VGND_c_337_n 0.0213669f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_118 N_A_288_74#_M1006_g N_A_405_138#_M1000_g 0.0312009f $X=2.66 $Y=2.34 $X2=0
+ $Y2=0
cc_119 N_A_288_74#_M1004_g N_A_405_138#_M1005_g 0.0198704f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_120 N_A_288_74#_M1004_g N_A_405_138#_c_216_n 0.0189992f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_121 N_A_288_74#_c_161_n N_A_405_138#_c_216_n 0.028346f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_122 N_A_288_74#_c_162_n N_A_405_138#_c_216_n 0.00668708f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_123 N_A_288_74#_M1006_g N_A_405_138#_c_222_n 0.0247695f $X=2.66 $Y=2.34 $X2=0
+ $Y2=0
cc_124 N_A_288_74#_c_161_n N_A_405_138#_c_222_n 0.0234159f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_125 N_A_288_74#_c_162_n N_A_405_138#_c_222_n 0.0042133f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_126 N_A_288_74#_M1004_g N_A_405_138#_c_217_n 0.00219888f $X=2.695 $Y=0.9
+ $X2=0 $Y2=0
cc_127 N_A_288_74#_c_161_n N_A_405_138#_c_217_n 0.0193923f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_128 N_A_288_74#_c_162_n N_A_405_138#_c_217_n 0.00410963f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_129 N_A_288_74#_M1006_g N_A_405_138#_c_218_n 0.00478601f $X=2.66 $Y=2.34
+ $X2=0 $Y2=0
cc_130 N_A_288_74#_M1004_g N_A_405_138#_c_219_n 0.0100145f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_131 N_A_288_74#_c_160_n N_A_405_138#_c_219_n 0.0301033f $X=1.597 $Y=1.38
+ $X2=0 $Y2=0
cc_132 N_A_288_74#_c_161_n N_A_405_138#_c_219_n 0.0290383f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_133 N_A_288_74#_c_162_n N_A_405_138#_c_219_n 0.00695677f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_134 N_A_288_74#_M1006_g N_A_405_138#_c_224_n 0.00802029f $X=2.66 $Y=2.34
+ $X2=0 $Y2=0
cc_135 N_A_288_74#_c_161_n N_A_405_138#_c_224_n 0.0237961f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_136 N_A_288_74#_c_162_n N_A_405_138#_c_224_n 0.0062457f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_137 N_A_288_74#_c_163_n N_A_405_138#_c_224_n 0.0219754f $X=1.567 $Y=2.395
+ $X2=0 $Y2=0
cc_138 N_A_288_74#_M1004_g N_A_405_138#_c_220_n 2.62551e-19 $X=2.695 $Y=0.9
+ $X2=0 $Y2=0
cc_139 N_A_288_74#_c_161_n N_A_405_138#_c_220_n 2.17534e-19 $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_140 N_A_288_74#_c_162_n N_A_405_138#_c_220_n 0.0213845f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_141 N_A_288_74#_c_166_n N_VPWR_c_275_n 0.0108408f $X=1.58 $Y=2.56 $X2=0 $Y2=0
cc_142 N_A_288_74#_M1006_g N_VPWR_c_276_n 0.00765051f $X=2.66 $Y=2.34 $X2=0
+ $Y2=0
cc_143 N_A_288_74#_M1006_g N_VPWR_c_277_n 0.00823417f $X=2.66 $Y=2.34 $X2=0
+ $Y2=0
cc_144 N_A_288_74#_c_166_n N_VPWR_c_277_n 0.00561205f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_145 N_A_288_74#_M1006_g N_VPWR_c_274_n 0.00847299f $X=2.66 $Y=2.34 $X2=0
+ $Y2=0
cc_146 N_A_288_74#_c_166_n N_VPWR_c_274_n 0.00918412f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_147 N_A_288_74#_c_159_n N_VGND_c_331_n 0.0111538f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_148 N_A_288_74#_M1004_g N_VGND_c_332_n 0.00468436f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_149 N_A_288_74#_M1004_g N_VGND_c_333_n 0.00459186f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_150 N_A_288_74#_c_159_n N_VGND_c_333_n 0.0163531f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_151 N_A_288_74#_M1004_g N_VGND_c_337_n 0.00542201f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_152 N_A_288_74#_c_159_n N_VGND_c_337_n 0.011395f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_153 N_A_405_138#_c_222_n N_VPWR_M1006_d 0.00246069f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_154 N_A_405_138#_M1000_g N_VPWR_c_276_n 0.0170272f $X=3.215 $Y=2.4 $X2=0
+ $Y2=0
cc_155 N_A_405_138#_c_222_n N_VPWR_c_276_n 0.022154f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_156 N_A_405_138#_c_220_n N_VPWR_c_276_n 3.71022e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_157 N_A_405_138#_M1000_g N_VPWR_c_280_n 0.00460063f $X=3.215 $Y=2.4 $X2=0
+ $Y2=0
cc_158 N_A_405_138#_M1000_g N_VPWR_c_274_n 0.00912647f $X=3.215 $Y=2.4 $X2=0
+ $Y2=0
cc_159 N_A_405_138#_M1000_g X 0.00311617f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_405_138#_M1005_g X 0.00260428f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_405_138#_c_217_n X 0.0327059f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_162 N_A_405_138#_c_218_n X 0.00709928f $X=3.032 $Y=1.825 $X2=0 $Y2=0
cc_163 N_A_405_138#_c_220_n X 0.00794767f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_164 N_A_405_138#_M1005_g N_X_c_310_n 0.00143568f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_405_138#_c_217_n X 0.0037592f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_166 N_A_405_138#_M1000_g N_X_c_314_n 0.00418785f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A_405_138#_c_222_n N_X_c_314_n 0.00776663f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_168 N_A_405_138#_c_218_n N_X_c_314_n 7.53343e-19 $X=3.032 $Y=1.825 $X2=0
+ $Y2=0
cc_169 N_A_405_138#_c_216_n N_VGND_M1004_d 7.12223e-19 $X=2.91 $Y=1.125 $X2=0
+ $Y2=0
cc_170 N_A_405_138#_c_217_n N_VGND_M1004_d 0.0018038f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_171 N_A_405_138#_M1005_g N_VGND_c_332_n 0.0156117f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_405_138#_c_216_n N_VGND_c_332_n 0.00549591f $X=2.91 $Y=1.125 $X2=0
+ $Y2=0
cc_173 N_A_405_138#_c_217_n N_VGND_c_332_n 0.016728f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_174 N_A_405_138#_c_220_n N_VGND_c_332_n 4.7706e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_175 N_A_405_138#_c_219_n N_VGND_c_333_n 0.00580898f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_176 N_A_405_138#_M1005_g N_VGND_c_336_n 0.00383152f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_405_138#_M1005_g N_VGND_c_337_n 0.00761589f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_405_138#_c_219_n N_VGND_c_337_n 0.0101265f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_276_n X 0.0378465f $X=2.99 $Y=2.27 $X2=0 $Y2=0
cc_180 N_VPWR_c_280_n X 0.0270407f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_274_n X 0.0159412f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_182 N_X_c_310_n N_VGND_c_332_n 0.019927f $X=3.42 $Y=0.52 $X2=0 $Y2=0
cc_183 N_X_c_310_n N_VGND_c_336_n 0.0180659f $X=3.42 $Y=0.52 $X2=0 $Y2=0
cc_184 N_X_c_310_n N_VGND_c_337_n 0.0152075f $X=3.42 $Y=0.52 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__nor4b_2.pxi.spice
* Created: Wed Sep  2 12:17:03 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4B_2%D_N N_D_N_M1001_g N_D_N_M1000_g D_N N_D_N_c_97_n
+ PM_SKY130_FD_SC_MS__NOR4B_2%D_N
x_PM_SKY130_FD_SC_MS__NOR4B_2%A_27_392# N_A_27_392#_M1000_s N_A_27_392#_M1001_s
+ N_A_27_392#_c_129_n N_A_27_392#_M1006_g N_A_27_392#_M1012_g
+ N_A_27_392#_c_131_n N_A_27_392#_M1009_g N_A_27_392#_M1014_g
+ N_A_27_392#_c_133_n N_A_27_392#_c_134_n N_A_27_392#_c_135_n
+ N_A_27_392#_c_136_n N_A_27_392#_c_137_n N_A_27_392#_c_138_n
+ PM_SKY130_FD_SC_MS__NOR4B_2%A_27_392#
x_PM_SKY130_FD_SC_MS__NOR4B_2%C N_C_M1010_g N_C_M1015_g N_C_M1017_g N_C_M1016_g
+ C C N_C_c_217_n PM_SKY130_FD_SC_MS__NOR4B_2%C
x_PM_SKY130_FD_SC_MS__NOR4B_2%B N_B_M1002_g N_B_c_272_n N_B_c_273_n N_B_M1005_g
+ N_B_M1011_g N_B_c_275_n N_B_M1007_g B B N_B_c_277_n
+ PM_SKY130_FD_SC_MS__NOR4B_2%B
x_PM_SKY130_FD_SC_MS__NOR4B_2%A N_A_M1003_g N_A_M1004_g N_A_M1008_g N_A_M1013_g
+ A A A N_A_c_334_n PM_SKY130_FD_SC_MS__NOR4B_2%A
x_PM_SKY130_FD_SC_MS__NOR4B_2%VPWR N_VPWR_M1001_d N_VPWR_M1003_s N_VPWR_c_375_n
+ N_VPWR_c_376_n VPWR N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n
+ N_VPWR_c_374_n N_VPWR_c_381_n N_VPWR_c_382_n PM_SKY130_FD_SC_MS__NOR4B_2%VPWR
x_PM_SKY130_FD_SC_MS__NOR4B_2%A_229_368# N_A_229_368#_M1012_s
+ N_A_229_368#_M1014_s N_A_229_368#_M1016_s N_A_229_368#_c_431_n
+ N_A_229_368#_c_432_n N_A_229_368#_c_433_n N_A_229_368#_c_445_n
+ N_A_229_368#_c_446_n N_A_229_368#_c_434_n N_A_229_368#_c_435_n
+ PM_SKY130_FD_SC_MS__NOR4B_2%A_229_368#
x_PM_SKY130_FD_SC_MS__NOR4B_2%Y N_Y_M1006_s N_Y_M1010_s N_Y_M1002_d N_Y_M1004_s
+ N_Y_M1012_d N_Y_c_473_n N_Y_c_486_n N_Y_c_489_n N_Y_c_482_n N_Y_c_540_n
+ N_Y_c_495_n N_Y_c_474_n N_Y_c_475_n N_Y_c_476_n N_Y_c_477_n N_Y_c_478_n
+ N_Y_c_479_n Y Y N_Y_c_481_n PM_SKY130_FD_SC_MS__NOR4B_2%Y
x_PM_SKY130_FD_SC_MS__NOR4B_2%A_501_368# N_A_501_368#_M1015_d
+ N_A_501_368#_M1005_d N_A_501_368#_c_573_n N_A_501_368#_c_580_n
+ N_A_501_368#_c_574_n PM_SKY130_FD_SC_MS__NOR4B_2%A_501_368#
x_PM_SKY130_FD_SC_MS__NOR4B_2%A_701_368# N_A_701_368#_M1005_s
+ N_A_701_368#_M1007_s N_A_701_368#_M1008_d N_A_701_368#_c_600_n
+ N_A_701_368#_c_601_n N_A_701_368#_c_609_n N_A_701_368#_c_602_n
+ N_A_701_368#_c_613_n N_A_701_368#_c_603_n N_A_701_368#_c_604_n
+ N_A_701_368#_c_619_n PM_SKY130_FD_SC_MS__NOR4B_2%A_701_368#
x_PM_SKY130_FD_SC_MS__NOR4B_2%VGND N_VGND_M1000_d N_VGND_M1009_d N_VGND_M1017_d
+ N_VGND_M1011_s N_VGND_M1013_d N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n VGND N_VGND_c_642_n
+ N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n
+ N_VGND_c_648_n PM_SKY130_FD_SC_MS__NOR4B_2%VGND
cc_1 VNB N_D_N_M1000_g 0.0450381f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_2 VNB D_N 0.00165062f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_N_c_97_n 0.0264696f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.635
cc_4 VNB N_A_27_392#_c_129_n 0.0182324f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_5 VNB N_A_27_392#_M1012_g 0.00699685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_392#_c_131_n 0.0183095f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.635
cc_7 VNB N_A_27_392#_M1014_g 0.00530441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_392#_c_133_n 0.0390192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_392#_c_134_n 0.0189495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_392#_c_135_n 0.0120801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_136_n 0.0081778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_392#_c_137_n 0.014353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_392#_c_138_n 0.0684587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C_M1010_g 0.0257645f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_15 VNB N_C_M1017_g 0.0249557f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.635
cc_16 VNB C 0.00340543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_c_217_n 0.0338177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_M1002_g 0.026244f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_19 VNB N_B_c_272_n 0.0157093f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.47
cc_20 VNB N_B_c_273_n 0.00974905f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_21 VNB N_B_M1011_g 0.0318253f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.635
cc_22 VNB N_B_c_275_n 0.0215786f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.635
cc_23 VNB B 0.00579351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_277_n 0.0101463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_M1004_g 0.0305489f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_26 VNB N_A_M1013_g 0.0326296f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.635
cc_27 VNB A 0.0218856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_c_334_n 0.0413018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_374_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_473_n 0.00291634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_474_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_475_n 0.00517051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_476_n 0.00687852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_477_n 0.00263681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_478_n 0.0117419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_479_n 0.0028038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB Y 0.00299091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_481_n 0.00245684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_636_n 0.00894653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_637_n 0.00830481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_638_n 0.0120411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_639_n 0.0421046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_640_n 0.0223929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_641_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_642_n 0.0184653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_643_n 0.0187266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_644_n 0.041024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_645_n 0.0185686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_646_n 0.0169675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_647_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_648_n 0.313921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_D_N_M1001_g 0.029246f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_53 VPB D_N 0.00249009f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_54 VPB N_D_N_c_97_n 0.021776f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_55 VPB N_A_27_392#_M1012_g 0.0259483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_392#_M1014_g 0.0212092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_392#_c_134_n 0.0556684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_C_M1015_g 0.0204354f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_59 VPB N_C_M1016_g 0.0244601f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_60 VPB C 0.0054379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_C_c_217_n 0.00477627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B_c_272_n 0.0103731f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.47
cc_63 VPB N_B_c_273_n 0.00491078f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_64 VPB N_B_M1005_g 0.0243443f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_65 VPB N_B_c_275_n 0.00389087f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_66 VPB N_B_M1007_g 0.0214081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB B 0.0137607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_B_c_277_n 3.82064e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_M1003_g 0.0203638f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_70 VPB N_A_M1008_g 0.0269566f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.635
cc_71 VPB A 0.0143682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_c_334_n 0.00594104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_375_n 0.0154162f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_74 VPB N_VPWR_c_376_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_75 VPB N_VPWR_c_377_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_378_n 0.0953538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_379_n 0.018982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_374_n 0.0875314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_381_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_382_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_229_368#_c_431_n 0.0128248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_229_368#_c_432_n 0.00439642f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_83 VPB N_A_229_368#_c_433_n 0.00413156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_229_368#_c_434_n 0.00225721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_229_368#_c_435_n 0.00256399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_Y_c_482_n 0.00312122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_Y_c_475_n 0.00185475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_501_368#_c_573_n 0.0187146f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_89 VPB N_A_501_368#_c_574_n 0.00195131f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_90 VPB N_A_701_368#_c_600_n 0.00196801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_701_368#_c_601_n 0.00650336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_701_368#_c_602_n 0.00179576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_701_368#_c_603_n 0.00723723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_701_368#_c_604_n 0.0339608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 N_D_N_M1000_g N_A_27_392#_c_129_n 0.0211411f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_96 D_N N_A_27_392#_M1012_g 0.0013121f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_97 N_D_N_c_97_n N_A_27_392#_M1012_g 0.00608659f $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_98 N_D_N_M1000_g N_A_27_392#_c_133_n 0.0131116f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_99 N_D_N_M1000_g N_A_27_392#_c_134_n 0.00592896f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_100 D_N N_A_27_392#_c_134_n 0.025547f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_101 N_D_N_c_97_n N_A_27_392#_c_134_n 0.0162755f $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_102 N_D_N_M1000_g N_A_27_392#_c_135_n 0.00449144f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_103 D_N N_A_27_392#_c_135_n 0.00361618f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_104 N_D_N_c_97_n N_A_27_392#_c_135_n 0.00600323f $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_105 N_D_N_M1000_g N_A_27_392#_c_136_n 9.66795e-19 $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_106 D_N N_A_27_392#_c_136_n 0.00477495f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_107 N_D_N_c_97_n N_A_27_392#_c_136_n 3.08012e-19 $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_108 N_D_N_M1000_g N_A_27_392#_c_137_n 0.0117536f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_109 D_N N_A_27_392#_c_137_n 0.0209481f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_110 N_D_N_c_97_n N_A_27_392#_c_137_n 0.00112087f $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_111 N_D_N_M1000_g N_A_27_392#_c_138_n 0.00670227f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_112 N_D_N_c_97_n N_A_27_392#_c_138_n 0.00440373f $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_113 N_D_N_M1001_g N_VPWR_c_375_n 0.020999f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_114 D_N N_VPWR_c_375_n 0.0220408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_115 N_D_N_c_97_n N_VPWR_c_375_n 0.00194594f $X=0.7 $Y=1.635 $X2=0 $Y2=0
cc_116 N_D_N_M1001_g N_VPWR_c_377_n 0.00460063f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_117 N_D_N_M1001_g N_VPWR_c_374_n 0.00912296f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_118 N_D_N_M1001_g N_A_229_368#_c_431_n 0.00377212f $X=0.505 $Y=2.46 $X2=0
+ $Y2=0
cc_119 N_D_N_M1001_g N_A_229_368#_c_433_n 6.08298e-19 $X=0.505 $Y=2.46 $X2=0
+ $Y2=0
cc_120 N_D_N_M1000_g N_VGND_c_636_n 0.00695483f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_121 N_D_N_M1000_g N_VGND_c_640_n 0.00434272f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_122 N_D_N_M1000_g N_VGND_c_648_n 0.0082535f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_123 N_A_27_392#_c_131_n N_C_M1010_g 0.0180513f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_124 N_A_27_392#_c_136_n N_C_M1010_g 8.7155e-19 $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A_27_392#_c_138_n N_C_M1010_g 0.0120031f $X=1.965 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_27_392#_M1014_g N_C_M1015_g 0.0340084f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_27_392#_M1012_g C 0.00103715f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_27_392#_M1014_g C 0.0070915f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_27_392#_c_136_n C 0.0115655f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_130 N_A_27_392#_c_138_n C 0.00624784f $X=1.965 $Y=1.385 $X2=0 $Y2=0
cc_131 N_A_27_392#_M1014_g N_C_c_217_n 0.0120031f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_27_392#_M1012_g N_VPWR_c_375_n 0.00263089f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_133 N_A_27_392#_c_134_n N_VPWR_c_375_n 0.0339508f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_134 N_A_27_392#_c_137_n N_VPWR_c_375_n 9.48018e-19 $X=1.105 $Y=1.34 $X2=0
+ $Y2=0
cc_135 N_A_27_392#_c_134_n N_VPWR_c_377_n 0.011066f $X=0.28 $Y=2.105 $X2=0 $Y2=0
cc_136 N_A_27_392#_M1012_g N_VPWR_c_378_n 0.00333896f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_137 N_A_27_392#_M1014_g N_VPWR_c_378_n 0.00333896f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_138 N_A_27_392#_M1012_g N_VPWR_c_374_n 0.00427818f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_139 N_A_27_392#_M1014_g N_VPWR_c_374_n 0.00422796f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_140 N_A_27_392#_c_134_n N_VPWR_c_374_n 0.00915947f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_141 N_A_27_392#_M1012_g N_A_229_368#_c_431_n 0.0160206f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_27_392#_M1014_g N_A_229_368#_c_431_n 6.27116e-19 $X=1.965 $Y=2.4
+ $X2=0 $Y2=0
cc_143 N_A_27_392#_c_136_n N_A_229_368#_c_431_n 0.0197823f $X=1.61 $Y=1.385
+ $X2=0 $Y2=0
cc_144 N_A_27_392#_c_138_n N_A_229_368#_c_431_n 0.00743382f $X=1.965 $Y=1.385
+ $X2=0 $Y2=0
cc_145 N_A_27_392#_M1012_g N_A_229_368#_c_432_n 0.0115958f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_146 N_A_27_392#_M1014_g N_A_229_368#_c_432_n 0.0132535f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_147 N_A_27_392#_M1012_g N_A_229_368#_c_433_n 0.00291744f $X=1.515 $Y=2.4
+ $X2=0 $Y2=0
cc_148 N_A_27_392#_M1014_g N_A_229_368#_c_445_n 0.00244698f $X=1.965 $Y=2.4
+ $X2=0 $Y2=0
cc_149 N_A_27_392#_M1012_g N_A_229_368#_c_446_n 5.20536e-19 $X=1.515 $Y=2.4
+ $X2=0 $Y2=0
cc_150 N_A_27_392#_M1014_g N_A_229_368#_c_446_n 0.00649085f $X=1.965 $Y=2.4
+ $X2=0 $Y2=0
cc_151 N_A_27_392#_c_129_n N_Y_c_473_n 0.0054187f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_152 N_A_27_392#_c_131_n N_Y_c_473_n 0.00252693f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_153 N_A_27_392#_c_131_n N_Y_c_486_n 0.0130155f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A_27_392#_c_136_n N_Y_c_486_n 0.0128666f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_155 N_A_27_392#_c_138_n N_Y_c_486_n 0.00950085f $X=1.965 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A_27_392#_c_129_n N_Y_c_489_n 0.00209321f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A_27_392#_c_136_n N_Y_c_489_n 0.0256756f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_158 N_A_27_392#_c_138_n N_Y_c_489_n 0.00105099f $X=1.965 $Y=1.385 $X2=0 $Y2=0
cc_159 N_A_27_392#_M1014_g N_Y_c_482_n 4.63009e-19 $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_27_392#_c_136_n N_Y_c_482_n 0.00728815f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_161 N_A_27_392#_c_138_n N_Y_c_482_n 0.00244512f $X=1.965 $Y=1.385 $X2=0 $Y2=0
cc_162 N_A_27_392#_M1014_g N_Y_c_495_n 0.0193484f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_27_392#_c_131_n N_Y_c_474_n 9.57264e-19 $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_27_392#_c_131_n N_Y_c_477_n 7.73117e-19 $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_27_392#_c_136_n N_Y_c_477_n 0.00131831f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_166 N_A_27_392#_c_129_n N_VGND_c_636_n 0.0054296f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_167 N_A_27_392#_c_133_n N_VGND_c_636_n 0.0249119f $X=0.415 $Y=0.515 $X2=0
+ $Y2=0
cc_168 N_A_27_392#_c_137_n N_VGND_c_636_n 0.0261348f $X=1.105 $Y=1.34 $X2=0
+ $Y2=0
cc_169 N_A_27_392#_c_133_n N_VGND_c_640_n 0.0205877f $X=0.415 $Y=0.515 $X2=0
+ $Y2=0
cc_170 N_A_27_392#_c_129_n N_VGND_c_642_n 0.00433834f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A_27_392#_c_131_n N_VGND_c_642_n 0.00384553f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A_27_392#_c_129_n N_VGND_c_646_n 3.64777e-19 $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_173 N_A_27_392#_c_131_n N_VGND_c_646_n 0.0117177f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A_27_392#_c_129_n N_VGND_c_648_n 0.00821665f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_27_392#_c_131_n N_VGND_c_648_n 0.00374134f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_176 N_A_27_392#_c_133_n N_VGND_c_648_n 0.0169844f $X=0.415 $Y=0.515 $X2=0
+ $Y2=0
cc_177 N_C_M1017_g N_B_M1002_g 0.0210645f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_178 N_C_c_217_n N_B_c_273_n 0.0116958f $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_179 N_C_M1016_g B 5.62894e-19 $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_180 N_C_c_217_n B 3.33564e-19 $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_181 N_C_M1015_g N_VPWR_c_378_n 0.00518311f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_182 N_C_M1016_g N_VPWR_c_378_n 0.00335119f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_183 N_C_M1015_g N_VPWR_c_374_n 0.00982392f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_184 N_C_M1016_g N_VPWR_c_374_n 0.00426909f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_185 N_C_M1015_g N_A_229_368#_c_432_n 0.00101073f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_186 N_C_M1015_g N_A_229_368#_c_434_n 0.0140196f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_187 N_C_M1016_g N_A_229_368#_c_434_n 0.0115668f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_188 N_C_M1010_g N_Y_c_486_n 0.0104376f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_189 C N_Y_c_486_n 0.0154053f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_190 N_C_M1015_g N_Y_c_495_n 0.0115861f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_191 N_C_M1016_g N_Y_c_495_n 0.0166954f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_192 C N_Y_c_495_n 0.0477277f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_193 N_C_c_217_n N_Y_c_495_n 4.88651e-19 $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_194 N_C_M1010_g N_Y_c_474_n 0.00798642f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_195 N_C_M1017_g N_Y_c_474_n 0.00570416f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_196 N_C_M1015_g N_Y_c_475_n 8.87005e-19 $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_197 N_C_M1017_g N_Y_c_475_n 0.00443118f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_198 N_C_M1016_g N_Y_c_475_n 0.00874477f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_199 C N_Y_c_475_n 0.0331353f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_200 N_C_c_217_n N_Y_c_475_n 0.00877689f $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_201 N_C_M1010_g N_Y_c_477_n 0.00661837f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_202 N_C_M1017_g N_Y_c_477_n 0.0217824f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_203 C N_Y_c_477_n 0.0269015f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_204 N_C_c_217_n N_Y_c_477_n 0.00373527f $X=2.865 $Y=1.515 $X2=0 $Y2=0
cc_205 N_C_M1017_g Y 6.11074e-19 $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_206 N_C_M1016_g N_A_501_368#_c_573_n 0.0116469f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_207 N_C_M1015_g N_A_501_368#_c_574_n 0.00714033f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_208 N_C_M1016_g N_A_501_368#_c_574_n 0.0117081f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_209 N_C_M1016_g N_A_701_368#_c_600_n 9.47506e-19 $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_210 N_C_M1016_g N_A_701_368#_c_601_n 0.00459472f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_211 N_C_M1017_g N_VGND_c_637_n 0.00470005f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_212 N_C_M1010_g N_VGND_c_643_n 0.00434272f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_213 N_C_M1017_g N_VGND_c_643_n 0.00434272f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_214 N_C_M1010_g N_VGND_c_646_n 0.00400351f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_215 N_C_M1010_g N_VGND_c_648_n 0.00436462f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_216 N_C_M1017_g N_VGND_c_648_n 0.00821165f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B_M1007_g N_A_M1003_g 0.0131302f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_218 N_B_c_275_n A 0.00270252f $X=4.235 $Y=1.605 $X2=0 $Y2=0
cc_219 B A 0.0298391f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B_c_277_n A 5.80008e-19 $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_221 N_B_c_275_n N_A_c_334_n 0.00827036f $X=4.235 $Y=1.605 $X2=0 $Y2=0
cc_222 B N_A_c_334_n 7.03106e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_223 N_B_c_277_n N_A_c_334_n 0.0018393f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_224 N_B_M1007_g N_VPWR_c_376_n 5.80674e-19 $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_225 N_B_M1005_g N_VPWR_c_378_n 0.00333896f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_226 N_B_M1007_g N_VPWR_c_378_n 0.00517089f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_227 N_B_M1005_g N_VPWR_c_374_n 0.00427818f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_228 N_B_M1007_g N_VPWR_c_374_n 0.00978686f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B_M1002_g N_Y_c_475_n 0.00358729f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B_c_273_n N_Y_c_475_n 0.00111277f $X=3.445 $Y=1.515 $X2=0 $Y2=0
cc_231 N_B_M1005_g N_Y_c_475_n 0.00262327f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_232 B N_Y_c_475_n 0.0306983f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B_M1002_g N_Y_c_476_n 0.0131887f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_234 B N_Y_c_476_n 0.0105458f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_B_M1002_g N_Y_c_477_n 4.69564e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B_M1011_g N_Y_c_478_n 0.0169209f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B_c_275_n N_Y_c_478_n 0.00857091f $X=4.235 $Y=1.605 $X2=0 $Y2=0
cc_238 B N_Y_c_478_n 0.0329461f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B_M1002_g Y 0.00856724f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B_M1011_g Y 0.00366931f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B_M1002_g N_Y_c_481_n 0.00116959f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B_c_272_n N_Y_c_481_n 0.00442617f $X=3.785 $Y=1.515 $X2=0 $Y2=0
cc_243 B N_Y_c_481_n 0.028285f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_244 N_B_M1005_g N_A_501_368#_c_573_n 0.0156999f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B_M1007_g N_A_501_368#_c_573_n 0.0041969f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B_M1005_g N_A_501_368#_c_580_n 0.0134366f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B_M1007_g N_A_501_368#_c_580_n 0.0076969f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_248 N_B_c_272_n N_A_701_368#_c_600_n 0.00151925f $X=3.785 $Y=1.515 $X2=0
+ $Y2=0
cc_249 B N_A_701_368#_c_600_n 0.0218203f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B_M1005_g N_A_701_368#_c_609_n 0.0142562f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_251 N_B_c_275_n N_A_701_368#_c_609_n 4.9731e-19 $X=4.235 $Y=1.605 $X2=0 $Y2=0
cc_252 N_B_M1007_g N_A_701_368#_c_609_n 0.01917f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_253 B N_A_701_368#_c_609_n 0.0308985f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_254 N_B_M1002_g N_VGND_c_637_n 0.0027066f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B_M1002_g N_VGND_c_644_n 0.00504858f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B_M1011_g N_VGND_c_644_n 0.0159343f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B_M1002_g N_VGND_c_648_n 0.00891136f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B_M1011_g N_VGND_c_648_n 0.00758371f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_M1003_g N_VPWR_c_376_n 0.0128677f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_M1008_g N_VPWR_c_376_n 0.0151943f $X=5.235 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A_M1003_g N_VPWR_c_378_n 0.00460063f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_M1008_g N_VPWR_c_379_n 0.00490827f $X=5.235 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A_M1003_g N_VPWR_c_374_n 0.00908665f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_M1008_g N_VPWR_c_374_n 0.00972577f $X=5.235 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A_M1004_g N_Y_c_478_n 0.0147517f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_M1013_g N_Y_c_478_n 0.00185032f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_267 A N_Y_c_478_n 0.0570125f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_268 N_A_c_334_n N_Y_c_478_n 0.00463218f $X=5.25 $Y=1.515 $X2=0 $Y2=0
cc_269 N_A_M1004_g N_Y_c_479_n 0.0153465f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_M1013_g N_Y_c_479_n 4.79228e-19 $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_M1003_g N_A_501_368#_c_573_n 2.99783e-19 $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A_M1003_g N_A_701_368#_c_613_n 0.0142639f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_M1008_g N_A_701_368#_c_613_n 0.0146245f $X=5.235 $Y=2.4 $X2=0 $Y2=0
cc_274 A N_A_701_368#_c_613_n 0.0486946f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_275 N_A_c_334_n N_A_701_368#_c_613_n 5.45297e-19 $X=5.25 $Y=1.515 $X2=0 $Y2=0
cc_276 A N_A_701_368#_c_603_n 0.0218206f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_277 N_A_M1008_g N_A_701_368#_c_604_n 4.72217e-19 $X=5.235 $Y=2.4 $X2=0 $Y2=0
cc_278 A N_A_701_368#_c_619_n 0.0143992f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A_M1004_g N_VGND_c_639_n 5.65034e-19 $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_M1013_g N_VGND_c_639_n 0.0137863f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_281 A N_VGND_c_639_n 0.023911f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_282 N_A_M1004_g N_VGND_c_644_n 0.00509578f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A_M1004_g N_VGND_c_645_n 0.00434272f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A_M1013_g N_VGND_c_645_n 0.00429299f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_M1004_g N_VGND_c_648_n 0.00825583f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_M1013_g N_VGND_c_648_n 0.00848048f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_287 N_VPWR_c_375_n N_A_229_368#_c_431_n 0.0630024f $X=0.73 $Y=2.135 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_378_n N_A_229_368#_c_432_n 0.0536089f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_374_n N_A_229_368#_c_432_n 0.0296408f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_375_n N_A_229_368#_c_433_n 0.0121616f $X=0.73 $Y=2.135 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_378_n N_A_229_368#_c_433_n 0.0235512f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_374_n N_A_229_368#_c_433_n 0.0126924f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_376_n N_A_501_368#_c_573_n 0.00279016f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_294 N_VPWR_c_378_n N_A_501_368#_c_573_n 0.0953389f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_374_n N_A_501_368#_c_573_n 0.053672f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_c_378_n N_A_501_368#_c_574_n 0.0225872f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_374_n N_A_501_368#_c_574_n 0.0123496f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_376_n N_A_701_368#_c_602_n 0.0233699f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_299 N_VPWR_c_378_n N_A_701_368#_c_602_n 0.00749631f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_374_n N_A_701_368#_c_602_n 0.0062048f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_301 N_VPWR_M1003_s N_A_701_368#_c_613_n 0.00333697f $X=4.865 $Y=1.84 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_376_n N_A_701_368#_c_613_n 0.0170777f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_303 N_VPWR_c_376_n N_A_701_368#_c_604_n 0.0225174f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_304 N_VPWR_c_379_n N_A_701_368#_c_604_n 0.011066f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_305 N_VPWR_c_374_n N_A_701_368#_c_604_n 0.00915947f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_A_229_368#_c_432_n N_Y_M1012_d 0.00165831f $X=2.025 $Y=2.99 $X2=0 $Y2=0
cc_307 N_A_229_368#_c_431_n N_Y_c_482_n 0.0105642f $X=1.29 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_229_368#_c_432_n N_Y_c_540_n 0.0118736f $X=2.025 $Y=2.99 $X2=0 $Y2=0
cc_309 N_A_229_368#_M1014_s N_Y_c_495_n 0.00332066f $X=2.055 $Y=1.84 $X2=0 $Y2=0
cc_310 N_A_229_368#_M1016_s N_Y_c_495_n 0.00343534f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_311 N_A_229_368#_c_445_n N_Y_c_495_n 0.0149351f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_312 N_A_229_368#_c_434_n N_Y_c_495_n 0.043084f $X=3.005 $Y=2.375 $X2=0 $Y2=0
cc_313 N_A_229_368#_M1016_s N_Y_c_475_n 0.00196027f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_314 N_A_229_368#_c_434_n N_A_501_368#_M1015_d 0.00324075f $X=3.005 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_315 N_A_229_368#_M1016_s N_A_501_368#_c_573_n 0.00266942f $X=2.955 $Y=1.84
+ $X2=0 $Y2=0
cc_316 N_A_229_368#_c_434_n N_A_501_368#_c_573_n 0.00464895f $X=3.005 $Y=2.375
+ $X2=0 $Y2=0
cc_317 N_A_229_368#_c_435_n N_A_501_368#_c_573_n 0.0178873f $X=3.13 $Y=2.46
+ $X2=0 $Y2=0
cc_318 N_A_229_368#_c_432_n N_A_501_368#_c_574_n 0.0103602f $X=2.025 $Y=2.99
+ $X2=0 $Y2=0
cc_319 N_A_229_368#_c_434_n N_A_501_368#_c_574_n 0.0164517f $X=3.005 $Y=2.375
+ $X2=0 $Y2=0
cc_320 N_A_229_368#_c_434_n N_A_701_368#_c_601_n 0.011925f $X=3.005 $Y=2.375
+ $X2=0 $Y2=0
cc_321 N_A_229_368#_c_435_n N_A_701_368#_c_601_n 0.0177445f $X=3.13 $Y=2.46
+ $X2=0 $Y2=0
cc_322 N_Y_c_495_n N_A_501_368#_M1015_d 0.0031478f $X=2.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_323 N_Y_c_495_n N_A_701_368#_c_600_n 0.0086044f $X=2.925 $Y=2.035 $X2=0 $Y2=0
cc_324 N_Y_c_486_n N_VGND_M1009_d 0.0123139f $X=2.44 $Y=0.875 $X2=0 $Y2=0
cc_325 N_Y_c_476_n N_VGND_M1017_d 0.0016136f $X=3.44 $Y=1.095 $X2=0 $Y2=0
cc_326 N_Y_c_477_n N_VGND_M1017_d 0.00169317f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_327 N_Y_c_478_n N_VGND_M1011_s 0.00926984f $X=4.815 $Y=1.095 $X2=0 $Y2=0
cc_328 N_Y_c_473_n N_VGND_c_636_n 0.0188454f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_329 N_Y_c_474_n N_VGND_c_637_n 0.0172628f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_330 N_Y_c_476_n N_VGND_c_637_n 0.0115978f $X=3.44 $Y=1.095 $X2=0 $Y2=0
cc_331 N_Y_c_477_n N_VGND_c_637_n 0.0128931f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_332 Y N_VGND_c_637_n 0.0191764f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_333 N_Y_c_478_n N_VGND_c_639_n 0.00540983f $X=4.815 $Y=1.095 $X2=0 $Y2=0
cc_334 N_Y_c_479_n N_VGND_c_639_n 0.0255552f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_335 N_Y_c_473_n N_VGND_c_642_n 0.0157475f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_336 N_Y_c_474_n N_VGND_c_643_n 0.0144922f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_337 N_Y_c_478_n N_VGND_c_644_n 0.0424937f $X=4.815 $Y=1.095 $X2=0 $Y2=0
cc_338 N_Y_c_479_n N_VGND_c_644_n 0.0173963f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_339 Y N_VGND_c_644_n 0.0339549f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_340 N_Y_c_479_n N_VGND_c_645_n 0.0145639f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_341 N_Y_c_473_n N_VGND_c_646_n 0.0124832f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_342 N_Y_c_486_n N_VGND_c_646_n 0.0323939f $X=2.44 $Y=0.875 $X2=0 $Y2=0
cc_343 N_Y_c_474_n N_VGND_c_646_n 0.0102273f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_344 N_Y_c_473_n N_VGND_c_648_n 0.0121127f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_345 N_Y_c_486_n N_VGND_c_648_n 0.0123705f $X=2.44 $Y=0.875 $X2=0 $Y2=0
cc_346 N_Y_c_474_n N_VGND_c_648_n 0.0118826f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_347 N_Y_c_479_n N_VGND_c_648_n 0.0119984f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_348 Y N_VGND_c_648_n 0.0120948f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_349 N_A_501_368#_c_573_n N_A_701_368#_M1005_s 0.00266942f $X=3.935 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_350 N_A_501_368#_c_573_n N_A_701_368#_c_601_n 0.0184743f $X=3.935 $Y=2.99
+ $X2=0 $Y2=0
cc_351 N_A_501_368#_M1005_d N_A_701_368#_c_609_n 0.00314376f $X=3.965 $Y=1.84
+ $X2=0 $Y2=0
cc_352 N_A_501_368#_c_580_n N_A_701_368#_c_609_n 0.0170259f $X=4.1 $Y=2.455
+ $X2=0 $Y2=0
cc_353 N_A_501_368#_c_573_n N_A_701_368#_c_602_n 0.00341172f $X=3.935 $Y=2.99
+ $X2=0 $Y2=0

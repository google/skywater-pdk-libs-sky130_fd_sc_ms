* File: sky130_fd_sc_ms__a22oi_2.spice
* Created: Fri Aug 28 17:03:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a22oi_2.pex.spice"
.subckt sky130_fd_sc_ms__a22oi_2  VNB VPB A1 A2 B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A1_M1002_g N_A_148_74#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1001 N_A_148_74#_M1002_s N_A2_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_148_74#_M1004_d N_A2_M1004_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_148_74#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.1036 PD=1.28 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1005 N_A_558_74#_M1005_d N_B1_M1005_g N_Y_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1998 PD=1.13 PS=1.28 NRD=11.34 NRS=25.128 M=1 R=4.93333
+ SA=75002.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_B2_M1007_g N_A_558_74#_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1443 PD=1.02 PS=1.13 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75002.8
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1007_d N_B2_M1014_g N_A_558_74#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_558_74#_M1014_s N_B1_M1006_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_66_368#_M1000_d N_A1_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1009 N_A_66_368#_M1009_d N_A2_M1009_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1011 N_A_66_368#_M1009_d N_A2_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3248 PD=1.39 PS=1.7 NRD=0 NRS=26.3783 M=1 R=6.22222 SA=90001.1
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1008 N_A_66_368#_M1008_d N_A1_M1008_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3248 PD=1.39 PS=1.7 NRD=0 NRS=26.3783 M=1 R=6.22222 SA=90001.8
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_66_368#_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.168 AS=0.1512 PD=1.42 PS=1.39 NRD=1.7533 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1010 N_A_66_368#_M1010_d N_B2_M1010_g N_Y_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.168 PD=1.39 PS=1.42 NRD=0 NRS=1.7533 M=1 R=6.22222 SA=90002.8
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1012 N_A_66_368#_M1010_d N_B2_M1012_g N_Y_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1015 N_Y_M1012_s N_B1_M1015_g N_A_66_368#_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__a22oi_2.pxi.spice"
*
.ends
*
*

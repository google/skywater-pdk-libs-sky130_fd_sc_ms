* NGSPICE file created from sky130_fd_sc_ms__sedfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sedfxtp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_2660_508# a_1538_74# a_2474_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=2.962e+11p ps=2.72e+06u
M1001 a_2474_74# a_1538_74# a_2402_74# VNB nlowvt w=640000u l=150000u
+  ad=1.915e+11p pd=1.93e+06u as=1.344e+11p ps=1.7e+06u
M1002 a_693_113# a_663_87# a_1082_455# VPB pshort w=640000u l=180000u
+  ad=4.728e+11p pd=5.07e+06u as=1.536e+11p ps=1.76e+06u
M1003 a_1068_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.2744e+12p ps=1.998e+07u
M1004 a_1340_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VPWR DE a_180_290# VPB pshort w=640000u l=180000u
+  ad=2.92365e+12p pd=2.518e+07u as=1.792e+11p ps=1.84e+06u
M1006 VPWR SCE a_663_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1007 a_1736_97# a_1538_74# a_693_113# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1008 a_693_113# SCE a_1068_125# VNB nlowvt w=420000u l=150000u
+  ad=3.885e+11p pd=4.37e+06u as=0p ps=0u
M1009 a_548_87# a_2474_74# VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1010 Q a_2474_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1011 a_1939_508# a_1340_74# a_1736_97# VPB pshort w=420000u l=180000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1012 a_138_74# D a_40_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.982e+11p ps=3.1e+06u
M1013 a_1538_74# a_1340_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1014 a_1979_71# a_1736_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1015 VPWR a_548_87# a_2660_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_40_464# a_548_87# a_578_463# VPB pshort w=640000u l=180000u
+  ad=3.52e+11p pd=3.66e+06u as=1.344e+11p ps=1.7e+06u
M1017 Q a_2474_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1018 a_132_464# D a_40_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_693_113# SCE a_40_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1736_97# a_1340_74# a_693_113# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1021 VGND DE a_180_290# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1022 a_2360_392# a_1979_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.8e+11p pd=3.56e+06u as=0p ps=0u
M1023 a_500_113# a_180_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1024 VPWR a_1979_71# a_1939_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_2474_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1082_455# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1872_97# a_1538_74# a_1736_97# VNB nlowvt w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1028 a_1979_71# a_1736_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1029 VGND a_1979_71# a_1872_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_578_463# DE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2569_74# a_1340_74# a_2474_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1032 VGND a_548_87# a_2569_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_548_87# a_2474_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1034 a_1340_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1035 a_1538_74# a_1340_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1036 a_40_464# a_548_87# a_500_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_693_113# a_663_87# a_40_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_180_290# a_132_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND DE a_138_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND SCE a_663_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1041 VGND a_2474_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_2474_74# a_1340_74# a_2360_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_2402_74# a_1979_71# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__o41a_4.pxi.spice
* Created: Wed Sep  2 12:27:03 2020
* 
x_PM_SKY130_FD_SC_MS__O41A_4%A_110_48# N_A_110_48#_M1005_s N_A_110_48#_M1011_d
+ N_A_110_48#_M1019_d N_A_110_48#_M1010_g N_A_110_48#_M1003_g
+ N_A_110_48#_M1017_g N_A_110_48#_M1006_g N_A_110_48#_M1020_g
+ N_A_110_48#_M1007_g N_A_110_48#_M1024_g N_A_110_48#_M1009_g
+ N_A_110_48#_c_149_n N_A_110_48#_c_150_n N_A_110_48#_c_161_p
+ N_A_110_48#_c_151_n N_A_110_48#_c_157_n N_A_110_48#_c_158_n
+ N_A_110_48#_c_152_n PM_SKY130_FD_SC_MS__O41A_4%A_110_48#
x_PM_SKY130_FD_SC_MS__O41A_4%B1 N_B1_M1011_g N_B1_M1005_g N_B1_M1014_g
+ N_B1_M1016_g B1 B1 N_B1_c_276_n PM_SKY130_FD_SC_MS__O41A_4%B1
x_PM_SKY130_FD_SC_MS__O41A_4%A4 N_A4_M1019_g N_A4_c_327_n N_A4_M1000_g
+ N_A4_M1021_g N_A4_c_328_n N_A4_M1027_g A4 A4 N_A4_c_330_n
+ PM_SKY130_FD_SC_MS__O41A_4%A4
x_PM_SKY130_FD_SC_MS__O41A_4%A3 N_A3_M1004_g N_A3_c_377_n N_A3_M1015_g
+ N_A3_c_379_n N_A3_c_380_n N_A3_M1023_g N_A3_M1018_g A3 N_A3_c_383_n
+ N_A3_c_384_n PM_SKY130_FD_SC_MS__O41A_4%A3
x_PM_SKY130_FD_SC_MS__O41A_4%A1 N_A1_c_450_n N_A1_M1012_g N_A1_M1001_g
+ N_A1_c_451_n N_A1_M1013_g N_A1_M1026_g A1 A1 N_A1_c_453_n
+ PM_SKY130_FD_SC_MS__O41A_4%A1
x_PM_SKY130_FD_SC_MS__O41A_4%A2 N_A2_M1008_g N_A2_c_499_n N_A2_M1002_g
+ N_A2_c_501_n N_A2_c_502_n N_A2_M1022_g N_A2_M1025_g N_A2_c_505_n A2
+ PM_SKY130_FD_SC_MS__O41A_4%A2
x_PM_SKY130_FD_SC_MS__O41A_4%VPWR N_VPWR_M1003_s N_VPWR_M1006_s N_VPWR_M1009_s
+ N_VPWR_M1014_s N_VPWR_M1001_s N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n
+ N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n
+ N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n
+ N_VPWR_c_575_n N_VPWR_c_576_n VPWR N_VPWR_c_577_n N_VPWR_c_561_n
+ PM_SKY130_FD_SC_MS__O41A_4%VPWR
x_PM_SKY130_FD_SC_MS__O41A_4%X N_X_M1010_d N_X_M1020_d N_X_M1003_d N_X_M1007_d
+ N_X_c_658_n N_X_c_673_n N_X_c_659_n N_X_c_663_n N_X_c_660_n N_X_c_664_n
+ N_X_c_683_n N_X_c_665_n N_X_c_661_n N_X_c_666_n N_X_c_667_n N_X_c_699_n
+ N_X_c_668_n X X X PM_SKY130_FD_SC_MS__O41A_4%X
x_PM_SKY130_FD_SC_MS__O41A_4%A_762_368# N_A_762_368#_M1015_s
+ N_A_762_368#_M1023_s N_A_762_368#_M1025_d N_A_762_368#_c_743_n
+ N_A_762_368#_c_737_n N_A_762_368#_c_754_n N_A_762_368#_c_738_n
+ N_A_762_368#_c_739_n N_A_762_368#_c_740_n N_A_762_368#_c_741_n
+ PM_SKY130_FD_SC_MS__O41A_4%A_762_368#
x_PM_SKY130_FD_SC_MS__O41A_4%A_854_368# N_A_854_368#_M1015_d
+ N_A_854_368#_M1021_s N_A_854_368#_c_788_n
+ PM_SKY130_FD_SC_MS__O41A_4%A_854_368#
x_PM_SKY130_FD_SC_MS__O41A_4%A_1216_368# N_A_1216_368#_M1002_s
+ N_A_1216_368#_M1026_d N_A_1216_368#_c_804_n N_A_1216_368#_c_802_n
+ N_A_1216_368#_c_803_n PM_SKY130_FD_SC_MS__O41A_4%A_1216_368#
x_PM_SKY130_FD_SC_MS__O41A_4%VGND N_VGND_M1010_s N_VGND_M1017_s N_VGND_M1024_s
+ N_VGND_M1004_s N_VGND_M1027_s N_VGND_M1008_s N_VGND_M1013_s N_VGND_c_825_n
+ N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n
+ N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n VGND
+ N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n
+ N_VGND_c_845_n N_VGND_c_846_n PM_SKY130_FD_SC_MS__O41A_4%VGND
x_PM_SKY130_FD_SC_MS__O41A_4%A_523_124# N_A_523_124#_M1005_d
+ N_A_523_124#_M1016_d N_A_523_124#_M1000_d N_A_523_124#_M1018_d
+ N_A_523_124#_M1012_d N_A_523_124#_M1022_d N_A_523_124#_c_946_n
+ N_A_523_124#_c_947_n N_A_523_124#_c_948_n N_A_523_124#_c_949_n
+ N_A_523_124#_c_950_n N_A_523_124#_c_951_n N_A_523_124#_c_952_n
+ N_A_523_124#_c_953_n N_A_523_124#_c_954_n N_A_523_124#_c_955_n
+ N_A_523_124#_c_956_n N_A_523_124#_c_957_n N_A_523_124#_c_1008_n
+ N_A_523_124#_c_958_n N_A_523_124#_c_959_n N_A_523_124#_c_960_n
+ PM_SKY130_FD_SC_MS__O41A_4%A_523_124#
cc_1 VNB N_A_110_48#_M1010_g 0.021193f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_2 VNB N_A_110_48#_M1003_g 0.00377054f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_3 VNB N_A_110_48#_M1017_g 0.0198267f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_4 VNB N_A_110_48#_M1006_g 0.00313923f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_5 VNB N_A_110_48#_M1020_g 0.0203883f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.74
cc_6 VNB N_A_110_48#_M1007_g 0.00313923f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=2.4
cc_7 VNB N_A_110_48#_M1024_g 0.0257334f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_8 VNB N_A_110_48#_M1009_g 0.00342768f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=2.4
cc_9 VNB N_A_110_48#_c_149_n 0.0185991f $X=-0.19 $Y=-0.245 $X2=2.78 $Y2=1.435
cc_10 VNB N_A_110_48#_c_150_n 0.00727972f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=1.6
cc_11 VNB N_A_110_48#_c_151_n 0.00170949f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=0.765
cc_12 VNB N_A_110_48#_c_152_n 0.103391f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.435
cc_13 VNB N_B1_M1011_g 0.00366516f $X=-0.19 $Y=-0.245 $X2=4.72 $Y2=1.84
cc_14 VNB N_B1_M1005_g 0.0213334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1016_g 0.020157f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_16 VNB B1 0.00226907f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.27
cc_17 VNB N_B1_c_276_n 0.0427953f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_18 VNB N_A4_c_327_n 0.0175218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A4_c_328_n 0.0139587f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_20 VNB A4 0.00518079f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_21 VNB N_A4_c_330_n 0.0351577f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.27
cc_22 VNB N_A3_M1004_g 0.00753503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A3_c_377_n 0.0256922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A3_M1015_g 0.00980353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_c_379_n 0.0989471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A3_c_380_n 0.0058681f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_27 VNB N_A3_M1023_g 0.0144043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A3_M1018_g 0.0235342f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.27
cc_29 VNB N_A3_c_383_n 0.0503978f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.27
cc_30 VNB N_A3_c_384_n 7.54705e-19 $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.6
cc_31 VNB N_A1_c_450_n 0.0147706f $X=-0.19 $Y=-0.245 $X2=3.05 $Y2=0.62
cc_32 VNB N_A1_c_451_n 0.0146138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB A1 0.00730714f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_34 VNB N_A1_c_453_n 0.0357709f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_35 VNB N_A2_M1008_g 0.0235707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_c_499_n 0.00579793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A2_M1002_g 0.0142072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A2_c_501_n 0.137982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A2_c_502_n 0.00954688f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.27
cc_40 VNB N_A2_M1022_g 0.01277f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.6
cc_41 VNB N_A2_M1025_g 0.0158535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A2_c_505_n 0.0202403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB A2 0.0401964f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.6
cc_44 VNB N_VPWR_c_561_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_658_n 0.0274757f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.6
cc_46 VNB N_X_c_659_n 0.00961898f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.4
cc_47 VNB N_X_c_660_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_X_c_661_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_49 VNB N_VGND_c_825_n 0.0141307f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.6
cc_50 VNB N_VGND_c_826_n 0.0274339f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_51 VNB N_VGND_c_827_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.74
cc_52 VNB N_VGND_c_828_n 0.0143472f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=2.4
cc_53 VNB N_VGND_c_829_n 0.00781633f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_54 VNB N_VGND_c_830_n 0.00341672f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=2.4
cc_55 VNB N_VGND_c_831_n 0.00469205f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.435
cc_56 VNB N_VGND_c_832_n 0.0160886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_833_n 0.0061168f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=1.6
cc_58 VNB N_VGND_c_834_n 0.0492942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_835_n 0.00229531f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.1
cc_60 VNB N_VGND_c_836_n 0.0160886f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=0.765
cc_61 VNB N_VGND_c_837_n 0.00445561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_838_n 0.0142087f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=2.035
cc_63 VNB N_VGND_c_839_n 0.00337546f $X=-0.19 $Y=-0.245 $X2=4.86 $Y2=2.035
cc_64 VNB N_VGND_c_840_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=3.027 $Y2=1.435
cc_65 VNB N_VGND_c_841_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.435
cc_66 VNB N_VGND_c_842_n 0.0272543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_843_n 0.437198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_844_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_845_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_846_n 0.00337546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_523_124#_c_946_n 0.00615577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_523_124#_c_947_n 0.0156685f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_73 VNB N_A_523_124#_c_948_n 0.00497327f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.4
cc_74 VNB N_A_523_124#_c_949_n 0.00215445f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.74
cc_75 VNB N_A_523_124#_c_950_n 0.00737922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_523_124#_c_951_n 0.00178935f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.6
cc_77 VNB N_A_523_124#_c_952_n 0.001978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_523_124#_c_953_n 0.0112124f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.74
cc_79 VNB N_A_523_124#_c_954_n 0.00254618f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=2.4
cc_80 VNB N_A_523_124#_c_955_n 0.0105793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_523_124#_c_956_n 0.00197771f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.435
cc_82 VNB N_A_523_124#_c_957_n 0.00525165f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=1.435
cc_83 VNB N_A_523_124#_c_958_n 0.00176133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_523_124#_c_959_n 0.00322493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_523_124#_c_960_n 0.00176197f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.1
cc_86 VPB N_A_110_48#_M1003_g 0.0247573f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.4
cc_87 VPB N_A_110_48#_M1006_g 0.0218093f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_88 VPB N_A_110_48#_M1007_g 0.0218093f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=2.4
cc_89 VPB N_A_110_48#_M1009_g 0.0237231f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.4
cc_90 VPB N_A_110_48#_c_157_n 0.0122307f $X=-0.19 $Y=1.66 $X2=4.86 $Y2=2.035
cc_91 VPB N_A_110_48#_c_158_n 0.00314017f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=2.075
cc_92 VPB N_B1_M1011_g 0.0272447f $X=-0.19 $Y=1.66 $X2=4.72 $Y2=1.84
cc_93 VPB N_B1_M1014_g 0.0252141f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=0.74
cc_94 VPB B1 0.0080897f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.27
cc_95 VPB N_B1_c_276_n 0.0197195f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_96 VPB N_A4_M1019_g 0.0208719f $X=-0.19 $Y=1.66 $X2=4.72 $Y2=1.84
cc_97 VPB N_A4_M1021_g 0.0208711f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.27
cc_98 VPB A4 0.00577f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.4
cc_99 VPB N_A4_c_330_n 0.00562645f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.27
cc_100 VPB N_A3_M1015_g 0.0267321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A3_M1023_g 0.023535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A1_M1001_g 0.0212756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A1_M1026_g 0.0212694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB A1 0.00647886f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.4
cc_105 VPB N_A1_c_453_n 0.00628559f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=2.4
cc_106 VPB N_A2_M1002_g 0.0234902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A2_M1025_g 0.0320291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_562_n 0.0111983f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.27
cc_109 VPB N_VPWR_c_563_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=1.6
cc_110 VPB N_VPWR_c_564_n 0.0163342f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.27
cc_111 VPB N_VPWR_c_565_n 0.023747f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=1.6
cc_112 VPB N_VPWR_c_566_n 0.00598808f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=1.27
cc_113 VPB N_VPWR_c_567_n 0.0173573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_568_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=1.6
cc_115 VPB N_VPWR_c_569_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.4
cc_116 VPB N_VPWR_c_570_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_571_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.435
cc_118 VPB N_VPWR_c_572_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.435
cc_119 VPB N_VPWR_c_573_n 0.0215627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_574_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_121 VPB N_VPWR_c_575_n 0.0805589f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_122 VPB N_VPWR_c_576_n 0.00535801f $X=-0.19 $Y=1.66 $X2=2.945 $Y2=1.6
cc_123 VPB N_VPWR_c_577_n 0.037911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_561_n 0.123341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_X_c_658_n 0.00575776f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.6
cc_126 VPB N_X_c_663_n 0.00885417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_X_c_664_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_X_c_665_n 0.00443716f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=2.4
cc_129 VPB N_X_c_666_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.4
cc_130 VPB N_X_c_667_n 0.00928121f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.435
cc_131 VPB N_X_c_668_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB X 0.0509563f $X=-0.19 $Y=1.66 $X2=2.11 $Y2=1.435
cc_133 VPB N_A_762_368#_c_737_n 0.00307266f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.6
cc_134 VPB N_A_762_368#_c_738_n 0.0233424f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_135 VPB N_A_762_368#_c_739_n 0.0357634f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=1.6
cc_136 VPB N_A_762_368#_c_740_n 0.00884675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_762_368#_c_741_n 0.00178969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_854_368#_c_788_n 0.00695998f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=0.74
cc_139 VPB N_A_1216_368#_c_802_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.6
cc_140 VPB N_A_1216_368#_c_803_n 0.00275743f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.4
cc_141 N_A_110_48#_M1009_g N_B1_M1011_g 0.0155799f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_110_48#_c_149_n N_B1_M1011_g 0.00734048f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_143 N_A_110_48#_c_161_p N_B1_M1011_g 0.0106664f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_144 N_A_110_48#_c_158_n N_B1_M1011_g 0.0127095f $X=2.945 $Y=2.075 $X2=0 $Y2=0
cc_145 N_A_110_48#_c_150_n N_B1_M1005_g 0.0194369f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_146 N_A_110_48#_c_152_n N_B1_M1005_g 0.00213441f $X=2.185 $Y=1.435 $X2=0
+ $Y2=0
cc_147 N_A_110_48#_c_161_p N_B1_M1014_g 0.00943938f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_148 N_A_110_48#_c_157_n N_B1_M1014_g 0.0193664f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_149 N_A_110_48#_c_158_n N_B1_M1014_g 0.0166896f $X=2.945 $Y=2.075 $X2=0 $Y2=0
cc_150 N_A_110_48#_c_150_n N_B1_M1016_g 0.00448353f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_151 N_A_110_48#_c_150_n B1 0.0134595f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_152 N_A_110_48#_c_161_p B1 0.0142537f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_153 N_A_110_48#_c_157_n B1 0.0677548f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_154 N_A_110_48#_c_149_n N_B1_c_276_n 0.00691491f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_155 N_A_110_48#_c_150_n N_B1_c_276_n 0.0162985f $X=2.945 $Y=1.6 $X2=0 $Y2=0
cc_156 N_A_110_48#_c_161_p N_B1_c_276_n 0.00479112f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_157 N_A_110_48#_c_157_n N_B1_c_276_n 0.00216518f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_158 N_A_110_48#_c_152_n N_B1_c_276_n 0.0155799f $X=2.185 $Y=1.435 $X2=0 $Y2=0
cc_159 N_A_110_48#_c_157_n N_A4_M1019_g 0.00963748f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_160 N_A_110_48#_c_157_n N_A4_M1021_g 0.00421605f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_161 N_A_110_48#_c_157_n A4 0.0382125f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_162 N_A_110_48#_c_157_n N_A4_c_330_n 5.43181e-19 $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_163 N_A_110_48#_c_157_n N_A3_c_377_n 8.11334e-19 $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_164 N_A_110_48#_c_157_n N_A3_M1015_g 0.0159132f $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_165 N_A_110_48#_c_157_n N_A3_M1023_g 5.03893e-19 $X=4.86 $Y=2.035 $X2=0 $Y2=0
cc_166 N_A_110_48#_c_157_n N_VPWR_M1014_s 0.00517312f $X=4.86 $Y=2.035 $X2=0
+ $Y2=0
cc_167 N_A_110_48#_M1003_g N_VPWR_c_562_n 0.00782815f $X=0.835 $Y=2.4 $X2=0
+ $Y2=0
cc_168 N_A_110_48#_M1006_g N_VPWR_c_563_n 0.00342026f $X=1.285 $Y=2.4 $X2=0
+ $Y2=0
cc_169 N_A_110_48#_M1007_g N_VPWR_c_563_n 0.00342026f $X=1.735 $Y=2.4 $X2=0
+ $Y2=0
cc_170 N_A_110_48#_M1009_g N_VPWR_c_564_n 0.00753041f $X=2.185 $Y=2.4 $X2=0
+ $Y2=0
cc_171 N_A_110_48#_c_149_n N_VPWR_c_564_n 0.013831f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_172 N_A_110_48#_c_161_p N_VPWR_c_564_n 0.00192425f $X=2.945 $Y=1.95 $X2=0
+ $Y2=0
cc_173 N_A_110_48#_c_158_n N_VPWR_c_564_n 0.0222747f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_174 N_A_110_48#_c_157_n N_VPWR_c_565_n 0.0197477f $X=4.86 $Y=2.035 $X2=0
+ $Y2=0
cc_175 N_A_110_48#_c_158_n N_VPWR_c_565_n 0.0171487f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_176 N_A_110_48#_M1003_g N_VPWR_c_569_n 0.005209f $X=0.835 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_110_48#_M1006_g N_VPWR_c_569_n 0.005209f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A_110_48#_M1007_g N_VPWR_c_571_n 0.005209f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_110_48#_M1009_g N_VPWR_c_571_n 0.005209f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_110_48#_c_158_n N_VPWR_c_573_n 0.00806582f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_181 N_A_110_48#_M1003_g N_VPWR_c_561_n 0.00987399f $X=0.835 $Y=2.4 $X2=0
+ $Y2=0
cc_182 N_A_110_48#_M1006_g N_VPWR_c_561_n 0.00982266f $X=1.285 $Y=2.4 $X2=0
+ $Y2=0
cc_183 N_A_110_48#_M1007_g N_VPWR_c_561_n 0.00982266f $X=1.735 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A_110_48#_M1009_g N_VPWR_c_561_n 0.00987399f $X=2.185 $Y=2.4 $X2=0
+ $Y2=0
cc_185 N_A_110_48#_c_158_n N_VPWR_c_561_n 0.0106017f $X=2.945 $Y=2.075 $X2=0
+ $Y2=0
cc_186 N_A_110_48#_M1010_g N_X_c_658_n 0.0135824f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_110_48#_M1003_g N_X_c_658_n 0.00439804f $X=0.835 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_110_48#_c_149_n N_X_c_658_n 0.0175348f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_189 N_A_110_48#_M1010_g N_X_c_673_n 0.0132299f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_110_48#_c_149_n N_X_c_673_n 0.00639324f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_191 N_A_110_48#_M1003_g N_X_c_663_n 0.0148618f $X=0.835 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_110_48#_c_149_n N_X_c_663_n 0.0227031f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_193 N_A_110_48#_c_152_n N_X_c_663_n 0.00531264f $X=2.185 $Y=1.435 $X2=0 $Y2=0
cc_194 N_A_110_48#_M1010_g N_X_c_660_n 0.0121547f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_110_48#_M1017_g N_X_c_660_n 2.71222e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_110_48#_M1003_g N_X_c_664_n 0.0154931f $X=0.835 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_110_48#_M1006_g N_X_c_664_n 0.014659f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_110_48#_M1007_g N_X_c_664_n 7.07432e-19 $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_110_48#_M1017_g N_X_c_683_n 0.012639f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_110_48#_M1020_g N_X_c_683_n 0.0122754f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_110_48#_c_149_n N_X_c_683_n 0.061224f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_202 N_A_110_48#_c_152_n N_X_c_683_n 0.00720526f $X=2.185 $Y=1.435 $X2=0 $Y2=0
cc_203 N_A_110_48#_M1006_g N_X_c_665_n 0.012931f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_110_48#_M1007_g N_X_c_665_n 0.0146352f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_110_48#_M1009_g N_X_c_665_n 0.00453707f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_110_48#_c_149_n N_X_c_665_n 0.0692143f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_207 N_A_110_48#_c_161_p N_X_c_665_n 0.00361447f $X=2.945 $Y=1.95 $X2=0 $Y2=0
cc_208 N_A_110_48#_c_152_n N_X_c_665_n 0.00482403f $X=2.185 $Y=1.435 $X2=0 $Y2=0
cc_209 N_A_110_48#_M1017_g N_X_c_661_n 9.1509e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_110_48#_M1020_g N_X_c_661_n 0.00804372f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_110_48#_M1024_g N_X_c_661_n 2.71222e-19 $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_110_48#_M1006_g N_X_c_666_n 7.07432e-19 $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A_110_48#_M1007_g N_X_c_666_n 0.014659f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_110_48#_M1009_g N_X_c_666_n 0.0136331f $X=2.185 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_110_48#_M1010_g N_X_c_699_n 7.32094e-19 $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_110_48#_c_149_n N_X_c_699_n 0.0178863f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_217 N_A_110_48#_c_152_n N_X_c_699_n 0.00272398f $X=2.185 $Y=1.435 $X2=0 $Y2=0
cc_218 N_A_110_48#_M1003_g N_X_c_668_n 0.00170419f $X=0.835 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_110_48#_M1006_g N_X_c_668_n 0.00170419f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_110_48#_c_149_n N_X_c_668_n 0.0275631f $X=2.78 $Y=1.435 $X2=0 $Y2=0
cc_221 N_A_110_48#_c_152_n N_X_c_668_n 0.00245159f $X=2.185 $Y=1.435 $X2=0 $Y2=0
cc_222 N_A_110_48#_M1003_g X 0.00389973f $X=0.835 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_110_48#_c_157_n N_A_762_368#_M1015_s 0.00544004f $X=4.86 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_224 N_A_110_48#_M1019_d N_A_762_368#_c_743_n 0.00344903f $X=4.72 $Y=1.84
+ $X2=0 $Y2=0
cc_225 N_A_110_48#_c_157_n N_A_762_368#_c_743_n 0.0497206f $X=4.86 $Y=2.035
+ $X2=0 $Y2=0
cc_226 N_A_110_48#_c_157_n N_A_762_368#_c_740_n 0.0198558f $X=4.86 $Y=2.035
+ $X2=0 $Y2=0
cc_227 N_A_110_48#_c_157_n N_A_854_368#_M1015_d 0.00656964f $X=4.86 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_228 N_A_110_48#_M1019_d N_A_854_368#_c_788_n 0.00180867f $X=4.72 $Y=1.84
+ $X2=0 $Y2=0
cc_229 N_A_110_48#_M1010_g N_VGND_c_826_n 0.0111726f $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_230 N_A_110_48#_M1010_g N_VGND_c_827_n 4.80326e-19 $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_110_48#_M1017_g N_VGND_c_827_n 0.00877665f $X=1.055 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_110_48#_M1020_g N_VGND_c_827_n 0.00382194f $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_110_48#_M1020_g N_VGND_c_828_n 5.81525e-19 $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_110_48#_M1024_g N_VGND_c_828_n 0.0138071f $X=1.985 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_110_48#_c_149_n N_VGND_c_828_n 0.0248195f $X=2.78 $Y=1.435 $X2=0
+ $Y2=0
cc_236 N_A_110_48#_c_152_n N_VGND_c_828_n 0.00568288f $X=2.185 $Y=1.435 $X2=0
+ $Y2=0
cc_237 N_A_110_48#_M1010_g N_VGND_c_840_n 0.00434272f $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_110_48#_M1017_g N_VGND_c_840_n 0.00383152f $X=1.055 $Y=0.74 $X2=0
+ $Y2=0
cc_239 N_A_110_48#_M1020_g N_VGND_c_841_n 0.00434272f $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_110_48#_M1024_g N_VGND_c_841_n 0.00383152f $X=1.985 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_110_48#_M1010_g N_VGND_c_843_n 0.00824087f $X=0.625 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_110_48#_M1017_g N_VGND_c_843_n 0.0075754f $X=1.055 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_110_48#_M1020_g N_VGND_c_843_n 0.00820718f $X=1.555 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_110_48#_M1024_g N_VGND_c_843_n 0.0075754f $X=1.985 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_110_48#_M1024_g N_A_523_124#_c_946_n 9.31825e-19 $X=1.985 $Y=0.74
+ $X2=0 $Y2=0
cc_246 N_A_110_48#_c_149_n N_A_523_124#_c_946_n 0.00970275f $X=2.78 $Y=1.435
+ $X2=0 $Y2=0
cc_247 N_A_110_48#_c_150_n N_A_523_124#_c_946_n 0.0062953f $X=2.945 $Y=1.6 $X2=0
+ $Y2=0
cc_248 N_A_110_48#_c_151_n N_A_523_124#_c_946_n 0.0125142f $X=3.19 $Y=0.765
+ $X2=0 $Y2=0
cc_249 N_A_110_48#_c_150_n N_A_523_124#_c_947_n 0.00380631f $X=2.945 $Y=1.6
+ $X2=0 $Y2=0
cc_250 N_A_110_48#_c_151_n N_A_523_124#_c_947_n 0.0132727f $X=3.19 $Y=0.765
+ $X2=0 $Y2=0
cc_251 N_A_110_48#_M1024_g N_A_523_124#_c_948_n 5.9337e-19 $X=1.985 $Y=0.74
+ $X2=0 $Y2=0
cc_252 N_A_110_48#_c_151_n N_A_523_124#_c_949_n 0.0173112f $X=3.19 $Y=0.765
+ $X2=0 $Y2=0
cc_253 N_A_110_48#_c_150_n N_A_523_124#_c_951_n 0.00714719f $X=2.945 $Y=1.6
+ $X2=0 $Y2=0
cc_254 B1 A4 0.0225058f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_255 B1 N_A4_c_330_n 2.39067e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_256 B1 N_A3_c_377_n 0.0108947f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_257 N_B1_c_276_n N_A3_c_377_n 0.00250407f $X=3.405 $Y=1.605 $X2=0 $Y2=0
cc_258 B1 N_A3_M1015_g 0.0119079f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_259 N_B1_c_276_n N_A3_M1015_g 0.00591861f $X=3.405 $Y=1.605 $X2=0 $Y2=0
cc_260 N_B1_M1016_g N_A3_c_383_n 0.0197827f $X=3.405 $Y=0.94 $X2=0 $Y2=0
cc_261 N_B1_M1011_g N_VPWR_c_564_n 0.00783518f $X=2.72 $Y=2.35 $X2=0 $Y2=0
cc_262 N_B1_M1014_g N_VPWR_c_565_n 0.0068611f $X=3.17 $Y=2.35 $X2=0 $Y2=0
cc_263 N_B1_M1011_g N_VPWR_c_573_n 0.00520125f $X=2.72 $Y=2.35 $X2=0 $Y2=0
cc_264 N_B1_M1014_g N_VPWR_c_573_n 0.00520125f $X=3.17 $Y=2.35 $X2=0 $Y2=0
cc_265 N_B1_M1011_g N_VPWR_c_561_n 0.00585323f $X=2.72 $Y=2.35 $X2=0 $Y2=0
cc_266 N_B1_M1014_g N_VPWR_c_561_n 0.00585323f $X=3.17 $Y=2.35 $X2=0 $Y2=0
cc_267 N_B1_M1011_g N_X_c_665_n 4.37439e-19 $X=2.72 $Y=2.35 $X2=0 $Y2=0
cc_268 N_B1_M1005_g N_VGND_c_828_n 0.00500871f $X=2.975 $Y=0.94 $X2=0 $Y2=0
cc_269 N_B1_M1005_g N_VGND_c_834_n 2.27419e-19 $X=2.975 $Y=0.94 $X2=0 $Y2=0
cc_270 N_B1_M1016_g N_VGND_c_834_n 2.27419e-19 $X=3.405 $Y=0.94 $X2=0 $Y2=0
cc_271 N_B1_M1005_g N_A_523_124#_c_946_n 0.00888778f $X=2.975 $Y=0.94 $X2=0
+ $Y2=0
cc_272 N_B1_M1016_g N_A_523_124#_c_946_n 4.22299e-19 $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_273 N_B1_c_276_n N_A_523_124#_c_946_n 0.00125597f $X=3.405 $Y=1.605 $X2=0
+ $Y2=0
cc_274 N_B1_M1005_g N_A_523_124#_c_947_n 0.0046393f $X=2.975 $Y=0.94 $X2=0 $Y2=0
cc_275 N_B1_M1016_g N_A_523_124#_c_947_n 0.00582977f $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_276 N_B1_M1005_g N_A_523_124#_c_949_n 4.69875e-19 $X=2.975 $Y=0.94 $X2=0
+ $Y2=0
cc_277 N_B1_M1016_g N_A_523_124#_c_949_n 0.00880445f $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_278 B1 N_A_523_124#_c_950_n 0.03029f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_279 N_B1_M1016_g N_A_523_124#_c_951_n 0.00236422f $X=3.405 $Y=0.94 $X2=0
+ $Y2=0
cc_280 B1 N_A_523_124#_c_951_n 0.0213654f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_281 N_B1_c_276_n N_A_523_124#_c_951_n 0.00302844f $X=3.405 $Y=1.605 $X2=0
+ $Y2=0
cc_282 N_A4_c_327_n N_A3_M1004_g 0.00814159f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_283 N_A4_c_327_n N_A3_c_377_n 6.90332e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_284 A4 N_A3_c_377_n 0.00293696f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_285 N_A4_c_330_n N_A3_c_377_n 0.0184214f $X=5.105 $Y=1.515 $X2=0 $Y2=0
cc_286 N_A4_M1019_g N_A3_M1015_g 0.0530691f $X=4.63 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A4_c_327_n N_A3_c_379_n 0.0103098f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_288 N_A4_c_328_n N_A3_c_379_n 0.0103186f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_289 N_A4_c_328_n N_A3_c_380_n 0.0345239f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_290 A4 N_A3_M1023_g 0.00224638f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_291 N_A4_c_330_n N_A3_M1023_g 0.0345239f $X=5.105 $Y=1.515 $X2=0 $Y2=0
cc_292 N_A4_c_328_n N_A3_M1018_g 0.0226172f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_293 N_A4_c_327_n N_A3_c_383_n 9.14655e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_294 N_A4_M1019_g N_VPWR_c_575_n 0.00349978f $X=4.63 $Y=2.4 $X2=0 $Y2=0
cc_295 N_A4_M1021_g N_VPWR_c_575_n 0.00349978f $X=5.09 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A4_M1019_g N_VPWR_c_561_n 0.00429731f $X=4.63 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A4_M1021_g N_VPWR_c_561_n 0.00429731f $X=5.09 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A4_M1019_g N_A_762_368#_c_743_n 0.0116873f $X=4.63 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A4_M1021_g N_A_762_368#_c_743_n 0.0133888f $X=5.09 $Y=2.4 $X2=0 $Y2=0
cc_300 A4 N_A_762_368#_c_743_n 0.00439412f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_301 N_A4_M1019_g N_A_854_368#_c_788_n 0.014539f $X=4.63 $Y=2.4 $X2=0 $Y2=0
cc_302 N_A4_M1021_g N_A_854_368#_c_788_n 0.014539f $X=5.09 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A4_c_327_n N_VGND_c_829_n 0.00291089f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_304 N_A4_c_327_n N_VGND_c_830_n 4.43476e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_305 N_A4_c_328_n N_VGND_c_830_n 0.0075897f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_306 N_A4_c_327_n N_VGND_c_843_n 9.33152e-19 $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_307 N_A4_c_328_n N_VGND_c_843_n 7.83848e-19 $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_308 N_A4_c_327_n N_A_523_124#_c_950_n 0.0121471f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_309 A4 N_A_523_124#_c_950_n 0.0209304f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_310 N_A4_c_330_n N_A_523_124#_c_950_n 0.00246149f $X=5.105 $Y=1.515 $X2=0
+ $Y2=0
cc_311 N_A4_c_327_n N_A_523_124#_c_952_n 0.0112487f $X=4.675 $Y=1.35 $X2=0 $Y2=0
cc_312 N_A4_c_328_n N_A_523_124#_c_953_n 0.0121744f $X=5.105 $Y=1.35 $X2=0 $Y2=0
cc_313 A4 N_A_523_124#_c_953_n 0.0148952f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_314 N_A4_c_327_n N_A_523_124#_c_958_n 9.00612e-19 $X=4.675 $Y=1.35 $X2=0
+ $Y2=0
cc_315 A4 N_A_523_124#_c_958_n 0.0210654f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_316 N_A4_c_330_n N_A_523_124#_c_958_n 0.00267502f $X=5.105 $Y=1.515 $X2=0
+ $Y2=0
cc_317 N_A3_M1018_g N_A2_M1008_g 0.0120828f $X=5.535 $Y=0.92 $X2=0 $Y2=0
cc_318 N_A3_c_380_n N_A2_c_499_n 0.0177768f $X=5.54 $Y=1.405 $X2=0 $Y2=0
cc_319 N_A3_M1023_g N_A2_M1002_g 0.0177768f $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_320 N_A3_c_379_n N_A2_c_502_n 0.0120828f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_321 N_A3_M1015_g N_VPWR_c_565_n 0.00356525f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_322 N_A3_M1015_g N_VPWR_c_575_n 0.00519794f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_323 N_A3_M1023_g N_VPWR_c_575_n 0.00519794f $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_324 N_A3_M1015_g N_VPWR_c_561_n 0.0098496f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A3_M1023_g N_VPWR_c_561_n 0.00979937f $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_326 N_A3_M1015_g N_A_762_368#_c_743_n 0.0139531f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_327 N_A3_M1023_g N_A_762_368#_c_743_n 0.01942f $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_328 N_A3_M1023_g N_A_762_368#_c_737_n 4.63009e-19 $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_329 N_A3_M1015_g N_A_762_368#_c_740_n 4.8693e-19 $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_330 N_A3_M1023_g N_A_762_368#_c_741_n 2.71287e-19 $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_331 N_A3_M1015_g N_A_854_368#_c_788_n 0.00528582f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_332 N_A3_M1023_g N_A_854_368#_c_788_n 0.00506122f $X=5.54 $Y=2.4 $X2=0 $Y2=0
cc_333 N_A3_c_384_n N_VGND_M1004_s 0.00269695f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_334 N_A3_M1004_g N_VGND_c_829_n 0.00247081f $X=3.925 $Y=0.94 $X2=0 $Y2=0
cc_335 N_A3_c_379_n N_VGND_c_829_n 0.0160258f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_336 N_A3_c_383_n N_VGND_c_829_n 0.0050871f $X=4.027 $Y=0.185 $X2=0 $Y2=0
cc_337 N_A3_c_384_n N_VGND_c_829_n 0.0316618f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_338 N_A3_c_379_n N_VGND_c_830_n 0.02003f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_339 N_A3_M1018_g N_VGND_c_830_n 0.0151923f $X=5.535 $Y=0.92 $X2=0 $Y2=0
cc_340 N_A3_c_379_n N_VGND_c_831_n 0.00157927f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_341 N_A3_c_383_n N_VGND_c_834_n 0.0147334f $X=4.027 $Y=0.185 $X2=0 $Y2=0
cc_342 N_A3_c_384_n N_VGND_c_834_n 0.0215843f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_343 N_A3_c_379_n N_VGND_c_836_n 0.0185349f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_344 N_A3_c_379_n N_VGND_c_838_n 0.0048178f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_345 N_A3_c_379_n N_VGND_c_843_n 0.0382998f $X=5.46 $Y=0.185 $X2=0 $Y2=0
cc_346 N_A3_c_383_n N_VGND_c_843_n 0.0117598f $X=4.027 $Y=0.185 $X2=0 $Y2=0
cc_347 N_A3_c_384_n N_VGND_c_843_n 0.0110944f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_348 N_A3_c_383_n N_A_523_124#_c_947_n 0.0041408f $X=4.027 $Y=0.185 $X2=0
+ $Y2=0
cc_349 N_A3_c_384_n N_A_523_124#_c_947_n 0.0143361f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_350 N_A3_c_383_n N_A_523_124#_c_949_n 0.0100067f $X=4.027 $Y=0.185 $X2=0
+ $Y2=0
cc_351 N_A3_c_384_n N_A_523_124#_c_949_n 0.0184329f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_352 N_A3_M1004_g N_A_523_124#_c_950_n 0.0139445f $X=3.925 $Y=0.94 $X2=0 $Y2=0
cc_353 N_A3_c_377_n N_A_523_124#_c_950_n 0.00830231f $X=4.18 $Y=1.485 $X2=0
+ $Y2=0
cc_354 N_A3_c_383_n N_A_523_124#_c_950_n 7.57014e-19 $X=4.027 $Y=0.185 $X2=0
+ $Y2=0
cc_355 N_A3_c_384_n N_A_523_124#_c_950_n 0.0103418f $X=4.04 $Y=0.345 $X2=0 $Y2=0
cc_356 N_A3_M1004_g N_A_523_124#_c_951_n 3.89157e-19 $X=3.925 $Y=0.94 $X2=0
+ $Y2=0
cc_357 N_A3_c_379_n N_A_523_124#_c_952_n 0.00461056f $X=5.46 $Y=0.185 $X2=0
+ $Y2=0
cc_358 N_A3_c_380_n N_A_523_124#_c_953_n 0.00140384f $X=5.54 $Y=1.405 $X2=0
+ $Y2=0
cc_359 N_A3_M1018_g N_A_523_124#_c_953_n 0.0169653f $X=5.535 $Y=0.92 $X2=0 $Y2=0
cc_360 N_A1_c_450_n N_A2_M1008_g 0.0218812f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_361 N_A1_c_450_n N_A2_c_499_n 0.00954005f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_362 N_A1_M1001_g N_A2_M1002_g 0.0344063f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_363 A1 N_A2_M1002_g 0.00416122f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_364 N_A1_c_453_n N_A2_M1002_g 0.00954005f $X=6.835 $Y=1.515 $X2=0 $Y2=0
cc_365 N_A1_c_450_n N_A2_c_501_n 0.0103098f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_366 N_A1_c_451_n N_A2_c_501_n 0.024217f $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_367 N_A1_c_453_n N_A2_M1022_g 0.0138985f $X=6.835 $Y=1.515 $X2=0 $Y2=0
cc_368 A1 N_A2_M1025_g 0.00755752f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_369 N_A1_c_453_n N_A2_M1025_g 0.0346794f $X=6.835 $Y=1.515 $X2=0 $Y2=0
cc_370 A1 N_A2_c_505_n 0.00166919f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A1_M1001_g N_VPWR_c_566_n 0.00313311f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A1_M1026_g N_VPWR_c_566_n 0.00826381f $X=6.93 $Y=2.4 $X2=0 $Y2=0
cc_373 N_A1_M1001_g N_VPWR_c_575_n 0.005209f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_374 N_A1_M1026_g N_VPWR_c_577_n 0.00460063f $X=6.93 $Y=2.4 $X2=0 $Y2=0
cc_375 N_A1_M1001_g N_VPWR_c_561_n 0.00982771f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_376 N_A1_M1026_g N_VPWR_c_561_n 0.00909121f $X=6.93 $Y=2.4 $X2=0 $Y2=0
cc_377 N_A1_M1001_g N_A_762_368#_c_754_n 0.0118637f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_378 N_A1_M1026_g N_A_762_368#_c_754_n 0.0121509f $X=6.93 $Y=2.4 $X2=0 $Y2=0
cc_379 A1 N_A_762_368#_c_754_n 0.0492494f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_380 N_A1_c_453_n N_A_762_368#_c_754_n 7.03243e-19 $X=6.835 $Y=1.515 $X2=0
+ $Y2=0
cc_381 N_A1_M1001_g N_A_1216_368#_c_804_n 0.012936f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_382 N_A1_M1026_g N_A_1216_368#_c_804_n 0.0142833f $X=6.93 $Y=2.4 $X2=0 $Y2=0
cc_383 N_A1_M1001_g N_A_1216_368#_c_802_n 0.00923349f $X=6.44 $Y=2.4 $X2=0 $Y2=0
cc_384 N_A1_M1026_g N_A_1216_368#_c_802_n 6.16295e-19 $X=6.93 $Y=2.4 $X2=0 $Y2=0
cc_385 N_A1_c_450_n N_VGND_c_831_n 0.00159705f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_386 N_A1_c_450_n N_VGND_c_833_n 4.43355e-19 $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_387 N_A1_c_451_n N_VGND_c_833_n 0.00739822f $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_388 N_A1_c_450_n N_VGND_c_843_n 9.33152e-19 $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_389 N_A1_c_451_n N_VGND_c_843_n 7.83848e-19 $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_390 N_A1_c_450_n N_A_523_124#_c_955_n 0.0108924f $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_391 A1 N_A_523_124#_c_955_n 0.00895556f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_392 N_A1_c_450_n N_A_523_124#_c_956_n 0.00706136f $X=6.405 $Y=1.35 $X2=0
+ $Y2=0
cc_393 N_A1_c_451_n N_A_523_124#_c_957_n 0.0126082f $X=6.835 $Y=1.35 $X2=0 $Y2=0
cc_394 A1 N_A_523_124#_c_957_n 0.0279976f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_395 N_A1_c_453_n N_A_523_124#_c_957_n 5.78783e-19 $X=6.835 $Y=1.515 $X2=0
+ $Y2=0
cc_396 N_A1_c_451_n N_A_523_124#_c_1008_n 7.33515e-19 $X=6.835 $Y=1.35 $X2=0
+ $Y2=0
cc_397 N_A1_c_450_n N_A_523_124#_c_960_n 8.4031e-19 $X=6.405 $Y=1.35 $X2=0 $Y2=0
cc_398 A1 N_A_523_124#_c_960_n 0.0210731f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_399 N_A1_c_453_n N_A_523_124#_c_960_n 0.00274327f $X=6.835 $Y=1.515 $X2=0
+ $Y2=0
cc_400 N_A2_M1025_g N_VPWR_c_566_n 6.14206e-19 $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_401 N_A2_M1002_g N_VPWR_c_575_n 0.005209f $X=5.99 $Y=2.4 $X2=0 $Y2=0
cc_402 N_A2_M1025_g N_VPWR_c_577_n 0.005209f $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_403 N_A2_M1002_g N_VPWR_c_561_n 0.00983585f $X=5.99 $Y=2.4 $X2=0 $Y2=0
cc_404 N_A2_M1025_g N_VPWR_c_561_n 0.0098824f $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_405 N_A2_M1002_g N_A_762_368#_c_737_n 4.63009e-19 $X=5.99 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A2_M1002_g N_A_762_368#_c_754_n 0.0196074f $X=5.99 $Y=2.4 $X2=0 $Y2=0
cc_407 N_A2_M1025_g N_A_762_368#_c_754_n 0.017111f $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_408 N_A2_c_505_n N_A_762_368#_c_754_n 0.00170114f $X=7.39 $Y=1.48 $X2=0 $Y2=0
cc_409 N_A2_M1025_g N_A_762_368#_c_738_n 8.68874e-19 $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_410 N_A2_M1025_g N_A_762_368#_c_739_n 0.00151912f $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A2_M1002_g N_A_762_368#_c_741_n 2.55042e-19 $X=5.99 $Y=2.4 $X2=0 $Y2=0
cc_412 N_A2_M1002_g N_A_1216_368#_c_802_n 0.00906731f $X=5.99 $Y=2.4 $X2=0 $Y2=0
cc_413 N_A2_M1025_g N_A_1216_368#_c_803_n 0.00900685f $X=7.43 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A2_c_502_n N_VGND_c_830_n 0.00158425f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_415 N_A2_M1008_g N_VGND_c_831_n 0.0145213f $X=5.975 $Y=0.92 $X2=0 $Y2=0
cc_416 N_A2_c_501_n N_VGND_c_831_n 0.0134054f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_417 N_A2_c_502_n N_VGND_c_831_n 0.0024927f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_418 N_A2_c_501_n N_VGND_c_832_n 0.0185349f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_419 N_A2_c_501_n N_VGND_c_833_n 0.029736f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_420 A2 N_VGND_c_833_n 0.0250425f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_421 N_A2_c_502_n N_VGND_c_838_n 0.0048178f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_422 N_A2_c_501_n N_VGND_c_842_n 0.0138662f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_423 A2 N_VGND_c_842_n 0.0386817f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_424 N_A2_c_501_n N_VGND_c_843_n 0.0400235f $X=7.26 $Y=0.185 $X2=0 $Y2=0
cc_425 N_A2_c_502_n N_VGND_c_843_n 0.00839621f $X=6.05 $Y=0.185 $X2=0 $Y2=0
cc_426 A2 N_VGND_c_843_n 0.0254788f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_427 N_A2_M1008_g N_A_523_124#_c_955_n 0.0169048f $X=5.975 $Y=0.92 $X2=0 $Y2=0
cc_428 N_A2_c_499_n N_A_523_124#_c_955_n 0.00139614f $X=5.99 $Y=1.405 $X2=0
+ $Y2=0
cc_429 N_A2_M1008_g N_A_523_124#_c_956_n 5.60436e-19 $X=5.975 $Y=0.92 $X2=0
+ $Y2=0
cc_430 N_A2_c_501_n N_A_523_124#_c_956_n 0.00460834f $X=7.26 $Y=0.185 $X2=0
+ $Y2=0
cc_431 N_A2_M1022_g N_A_523_124#_c_957_n 0.0170722f $X=7.335 $Y=0.935 $X2=0
+ $Y2=0
cc_432 N_A2_c_505_n N_A_523_124#_c_957_n 0.00475534f $X=7.39 $Y=1.48 $X2=0 $Y2=0
cc_433 A2 N_A_523_124#_c_957_n 0.00203938f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_434 N_A2_c_501_n N_A_523_124#_c_1008_n 0.00157463f $X=7.26 $Y=0.185 $X2=0
+ $Y2=0
cc_435 N_A2_M1022_g N_A_523_124#_c_1008_n 0.0083412f $X=7.335 $Y=0.935 $X2=0
+ $Y2=0
cc_436 A2 N_A_523_124#_c_1008_n 0.0166591f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_437 N_VPWR_M1003_s N_X_c_663_n 0.00459755f $X=0.465 $Y=1.84 $X2=0 $Y2=0
cc_438 N_VPWR_c_562_n N_X_c_663_n 0.0131801f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_439 N_VPWR_c_562_n N_X_c_664_n 0.0293f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_440 N_VPWR_c_563_n N_X_c_664_n 0.0293f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_441 N_VPWR_c_569_n N_X_c_664_n 0.0144623f $X=1.425 $Y=3.33 $X2=0 $Y2=0
cc_442 N_VPWR_c_561_n N_X_c_664_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_443 N_VPWR_M1006_s N_X_c_665_n 0.00165831f $X=1.375 $Y=1.84 $X2=0 $Y2=0
cc_444 N_VPWR_c_563_n N_X_c_665_n 0.0126919f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_445 N_VPWR_c_563_n N_X_c_666_n 0.0293f $X=1.51 $Y=2.275 $X2=0 $Y2=0
cc_446 N_VPWR_c_564_n N_X_c_666_n 0.0349062f $X=2.41 $Y=2.075 $X2=0 $Y2=0
cc_447 N_VPWR_c_571_n N_X_c_666_n 0.0144623f $X=2.325 $Y=3.33 $X2=0 $Y2=0
cc_448 N_VPWR_c_561_n N_X_c_666_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_449 N_VPWR_c_562_n X 0.0590724f $X=0.61 $Y=2.275 $X2=0 $Y2=0
cc_450 N_VPWR_c_567_n X 0.00745548f $X=0.525 $Y=3.33 $X2=0 $Y2=0
cc_451 N_VPWR_c_561_n X 0.00794958f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_452 N_VPWR_M1001_s N_A_762_368#_c_754_n 0.00392167f $X=6.53 $Y=1.84 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_577_n N_A_762_368#_c_739_n 0.0146357f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_561_n N_A_762_368#_c_739_n 0.0121141f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_565_n N_A_762_368#_c_740_n 0.0455071f $X=3.395 $Y=2.54 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_575_n N_A_762_368#_c_740_n 0.0110778f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_561_n N_A_762_368#_c_740_n 0.00916405f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_575_n N_A_762_368#_c_741_n 0.00749631f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_561_n N_A_762_368#_c_741_n 0.0062048f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_575_n N_A_854_368#_c_788_n 0.0513994f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_561_n N_A_854_368#_c_788_n 0.042767f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_462 N_VPWR_M1001_s N_A_1216_368#_c_804_n 0.00415741f $X=6.53 $Y=1.84 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_566_n N_A_1216_368#_c_804_n 0.0166568f $X=6.685 $Y=2.815 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_566_n N_A_1216_368#_c_802_n 0.0115634f $X=6.685 $Y=2.815 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_575_n N_A_1216_368#_c_802_n 0.0144776f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_561_n N_A_1216_368#_c_802_n 0.0118404f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_566_n N_A_1216_368#_c_803_n 0.0129302f $X=6.685 $Y=2.815 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_577_n N_A_1216_368#_c_803_n 0.0145644f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_561_n N_A_1216_368#_c_803_n 0.0119803f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_470 N_X_c_673_n N_VGND_M1010_s 0.00672868f $X=0.675 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_471 N_X_c_659_n N_VGND_M1010_s 0.00204758f $X=0.295 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_472 N_X_c_683_n N_VGND_M1017_s 0.00463478f $X=1.605 $Y=1.015 $X2=0 $Y2=0
cc_473 N_X_c_673_n N_VGND_c_826_n 0.0160725f $X=0.675 $Y=1.015 $X2=0 $Y2=0
cc_474 N_X_c_659_n N_VGND_c_826_n 0.0107964f $X=0.295 $Y=1.015 $X2=0 $Y2=0
cc_475 N_X_c_660_n N_VGND_c_826_n 0.0155339f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_476 N_X_c_660_n N_VGND_c_827_n 0.0154229f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_477 N_X_c_683_n N_VGND_c_827_n 0.0210288f $X=1.605 $Y=1.015 $X2=0 $Y2=0
cc_478 N_X_c_661_n N_VGND_c_827_n 0.0155339f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_479 N_X_c_661_n N_VGND_c_828_n 0.0215159f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_480 N_X_c_660_n N_VGND_c_840_n 0.0109942f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_481 N_X_c_661_n N_VGND_c_841_n 0.0109942f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_482 N_X_c_660_n N_VGND_c_843_n 0.00904371f $X=0.84 $Y=0.515 $X2=0 $Y2=0
cc_483 N_X_c_661_n N_VGND_c_843_n 0.00904371f $X=1.77 $Y=0.515 $X2=0 $Y2=0
cc_484 N_A_762_368#_c_743_n N_A_854_368#_M1015_d 0.00332471f $X=5.68 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_485 N_A_762_368#_c_743_n N_A_854_368#_M1021_s 0.00761462f $X=5.68 $Y=2.375
+ $X2=0 $Y2=0
cc_486 N_A_762_368#_c_743_n N_A_854_368#_c_788_n 0.0666831f $X=5.68 $Y=2.375
+ $X2=0 $Y2=0
cc_487 N_A_762_368#_c_740_n N_A_854_368#_c_788_n 0.0135043f $X=3.955 $Y=2.455
+ $X2=0 $Y2=0
cc_488 N_A_762_368#_c_741_n N_A_854_368#_c_788_n 0.0134678f $X=5.765 $Y=2.4
+ $X2=0 $Y2=0
cc_489 N_A_762_368#_c_754_n N_A_1216_368#_M1002_s 0.00761058f $X=7.54 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_490 N_A_762_368#_c_754_n N_A_1216_368#_M1026_d 0.0095173f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_491 N_A_762_368#_c_754_n N_A_1216_368#_c_804_n 0.0365359f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_492 N_A_762_368#_c_754_n N_A_1216_368#_c_802_n 0.0171986f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_493 N_A_762_368#_c_741_n N_A_1216_368#_c_802_n 0.0177362f $X=5.765 $Y=2.4
+ $X2=0 $Y2=0
cc_494 N_A_762_368#_c_754_n N_A_1216_368#_c_803_n 0.0190257f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_495 N_A_762_368#_c_739_n N_A_1216_368#_c_803_n 0.0202646f $X=7.705 $Y=2.4
+ $X2=0 $Y2=0
cc_496 N_A_762_368#_c_754_n N_A_523_124#_c_957_n 0.00281217f $X=7.54 $Y=2.035
+ $X2=0 $Y2=0
cc_497 N_A_762_368#_c_738_n N_A_523_124#_c_957_n 0.00391062f $X=7.705 $Y=2.12
+ $X2=0 $Y2=0
cc_498 N_A_762_368#_c_737_n N_A_523_124#_c_959_n 0.00667642f $X=5.765 $Y=2.12
+ $X2=0 $Y2=0
cc_499 N_VGND_c_828_n N_A_523_124#_c_946_n 0.0336756f $X=2.2 $Y=0.515 $X2=0
+ $Y2=0
cc_500 N_VGND_c_834_n N_A_523_124#_c_947_n 0.0504256f $X=4.375 $Y=0 $X2=0 $Y2=0
cc_501 N_VGND_c_843_n N_A_523_124#_c_947_n 0.0295559f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_c_828_n N_A_523_124#_c_948_n 0.0121618f $X=2.2 $Y=0.515 $X2=0
+ $Y2=0
cc_503 N_VGND_c_834_n N_A_523_124#_c_948_n 0.0229068f $X=4.375 $Y=0 $X2=0 $Y2=0
cc_504 N_VGND_c_843_n N_A_523_124#_c_948_n 0.0127944f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_505 N_VGND_c_829_n N_A_523_124#_c_949_n 0.00647753f $X=4.46 $Y=0.75 $X2=0
+ $Y2=0
cc_506 N_VGND_M1004_s N_A_523_124#_c_950_n 0.0143195f $X=4 $Y=0.62 $X2=0 $Y2=0
cc_507 N_VGND_c_829_n N_A_523_124#_c_950_n 0.0135869f $X=4.46 $Y=0.75 $X2=0
+ $Y2=0
cc_508 N_VGND_c_829_n N_A_523_124#_c_952_n 0.0121933f $X=4.46 $Y=0.75 $X2=0
+ $Y2=0
cc_509 N_VGND_c_830_n N_A_523_124#_c_952_n 0.0127348f $X=5.32 $Y=0.745 $X2=0
+ $Y2=0
cc_510 N_VGND_c_836_n N_A_523_124#_c_952_n 0.00558557f $X=5.155 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_843_n N_A_523_124#_c_952_n 0.0068223f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_M1027_s N_A_523_124#_c_953_n 0.00176461f $X=5.18 $Y=0.6 $X2=0
+ $Y2=0
cc_513 N_VGND_c_830_n N_A_523_124#_c_953_n 0.0170777f $X=5.32 $Y=0.745 $X2=0
+ $Y2=0
cc_514 N_VGND_c_830_n N_A_523_124#_c_954_n 0.0126994f $X=5.32 $Y=0.745 $X2=0
+ $Y2=0
cc_515 N_VGND_c_831_n N_A_523_124#_c_954_n 0.0120275f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_516 N_VGND_c_838_n N_A_523_124#_c_954_n 0.00405637f $X=6.025 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_843_n N_A_523_124#_c_954_n 0.00562174f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_M1008_s N_A_523_124#_c_955_n 0.00176461f $X=6.05 $Y=0.6 $X2=0
+ $Y2=0
cc_519 N_VGND_c_831_n N_A_523_124#_c_955_n 0.0152916f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_520 N_VGND_c_831_n N_A_523_124#_c_956_n 0.0120629f $X=6.19 $Y=0.745 $X2=0
+ $Y2=0
cc_521 N_VGND_c_832_n N_A_523_124#_c_956_n 0.00558247f $X=6.885 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_833_n N_A_523_124#_c_956_n 0.0120629f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
cc_523 N_VGND_c_843_n N_A_523_124#_c_956_n 0.00681968f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_M1013_s N_A_523_124#_c_957_n 0.00996523f $X=6.91 $Y=0.6 $X2=0
+ $Y2=0
cc_525 N_VGND_c_833_n N_A_523_124#_c_957_n 0.015373f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0
cc_526 N_VGND_c_833_n N_A_523_124#_c_1008_n 0.0130127f $X=7.05 $Y=0.745 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__dlrtp_4.pex.spice
* Created: Wed Sep  2 12:05:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRTP_4%D 3 7 9 12 13
c29 3 0 1.88806e-19 $X=0.505 $Y=2.39
r30 12 15 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.78
r31 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.45
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r33 9 13 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r34 7 14 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.495 $Y=0.905
+ $X2=0.495 $Y2=1.45
r35 3 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.505 $Y=2.39
+ $X2=0.505 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%GATE 3 7 9 12
c37 7 0 3.6533e-19 $X=1.19 $Y=0.81
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.615
+ $X2=1.165 $Y2=1.78
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.615
+ $X2=1.165 $Y2=1.45
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.615 $X2=1.165 $Y2=1.615
r41 7 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.19 $Y=0.81 $X2=1.19
+ $Y2=1.45
r42 3 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.125 $Y=2.39
+ $X2=1.125 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%A_243_394# 1 2 9 11 13 14 16 17 18 21 23 24
+ 25 30 32 33 36 37 38 42 49 53 54 55
c147 54 0 1.30138e-19 $X=3.985 $Y=1.39
c148 38 0 5.47968e-20 $X=3.005 $Y=0.34
c149 33 0 1.82632e-19 $X=2.835 $Y=0.855
c150 25 0 1.88806e-19 $X=1.46 $Y=2.075
c151 18 0 2.60199e-19 $X=3.215 $Y=1.765
c152 14 0 1.99356e-19 $X=3.125 $Y=1.84
r153 53 55 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=1.39 $X2=4
+ $Y2=1.225
r154 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.985
+ $Y=1.39 $X2=3.985 $Y2=1.39
r155 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.615 $X2=1.735 $Y2=1.615
r156 46 49 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.545 $Y=1.615
+ $X2=1.735 $Y2=1.615
r157 44 45 13.9266 $w=3.88e-07 $l=3.45e-07 $layer=LI1_cond $X=1.435 $Y=0.855
+ $X2=1.435 $Y2=1.2
r158 42 44 7.97845 $w=3.88e-07 $l=2.7e-07 $layer=LI1_cond $X=1.435 $Y=0.585
+ $X2=1.435 $Y2=0.855
r159 39 55 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.935 $Y=0.425
+ $X2=3.935 $Y2=1.225
r160 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.85 $Y=0.34
+ $X2=3.935 $Y2=0.425
r161 37 38 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.85 $Y=0.34
+ $X2=3.005 $Y2=0.34
r162 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.92 $Y=0.425
+ $X2=3.005 $Y2=0.34
r163 35 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.92 $Y=0.425
+ $X2=2.92 $Y2=0.77
r164 34 44 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.63 $Y=0.855
+ $X2=1.435 $Y2=0.855
r165 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.835 $Y=0.855
+ $X2=2.92 $Y2=0.77
r166 33 34 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=2.835 $Y=0.855
+ $X2=1.63 $Y2=0.855
r167 31 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.78
+ $X2=1.545 $Y2=1.615
r168 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.545 $Y=1.78
+ $X2=1.545 $Y2=1.95
r169 30 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.45
+ $X2=1.545 $Y2=1.615
r170 30 45 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.545 $Y=1.45
+ $X2=1.545 $Y2=1.2
r171 25 32 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.46 $Y=2.075
+ $X2=1.545 $Y2=1.95
r172 25 27 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=2.075
+ $X2=1.375 $Y2=2.075
r173 23 50 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.1 $Y=1.615
+ $X2=1.735 $Y2=1.615
r174 23 24 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.1 $Y=1.615 $X2=2.19
+ $Y2=1.615
r175 19 54 38.7956 $w=3.51e-07 $l=2.56562e-07 $layer=POLY_cond $X=3.7 $Y=1.225
+ $X2=3.887 $Y2=1.39
r176 19 21 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.7 $Y=1.225
+ $X2=3.7 $Y2=0.58
r177 17 54 51.4957 $w=3.51e-07 $l=4.88748e-07 $layer=POLY_cond $X=3.625 $Y=1.765
+ $X2=3.887 $Y2=1.39
r178 17 18 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.625 $Y=1.765
+ $X2=3.215 $Y2=1.765
r179 14 18 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.125 $Y=1.84
+ $X2=3.215 $Y2=1.765
r180 14 16 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.125 $Y=1.84
+ $X2=3.125 $Y2=2.46
r181 11 24 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.205 $Y=1.45
+ $X2=2.19 $Y2=1.615
r182 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.205 $Y=1.45
+ $X2=2.205 $Y2=0.97
r183 7 24 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.78
+ $X2=2.19 $Y2=1.615
r184 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=2.19 $Y=1.78 $X2=2.19
+ $Y2=2.38
r185 2 27 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.97 $X2=1.375 $Y2=2.115
r186 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.265
+ $Y=0.44 $X2=1.405 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%A_27_126# 1 2 9 13 17 19 20 22 23 26 28 31
+ 32
c91 31 0 1.08744e-19 $X=2.66 $Y=1.635
c92 26 0 4.0055e-19 $X=2.58 $Y=2.37
c93 13 0 1.75109e-19 $X=2.735 $Y=2.46
c94 9 0 1.68329e-19 $X=2.72 $Y=0.69
r95 32 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.635
+ $X2=2.66 $Y2=1.8
r96 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.635
+ $X2=2.66 $Y2=1.47
r97 31 34 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.635
+ $X2=2.64 $Y2=1.8
r98 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.635 $X2=2.66 $Y2=1.635
r99 28 29 6.86755 $w=6.04e-07 $l=3.4e-07 $layer=LI1_cond $X=0.485 $Y=2.115
+ $X2=0.485 $Y2=2.455
r100 26 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.58 $Y=2.37
+ $X2=2.58 $Y2=1.8
r101 24 29 8.35964 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.855 $Y=2.455
+ $X2=0.485 $Y2=2.455
r102 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.495 $Y=2.455
+ $X2=2.58 $Y2=2.37
r103 23 24 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=2.495 $Y=2.455
+ $X2=0.855 $Y2=2.455
r104 22 28 10.3858 $w=6.04e-07 $l=3.5812e-07 $layer=LI1_cond $X=0.77 $Y=1.95
+ $X2=0.485 $Y2=2.115
r105 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.77 $Y=1.28
+ $X2=0.77 $Y2=1.95
r106 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.77 $Y2=1.28
r107 19 20 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.445 $Y2=1.195
r108 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.445 $Y2=1.195
r109 15 17 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.28 $Y2=0.905
r110 13 37 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=1.8
r111 9 36 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.72 $Y=0.69
+ $X2=2.72 $Y2=1.47
r112 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.97 $X2=0.28 $Y2=2.115
r113 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.63 $X2=0.28 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%A_364_120# 1 2 9 12 15 16 17 19 21 22 23 26
+ 27 36 40 46 49
c109 36 0 1.75109e-19 $X=2.155 $Y=2.11
c110 26 0 1.30138e-19 $X=3.82 $Y=2.215
c111 21 0 1.67587e-19 $X=3.04 $Y=1.97
c112 17 0 1.82698e-19 $X=2.24 $Y=1.195
c113 12 0 9.02322e-20 $X=3.66 $Y=2.75
r114 46 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.285
+ $X2=3.2 $Y2=1.12
r115 45 47 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.147 $Y=1.285
+ $X2=3.147 $Y2=1.45
r116 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.285 $X2=3.2 $Y2=1.285
r117 38 40 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.93 $Y=2.055
+ $X2=3.04 $Y2=2.055
r118 34 36 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=1.965 $Y=2.11
+ $X2=2.155 $Y2=2.11
r119 30 32 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.975 $Y=1.195
+ $X2=2.155 $Y2=1.195
r120 27 51 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.82 $Y=2.215
+ $X2=3.66 $Y2=2.215
r121 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.82
+ $Y=2.215 $X2=3.82 $Y2=2.215
r122 24 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.82 $Y=2.905
+ $X2=3.82 $Y2=2.215
r123 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.655 $Y=2.99
+ $X2=3.82 $Y2=2.905
r124 22 23 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.655 $Y=2.99
+ $X2=3.015 $Y2=2.99
r125 21 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=1.97
+ $X2=3.04 $Y2=2.055
r126 21 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.04 $Y=1.97
+ $X2=3.04 $Y2=1.45
r127 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.93 $Y=2.905
+ $X2=3.015 $Y2=2.99
r128 18 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=2.14
+ $X2=2.93 $Y2=2.055
r129 18 19 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.93 $Y=2.14
+ $X2=2.93 $Y2=2.905
r130 17 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=1.195
+ $X2=2.155 $Y2=1.195
r131 16 45 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=3.147 $Y=1.195
+ $X2=3.147 $Y2=1.285
r132 16 17 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.955 $Y=1.195
+ $X2=2.24 $Y2=1.195
r133 15 36 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.155 $Y=2.02
+ $X2=2.155 $Y2=2.11
r134 14 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.28
+ $X2=2.155 $Y2=1.195
r135 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.155 $Y=1.28
+ $X2=2.155 $Y2=2.02
r136 10 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=2.38
+ $X2=3.66 $Y2=2.215
r137 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.66 $Y=2.38
+ $X2=3.66 $Y2=2.75
r138 9 49 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.125 $Y=0.69
+ $X2=3.125 $Y2=1.12
r139 2 34 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=1.96 $X2=1.965 $Y2=2.11
r140 1 30 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.6 $X2=1.975 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%A_797_48# 1 2 3 10 12 13 14 17 23 27 31 35
+ 39 43 47 51 53 56 59 63 64 68 77 86 89 90 91 92 94 104
c197 53 0 1.98009e-19 $X=5.11 $Y=2.272
c198 14 0 7.47035e-20 $X=4.135 $Y=0.94
r199 101 102 31.7304 $w=3.19e-07 $l=2.1e-07 $layer=POLY_cond $X=7.985 $Y=1.465
+ $X2=8.195 $Y2=1.465
r200 100 101 33.2414 $w=3.19e-07 $l=2.2e-07 $layer=POLY_cond $X=7.765 $Y=1.465
+ $X2=7.985 $Y2=1.465
r201 99 100 42.3072 $w=3.19e-07 $l=2.8e-07 $layer=POLY_cond $X=7.485 $Y=1.465
+ $X2=7.765 $Y2=1.465
r202 96 97 45.3292 $w=3.19e-07 $l=3e-07 $layer=POLY_cond $X=7.035 $Y=1.465
+ $X2=7.335 $Y2=1.465
r203 91 92 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.765 $Y=1.545
+ $X2=6.935 $Y2=1.545
r204 86 88 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=0.785
+ $X2=5.27 $Y2=0.95
r205 78 104 11.3323 $w=3.19e-07 $l=7.5e-08 $layer=POLY_cond $X=8.43 $Y=1.465
+ $X2=8.505 $Y2=1.465
r206 78 102 35.5078 $w=3.19e-07 $l=2.35e-07 $layer=POLY_cond $X=8.43 $Y=1.465
+ $X2=8.195 $Y2=1.465
r207 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.43
+ $Y=1.465 $X2=8.43 $Y2=1.465
r208 75 99 11.3323 $w=3.19e-07 $l=7.5e-08 $layer=POLY_cond $X=7.41 $Y=1.465
+ $X2=7.485 $Y2=1.465
r209 75 97 11.3323 $w=3.19e-07 $l=7.5e-08 $layer=POLY_cond $X=7.41 $Y=1.465
+ $X2=7.335 $Y2=1.465
r210 74 77 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=7.41 $Y=1.465
+ $X2=8.43 $Y2=1.465
r211 74 92 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=7.41 $Y=1.465
+ $X2=6.935 $Y2=1.465
r212 74 75 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.41
+ $Y=1.465 $X2=7.41 $Y2=1.465
r213 71 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.44 $Y=1.705
+ $X2=6.275 $Y2=1.705
r214 71 91 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.44 $Y=1.705
+ $X2=6.765 $Y2=1.705
r215 66 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=1.79
+ $X2=6.275 $Y2=1.705
r216 66 68 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.275 $Y=1.79
+ $X2=6.275 $Y2=1.985
r217 65 89 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.44 $Y=1.705
+ $X2=5.315 $Y2=1.705
r218 64 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.11 $Y=1.705
+ $X2=6.275 $Y2=1.705
r219 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.11 $Y=1.705
+ $X2=5.44 $Y2=1.705
r220 63 81 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=5.315 $Y=1.965
+ $X2=5.315 $Y2=2.065
r221 60 89 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=1.79
+ $X2=5.315 $Y2=1.705
r222 60 63 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=5.315 $Y=1.79
+ $X2=5.315 $Y2=1.965
r223 59 89 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.275 $Y=1.62
+ $X2=5.315 $Y2=1.705
r224 59 88 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.275 $Y=1.62
+ $X2=5.275 $Y2=0.95
r225 56 95 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=2.215
+ $X2=4.36 $Y2=2.38
r226 56 94 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=2.215
+ $X2=4.36 $Y2=2.05
r227 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=2.215 $X2=4.36 $Y2=2.215
r228 53 83 9.18462 $w=3.28e-07 $l=2.63e-07 $layer=LI1_cond $X=5.275 $Y=2.272
+ $X2=5.275 $Y2=2.535
r229 53 81 7.93363 $w=3.28e-07 $l=2.07e-07 $layer=LI1_cond $X=5.275 $Y=2.272
+ $X2=5.275 $Y2=2.065
r230 53 55 20.8273 $w=4.13e-07 $l=7.5e-07 $layer=LI1_cond $X=5.11 $Y=2.272
+ $X2=4.36 $Y2=2.272
r231 49 104 18.1317 $w=3.19e-07 $l=2.16852e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.505 $Y2=1.465
r232 49 51 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=0.74
r233 45 104 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.505 $Y=1.63
+ $X2=8.505 $Y2=1.465
r234 45 47 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.505 $Y=1.63
+ $X2=8.505 $Y2=2.4
r235 41 102 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=1.465
r236 41 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=0.74
r237 37 101 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.985 $Y=1.63
+ $X2=7.985 $Y2=1.465
r238 37 39 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.985 $Y=1.63
+ $X2=7.985 $Y2=2.4
r239 33 100 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=1.465
r240 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=0.74
r241 29 99 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.485 $Y=1.63
+ $X2=7.485 $Y2=1.465
r242 29 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.485 $Y=1.63
+ $X2=7.485 $Y2=2.4
r243 25 97 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.335 $Y=1.3
+ $X2=7.335 $Y2=1.465
r244 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.335 $Y=1.3
+ $X2=7.335 $Y2=0.74
r245 21 96 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.035 $Y=1.63
+ $X2=7.035 $Y2=1.465
r246 21 23 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.035 $Y=1.63
+ $X2=7.035 $Y2=2.4
r247 19 94 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=4.435 $Y=1.015
+ $X2=4.435 $Y2=2.05
r248 17 95 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.285 $Y=2.75
+ $X2=4.285 $Y2=2.38
r249 13 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.36 $Y=0.94
+ $X2=4.435 $Y2=1.015
r250 13 14 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.36 $Y=0.94
+ $X2=4.135 $Y2=0.94
r251 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.06 $Y=0.865
+ $X2=4.135 $Y2=0.94
r252 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.06 $Y=0.865
+ $X2=4.06 $Y2=0.58
r253 3 68 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=6.09
+ $Y=1.84 $X2=6.275 $Y2=1.985
r254 2 83 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=1.84 $X2=5.275 $Y2=2.535
r255 2 63 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=1.84 $X2=5.275 $Y2=1.965
r256 1 86 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.37 $X2=5.265 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%A_640_74# 1 2 9 13 15 19 23 25 27 34 35 36
+ 39 43 44 52
c109 44 0 4.97389e-20 $X=3.325 $Y=2.405
c110 34 0 7.47035e-20 $X=3.595 $Y=1.725
c111 27 0 1.68329e-19 $X=3.51 $Y=0.76
c112 23 0 1.07777e-19 $X=5.5 $Y=2.26
r113 51 52 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.05 $Y=1.515
+ $X2=5.14 $Y2=1.515
r114 46 48 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.38 $Y=1.81
+ $X2=3.595 $Y2=1.81
r115 43 44 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=2.57
+ $X2=3.325 $Y2=2.405
r116 40 51 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.885 $Y=1.515
+ $X2=5.05 $Y2=1.515
r117 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.885
+ $Y=1.515 $X2=4.885 $Y2=1.515
r118 37 39 8.0671 $w=2.98e-07 $l=2.1e-07 $layer=LI1_cond $X=4.87 $Y=1.725
+ $X2=4.87 $Y2=1.515
r119 36 48 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.81
+ $X2=3.595 $Y2=1.81
r120 35 37 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.72 $Y=1.81
+ $X2=4.87 $Y2=1.725
r121 35 36 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.72 $Y=1.81
+ $X2=3.68 $Y2=1.81
r122 34 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=1.725
+ $X2=3.595 $Y2=1.81
r123 33 34 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.595 $Y=0.925
+ $X2=3.595 $Y2=1.725
r124 31 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=1.895
+ $X2=3.38 $Y2=1.81
r125 31 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.38 $Y=1.895
+ $X2=3.38 $Y2=2.405
r126 27 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.51 $Y=0.76
+ $X2=3.595 $Y2=0.925
r127 27 29 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.51 $Y=0.76
+ $X2=3.37 $Y2=0.76
r128 25 26 89.6095 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=5.5 $Y=1.425
+ $X2=5.5 $Y2=1.2
r129 21 25 29.1532 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.5 $Y=1.5 $X2=5.5
+ $Y2=1.425
r130 21 23 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=5.5 $Y=1.5 $X2=5.5
+ $Y2=2.26
r131 19 26 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.485 $Y=0.69
+ $X2=5.485 $Y2=1.2
r132 15 25 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.41 $Y=1.425 $X2=5.5
+ $Y2=1.425
r133 15 52 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.41 $Y=1.425
+ $X2=5.14 $Y2=1.425
r134 11 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.35
+ $X2=5.05 $Y2=1.515
r135 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.35
+ $X2=5.05 $Y2=0.69
r136 7 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.68
+ $X2=5.05 $Y2=1.515
r137 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=5.05 $Y=1.68 $X2=5.05
+ $Y2=2.26
r138 2 43 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.96 $X2=3.35 $Y2=2.57
r139 1 29 182 $w=1.7e-07 $l=4.67333e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.37 $X2=3.37 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%RESET_B 1 3 6 8 10 13 15 16 26
c57 26 0 3.8972e-20 $X=6.5 $Y=1.285
r58 24 26 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.39 $Y=1.285
+ $X2=6.5 $Y2=1.285
r59 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.39
+ $Y=1.285 $X2=6.39 $Y2=1.285
r60 22 24 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.345 $Y=1.285
+ $X2=6.39 $Y2=1.285
r61 21 22 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=6 $Y=1.285
+ $X2=6.345 $Y2=1.285
r62 19 21 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.915 $Y=1.285 $X2=6
+ $Y2=1.285
r63 16 25 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.48 $Y=1.285 $X2=6.39
+ $Y2=1.285
r64 15 25 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6 $Y=1.285 $X2=6.39
+ $Y2=1.285
r65 11 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=1.285
r66 11 13 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=2.26
r67 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.12
+ $X2=6.345 $Y2=1.285
r68 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.345 $Y=1.12
+ $X2=6.345 $Y2=0.69
r69 4 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6 $Y=1.45 $X2=6
+ $Y2=1.285
r70 4 6 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=6 $Y=1.45 $X2=6
+ $Y2=2.26
r71 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.12
+ $X2=5.915 $Y2=1.285
r72 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.915 $Y=1.12
+ $X2=5.915 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%VPWR 1 2 3 4 5 6 7 26 30 34 38 42 48 50 52
+ 55 56 58 59 61 62 63 65 73 88 93 96 99 103
r113 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 91 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r118 88 102 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.857 $Y2=3.33
r119 88 90 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.4 $Y2=3.33
r120 87 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r125 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 78 99 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.625 $Y2=3.33
r127 78 80 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 77 97 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 74 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=2.5 $Y2=3.33
r131 74 76 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 73 99 12.0744 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.625 $Y2=3.33
r133 73 76 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 72 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r139 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 66 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r141 66 68 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 65 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.5 $Y2=3.33
r143 65 71 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.16 $Y2=3.33
r144 63 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r145 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r146 63 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r147 61 86 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.44 $Y2=3.33
r148 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.76 $Y2=3.33
r149 60 90 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=8.4 $Y2=3.33
r150 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=7.76 $Y2=3.33
r151 58 83 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.81 $Y2=3.33
r153 57 86 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=6.81 $Y2=3.33
r155 55 80 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.61 $Y=3.33 $X2=5.52
+ $Y2=3.33
r156 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=3.33
+ $X2=5.775 $Y2=3.33
r157 54 83 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=6.48 $Y2=3.33
r158 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=5.775 $Y2=3.33
r159 50 102 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.857 $Y2=3.33
r160 50 52 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.76 $Y2=2.225
r161 46 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=3.245
+ $X2=7.76 $Y2=3.33
r162 46 48 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=7.76 $Y=3.245
+ $X2=7.76 $Y2=2.225
r163 42 45 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.81 $Y=2.045
+ $X2=6.81 $Y2=2.815
r164 40 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=3.245
+ $X2=6.81 $Y2=3.33
r165 40 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.81 $Y=3.245
+ $X2=6.81 $Y2=2.815
r166 36 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=3.245
+ $X2=5.775 $Y2=3.33
r167 36 38 41.034 $w=3.28e-07 $l=1.175e-06 $layer=LI1_cond $X=5.775 $Y=3.245
+ $X2=5.775 $Y2=2.07
r168 32 99 2.35715 $w=5.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r169 32 34 9.18417 $w=5.58e-07 $l=4.3e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.815
r170 28 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=3.245 $X2=2.5
+ $Y2=3.33
r171 28 30 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.5 $Y=3.245
+ $X2=2.5 $Y2=2.805
r172 24 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r173 24 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.875
r174 7 52 300 $w=1.7e-07 $l=4.60163e-07 $layer=licon1_PDIFF $count=2 $X=8.595
+ $Y=1.84 $X2=8.76 $Y2=2.225
r175 6 48 300 $w=1.7e-07 $l=4.68455e-07 $layer=licon1_PDIFF $count=2 $X=7.575
+ $Y=1.84 $X2=7.76 $Y2=2.225
r176 5 45 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=6.59
+ $Y=1.84 $X2=6.81 $Y2=2.815
r177 5 42 300 $w=1.7e-07 $l=3.05778e-07 $layer=licon1_PDIFF $count=2 $X=6.59
+ $Y=1.84 $X2=6.81 $Y2=2.045
r178 4 38 300 $w=1.7e-07 $l=3.0895e-07 $layer=licon1_PDIFF $count=2 $X=5.59
+ $Y=1.84 $X2=5.775 $Y2=2.07
r179 3 34 600 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=2.54 $X2=4.625 $Y2=2.815
r180 2 30 600 $w=1.7e-07 $l=9.48644e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.96 $X2=2.5 $Y2=2.805
r181 1 26 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.97 $X2=0.815 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%Q 1 2 3 4 15 19 21 23 24 25 29 35 37 39 43
+ 45 48 49
r76 48 49 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.665
r77 47 49 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.88 $Y=1.8
+ $X2=8.88 $Y2=1.665
r78 46 48 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=1.13
+ $X2=8.88 $Y2=1.295
r79 40 45 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=8.505 $Y=1.005
+ $X2=8.41 $Y2=1.005
r80 39 46 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=8.765 $Y=1.005
+ $X2=8.88 $Y2=1.13
r81 39 40 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=8.765 $Y=1.005
+ $X2=8.505 $Y2=1.005
r82 38 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.425 $Y=1.885
+ $X2=8.26 $Y2=1.885
r83 37 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.765 $Y=1.885
+ $X2=8.88 $Y2=1.8
r84 37 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.765 $Y=1.885
+ $X2=8.425 $Y2=1.885
r85 33 45 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=8.41 $Y=0.88
+ $X2=8.41 $Y2=1.005
r86 33 35 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=8.41 $Y=0.88
+ $X2=8.41 $Y2=0.53
r87 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.26 $Y=1.985
+ $X2=8.26 $Y2=2.815
r88 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.26 $Y=1.97 $X2=8.26
+ $Y2=1.885
r89 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.26 $Y=1.97
+ $X2=8.26 $Y2=1.985
r90 26 42 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=7.645 $Y=1.005
+ $X2=7.515 $Y2=1.005
r91 25 45 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=8.315 $Y=1.005
+ $X2=8.41 $Y2=1.005
r92 25 26 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=8.315 $Y=1.005
+ $X2=7.645 $Y2=1.005
r93 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=1.885
+ $X2=8.26 $Y2=1.885
r94 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.095 $Y=1.885
+ $X2=7.425 $Y2=1.885
r95 19 42 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=0.88
+ $X2=7.515 $Y2=1.005
r96 19 21 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=7.515 $Y=0.88
+ $X2=7.515 $Y2=0.53
r97 15 17 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.3 $Y=1.985 $X2=7.3
+ $Y2=2.815
r98 13 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.3 $Y=1.97
+ $X2=7.425 $Y2=1.885
r99 13 15 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=7.3 $Y=1.97 $X2=7.3
+ $Y2=1.985
r100 4 31 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=8.075
+ $Y=1.84 $X2=8.26 $Y2=2.815
r101 4 29 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=8.075
+ $Y=1.84 $X2=8.26 $Y2=1.985
r102 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.125
+ $Y=1.84 $X2=7.26 $Y2=2.815
r103 3 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.125
+ $Y=1.84 $X2=7.26 $Y2=1.985
r104 2 45 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.965
r105 2 35 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.53
r106 1 42 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.37 $X2=7.55 $Y2=0.965
r107 1 21 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.37 $X2=7.55 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%VGND 1 2 3 4 5 6 7 26 30 34 38 40 44 48 50
+ 52 55 56 57 59 71 75 80 86 89 92 95 98 102
c122 44 0 3.8972e-20 $X=7.12 $Y=0.53
r123 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r124 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r125 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r126 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r127 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r128 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r129 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r130 84 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r131 84 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r132 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r133 81 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.145 $Y=0 $X2=7.98
+ $Y2=0
r134 81 83 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.145 $Y=0 $X2=8.4
+ $Y2=0
r135 80 101 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r136 80 83 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r137 79 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r138 79 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r139 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r140 76 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.215 $Y=0 $X2=7.085
+ $Y2=0
r141 76 78 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.215 $Y=0
+ $X2=7.44 $Y2=0
r142 75 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=0 $X2=7.98
+ $Y2=0
r143 75 78 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.815 $Y=0
+ $X2=7.44 $Y2=0
r144 71 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=0 $X2=6.13
+ $Y2=0
r145 71 73 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=4.56 $Y2=0
r146 70 90 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r147 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r148 67 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=0 $X2=2.5
+ $Y2=0
r149 67 69 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.665 $Y=0
+ $X2=4.08 $Y2=0
r150 66 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r151 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r152 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r153 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r154 62 65 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r155 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r156 60 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.845
+ $Y2=0
r157 60 62 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.2
+ $Y2=0
r158 59 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.5
+ $Y2=0
r159 59 65 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=0
+ $X2=2.16 $Y2=0
r160 57 93 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r161 57 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r162 57 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r163 55 69 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.08
+ $Y2=0
r164 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.315
+ $Y2=0
r165 54 73 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.56
+ $Y2=0
r166 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.315
+ $Y2=0
r167 50 101 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.897 $Y2=0
r168 50 52 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.84 $Y2=0.53
r169 46 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0
r170 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0.53
r171 42 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.085 $Y=0.085
+ $X2=7.085 $Y2=0
r172 42 44 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=7.085 $Y=0.085
+ $X2=7.085 $Y2=0.53
r173 41 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r174 40 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.955 $Y=0 $X2=7.085
+ $Y2=0
r175 40 41 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.955 $Y=0
+ $X2=6.295 $Y2=0
r176 36 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0
r177 36 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0.515
r178 32 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=0.085
+ $X2=4.315 $Y2=0
r179 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.315 $Y=0.085
+ $X2=4.315 $Y2=0.58
r180 28 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=0.085 $X2=2.5
+ $Y2=0
r181 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.5 $Y=0.085
+ $X2=2.5 $Y2=0.515
r182 24 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0
r183 24 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0.775
r184 7 52 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.53
r185 6 48 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.84
+ $Y=0.37 $X2=7.98 $Y2=0.53
r186 5 44 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=6.975
+ $Y=0.37 $X2=7.12 $Y2=0.53
r187 4 38 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.37 $X2=6.13 $Y2=0.515
r188 3 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.135
+ $Y=0.37 $X2=4.275 $Y2=0.58
r189 2 30 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.6 $X2=2.5 $Y2=0.515
r190 1 26 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.63 $X2=0.845 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_4%A_938_74# 1 2 3 12 14 15 17 19 20 22 24
r47 22 29 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=6.595 $Y=0.77 $X2=6.595
+ $Y2=0.86
r48 22 24 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=6.595 $Y=0.77
+ $X2=6.595 $Y2=0.51
r49 21 27 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=5.785 $Y=0.86
+ $X2=5.66 $Y2=0.86
r50 20 29 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=6.465 $Y=0.86
+ $X2=6.595 $Y2=0.86
r51 20 21 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.465 $Y=0.86
+ $X2=5.785 $Y2=0.86
r52 17 27 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.66 $Y=0.77 $X2=5.66
+ $Y2=0.86
r53 17 19 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.66 $Y=0.77
+ $X2=5.66 $Y2=0.495
r54 16 19 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=5.66 $Y=0.45 $X2=5.66
+ $Y2=0.495
r55 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.535 $Y=0.365
+ $X2=5.66 $Y2=0.45
r56 14 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.535 $Y=0.365
+ $X2=5 $Y2=0.365
r57 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.835 $Y=0.45
+ $X2=5 $Y2=0.365
r58 10 12 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=4.835 $Y=0.45
+ $X2=4.835 $Y2=0.515
r59 3 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.42
+ $Y=0.37 $X2=6.56 $Y2=0.86
r60 3 24 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=6.42
+ $Y=0.37 $X2=6.56 $Y2=0.51
r61 2 27 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.37 $X2=5.7 $Y2=0.855
r62 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.37 $X2=5.7 $Y2=0.495
r63 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.69
+ $Y=0.37 $X2=4.835 $Y2=0.515
.ends


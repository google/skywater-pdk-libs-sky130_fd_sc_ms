# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__nand4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.835000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.130000 1.430000 4.140000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 7.555000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.300000 9.015000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.665600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.880000 2.725000 1.090000 ;
        RECT 1.535000 1.090000 4.675000 1.130000 ;
        RECT 2.050000 1.850000 2.680000 1.950000 ;
        RECT 2.050000 1.950000 8.505000 2.120000 ;
        RECT 2.050000 2.120000 2.670000 2.980000 ;
        RECT 2.395000 0.595000 2.725000 0.880000 ;
        RECT 2.395000 1.130000 4.675000 1.260000 ;
        RECT 4.310000 1.820000 4.675000 1.950000 ;
        RECT 4.370000 2.120000 4.590000 2.980000 ;
        RECT 4.445000 1.260000 4.675000 1.820000 ;
        RECT 6.065000 2.120000 6.660000 2.980000 ;
        RECT 8.215000 2.120000 8.505000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  0.770000 0.445000 0.960000 ;
      RECT 0.115000  0.960000 1.335000 1.130000 ;
      RECT 0.505000  1.950000 0.835000 3.245000 ;
      RECT 0.545000  0.085000 0.875000 0.600000 ;
      RECT 1.005000  1.130000 1.335000 1.430000 ;
      RECT 1.005000  1.430000 2.850000 1.680000 ;
      RECT 1.005000  1.680000 1.335000 2.700000 ;
      RECT 1.105000  0.255000 3.075000 0.425000 ;
      RECT 1.105000  0.425000 1.435000 0.710000 ;
      RECT 1.540000  1.850000 1.870000 3.245000 ;
      RECT 1.965000  0.425000 2.215000 0.710000 ;
      RECT 2.850000  2.290000 4.190000 3.245000 ;
      RECT 2.905000  0.425000 3.075000 0.750000 ;
      RECT 2.905000  0.750000 4.875000 0.920000 ;
      RECT 3.255000  0.330000 6.725000 0.580000 ;
      RECT 4.760000  2.290000 5.885000 3.245000 ;
      RECT 5.105000  0.770000 5.435000 0.960000 ;
      RECT 5.105000  0.960000 6.215000 1.010000 ;
      RECT 5.105000  1.010000 9.005000 1.130000 ;
      RECT 5.535000  0.580000 6.725000 0.600000 ;
      RECT 5.605000  0.600000 5.795000 0.710000 ;
      RECT 5.965000  0.770000 6.215000 0.960000 ;
      RECT 5.965000  1.130000 7.170000 1.180000 ;
      RECT 6.395000  0.600000 6.725000 0.840000 ;
      RECT 6.835000  2.290000 8.035000 3.245000 ;
      RECT 6.920000  0.350000 7.100000 0.960000 ;
      RECT 6.920000  0.960000 9.005000 1.010000 ;
      RECT 7.270000  0.085000 7.600000 0.780000 ;
      RECT 7.770000  0.350000 7.960000 0.960000 ;
      RECT 8.130000  0.085000 8.505000 0.780000 ;
      RECT 8.675000  0.350000 9.005000 0.960000 ;
      RECT 8.675000  1.950000 8.955000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_ms__nand4b_4

* File: sky130_fd_sc_ms__dlxbp_1.pex.spice
* Created: Wed Sep  2 12:06:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLXBP_1%D 2 5 9 10 11 14 16
c38 10 0 1.56139e-19 $X=0.587 $Y=1.89
r39 14 16 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.385
+ $X2=0.587 $Y2=1.22
r40 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r41 11 15 2.14223 $w=6.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.555
+ $X2=0.6 $Y2=1.555
r42 9 16 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.5 $Y=0.835 $X2=0.5
+ $Y2=1.22
r43 5 10 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=0.5 $Y=2.485 $X2=0.5
+ $Y2=1.89
r44 2 10 42.7652 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.587 $Y=1.713
+ $X2=0.587 $Y2=1.89
r45 1 14 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.587 $Y=1.397
+ $X2=0.587 $Y2=1.385
r46 1 2 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.587 $Y=1.397
+ $X2=0.587 $Y2=1.713
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%GATE 3 6 8 11 13
c38 13 0 3.53875e-20 $X=1.17 $Y=1.22
c39 8 0 7.84293e-20 $X=1.2 $Y=1.295
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.385
+ $X2=1.17 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.385
+ $X2=1.17 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.385 $X2=1.17 $Y2=1.385
r43 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=1.295 $X2=1.17
+ $Y2=1.385
r44 6 14 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=1.11 $Y=2.485
+ $X2=1.11 $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.08 $Y=0.74 $X2=1.08
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%A_231_74# 1 2 11 15 17 19 20 21 25 28 31 32
+ 34 36 37 39 41 42 45
c132 41 0 6.89381e-20 $X=3.91 $Y=0.345
c133 37 0 7.84293e-20 $X=2.165 $Y=1.635
c134 36 0 8.26417e-20 $X=2.165 $Y=1.635
c135 34 0 1.56139e-19 $X=1.675 $Y=1.68
c136 32 0 3.53875e-20 $X=2.91 $Y=0.665
c137 20 0 1.49705e-19 $X=3.925 $Y=1.765
c138 17 0 1.53417e-19 $X=3.245 $Y=1.84
r139 49 50 14.1693 $w=2.54e-07 $l=2.95e-07 $layer=LI1_cond $X=1.295 $Y=1.72
+ $X2=1.59 $Y2=1.72
r140 47 48 13.7503 $w=5.43e-07 $l=3.45e-07 $layer=LI1_cond $X=1.402 $Y=0.665
+ $X2=1.402 $Y2=1.01
r141 45 47 3.18223 $w=5.43e-07 $l=1.45e-07 $layer=LI1_cond $X=1.402 $Y=0.52
+ $X2=1.402 $Y2=0.665
r142 42 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=0.345
+ $X2=3.91 $Y2=0.51
r143 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=0.345 $X2=3.91 $Y2=0.345
r144 39 53 18.4631 $w=1.68e-07 $l=2.83e-07 $layer=LI1_cond $X=2.995 $Y=0.382
+ $X2=2.995 $Y2=0.665
r145 39 41 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=3.08 $Y=0.382
+ $X2=3.91 $Y2=0.382
r146 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.165
+ $Y=1.635 $X2=2.165 $Y2=1.635
r147 34 50 4.36065 $w=4.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.675 $Y=1.68
+ $X2=1.59 $Y2=1.72
r148 34 36 13.4452 $w=4.18e-07 $l=4.9e-07 $layer=LI1_cond $X=1.675 $Y=1.68
+ $X2=2.165 $Y2=1.68
r149 33 47 7.70116 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=1.675 $Y=0.665
+ $X2=1.402 $Y2=0.665
r150 32 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0.665
+ $X2=2.995 $Y2=0.665
r151 32 33 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.91 $Y=0.665
+ $X2=1.675 $Y2=0.665
r152 31 50 3.08766 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.59 $Y=1.47
+ $X2=1.59 $Y2=1.72
r153 31 48 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.59 $Y=1.47
+ $X2=1.59 $Y2=1.01
r154 26 49 0.813113 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=1.295 $Y=1.89
+ $X2=1.295 $Y2=1.72
r155 26 28 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=1.295 $Y=1.89
+ $X2=1.295 $Y2=2.21
r156 25 58 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4 $Y=0.83 $X2=4
+ $Y2=0.51
r157 23 25 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4 $Y=1.69 $X2=4
+ $Y2=0.83
r158 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.925 $Y=1.765
+ $X2=4 $Y2=1.69
r159 20 21 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.925 $Y=1.765
+ $X2=3.335 $Y2=1.765
r160 17 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.245 $Y=1.84
+ $X2=3.335 $Y2=1.765
r161 17 19 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.245 $Y=1.84
+ $X2=3.245 $Y2=2.46
r162 13 37 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.8
+ $X2=2.24 $Y2=1.635
r163 13 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.24 $Y=1.8
+ $X2=2.24 $Y2=2.38
r164 9 37 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.225 $Y=1.47
+ $X2=2.24 $Y2=1.635
r165 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.225 $Y=1.47
+ $X2=2.225 $Y2=0.78
r166 2 28 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.065 $X2=1.335 $Y2=2.21
r167 1 45 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.295 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%A_27_413# 1 2 9 13 18 19 20 22 23 24 27 28
+ 31 35 36
c96 27 0 8.79278e-21 $X=2.71 $Y=1.635
c97 23 0 1.53417e-19 $X=2.545 $Y=2.145
c98 9 0 8.26417e-20 $X=2.855 $Y=2.46
r99 35 36 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.267 $Y=2.225
+ $X2=0.267 $Y2=2.06
r100 33 36 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.18 $Y=1.05
+ $X2=0.18 $Y2=2.06
r101 31 33 11.4207 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.272 $Y=0.795
+ $X2=0.272 $Y2=1.05
r102 28 39 39.9775 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.635
+ $X2=2.745 $Y2=1.8
r103 28 38 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.635
+ $X2=2.745 $Y2=1.47
r104 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.635 $X2=2.71 $Y2=1.635
r105 25 27 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.71 $Y=2.06
+ $X2=2.71 $Y2=1.635
r106 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.545 $Y=2.145
+ $X2=2.71 $Y2=2.06
r107 23 24 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.545 $Y=2.145
+ $X2=1.76 $Y2=2.145
r108 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.675 $Y=2.23
+ $X2=1.76 $Y2=2.145
r109 21 22 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.675 $Y=2.23
+ $X2=1.675 $Y2=2.545
r110 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.59 $Y=2.63
+ $X2=1.675 $Y2=2.545
r111 19 20 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=1.59 $Y=2.63
+ $X2=0.44 $Y2=2.63
r112 18 20 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.267 $Y=2.545
+ $X2=0.44 $Y2=2.63
r113 17 35 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=0.267 $Y=2.232
+ $X2=0.267 $Y2=2.225
r114 17 18 10.4555 $w=3.43e-07 $l=3.13e-07 $layer=LI1_cond $X=0.267 $Y=2.232
+ $X2=0.267 $Y2=2.545
r115 13 38 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.87 $Y=0.72
+ $X2=2.87 $Y2=1.47
r116 9 39 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.855 $Y=2.46
+ $X2=2.855 $Y2=1.8
r117 2 35 300 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.065 $X2=0.275 $Y2=2.225
r118 1 31 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.56 $X2=0.285 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%A_373_82# 1 2 9 12 14 16 19 20 24 25 28 32
+ 37 41 43 45
c117 41 0 8.79278e-21 $X=3.35 $Y=1.315
c118 37 0 1.49705e-19 $X=3.28 $Y=1.105
r119 41 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.315
+ $X2=3.35 $Y2=1.15
r120 40 42 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=1.315
+ $X2=3.28 $Y2=1.48
r121 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.315 $X2=3.35 $Y2=1.315
r122 37 40 5.34418 $w=4.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.28 $Y=1.105
+ $X2=3.28 $Y2=1.315
r123 32 35 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.525
+ $X2=2.055 $Y2=2.61
r124 28 30 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.01 $Y=1.005
+ $X2=2.01 $Y2=1.105
r125 25 47 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.935 $Y=2.215
+ $X2=3.775 $Y2=2.215
r126 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.935
+ $Y=2.215 $X2=3.935 $Y2=2.215
r127 22 24 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.935 $Y=2.44
+ $X2=3.935 $Y2=2.215
r128 21 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.525
+ $X2=3.13 $Y2=2.525
r129 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.77 $Y=2.525
+ $X2=3.935 $Y2=2.44
r130 20 21 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.77 $Y=2.525
+ $X2=3.215 $Y2=2.525
r131 19 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=2.44
+ $X2=3.13 $Y2=2.525
r132 19 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.13 $Y=2.44
+ $X2=3.13 $Y2=1.48
r133 17 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.18 $Y=2.525
+ $X2=2.055 $Y2=2.525
r134 16 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=2.525
+ $X2=3.13 $Y2=2.525
r135 16 17 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.045 $Y=2.525
+ $X2=2.18 $Y2=2.525
r136 15 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.105
+ $X2=2.01 $Y2=1.105
r137 14 37 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.045 $Y=1.105
+ $X2=3.28 $Y2=1.105
r138 14 15 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.045 $Y=1.105
+ $X2=2.175 $Y2=1.105
r139 10 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=2.38
+ $X2=3.775 $Y2=2.215
r140 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.775 $Y=2.38
+ $X2=3.775 $Y2=2.75
r141 9 45 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.26 $Y=0.72
+ $X2=3.26 $Y2=1.15
r142 2 35 600 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.96 $X2=2.015 $Y2=2.61
r143 1 28 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.41 $X2=2.01 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%A_863_98# 1 2 9 11 15 19 23 27 31 34 38 40
+ 43 47 50 54 57 59 64 67 71
c118 50 0 1.86828e-19 $X=5.29 $Y=1.32
c119 38 0 1.82849e-19 $X=6.675 $Y=1.485
c120 34 0 1.77373e-19 $X=6.065 $Y=1.485
c121 9 0 6.89381e-20 $X=4.39 $Y=0.83
r122 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.61
+ $Y=1.485 $X2=5.61 $Y2=1.485
r123 62 64 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.37 $Y=1.485
+ $X2=5.61 $Y2=1.485
r124 60 62 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.29 $Y=1.485 $X2=5.37
+ $Y2=1.485
r125 55 67 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=2.32
+ $X2=5.37 $Y2=2.155
r126 55 57 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.37 $Y=2.32
+ $X2=5.37 $Y2=2.815
r127 52 67 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=1.99
+ $X2=5.37 $Y2=2.155
r128 52 54 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=5.37 $Y=1.99
+ $X2=5.37 $Y2=1.985
r129 51 62 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=1.65
+ $X2=5.37 $Y2=1.485
r130 51 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.37 $Y=1.65
+ $X2=5.37 $Y2=1.985
r131 50 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=1.32
+ $X2=5.29 $Y2=1.485
r132 50 59 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.29 $Y=1.32
+ $X2=5.29 $Y2=1.07
r133 45 59 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=5.197 $Y=0.893
+ $X2=5.197 $Y2=1.07
r134 45 47 12.2711 $w=3.53e-07 $l=3.78e-07 $layer=LI1_cond $X=5.197 $Y=0.893
+ $X2=5.197 $Y2=0.515
r135 43 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=2.155
+ $X2=4.48 $Y2=2.32
r136 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.48
+ $Y=2.155 $X2=4.48 $Y2=2.155
r137 40 67 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=2.155
+ $X2=5.37 $Y2=2.155
r138 40 42 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=5.205 $Y=2.155
+ $X2=4.48 $Y2=2.155
r139 37 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.66 $Y=1.485
+ $X2=6.675 $Y2=1.485
r140 36 37 84.8077 $w=3.3e-07 $l=4.85e-07 $layer=POLY_cond $X=6.175 $Y=1.485
+ $X2=6.66 $Y2=1.485
r141 35 36 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.155 $Y=1.485
+ $X2=6.175 $Y2=1.485
r142 34 65 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=6.065 $Y=1.485
+ $X2=5.61 $Y2=1.485
r143 34 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.065 $Y=1.485
+ $X2=6.155 $Y2=1.485
r144 29 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.675 $Y=1.32
+ $X2=6.675 $Y2=1.485
r145 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.675 $Y=1.32
+ $X2=6.675 $Y2=0.855
r146 25 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.65
+ $X2=6.66 $Y2=1.485
r147 25 27 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=6.66 $Y=1.65
+ $X2=6.66 $Y2=2.54
r148 21 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.175 $Y=1.32
+ $X2=6.175 $Y2=1.485
r149 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.175 $Y=1.32
+ $X2=6.175 $Y2=0.76
r150 17 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.65
+ $X2=6.155 $Y2=1.485
r151 17 19 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.155 $Y=1.65
+ $X2=6.155 $Y2=2.4
r152 15 71 167.145 $w=1.8e-07 $l=4.3e-07 $layer=POLY_cond $X=4.43 $Y=2.75
+ $X2=4.43 $Y2=2.32
r153 11 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=1.975
+ $X2=4.48 $Y2=1.81
r154 11 43 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.48 $Y=1.975
+ $X2=4.48 $Y2=2.155
r155 9 33 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.39 $Y=0.83
+ $X2=4.39 $Y2=1.81
r156 2 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.84 $X2=5.37 $Y2=2.815
r157 2 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.84 $X2=5.37 $Y2=1.985
r158 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.045
+ $Y=0.37 $X2=5.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%A_667_80# 1 2 9 13 15 21 23 24 26 27 31 34
+ 36
c88 36 0 1.86828e-19 $X=4.97 $Y=1.405
c89 31 0 1.77373e-19 $X=4.87 $Y=1.405
r90 32 36 18.1887 $w=2.65e-07 $l=1e-07 $layer=POLY_cond $X=4.87 $Y=1.405
+ $X2=4.97 $Y2=1.405
r91 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.87
+ $Y=1.405 $X2=4.87 $Y2=1.405
r92 29 31 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=4.87 $Y=1.65
+ $X2=4.87 $Y2=1.405
r93 28 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=1.735
+ $X2=3.865 $Y2=1.735
r94 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.705 $Y=1.735
+ $X2=4.87 $Y2=1.65
r95 27 28 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.705 $Y=1.735
+ $X2=3.95 $Y2=1.735
r96 26 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=1.65
+ $X2=3.865 $Y2=1.735
r97 25 26 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.865 $Y=0.85
+ $X2=3.865 $Y2=1.65
r98 23 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=1.735
+ $X2=3.865 $Y2=1.735
r99 23 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.78 $Y=1.735
+ $X2=3.555 $Y2=1.735
r100 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=1.82
+ $X2=3.555 $Y2=1.735
r101 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.47 $Y=1.82
+ $X2=3.47 $Y2=2.105
r102 15 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.78 $Y=0.765
+ $X2=3.865 $Y2=0.85
r103 15 17 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.78 $Y=0.765
+ $X2=3.63 $Y2=0.765
r104 11 36 31.8302 $w=2.65e-07 $l=2.43926e-07 $layer=POLY_cond $X=5.145 $Y=1.57
+ $X2=4.97 $Y2=1.405
r105 11 13 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=5.145 $Y=1.57
+ $X2=5.145 $Y2=2.4
r106 7 36 16.0701 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.24
+ $X2=4.97 $Y2=1.405
r107 7 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=4.97 $Y=1.24 $X2=4.97
+ $Y2=0.74
r108 2 21 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.96 $X2=3.47 $Y2=2.105
r109 1 17 182 $w=1.7e-07 $l=4.90816e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.4 $X2=3.63 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%A_1350_116# 1 2 9 13 15 16 19 23 29
c42 23 0 9.14246e-20 $X=6.885 $Y=2.265
c43 19 0 9.14246e-20 $X=6.89 $Y=0.855
r44 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.155
+ $Y=1.485 $X2=7.155 $Y2=1.485
r45 27 29 9.35923 $w=3.28e-07 $l=2.68e-07 $layer=LI1_cond $X=6.887 $Y=1.485
+ $X2=7.155 $Y2=1.485
r46 25 27 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=6.885 $Y=1.485
+ $X2=6.887 $Y2=1.485
r47 21 25 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.885 $Y=1.65
+ $X2=6.885 $Y2=1.485
r48 21 23 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=6.885 $Y=1.65
+ $X2=6.885 $Y2=2.265
r49 17 27 0.643053 $w=3.35e-07 $l=1.65e-07 $layer=LI1_cond $X=6.887 $Y=1.32
+ $X2=6.887 $Y2=1.485
r50 17 19 15.9966 $w=3.33e-07 $l=4.65e-07 $layer=LI1_cond $X=6.887 $Y=1.32
+ $X2=6.887 $Y2=0.855
r51 15 30 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=7.57 $Y=1.485
+ $X2=7.155 $Y2=1.485
r52 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.57 $Y=1.485 $X2=7.66
+ $Y2=1.485
r53 11 16 34.7346 $w=1.65e-07 $l=1.67481e-07 $layer=POLY_cond $X=7.665 $Y=1.32
+ $X2=7.66 $Y2=1.485
r54 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.665 $Y=1.32
+ $X2=7.665 $Y2=0.74
r55 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=7.66 $Y=1.65
+ $X2=7.66 $Y2=1.485
r56 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.66 $Y=1.65 $X2=7.66
+ $Y2=2.4
r57 2 23 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.12 $X2=6.885 $Y2=2.265
r58 1 19 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=6.75
+ $Y=0.58 $X2=6.89 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%VPWR 1 2 3 4 5 20 24 26 30 34 38 43 44 46 47
+ 48 50 69 70 73 76 79
r92 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r96 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r97 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r98 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r99 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r100 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r101 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r103 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 58 79 11.8853 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.762 $Y2=3.33
r105 58 60 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r111 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r113 51 53 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r115 50 56 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 48 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 48 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 46 66 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.27 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.27 $Y=3.33
+ $X2=7.395 $Y2=3.33
r120 45 69 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.52 $Y=3.33 $X2=7.92
+ $Y2=3.33
r121 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.52 $Y=3.33
+ $X2=7.395 $Y2=3.33
r122 43 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.295 $Y=3.33 $X2=6
+ $Y2=3.33
r123 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=3.33
+ $X2=6.42 $Y2=3.33
r124 42 66 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.42 $Y2=3.33
r126 38 41 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.395 $Y=1.985
+ $X2=7.395 $Y2=2.815
r127 36 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.395 $Y=3.245
+ $X2=7.395 $Y2=3.33
r128 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.395 $Y=3.245
+ $X2=7.395 $Y2=2.815
r129 32 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=3.33
r130 32 34 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=2.265
r131 28 79 2.29102 $w=5.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.762 $Y=3.245
+ $X2=4.762 $Y2=3.33
r132 28 30 11.7413 $w=5.43e-07 $l=5.35e-07 $layer=LI1_cond $X=4.762 $Y=3.245
+ $X2=4.762 $Y2=2.71
r133 27 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r134 26 79 11.8853 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=4.762 $Y2=3.33
r135 26 27 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=2.71 $Y2=3.33
r136 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r137 22 24 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=2.945
r138 18 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r139 18 20 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.05
r140 5 41 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.435 $Y2=2.815
r141 5 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.435 $Y2=1.985
r142 4 34 300 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_PDIFF $count=2 $X=6.245
+ $Y=1.84 $X2=6.38 $Y2=2.265
r143 3 30 600 $w=1.7e-07 $l=3.13688e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=2.54 $X2=4.76 $Y2=2.71
r144 2 24 600 $w=1.7e-07 $l=1.0872e-06 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=1.96 $X2=2.545 $Y2=2.945
r145 1 20 600 $w=1.7e-07 $l=1.0872e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=2.065 $X2=0.805 $Y2=3.05
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%Q 1 2 9 14 15 16 17 28
r37 21 28 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=5.96 $Y=0.985 $X2=5.96
+ $Y2=0.925
r38 17 30 8.04311 $w=3.28e-07 $l=1.53e-07 $layer=LI1_cond $X=5.96 $Y=0.997
+ $X2=5.96 $Y2=1.15
r39 17 21 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=5.96 $Y=0.997
+ $X2=5.96 $Y2=0.985
r40 17 28 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=5.96 $Y=0.912
+ $X2=5.96 $Y2=0.925
r41 16 17 13.1658 $w=3.28e-07 $l=3.77e-07 $layer=LI1_cond $X=5.96 $Y=0.535
+ $X2=5.96 $Y2=0.912
r42 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.04 $Y=1.82
+ $X2=6.04 $Y2=1.15
r43 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.945 $Y=1.985
+ $X2=5.945 $Y2=1.82
r44 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.945 $Y=2 $X2=5.945
+ $Y2=1.985
r45 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=5.945 $Y=2 $X2=5.945
+ $Y2=2.815
r46 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.93 $Y2=1.985
r47 2 9 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.93 $Y2=2.815
r48 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.39 $X2=5.96 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%Q_N 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=2.405
+ $X2=7.882 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.882 $Y=1.985
+ $X2=7.882 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=7.882 $Y=1.665
+ $X2=7.882 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=1.295
+ $X2=7.882 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=0.925
+ $X2=7.882 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=7.882 $Y=0.515
+ $X2=7.882 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=1.84 $X2=7.885 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=1.84 $X2=7.885 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.37 $X2=7.88 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBP_1%VGND 1 2 3 4 5 18 22 26 30 33 34 35 37 42 50
+ 62 68 69 72 82 85
r85 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r86 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r87 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r88 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r89 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r90 66 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.41
+ $Y2=0
r91 66 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.92
+ $Y2=0
r92 65 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r93 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r94 62 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.285 $Y=0 $X2=7.41
+ $Y2=0
r95 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.285 $Y=0 $X2=6.96
+ $Y2=0
r96 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r97 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r98 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r99 58 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r100 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r101 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 55 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=4.685
+ $Y2=0
r103 55 57 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.85 $Y=0 $X2=5.04
+ $Y2=0
r104 54 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r105 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r106 51 53 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=3.12
+ $Y2=0
r107 50 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=0 $X2=4.685
+ $Y2=0
r108 50 53 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=4.52 $Y=0 $X2=3.12
+ $Y2=0
r109 49 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r110 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r111 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r112 46 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r113 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r114 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r115 43 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r116 43 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r117 42 79 9.72841 $w=3.83e-07 $l=3.25e-07 $layer=LI1_cond $X=2.547 $Y=0
+ $X2=2.547 $Y2=0.325
r118 42 51 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.547 $Y=0 $X2=2.74
+ $Y2=0
r119 42 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r120 42 48 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.16 $Y2=0
r121 40 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 37 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.795
+ $Y2=0
r124 37 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r125 35 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r126 35 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r127 33 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6
+ $Y2=0
r128 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.42
+ $Y2=0
r129 32 64 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.96 $Y2=0
r130 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=0 $X2=6.42
+ $Y2=0
r131 28 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0
r132 28 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0.515
r133 24 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r134 24 26 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.855
r135 20 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0
r136 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0.515
r137 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r138 16 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.52
r139 5 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.305
+ $Y=0.37 $X2=7.45 $Y2=0.515
r140 4 26 182 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.39 $X2=6.425 $Y2=0.855
r141 3 22 91 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_NDIFF $count=2 $X=4.465
+ $Y=0.62 $X2=4.685 $Y2=0.515
r142 2 79 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.41 $X2=2.545 $Y2=0.325
r143 1 18 91 $w=1.7e-07 $l=2.39165e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.52
.ends


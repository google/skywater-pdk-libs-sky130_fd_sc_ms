* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
M1000 VGND C2 a_119_74# VNB nlowvt w=640000u l=150000u
+  ad=9.082e+11p pd=5.52e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_32_74# C1 a_27_390# VPB pshort w=1e+06u l=180000u
+  ad=4.25e+11p pd=2.85e+06u as=8.8e+11p ps=7.76e+06u
M1002 X a_32_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 VGND A2 a_651_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1004 a_651_74# A1 a_32_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.848e+11p ps=4.7e+06u
M1005 a_119_74# C1 a_32_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_386_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1007 a_32_74# B1 a_386_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_340_390# B2 a_27_390# VPB pshort w=1e+06u l=180000u
+  ad=6.8e+11p pd=5.36e+06u as=0p ps=0u
M1009 a_27_390# C2 a_32_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_390# B1 a_340_390# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_340_390# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.686e+11p ps=5.71e+06u
M1012 VPWR A2 a_340_390# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_32_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__a31o_4.pxi.spice
* Created: Wed Sep  2 11:55:15 2020
* 
x_PM_SKY130_FD_SC_MS__A31O_4%A_83_274# N_A_83_274#_M1002_d N_A_83_274#_M1007_d
+ N_A_83_274#_M1015_d N_A_83_274#_M1010_d N_A_83_274#_M1001_g
+ N_A_83_274#_c_131_n N_A_83_274#_M1012_g N_A_83_274#_M1005_g
+ N_A_83_274#_c_133_n N_A_83_274#_M1013_g N_A_83_274#_c_134_n
+ N_A_83_274#_M1018_g N_A_83_274#_M1008_g N_A_83_274#_c_136_n
+ N_A_83_274#_M1019_g N_A_83_274#_M1009_g N_A_83_274#_c_211_p
+ N_A_83_274#_c_138_n N_A_83_274#_c_139_n N_A_83_274#_c_140_n
+ N_A_83_274#_c_141_n N_A_83_274#_c_142_n N_A_83_274#_c_143_n
+ N_A_83_274#_c_163_p N_A_83_274#_c_144_n N_A_83_274#_c_145_n
+ N_A_83_274#_c_146_n PM_SKY130_FD_SC_MS__A31O_4%A_83_274#
x_PM_SKY130_FD_SC_MS__A31O_4%B1 N_B1_M1002_g N_B1_M1010_g N_B1_M1007_g
+ N_B1_M1011_g B1 N_B1_c_274_n PM_SKY130_FD_SC_MS__A31O_4%B1
x_PM_SKY130_FD_SC_MS__A31O_4%A1 N_A1_c_332_n N_A1_M1014_g N_A1_c_333_n
+ N_A1_c_334_n N_A1_c_335_n N_A1_M1000_g N_A1_c_336_n N_A1_M1015_g N_A1_M1022_g
+ N_A1_c_337_n A1 A1 N_A1_c_339_n PM_SKY130_FD_SC_MS__A31O_4%A1
x_PM_SKY130_FD_SC_MS__A31O_4%A2 N_A2_M1004_g N_A2_c_399_n N_A2_c_400_n
+ N_A2_c_401_n N_A2_M1006_g N_A2_M1023_g N_A2_M1017_g N_A2_c_403_n N_A2_c_404_n
+ A2 A2 N_A2_c_405_n N_A2_c_406_n PM_SKY130_FD_SC_MS__A31O_4%A2
x_PM_SKY130_FD_SC_MS__A31O_4%A3 N_A3_M1020_g N_A3_M1003_g N_A3_M1016_g
+ N_A3_M1021_g A3 A3 N_A3_c_470_n PM_SKY130_FD_SC_MS__A31O_4%A3
x_PM_SKY130_FD_SC_MS__A31O_4%VPWR N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_M1009_s
+ N_VPWR_M1000_d N_VPWR_M1004_d N_VPWR_M1020_s N_VPWR_c_509_n N_VPWR_c_510_n
+ N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_515_n
+ N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n VPWR
+ N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n N_VPWR_c_508_n
+ N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n PM_SKY130_FD_SC_MS__A31O_4%VPWR
x_PM_SKY130_FD_SC_MS__A31O_4%X N_X_M1012_d N_X_M1018_d N_X_M1001_d N_X_M1008_d
+ N_X_c_603_n N_X_c_611_n N_X_c_606_n N_X_c_604_n N_X_c_607_n X X X X
+ N_X_c_605_n PM_SKY130_FD_SC_MS__A31O_4%X
x_PM_SKY130_FD_SC_MS__A31O_4%A_529_392# N_A_529_392#_M1010_s
+ N_A_529_392#_M1011_s N_A_529_392#_M1022_s N_A_529_392#_M1023_s
+ N_A_529_392#_M1021_d N_A_529_392#_c_660_n N_A_529_392#_c_661_n
+ N_A_529_392#_c_662_n N_A_529_392#_c_663_n N_A_529_392#_c_664_n
+ N_A_529_392#_c_665_n N_A_529_392#_c_666_n N_A_529_392#_c_667_n
+ N_A_529_392#_c_668_n N_A_529_392#_c_669_n N_A_529_392#_c_670_n
+ N_A_529_392#_c_671_n N_A_529_392#_c_672_n N_A_529_392#_c_673_n
+ PM_SKY130_FD_SC_MS__A31O_4%A_529_392#
x_PM_SKY130_FD_SC_MS__A31O_4%VGND N_VGND_M1012_s N_VGND_M1013_s N_VGND_M1019_s
+ N_VGND_M1002_s N_VGND_M1003_d N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n
+ N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n VGND N_VGND_c_756_n
+ N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n
+ N_VGND_c_762_n N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n
+ PM_SKY130_FD_SC_MS__A31O_4%VGND
x_PM_SKY130_FD_SC_MS__A31O_4%A_775_74# N_A_775_74#_M1014_s N_A_775_74#_M1006_d
+ N_A_775_74#_c_842_n N_A_775_74#_c_840_n N_A_775_74#_c_841_n
+ N_A_775_74#_c_854_n PM_SKY130_FD_SC_MS__A31O_4%A_775_74#
x_PM_SKY130_FD_SC_MS__A31O_4%A_1000_74# N_A_1000_74#_M1006_s
+ N_A_1000_74#_M1017_s N_A_1000_74#_M1016_s N_A_1000_74#_c_867_n
+ N_A_1000_74#_c_868_n N_A_1000_74#_c_869_n N_A_1000_74#_c_870_n
+ N_A_1000_74#_c_871_n N_A_1000_74#_c_872_n N_A_1000_74#_c_873_n
+ PM_SKY130_FD_SC_MS__A31O_4%A_1000_74#
cc_1 VNB N_A_83_274#_M1001_g 0.00871317f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_274#_c_131_n 0.0208118f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_3 VNB N_A_83_274#_M1005_g 0.00577081f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_4 VNB N_A_83_274#_c_133_n 0.0168814f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_5 VNB N_A_83_274#_c_134_n 0.0167202f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.22
cc_6 VNB N_A_83_274#_M1008_g 0.00621938f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_7 VNB N_A_83_274#_c_136_n 0.0199378f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.22
cc_8 VNB N_A_83_274#_M1009_g 0.00688285f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_9 VNB N_A_83_274#_c_138_n 0.0117524f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=0.515
cc_10 VNB N_A_83_274#_c_139_n 0.00958212f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.215
cc_11 VNB N_A_83_274#_c_140_n 0.0268008f $X=-0.19 $Y=-0.245 $X2=2.74 $Y2=1.215
cc_12 VNB N_A_83_274#_c_141_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=0.515
cc_13 VNB N_A_83_274#_c_142_n 0.0107873f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=1.195
cc_14 VNB N_A_83_274#_c_143_n 0.00616633f $X=-0.19 $Y=-0.245 $X2=4.585 $Y2=0.76
cc_15 VNB N_A_83_274#_c_144_n 0.00376476f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=1.97
cc_16 VNB N_A_83_274#_c_145_n 0.00593555f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.13
cc_17 VNB N_A_83_274#_c_146_n 0.130207f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.385
cc_18 VNB N_B1_M1002_g 0.0393688f $X=-0.19 $Y=-0.245 $X2=4.375 $Y2=0.37
cc_19 VNB N_B1_M1007_g 0.0360572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.00224847f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_21 VNB N_B1_c_274_n 0.0404856f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_22 VNB N_A1_c_332_n 0.0156956f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=0.37
cc_23 VNB N_A1_c_333_n 0.00921382f $X=-0.19 $Y=-0.245 $X2=3.105 $Y2=1.96
cc_24 VNB N_A1_c_334_n 0.00862272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_c_335_n 0.0199174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_c_336_n 0.0174223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_337_n 0.0112882f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_28 VNB A1 0.00258642f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_29 VNB N_A1_c_339_n 0.0360126f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.55
cc_30 VNB N_A2_c_399_n 0.0108595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_400_n 0.0144295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_401_n 0.0168779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_M1017_g 0.0376337f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_34 VNB N_A2_c_403_n 0.00726442f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.55
cc_35 VNB N_A2_c_404_n 0.0211715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_c_405_n 0.00873674f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.55
cc_37 VNB N_A2_c_406_n 0.00587819f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_38 VNB N_A3_M1003_g 0.0324872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A3_M1016_g 0.0431332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB A3 0.0133116f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_41 VNB N_A3_c_470_n 0.0299617f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_42 VNB N_VPWR_c_508_n 0.302998f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.385
cc_43 VNB N_X_c_603_n 0.00253236f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_44 VNB N_X_c_604_n 0.00211712f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_45 VNB N_X_c_605_n 0.002f $X=-0.19 $Y=-0.245 $X2=2.74 $Y2=1.215
cc_46 VNB N_VGND_c_750_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_751_n 0.0542158f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_48 VNB N_VGND_c_752_n 0.00263668f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_49 VNB N_VGND_c_753_n 0.0107234f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_50 VNB N_VGND_c_754_n 0.00583463f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.55
cc_51 VNB N_VGND_c_755_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.22
cc_52 VNB N_VGND_c_756_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_53 VNB N_VGND_c_757_n 0.0159167f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.385
cc_54 VNB N_VGND_c_758_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.385
cc_55 VNB N_VGND_c_759_n 0.0744736f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.215
cc_56 VNB N_VGND_c_760_n 0.0191411f $X=-0.19 $Y=-0.245 $X2=4.585 $Y2=1.11
cc_57 VNB N_VGND_c_761_n 0.400335f $X=-0.19 $Y=-0.245 $X2=4.585 $Y2=0.76
cc_58 VNB N_VGND_c_762_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.13
cc_59 VNB N_VGND_c_763_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=1.97
cc_60 VNB N_VGND_c_764_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_61 VNB N_VGND_c_765_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.385
cc_62 VNB N_A_775_74#_c_840_n 0.0196946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_775_74#_c_841_n 0.00374971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1000_74#_c_867_n 0.00537913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1000_74#_c_868_n 0.00878949f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_66 VNB N_A_1000_74#_c_869_n 0.00222615f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_67 VNB N_A_1000_74#_c_870_n 0.00356893f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_68 VNB N_A_1000_74#_c_871_n 0.0193916f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.55
cc_69 VNB N_A_1000_74#_c_872_n 0.0316008f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_70 VNB N_A_1000_74#_c_873_n 0.00294697f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_71 VPB N_A_83_274#_M1001_g 0.0274205f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_72 VPB N_A_83_274#_M1005_g 0.0222985f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_73 VPB N_A_83_274#_M1008_g 0.0225445f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_74 VPB N_A_83_274#_M1009_g 0.0246942f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_75 VPB N_A_83_274#_c_144_n 0.0016955f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=1.97
cc_76 VPB N_B1_M1010_g 0.0260324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_B1_M1011_g 0.0233607f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_78 VPB B1 0.0019221f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_79 VPB N_B1_c_274_n 0.0368653f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.22
cc_80 VPB N_A1_M1000_g 0.0255432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A1_M1022_g 0.0239355f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_82 VPB A1 0.00182137f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_83 VPB N_A1_c_339_n 0.0184685f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.55
cc_84 VPB N_A2_M1004_g 0.0240433f $X=-0.19 $Y=1.66 $X2=4.375 $Y2=0.37
cc_85 VPB N_A2_c_400_n 0.00964737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A2_M1023_g 0.0246231f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_87 VPB N_A2_c_403_n 0.00382585f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.55
cc_88 VPB N_A2_c_405_n 0.00678093f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.55
cc_89 VPB N_A2_c_406_n 0.00279107f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_90 VPB N_A3_M1020_g 0.0234013f $X=-0.19 $Y=1.66 $X2=4.375 $Y2=0.37
cc_91 VPB N_A3_M1021_g 0.0318882f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_92 VPB A3 0.00802022f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_93 VPB N_A3_c_470_n 0.017688f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_94 VPB N_VPWR_c_509_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_95 VPB N_VPWR_c_510_n 0.0645583f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_96 VPB N_VPWR_c_511_n 0.00899828f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.22
cc_97 VPB N_VPWR_c_512_n 0.0237727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_513_n 0.00898491f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_99 VPB N_VPWR_c_514_n 0.00906077f $X=-0.19 $Y=1.66 $X2=1.15 $Y2=1.385
cc_100 VPB N_VPWR_c_515_n 0.00635773f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.385
cc_101 VPB N_VPWR_c_516_n 0.0474919f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.515
cc_102 VPB N_VPWR_c_517_n 0.00632158f $X=-0.19 $Y=1.66 $X2=2.655 $Y2=0.515
cc_103 VPB N_VPWR_c_518_n 0.0186948f $X=-0.19 $Y=1.66 $X2=3.405 $Y2=1.215
cc_104 VPB N_VPWR_c_519_n 0.00632158f $X=-0.19 $Y=1.66 $X2=2.74 $Y2=1.215
cc_105 VPB N_VPWR_c_520_n 0.0196495f $X=-0.19 $Y=1.66 $X2=3.585 $Y2=1.11
cc_106 VPB N_VPWR_c_521_n 0.0186948f $X=-0.19 $Y=1.66 $X2=3.75 $Y2=1.195
cc_107 VPB N_VPWR_c_522_n 0.018855f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_108 VPB N_VPWR_c_523_n 0.0191515f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.385
cc_109 VPB N_VPWR_c_508_n 0.0837558f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.385
cc_110 VPB N_VPWR_c_525_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_526_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_527_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_X_c_606_n 0.00558234f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_114 VPB N_X_c_607_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_115 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=0.74
cc_116 VPB N_A_529_392#_c_660_n 0.00420248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_529_392#_c_661_n 0.00767625f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_118 VPB N_A_529_392#_c_662_n 0.00384413f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.55
cc_119 VPB N_A_529_392#_c_663_n 0.00466903f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_120 VPB N_A_529_392#_c_664_n 0.00261786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_529_392#_c_665_n 0.00279507f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.22
cc_122 VPB N_A_529_392#_c_666_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_123 VPB N_A_529_392#_c_667_n 0.00285515f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.55
cc_124 VPB N_A_529_392#_c_668_n 0.00275675f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.22
cc_125 VPB N_A_529_392#_c_669_n 0.00274662f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=0.74
cc_126 VPB N_A_529_392#_c_670_n 0.0102169f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_127 VPB N_A_529_392#_c_671_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_529_392#_c_672_n 0.00723598f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=1.13
cc_129 VPB N_A_529_392#_c_673_n 0.00430557f $X=-0.19 $Y=1.66 $X2=2.655 $Y2=0.515
cc_130 N_A_83_274#_c_138_n N_B1_M1002_g 0.00527749f $X=2.655 $Y=0.515 $X2=0
+ $Y2=0
cc_131 N_A_83_274#_c_139_n N_B1_M1002_g 0.0161307f $X=3.405 $Y=1.215 $X2=0 $Y2=0
cc_132 N_A_83_274#_c_140_n N_B1_M1002_g 9.26602e-19 $X=2.74 $Y=1.215 $X2=0 $Y2=0
cc_133 N_A_83_274#_c_141_n N_B1_M1002_g 7.42424e-19 $X=3.585 $Y=0.515 $X2=0
+ $Y2=0
cc_134 N_A_83_274#_c_144_n N_B1_M1002_g 8.24452e-19 $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_135 N_A_83_274#_c_146_n N_B1_M1002_g 0.00546699f $X=1.955 $Y=1.385 $X2=0
+ $Y2=0
cc_136 N_A_83_274#_c_144_n N_B1_M1010_g 0.00291431f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_137 N_A_83_274#_c_139_n N_B1_M1007_g 0.0118906f $X=3.405 $Y=1.215 $X2=0 $Y2=0
cc_138 N_A_83_274#_c_141_n N_B1_M1007_g 0.0107217f $X=3.585 $Y=0.515 $X2=0 $Y2=0
cc_139 N_A_83_274#_c_144_n N_B1_M1007_g 0.00531551f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_140 N_A_83_274#_c_145_n N_B1_M1007_g 0.00442223f $X=3.405 $Y=1.13 $X2=0 $Y2=0
cc_141 N_A_83_274#_c_163_p N_B1_M1011_g 0.0143936f $X=3.3 $Y=2.085 $X2=0 $Y2=0
cc_142 N_A_83_274#_c_144_n N_B1_M1011_g 0.00531948f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_143 N_A_83_274#_M1009_g B1 0.00122078f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_83_274#_c_139_n B1 0.0366052f $X=3.405 $Y=1.215 $X2=0 $Y2=0
cc_145 N_A_83_274#_c_140_n B1 0.0199912f $X=2.74 $Y=1.215 $X2=0 $Y2=0
cc_146 N_A_83_274#_c_163_p B1 0.00737847f $X=3.3 $Y=2.085 $X2=0 $Y2=0
cc_147 N_A_83_274#_c_144_n B1 0.0249544f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_148 N_A_83_274#_M1009_g N_B1_c_274_n 0.00459228f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_83_274#_c_139_n N_B1_c_274_n 0.00567282f $X=3.405 $Y=1.215 $X2=0
+ $Y2=0
cc_150 N_A_83_274#_c_140_n N_B1_c_274_n 0.00417566f $X=2.74 $Y=1.215 $X2=0 $Y2=0
cc_151 N_A_83_274#_c_163_p N_B1_c_274_n 0.00512322f $X=3.3 $Y=2.085 $X2=0 $Y2=0
cc_152 N_A_83_274#_c_144_n N_B1_c_274_n 0.014735f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_153 N_A_83_274#_c_145_n N_B1_c_274_n 0.00196877f $X=3.405 $Y=1.13 $X2=0 $Y2=0
cc_154 N_A_83_274#_c_146_n N_B1_c_274_n 0.00468439f $X=1.955 $Y=1.385 $X2=0
+ $Y2=0
cc_155 N_A_83_274#_c_141_n N_A1_c_332_n 0.010214f $X=3.585 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_83_274#_c_142_n N_A1_c_333_n 0.00749193f $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_157 N_A_83_274#_c_141_n N_A1_c_334_n 9.8511e-19 $X=3.585 $Y=0.515 $X2=0 $Y2=0
cc_158 N_A_83_274#_c_142_n N_A1_c_334_n 0.00877685f $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_159 N_A_83_274#_c_145_n N_A1_c_334_n 0.00215915f $X=3.405 $Y=1.13 $X2=0 $Y2=0
cc_160 N_A_83_274#_c_142_n N_A1_c_335_n 0.00746623f $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_161 N_A_83_274#_c_144_n N_A1_c_335_n 0.00257472f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_162 N_A_83_274#_c_145_n N_A1_c_335_n 4.51009e-19 $X=3.405 $Y=1.13 $X2=0 $Y2=0
cc_163 N_A_83_274#_c_141_n N_A1_c_336_n 4.36444e-19 $X=3.585 $Y=0.515 $X2=0
+ $Y2=0
cc_164 N_A_83_274#_c_143_n N_A1_c_336_n 0.010812f $X=4.585 $Y=0.76 $X2=0 $Y2=0
cc_165 N_A_83_274#_c_142_n N_A1_c_337_n 0.0137085f $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_166 N_A_83_274#_c_142_n A1 0.0547704f $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_167 N_A_83_274#_c_144_n A1 0.0151243f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_168 N_A_83_274#_c_142_n N_A1_c_339_n 0.0101596f $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_169 N_A_83_274#_c_144_n N_A1_c_339_n 0.00172043f $X=3.35 $Y=1.97 $X2=0 $Y2=0
cc_170 N_A_83_274#_c_142_n N_A2_c_404_n 7.12337e-19 $X=4.42 $Y=1.195 $X2=0 $Y2=0
cc_171 N_A_83_274#_M1001_g N_VPWR_c_510_n 0.00649215f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_172 N_A_83_274#_M1005_g N_VPWR_c_511_n 0.00343717f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_173 N_A_83_274#_M1008_g N_VPWR_c_511_n 0.00203999f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_174 N_A_83_274#_M1009_g N_VPWR_c_512_n 0.00546726f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_175 N_A_83_274#_c_140_n N_VPWR_c_512_n 0.0186821f $X=2.74 $Y=1.215 $X2=0
+ $Y2=0
cc_176 N_A_83_274#_c_146_n N_VPWR_c_512_n 0.0020126f $X=1.955 $Y=1.385 $X2=0
+ $Y2=0
cc_177 N_A_83_274#_M1001_g N_VPWR_c_520_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A_83_274#_M1005_g N_VPWR_c_520_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_83_274#_M1008_g N_VPWR_c_521_n 0.005209f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_83_274#_M1009_g N_VPWR_c_521_n 0.005209f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_83_274#_M1001_g N_VPWR_c_508_n 0.00986008f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_182 N_A_83_274#_M1005_g N_VPWR_c_508_n 0.00982526f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_183 N_A_83_274#_M1008_g N_VPWR_c_508_n 0.00982526f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A_83_274#_M1009_g N_VPWR_c_508_n 0.00986727f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_185 N_A_83_274#_c_131_n N_X_c_603_n 4.74419e-19 $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_186 N_A_83_274#_c_133_n N_X_c_603_n 4.44219e-19 $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_187 N_A_83_274#_c_133_n N_X_c_611_n 0.0139501f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_188 N_A_83_274#_c_134_n N_X_c_611_n 0.00988574f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_189 N_A_83_274#_c_211_p N_X_c_611_n 0.0355741f $X=1.895 $Y=1.385 $X2=0 $Y2=0
cc_190 N_A_83_274#_c_146_n N_X_c_611_n 0.00535312f $X=1.955 $Y=1.385 $X2=0 $Y2=0
cc_191 N_A_83_274#_M1005_g N_X_c_606_n 0.0191156f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_83_274#_M1008_g N_X_c_606_n 0.0157736f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_83_274#_M1009_g N_X_c_606_n 0.00538979f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_83_274#_c_211_p N_X_c_606_n 0.0645108f $X=1.895 $Y=1.385 $X2=0 $Y2=0
cc_195 N_A_83_274#_c_146_n N_X_c_606_n 0.00694776f $X=1.955 $Y=1.385 $X2=0 $Y2=0
cc_196 N_A_83_274#_c_134_n N_X_c_604_n 2.95615e-19 $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_197 N_A_83_274#_c_136_n N_X_c_604_n 0.00173245f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_198 N_A_83_274#_M1005_g N_X_c_607_n 4.58171e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_83_274#_M1008_g N_X_c_607_n 0.0151125f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_83_274#_M1009_g N_X_c_607_n 0.013879f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_83_274#_M1001_g X 0.0161078f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_83_274#_M1005_g X 0.00782078f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_83_274#_M1008_g X 0.00131515f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_83_274#_c_146_n X 0.0054939f $X=1.955 $Y=1.385 $X2=0 $Y2=0
cc_205 N_A_83_274#_M1001_g X 0.014728f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_83_274#_M1005_g X 0.0151125f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_83_274#_c_131_n N_X_c_605_n 0.00263346f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_208 N_A_83_274#_c_133_n N_X_c_605_n 0.00286407f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_209 N_A_83_274#_c_211_p N_X_c_605_n 0.0225199f $X=1.895 $Y=1.385 $X2=0 $Y2=0
cc_210 N_A_83_274#_c_146_n N_X_c_605_n 0.0295979f $X=1.955 $Y=1.385 $X2=0 $Y2=0
cc_211 N_A_83_274#_M1010_d N_A_529_392#_c_662_n 0.00240242f $X=3.105 $Y=1.96
+ $X2=0 $Y2=0
cc_212 N_A_83_274#_c_163_p N_A_529_392#_c_662_n 0.0268288f $X=3.3 $Y=2.085 $X2=0
+ $Y2=0
cc_213 N_A_83_274#_c_142_n N_A_529_392#_c_663_n 0.00693098f $X=4.42 $Y=1.195
+ $X2=0 $Y2=0
cc_214 N_A_83_274#_c_144_n N_A_529_392#_c_663_n 0.0142238f $X=3.35 $Y=1.97 $X2=0
+ $Y2=0
cc_215 N_A_83_274#_c_163_p N_A_529_392#_c_664_n 0.041273f $X=3.3 $Y=2.085 $X2=0
+ $Y2=0
cc_216 N_A_83_274#_c_142_n N_A_529_392#_c_665_n 0.00197378f $X=4.42 $Y=1.195
+ $X2=0 $Y2=0
cc_217 N_A_83_274#_c_131_n N_VGND_c_751_n 0.00551153f $X=0.52 $Y=1.22 $X2=0
+ $Y2=0
cc_218 N_A_83_274#_c_146_n N_VGND_c_751_n 0.00130153f $X=1.955 $Y=1.385 $X2=0
+ $Y2=0
cc_219 N_A_83_274#_c_131_n N_VGND_c_752_n 4.20062e-19 $X=0.52 $Y=1.22 $X2=0
+ $Y2=0
cc_220 N_A_83_274#_c_133_n N_VGND_c_752_n 0.00759271f $X=0.995 $Y=1.22 $X2=0
+ $Y2=0
cc_221 N_A_83_274#_c_134_n N_VGND_c_752_n 0.00739907f $X=1.425 $Y=1.22 $X2=0
+ $Y2=0
cc_222 N_A_83_274#_c_136_n N_VGND_c_752_n 3.63246e-19 $X=1.88 $Y=1.22 $X2=0
+ $Y2=0
cc_223 N_A_83_274#_c_134_n N_VGND_c_753_n 4.28983e-19 $X=1.425 $Y=1.22 $X2=0
+ $Y2=0
cc_224 N_A_83_274#_c_136_n N_VGND_c_753_n 0.0119292f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_225 N_A_83_274#_c_138_n N_VGND_c_753_n 0.0402788f $X=2.655 $Y=0.515 $X2=0
+ $Y2=0
cc_226 N_A_83_274#_c_140_n N_VGND_c_753_n 0.0263324f $X=2.74 $Y=1.215 $X2=0
+ $Y2=0
cc_227 N_A_83_274#_c_146_n N_VGND_c_753_n 0.00176127f $X=1.955 $Y=1.385 $X2=0
+ $Y2=0
cc_228 N_A_83_274#_c_138_n N_VGND_c_754_n 0.0225912f $X=2.655 $Y=0.515 $X2=0
+ $Y2=0
cc_229 N_A_83_274#_c_139_n N_VGND_c_754_n 0.0238718f $X=3.405 $Y=1.215 $X2=0
+ $Y2=0
cc_230 N_A_83_274#_c_141_n N_VGND_c_754_n 0.0236791f $X=3.585 $Y=0.515 $X2=0
+ $Y2=0
cc_231 N_A_83_274#_c_131_n N_VGND_c_756_n 0.00460063f $X=0.52 $Y=1.22 $X2=0
+ $Y2=0
cc_232 N_A_83_274#_c_133_n N_VGND_c_756_n 0.00383152f $X=0.995 $Y=1.22 $X2=0
+ $Y2=0
cc_233 N_A_83_274#_c_134_n N_VGND_c_757_n 0.00383152f $X=1.425 $Y=1.22 $X2=0
+ $Y2=0
cc_234 N_A_83_274#_c_136_n N_VGND_c_757_n 0.00383152f $X=1.88 $Y=1.22 $X2=0
+ $Y2=0
cc_235 N_A_83_274#_c_138_n N_VGND_c_758_n 0.011066f $X=2.655 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_A_83_274#_c_141_n N_VGND_c_759_n 0.0144922f $X=3.585 $Y=0.515 $X2=0
+ $Y2=0
cc_237 N_A_83_274#_c_131_n N_VGND_c_761_n 0.00911274f $X=0.52 $Y=1.22 $X2=0
+ $Y2=0
cc_238 N_A_83_274#_c_133_n N_VGND_c_761_n 0.00382307f $X=0.995 $Y=1.22 $X2=0
+ $Y2=0
cc_239 N_A_83_274#_c_134_n N_VGND_c_761_n 0.00382119f $X=1.425 $Y=1.22 $X2=0
+ $Y2=0
cc_240 N_A_83_274#_c_136_n N_VGND_c_761_n 0.00757785f $X=1.88 $Y=1.22 $X2=0
+ $Y2=0
cc_241 N_A_83_274#_c_138_n N_VGND_c_761_n 0.00915947f $X=2.655 $Y=0.515 $X2=0
+ $Y2=0
cc_242 N_A_83_274#_c_141_n N_VGND_c_761_n 0.0118826f $X=3.585 $Y=0.515 $X2=0
+ $Y2=0
cc_243 N_A_83_274#_c_142_n N_A_775_74#_c_842_n 0.0227079f $X=4.42 $Y=1.195 $X2=0
+ $Y2=0
cc_244 N_A_83_274#_M1015_d N_A_775_74#_c_840_n 0.00369086f $X=4.375 $Y=0.37
+ $X2=0 $Y2=0
cc_245 N_A_83_274#_c_143_n N_A_775_74#_c_840_n 0.0241965f $X=4.585 $Y=0.76 $X2=0
+ $Y2=0
cc_246 N_A_83_274#_c_141_n N_A_775_74#_c_841_n 0.00371332f $X=3.585 $Y=0.515
+ $X2=0 $Y2=0
cc_247 N_A_83_274#_c_143_n N_A_1000_74#_c_867_n 0.0339399f $X=4.585 $Y=0.76
+ $X2=0 $Y2=0
cc_248 N_A_83_274#_c_142_n N_A_1000_74#_c_869_n 0.012865f $X=4.42 $Y=1.195 $X2=0
+ $Y2=0
cc_249 N_B1_M1007_g N_A1_c_332_n 0.0157482f $X=3.37 $Y=0.69 $X2=-0.19 $Y2=-0.245
cc_250 N_B1_M1007_g N_A1_c_335_n 0.00291887f $X=3.37 $Y=0.69 $X2=0 $Y2=0
cc_251 N_B1_M1011_g N_A1_M1000_g 0.011669f $X=3.535 $Y=2.46 $X2=0 $Y2=0
cc_252 N_B1_M1007_g A1 8.09225e-19 $X=3.37 $Y=0.69 $X2=0 $Y2=0
cc_253 N_B1_c_274_n A1 0.001245f $X=3.37 $Y=1.635 $X2=0 $Y2=0
cc_254 N_B1_c_274_n N_A1_c_339_n 0.0145879f $X=3.37 $Y=1.635 $X2=0 $Y2=0
cc_255 N_B1_M1010_g N_VPWR_c_512_n 0.00838372f $X=3.015 $Y=2.46 $X2=0 $Y2=0
cc_256 N_B1_M1010_g N_VPWR_c_516_n 0.00349951f $X=3.015 $Y=2.46 $X2=0 $Y2=0
cc_257 N_B1_M1011_g N_VPWR_c_516_n 0.00349978f $X=3.535 $Y=2.46 $X2=0 $Y2=0
cc_258 N_B1_M1010_g N_VPWR_c_508_n 0.00435301f $X=3.015 $Y=2.46 $X2=0 $Y2=0
cc_259 N_B1_M1011_g N_VPWR_c_508_n 0.00431552f $X=3.535 $Y=2.46 $X2=0 $Y2=0
cc_260 B1 N_X_c_606_n 0.00210779f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_261 N_B1_M1010_g N_A_529_392#_c_660_n 0.00114413f $X=3.015 $Y=2.46 $X2=0
+ $Y2=0
cc_262 N_B1_M1010_g N_A_529_392#_c_661_n 0.0113795f $X=3.015 $Y=2.46 $X2=0 $Y2=0
cc_263 N_B1_M1011_g N_A_529_392#_c_661_n 8.03016e-19 $X=3.535 $Y=2.46 $X2=0
+ $Y2=0
cc_264 B1 N_A_529_392#_c_661_n 0.0244395f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_265 N_B1_c_274_n N_A_529_392#_c_661_n 0.00730446f $X=3.37 $Y=1.635 $X2=0
+ $Y2=0
cc_266 N_B1_M1010_g N_A_529_392#_c_662_n 0.0127709f $X=3.015 $Y=2.46 $X2=0 $Y2=0
cc_267 N_B1_M1011_g N_A_529_392#_c_662_n 0.013657f $X=3.535 $Y=2.46 $X2=0 $Y2=0
cc_268 N_B1_M1011_g N_A_529_392#_c_663_n 0.00150244f $X=3.535 $Y=2.46 $X2=0
+ $Y2=0
cc_269 N_B1_M1011_g N_A_529_392#_c_664_n 0.00883593f $X=3.535 $Y=2.46 $X2=0
+ $Y2=0
cc_270 N_B1_M1002_g N_VGND_c_753_n 0.00277984f $X=2.87 $Y=0.69 $X2=0 $Y2=0
cc_271 N_B1_M1002_g N_VGND_c_754_n 0.0114424f $X=2.87 $Y=0.69 $X2=0 $Y2=0
cc_272 N_B1_M1007_g N_VGND_c_754_n 0.00513027f $X=3.37 $Y=0.69 $X2=0 $Y2=0
cc_273 N_B1_M1002_g N_VGND_c_758_n 0.00383152f $X=2.87 $Y=0.69 $X2=0 $Y2=0
cc_274 N_B1_M1007_g N_VGND_c_759_n 0.00434272f $X=3.37 $Y=0.69 $X2=0 $Y2=0
cc_275 N_B1_M1002_g N_VGND_c_761_n 0.00762539f $X=2.87 $Y=0.69 $X2=0 $Y2=0
cc_276 N_B1_M1007_g N_VGND_c_761_n 0.00820816f $X=3.37 $Y=0.69 $X2=0 $Y2=0
cc_277 N_A1_M1022_g N_A2_M1004_g 0.0120715f $X=4.685 $Y=2.46 $X2=0 $Y2=0
cc_278 N_A1_c_335_n N_A2_c_399_n 0.00309966f $X=4.21 $Y=1.45 $X2=0 $Y2=0
cc_279 A1 N_A2_c_403_n 2.91215e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_280 N_A1_c_339_n N_A2_c_403_n 0.0183213f $X=4.685 $Y=1.615 $X2=0 $Y2=0
cc_281 N_A1_c_337_n N_A2_c_404_n 0.00309966f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_282 A1 N_A2_c_406_n 0.0219354f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_283 N_A1_c_339_n N_A2_c_406_n 0.00312586f $X=4.685 $Y=1.615 $X2=0 $Y2=0
cc_284 N_A1_M1000_g N_VPWR_c_513_n 0.00343682f $X=4.135 $Y=2.46 $X2=0 $Y2=0
cc_285 N_A1_M1022_g N_VPWR_c_513_n 0.00203999f $X=4.685 $Y=2.46 $X2=0 $Y2=0
cc_286 N_A1_M1000_g N_VPWR_c_516_n 0.00519767f $X=4.135 $Y=2.46 $X2=0 $Y2=0
cc_287 N_A1_M1022_g N_VPWR_c_518_n 0.005209f $X=4.685 $Y=2.46 $X2=0 $Y2=0
cc_288 N_A1_M1000_g N_VPWR_c_508_n 0.0098022f $X=4.135 $Y=2.46 $X2=0 $Y2=0
cc_289 N_A1_M1022_g N_VPWR_c_508_n 0.00982636f $X=4.685 $Y=2.46 $X2=0 $Y2=0
cc_290 N_A1_M1000_g N_A_529_392#_c_663_n 0.00101935f $X=4.135 $Y=2.46 $X2=0
+ $Y2=0
cc_291 A1 N_A_529_392#_c_663_n 0.00947167f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_292 N_A1_M1000_g N_A_529_392#_c_664_n 0.0120075f $X=4.135 $Y=2.46 $X2=0 $Y2=0
cc_293 N_A1_M1022_g N_A_529_392#_c_664_n 4.92553e-19 $X=4.685 $Y=2.46 $X2=0
+ $Y2=0
cc_294 N_A1_M1000_g N_A_529_392#_c_665_n 0.0134861f $X=4.135 $Y=2.46 $X2=0 $Y2=0
cc_295 N_A1_M1022_g N_A_529_392#_c_665_n 0.0143281f $X=4.685 $Y=2.46 $X2=0 $Y2=0
cc_296 A1 N_A_529_392#_c_665_n 0.0442019f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_297 N_A1_c_339_n N_A_529_392#_c_665_n 0.0044963f $X=4.685 $Y=1.615 $X2=0
+ $Y2=0
cc_298 N_A1_M1000_g N_A_529_392#_c_666_n 5.28651e-19 $X=4.135 $Y=2.46 $X2=0
+ $Y2=0
cc_299 N_A1_M1022_g N_A_529_392#_c_666_n 0.0119155f $X=4.685 $Y=2.46 $X2=0 $Y2=0
cc_300 N_A1_M1022_g N_A_529_392#_c_672_n 0.00191681f $X=4.685 $Y=2.46 $X2=0
+ $Y2=0
cc_301 N_A1_c_332_n N_VGND_c_759_n 0.00434272f $X=3.8 $Y=1.085 $X2=0 $Y2=0
cc_302 N_A1_c_336_n N_VGND_c_759_n 0.00278247f $X=4.3 $Y=1.085 $X2=0 $Y2=0
cc_303 N_A1_c_332_n N_VGND_c_761_n 0.00822026f $X=3.8 $Y=1.085 $X2=0 $Y2=0
cc_304 N_A1_c_336_n N_VGND_c_761_n 0.00359084f $X=4.3 $Y=1.085 $X2=0 $Y2=0
cc_305 N_A1_c_333_n N_A_775_74#_c_842_n 0.00414859f $X=4.045 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A1_c_336_n N_A_775_74#_c_842_n 0.0113332f $X=4.3 $Y=1.085 $X2=0 $Y2=0
cc_307 N_A1_c_336_n N_A_775_74#_c_840_n 0.0121116f $X=4.3 $Y=1.085 $X2=0 $Y2=0
cc_308 N_A1_c_332_n N_A_775_74#_c_841_n 0.00215418f $X=3.8 $Y=1.085 $X2=0 $Y2=0
cc_309 N_A1_c_336_n N_A_775_74#_c_841_n 0.00188363f $X=4.3 $Y=1.085 $X2=0 $Y2=0
cc_310 N_A1_c_337_n N_A_1000_74#_c_869_n 4.09982e-19 $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A2_M1023_g N_A3_M1020_g 0.0129282f $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_312 N_A2_M1017_g N_A3_M1003_g 0.0249921f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_313 N_A2_c_405_n A3 4.05423e-19 $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_314 N_A2_c_406_n A3 0.0203396f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_315 N_A2_c_405_n N_A3_c_470_n 0.0187073f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_316 N_A2_c_406_n N_A3_c_470_n 0.00139133f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_317 N_A2_M1004_g N_VPWR_c_514_n 0.0020575f $X=5.135 $Y=2.46 $X2=0 $Y2=0
cc_318 N_A2_M1023_g N_VPWR_c_514_n 0.00341126f $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_319 N_A2_M1023_g N_VPWR_c_515_n 6.9941e-19 $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_320 N_A2_M1004_g N_VPWR_c_518_n 0.005209f $X=5.135 $Y=2.46 $X2=0 $Y2=0
cc_321 N_A2_M1023_g N_VPWR_c_522_n 0.005209f $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_322 N_A2_M1004_g N_VPWR_c_508_n 0.0098272f $X=5.135 $Y=2.46 $X2=0 $Y2=0
cc_323 N_A2_M1023_g N_VPWR_c_508_n 0.009834f $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_324 N_A2_M1004_g N_A_529_392#_c_666_n 0.0118459f $X=5.135 $Y=2.46 $X2=0 $Y2=0
cc_325 N_A2_M1023_g N_A_529_392#_c_666_n 7.71767e-19 $X=5.695 $Y=2.46 $X2=0
+ $Y2=0
cc_326 N_A2_M1004_g N_A_529_392#_c_667_n 0.0135339f $X=5.135 $Y=2.46 $X2=0 $Y2=0
cc_327 N_A2_c_400_n N_A_529_392#_c_667_n 0.00448411f $X=5.605 $Y=1.615 $X2=0
+ $Y2=0
cc_328 N_A2_M1023_g N_A_529_392#_c_667_n 0.0135339f $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_329 N_A2_c_406_n N_A_529_392#_c_667_n 0.0498434f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_330 N_A2_M1004_g N_A_529_392#_c_668_n 7.79605e-19 $X=5.135 $Y=2.46 $X2=0
+ $Y2=0
cc_331 N_A2_M1023_g N_A_529_392#_c_668_n 0.0120093f $X=5.695 $Y=2.46 $X2=0 $Y2=0
cc_332 N_A2_M1004_g N_A_529_392#_c_672_n 0.00100213f $X=5.135 $Y=2.46 $X2=0
+ $Y2=0
cc_333 N_A2_c_406_n N_A_529_392#_c_672_n 0.0130101f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_334 N_A2_M1023_g N_A_529_392#_c_673_n 0.00101745f $X=5.695 $Y=2.46 $X2=0
+ $Y2=0
cc_335 N_A2_c_405_n N_A_529_392#_c_673_n 0.00217919f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_336 N_A2_c_406_n N_A_529_392#_c_673_n 0.00914141f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_337 N_A2_M1017_g N_VGND_c_755_n 5.42935e-19 $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_338 N_A2_c_401_n N_VGND_c_759_n 0.00278247f $X=5.36 $Y=1.085 $X2=0 $Y2=0
cc_339 N_A2_M1017_g N_VGND_c_759_n 0.00430908f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_340 N_A2_c_401_n N_VGND_c_761_n 0.00358425f $X=5.36 $Y=1.085 $X2=0 $Y2=0
cc_341 N_A2_M1017_g N_VGND_c_761_n 0.00816766f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_342 N_A2_c_401_n N_A_775_74#_c_840_n 0.0139866f $X=5.36 $Y=1.085 $X2=0 $Y2=0
cc_343 N_A2_M1017_g N_A_775_74#_c_840_n 0.00393174f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_344 N_A2_c_404_n N_A_775_74#_c_840_n 4.0436e-19 $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A2_c_401_n N_A_775_74#_c_854_n 0.0114072f $X=5.36 $Y=1.085 $X2=0 $Y2=0
cc_346 N_A2_M1017_g N_A_775_74#_c_854_n 0.00564547f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_347 N_A2_c_401_n N_A_1000_74#_c_867_n 0.00406074f $X=5.36 $Y=1.085 $X2=0
+ $Y2=0
cc_348 N_A2_c_404_n N_A_1000_74#_c_867_n 0.00442645f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A2_c_400_n N_A_1000_74#_c_868_n 0.00530999f $X=5.605 $Y=1.615 $X2=0
+ $Y2=0
cc_350 N_A2_M1017_g N_A_1000_74#_c_868_n 0.0148277f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_351 N_A2_c_404_n N_A_1000_74#_c_868_n 0.0133304f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A2_c_406_n N_A_1000_74#_c_868_n 0.0470905f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_353 N_A2_c_399_n N_A_1000_74#_c_869_n 0.00335202f $X=5.15 $Y=1.45 $X2=0 $Y2=0
cc_354 N_A2_c_404_n N_A_1000_74#_c_869_n 0.00347692f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_355 N_A2_c_406_n N_A_1000_74#_c_869_n 0.0207735f $X=5.7 $Y=1.615 $X2=0 $Y2=0
cc_356 N_A2_M1017_g N_A_1000_74#_c_870_n 0.00248673f $X=5.79 $Y=0.69 $X2=0 $Y2=0
cc_357 N_A3_M1020_g N_VPWR_c_515_n 0.0124389f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_358 N_A3_M1021_g N_VPWR_c_515_n 0.00334717f $X=6.695 $Y=2.46 $X2=0 $Y2=0
cc_359 N_A3_M1020_g N_VPWR_c_522_n 0.00460063f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_360 N_A3_M1021_g N_VPWR_c_523_n 0.005209f $X=6.695 $Y=2.46 $X2=0 $Y2=0
cc_361 N_A3_M1020_g N_VPWR_c_508_n 0.00909121f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_362 N_A3_M1021_g N_VPWR_c_508_n 0.00985824f $X=6.695 $Y=2.46 $X2=0 $Y2=0
cc_363 N_A3_M1020_g N_A_529_392#_c_669_n 0.0147935f $X=6.195 $Y=2.46 $X2=0 $Y2=0
cc_364 N_A3_M1021_g N_A_529_392#_c_669_n 0.0132272f $X=6.695 $Y=2.46 $X2=0 $Y2=0
cc_365 A3 N_A_529_392#_c_669_n 0.0468712f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_366 N_A3_c_470_n N_A_529_392#_c_669_n 0.00329647f $X=6.695 $Y=1.615 $X2=0
+ $Y2=0
cc_367 N_A3_M1021_g N_A_529_392#_c_670_n 0.00108119f $X=6.695 $Y=2.46 $X2=0
+ $Y2=0
cc_368 A3 N_A_529_392#_c_670_n 0.0280486f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_369 N_A3_M1020_g N_A_529_392#_c_671_n 5.59637e-19 $X=6.195 $Y=2.46 $X2=0
+ $Y2=0
cc_370 N_A3_M1021_g N_A_529_392#_c_671_n 0.0119802f $X=6.695 $Y=2.46 $X2=0 $Y2=0
cc_371 N_A3_M1003_g N_VGND_c_755_n 0.0104218f $X=6.22 $Y=0.69 $X2=0 $Y2=0
cc_372 N_A3_M1016_g N_VGND_c_755_n 0.013474f $X=6.65 $Y=0.69 $X2=0 $Y2=0
cc_373 N_A3_M1003_g N_VGND_c_759_n 0.00383152f $X=6.22 $Y=0.69 $X2=0 $Y2=0
cc_374 N_A3_M1016_g N_VGND_c_760_n 0.00383152f $X=6.65 $Y=0.69 $X2=0 $Y2=0
cc_375 N_A3_M1003_g N_VGND_c_761_n 0.00757637f $X=6.22 $Y=0.69 $X2=0 $Y2=0
cc_376 N_A3_M1016_g N_VGND_c_761_n 0.00761372f $X=6.65 $Y=0.69 $X2=0 $Y2=0
cc_377 N_A3_M1003_g N_A_775_74#_c_840_n 3.00542e-19 $X=6.22 $Y=0.69 $X2=0 $Y2=0
cc_378 N_A3_M1003_g N_A_1000_74#_c_870_n 0.00248702f $X=6.22 $Y=0.69 $X2=0 $Y2=0
cc_379 N_A3_M1003_g N_A_1000_74#_c_871_n 0.0142932f $X=6.22 $Y=0.69 $X2=0 $Y2=0
cc_380 N_A3_M1016_g N_A_1000_74#_c_871_n 0.0157274f $X=6.65 $Y=0.69 $X2=0 $Y2=0
cc_381 A3 N_A_1000_74#_c_871_n 0.070916f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_382 N_A3_c_470_n N_A_1000_74#_c_871_n 0.00492955f $X=6.695 $Y=1.615 $X2=0
+ $Y2=0
cc_383 N_A3_M1016_g N_A_1000_74#_c_872_n 0.00446473f $X=6.65 $Y=0.69 $X2=0 $Y2=0
cc_384 N_VPWR_M1005_s N_X_c_606_n 0.00274845f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_385 N_VPWR_c_511_n N_X_c_606_n 0.0208278f $X=1.23 $Y=2.145 $X2=0 $Y2=0
cc_386 N_VPWR_c_512_n N_X_c_606_n 0.00374248f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_387 N_VPWR_c_511_n N_X_c_607_n 0.0353111f $X=1.23 $Y=2.145 $X2=0 $Y2=0
cc_388 N_VPWR_c_512_n N_X_c_607_n 0.0416523f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_389 N_VPWR_c_521_n N_X_c_607_n 0.0144623f $X=2.065 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_c_508_n N_X_c_607_n 0.0118344f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_c_510_n X 0.0395357f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_392 N_VPWR_c_511_n X 0.0353111f $X=1.23 $Y=2.145 $X2=0 $Y2=0
cc_393 N_VPWR_c_520_n X 0.0144623f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_c_508_n X 0.0118344f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_c_512_n N_A_529_392#_c_660_n 0.0121617f $X=2.23 $Y=1.985 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_516_n N_A_529_392#_c_660_n 0.0146352f $X=4.245 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_508_n N_A_529_392#_c_660_n 0.0120433f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_512_n N_A_529_392#_c_661_n 0.0565981f $X=2.23 $Y=1.985 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_516_n N_A_529_392#_c_662_n 0.0310297f $X=4.245 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_508_n N_A_529_392#_c_662_n 0.0263528f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_513_n N_A_529_392#_c_664_n 0.0079549f $X=4.41 $Y=2.425 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_516_n N_A_529_392#_c_664_n 0.0146352f $X=4.245 $Y=3.33 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_508_n N_A_529_392#_c_664_n 0.0120433f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_M1000_d N_A_529_392#_c_665_n 0.00280934f $X=4.225 $Y=1.96 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_513_n N_A_529_392#_c_665_n 0.0208278f $X=4.41 $Y=2.425 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_513_n N_A_529_392#_c_666_n 0.0266809f $X=4.41 $Y=2.425 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_514_n N_A_529_392#_c_666_n 0.0266809f $X=5.41 $Y=2.425 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_518_n N_A_529_392#_c_666_n 0.0144623f $X=5.245 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_508_n N_A_529_392#_c_666_n 0.0118344f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_M1004_d N_A_529_392#_c_667_n 0.00300365f $X=5.225 $Y=1.96 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_514_n N_A_529_392#_c_667_n 0.0216414f $X=5.41 $Y=2.425 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_514_n N_A_529_392#_c_668_n 0.0254897f $X=5.41 $Y=2.425 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_515_n N_A_529_392#_c_668_n 0.0266809f $X=6.42 $Y=2.425 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_522_n N_A_529_392#_c_668_n 0.014549f $X=6.255 $Y=3.33 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_508_n N_A_529_392#_c_668_n 0.0119743f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_416 N_VPWR_M1020_s N_A_529_392#_c_669_n 0.00218982f $X=6.285 $Y=1.96 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_515_n N_A_529_392#_c_669_n 0.0189268f $X=6.42 $Y=2.425 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_515_n N_A_529_392#_c_671_n 0.0266809f $X=6.42 $Y=2.425 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_523_n N_A_529_392#_c_671_n 0.014549f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_508_n N_A_529_392#_c_671_n 0.0119743f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_X_c_611_n N_VGND_M1013_s 0.00346908f $X=1.555 $Y=0.915 $X2=0 $Y2=0
cc_422 N_X_c_603_n N_VGND_c_751_n 0.01819f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_423 N_X_c_605_n N_VGND_c_751_n 0.00612485f $X=0.73 $Y=1.55 $X2=0 $Y2=0
cc_424 N_X_c_603_n N_VGND_c_752_n 0.0118388f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_425 N_X_c_611_n N_VGND_c_752_n 0.0166873f $X=1.555 $Y=0.915 $X2=0 $Y2=0
cc_426 N_X_c_604_n N_VGND_c_752_n 0.0132369f $X=1.64 $Y=0.495 $X2=0 $Y2=0
cc_427 N_X_c_611_n N_VGND_c_753_n 0.0092903f $X=1.555 $Y=0.915 $X2=0 $Y2=0
cc_428 N_X_c_604_n N_VGND_c_753_n 0.0319798f $X=1.64 $Y=0.495 $X2=0 $Y2=0
cc_429 N_X_c_603_n N_VGND_c_756_n 0.011066f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_430 N_X_c_604_n N_VGND_c_757_n 0.00814007f $X=1.64 $Y=0.495 $X2=0 $Y2=0
cc_431 N_X_c_603_n N_VGND_c_761_n 0.00915947f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_432 N_X_c_611_n N_VGND_c_761_n 0.0117746f $X=1.555 $Y=0.915 $X2=0 $Y2=0
cc_433 N_X_c_604_n N_VGND_c_761_n 0.00627537f $X=1.64 $Y=0.495 $X2=0 $Y2=0
cc_434 N_A_529_392#_c_673_n N_A_1000_74#_c_868_n 0.00176228f $X=5.92 $Y=2.115
+ $X2=0 $Y2=0
cc_435 N_A_529_392#_c_669_n N_A_1000_74#_c_871_n 6.68628e-19 $X=6.755 $Y=2.035
+ $X2=0 $Y2=0
cc_436 N_A_529_392#_c_673_n N_A_1000_74#_c_873_n 0.00589499f $X=5.92 $Y=2.115
+ $X2=0 $Y2=0
cc_437 N_VGND_c_755_n N_A_775_74#_c_840_n 0.0029789f $X=6.435 $Y=0.495 $X2=0
+ $Y2=0
cc_438 N_VGND_c_759_n N_A_775_74#_c_840_n 0.0974389f $X=6.27 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_761_n N_A_775_74#_c_840_n 0.0550722f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_754_n N_A_775_74#_c_841_n 0.00314463f $X=3.085 $Y=0.495 $X2=0
+ $Y2=0
cc_441 N_VGND_c_759_n N_A_775_74#_c_841_n 0.0235818f $X=6.27 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_c_761_n N_A_775_74#_c_841_n 0.0127177f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_755_n N_A_1000_74#_c_870_n 0.0218329f $X=6.435 $Y=0.495 $X2=0
+ $Y2=0
cc_444 N_VGND_c_759_n N_A_1000_74#_c_870_n 0.00749631f $X=6.27 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_761_n N_A_1000_74#_c_870_n 0.0062048f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_755_n N_A_1000_74#_c_871_n 0.0216087f $X=6.435 $Y=0.495 $X2=0
+ $Y2=0
cc_447 N_VGND_c_755_n N_A_1000_74#_c_872_n 0.0218743f $X=6.435 $Y=0.495 $X2=0
+ $Y2=0
cc_448 N_VGND_c_760_n N_A_1000_74#_c_872_n 0.011066f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_761_n N_A_1000_74#_c_872_n 0.00915947f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_450 N_A_775_74#_c_840_n N_A_1000_74#_M1006_s 0.00261961f $X=5.41 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_451 N_A_775_74#_c_840_n N_A_1000_74#_c_867_n 0.0188656f $X=5.41 $Y=0.34 $X2=0
+ $Y2=0
cc_452 N_A_775_74#_c_854_n N_A_1000_74#_c_868_n 0.021619f $X=5.575 $Y=0.495
+ $X2=0 $Y2=0
cc_453 N_A_775_74#_c_840_n N_A_1000_74#_c_870_n 0.00370621f $X=5.41 $Y=0.34
+ $X2=0 $Y2=0

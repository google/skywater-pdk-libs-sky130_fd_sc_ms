* NGSPICE file created from sky130_fd_sc_ms__a2bb2oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_126_112# A1_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=8.322e+11p ps=6.72e+06u
M1001 Y a_126_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1002 a_126_112# A2_N a_120_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1003 VGND B1 a_488_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1004 a_402_368# a_126_112# Y VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=2.912e+11p ps=2.76e+06u
M1005 a_402_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.96e+11p ps=5.36e+06u
M1006 VPWR B2 a_402_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_488_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_120_392# A1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2_N a_126_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


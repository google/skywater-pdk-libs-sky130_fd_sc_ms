* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor3_1 A B C VGND VNB VPB VPWR X
M1000 a_81_268# C a_363_394# VPB pshort w=840000u l=180000u
+  ad=3.9275e+11p pd=2.79e+06u as=5.184e+11p ps=4.63e+06u
M1001 a_786_100# B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.0267e+12p ps=7.95e+06u
M1002 a_786_100# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.212e+12p ps=9e+06u
M1003 VGND a_81_268# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1004 a_1116_383# B a_371_74# VNB nlowvt w=640000u l=150000u
+  ad=4.096e+11p pd=3.95e+06u as=4.48e+11p ps=3.96e+06u
M1005 a_1116_383# a_897_54# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_363_394# a_232_162# a_81_268# VNB nlowvt w=640000u l=150000u
+  ad=4.271e+11p pd=3.96e+06u as=2.24e+11p ps=1.98e+06u
M1007 a_371_74# a_786_100# a_897_54# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.95425e+11p ps=4.74e+06u
M1008 a_81_268# C a_371_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_363_394# a_786_100# a_897_54# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=6.9725e+11p ps=5.56e+06u
M1010 a_1116_383# B a_363_394# VPB pshort w=640000u l=180000u
+  ad=4.578e+11p pd=4.39e+06u as=0p ps=0u
M1011 a_1116_383# a_897_54# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_371_74# a_786_100# a_1116_383# VPB pshort w=640000u l=180000u
+  ad=5.792e+11p pd=4.82e+06u as=0p ps=0u
M1013 a_232_162# C VGND VNB nlowvt w=420000u l=150000u
+  ad=1.575e+11p pd=1.59e+06u as=0p ps=0u
M1014 a_897_54# B a_363_394# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_897_54# B a_371_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_81_268# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1017 VGND A a_897_54# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_232_162# C VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1019 a_371_74# a_232_162# a_81_268# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_897_54# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_363_394# a_786_100# a_1116_383# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__a311oi_1.pxi.spice
* Created: Wed Sep  2 11:54:42 2020
* 
x_PM_SKY130_FD_SC_MS__A311OI_1%A3 N_A3_M1007_g N_A3_c_62_n N_A3_M1005_g
+ N_A3_c_63_n N_A3_c_64_n A3 A3 PM_SKY130_FD_SC_MS__A311OI_1%A3
x_PM_SKY130_FD_SC_MS__A311OI_1%A2 N_A2_M1001_g N_A2_M1008_g A2 N_A2_c_91_n
+ N_A2_c_92_n PM_SKY130_FD_SC_MS__A311OI_1%A2
x_PM_SKY130_FD_SC_MS__A311OI_1%A1 N_A1_M1006_g N_A1_M1000_g A1 N_A1_c_129_n
+ N_A1_c_130_n PM_SKY130_FD_SC_MS__A311OI_1%A1
x_PM_SKY130_FD_SC_MS__A311OI_1%B1 N_B1_M1009_g N_B1_M1003_g B1 B1 N_B1_c_165_n
+ PM_SKY130_FD_SC_MS__A311OI_1%B1
x_PM_SKY130_FD_SC_MS__A311OI_1%C1 N_C1_M1004_g N_C1_M1002_g N_C1_c_197_n C1
+ N_C1_c_198_n N_C1_c_199_n PM_SKY130_FD_SC_MS__A311OI_1%C1
x_PM_SKY130_FD_SC_MS__A311OI_1%VPWR N_VPWR_M1007_s N_VPWR_M1008_d N_VPWR_c_227_n
+ N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_232_n
+ VPWR N_VPWR_c_233_n N_VPWR_c_226_n PM_SKY130_FD_SC_MS__A311OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A311OI_1%A_159_368# N_A_159_368#_M1007_d
+ N_A_159_368#_M1000_d N_A_159_368#_c_264_n N_A_159_368#_c_261_n
+ N_A_159_368#_c_262_n PM_SKY130_FD_SC_MS__A311OI_1%A_159_368#
x_PM_SKY130_FD_SC_MS__A311OI_1%Y N_Y_M1006_d N_Y_M1004_d N_Y_M1002_d N_Y_c_289_n
+ N_Y_c_301_n N_Y_c_307_n N_Y_c_302_n N_Y_c_290_n N_Y_c_291_n N_Y_c_295_n
+ N_Y_c_296_n Y Y N_Y_c_292_n N_Y_c_293_n PM_SKY130_FD_SC_MS__A311OI_1%Y
x_PM_SKY130_FD_SC_MS__A311OI_1%VGND N_VGND_M1005_s N_VGND_M1009_d N_VGND_c_361_n
+ N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n
+ VGND N_VGND_c_367_n N_VGND_c_368_n PM_SKY130_FD_SC_MS__A311OI_1%VGND
cc_1 VNB N_A3_M1007_g 0.00560732f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_2 VNB N_A3_c_62_n 0.0197654f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.22
cc_3 VNB N_A3_c_63_n 0.0534421f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_4 VNB N_A3_c_64_n 0.0105651f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_5 VNB A3 0.0295507f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A2_M1001_g 0.0244269f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_7 VNB N_A2_c_91_n 0.026255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_92_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_M1006_g 0.0268314f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_10 VNB N_A1_c_129_n 0.0262338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_130_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1009_g 0.0261863f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_13 VNB B1 0.00423229f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_B1_c_165_n 0.0216755f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_15 VNB N_C1_M1004_g 0.0345407f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_16 VNB N_C1_c_197_n 0.00984469f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_C1_c_198_n 0.0439496f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_18 VNB N_C1_c_199_n 0.00813406f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_19 VNB N_VPWR_c_226_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_289_n 0.00348446f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_Y_c_290_n 0.0134556f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_22 VNB N_Y_c_291_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_292_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_293_n 0.0242391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_361_n 0.0285265f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_26 VNB N_VGND_c_362_n 0.00685406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_363_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.385
cc_28 VNB N_VGND_c_364_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_365_n 0.0411805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_366_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_367_n 0.0244021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_368_n 0.225214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A3_M1007_g 0.0249909f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_34 VPB A3 0.0162107f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_35 VPB N_A2_M1008_g 0.0228477f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_36 VPB N_A2_c_91_n 0.0055922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A2_c_92_n 0.00271794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A1_M1000_g 0.0234277f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_39 VPB N_A1_c_129_n 0.00561629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A1_c_130_n 0.00208354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_B1_M1003_g 0.0215351f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_42 VPB B1 0.00446509f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB N_B1_c_165_n 0.00539277f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_44 VPB N_C1_M1002_g 0.0276459f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_45 VPB N_C1_c_197_n 5.8517e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_46 VPB N_C1_c_198_n 0.0145157f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_47 VPB N_C1_c_199_n 0.0117191f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_48 VPB N_VPWR_c_227_n 0.0379948f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.385
cc_49 VPB N_VPWR_c_228_n 0.0105998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_229_n 0.0121672f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_51 VPB N_VPWR_c_230_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_231_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_232_n 0.00786036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_233_n 0.0506387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_226_n 0.0814749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_159_368#_c_261_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_57 VPB N_A_159_368#_c_262_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.385
cc_58 VPB N_Y_c_289_n 0.00133119f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_59 VPB N_Y_c_295_n 0.00743317f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_60 VPB N_Y_c_296_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_A3_c_62_n N_A2_M1001_g 0.0431007f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A3_M1007_g N_A2_M1008_g 0.0319382f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A3_c_64_n N_A2_c_91_n 0.0431007f $X=0.705 $Y=1.385 $X2=0 $Y2=0
cc_64 N_A3_M1007_g N_A2_c_92_n 3.16626e-19 $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_65 N_A3_c_64_n N_A2_c_92_n 3.7927e-19 $X=0.705 $Y=1.385 $X2=0 $Y2=0
cc_66 N_A3_M1007_g N_VPWR_c_227_n 0.00501904f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_67 A3 N_VPWR_c_227_n 0.00741364f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A3_M1007_g N_VPWR_c_231_n 0.005209f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A3_M1007_g N_VPWR_c_226_n 0.00986641f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A3_M1007_g N_A_159_368#_c_261_n 0.00971514f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_71 N_A3_M1007_g N_Y_c_289_n 0.0139572f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A3_c_62_n N_Y_c_289_n 7.61601e-19 $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_73 N_A3_c_64_n N_Y_c_289_n 0.0093363f $X=0.705 $Y=1.385 $X2=0 $Y2=0
cc_74 A3 N_Y_c_289_n 0.0442649f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A3_c_62_n N_Y_c_301_n 0.0174993f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_76 N_A3_M1007_g N_Y_c_302_n 0.0170159f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A3_c_62_n N_Y_c_293_n 0.00235309f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_78 N_A3_c_62_n N_VGND_c_361_n 0.0158743f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_79 N_A3_c_63_n N_VGND_c_361_n 0.00537271f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_80 A3 N_VGND_c_361_n 0.0085354f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A3_c_62_n N_VGND_c_365_n 0.00383152f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_82 N_A3_c_62_n N_VGND_c_368_n 0.0075694f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A2_M1001_g N_A1_M1006_g 0.0343434f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A2_M1008_g N_A1_M1000_g 0.0338588f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A2_c_92_n N_A1_M1000_g 2.93655e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A2_c_91_n N_A1_c_129_n 0.0201104f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A2_c_92_n N_A1_c_129_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A2_M1008_g N_A1_c_130_n 3.33652e-19 $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A2_c_91_n N_A1_c_130_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_90 N_A2_c_92_n N_A1_c_130_n 0.0280927f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A2_M1008_g N_VPWR_c_228_n 0.00603141f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A2_M1008_g N_VPWR_c_231_n 0.005209f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A2_M1008_g N_VPWR_c_226_n 0.00983279f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A2_M1008_g N_A_159_368#_c_264_n 0.0135335f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A2_M1008_g N_A_159_368#_c_261_n 0.0092369f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A2_M1008_g N_A_159_368#_c_262_n 8.09876e-19 $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A2_M1001_g N_Y_c_289_n 0.0051053f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A2_M1008_g N_Y_c_289_n 0.00173837f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A2_c_92_n N_Y_c_289_n 0.0327278f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A2_M1008_g N_Y_c_307_n 0.0124538f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A2_c_91_n N_Y_c_307_n 5.96642e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A2_c_92_n N_Y_c_307_n 0.0208858f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A2_M1001_g N_Y_c_292_n 0.00731318f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A2_c_92_n N_Y_c_292_n 0.0268379f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A2_M1001_g N_Y_c_293_n 0.0279819f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A2_c_91_n N_Y_c_293_n 0.00140716f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A2_M1001_g N_VGND_c_361_n 0.00186934f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A2_M1001_g N_VGND_c_365_n 0.00382217f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A2_M1001_g N_VGND_c_368_n 0.00652989f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A1_M1006_g N_B1_M1009_g 0.0215861f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A1_M1000_g N_B1_M1003_g 0.0337279f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A1_c_129_n B1 0.00264603f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_113 N_A1_c_130_n B1 0.0361869f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A1_c_129_n N_B1_c_165_n 0.0206382f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A1_c_130_n N_B1_c_165_n 3.7859e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A1_M1000_g N_VPWR_c_228_n 0.00603141f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A1_M1000_g N_VPWR_c_233_n 0.005209f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A1_M1000_g N_VPWR_c_226_n 0.00983279f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A1_M1000_g N_A_159_368#_c_264_n 0.0135335f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A1_M1000_g N_A_159_368#_c_261_n 8.09876e-19 $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A1_M1000_g N_A_159_368#_c_262_n 0.00922705f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A1_M1000_g N_Y_c_307_n 0.0124265f $X=1.785 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A1_c_129_n N_Y_c_307_n 6.98124e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A1_c_130_n N_Y_c_307_n 0.0229716f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A1_M1006_g N_Y_c_293_n 0.0297967f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A1_c_129_n N_Y_c_293_n 0.00139878f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A1_c_130_n N_Y_c_293_n 0.0275097f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A1_M1006_g N_VGND_c_362_n 6.64319e-19 $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A1_M1006_g N_VGND_c_365_n 0.00291649f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A1_M1006_g N_VGND_c_368_n 0.00361179f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B1_M1009_g N_C1_M1004_g 0.0254529f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B1_M1003_g N_C1_M1002_g 0.0590827f $X=2.235 $Y=2.4 $X2=0 $Y2=0
cc_133 B1 N_C1_M1002_g 0.00488713f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_134 B1 N_C1_c_197_n 0.0136716f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_135 N_B1_c_165_n N_C1_c_197_n 0.021497f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_136 B1 N_C1_c_199_n 0.0346458f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_137 N_B1_M1003_g N_VPWR_c_233_n 0.005209f $X=2.235 $Y=2.4 $X2=0 $Y2=0
cc_138 N_B1_M1003_g N_VPWR_c_226_n 0.00983863f $X=2.235 $Y=2.4 $X2=0 $Y2=0
cc_139 N_B1_M1003_g N_A_159_368#_c_262_n 0.0147202f $X=2.235 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B1_M1003_g N_Y_c_307_n 0.0163421f $X=2.235 $Y=2.4 $X2=0 $Y2=0
cc_141 B1 N_Y_c_307_n 0.0482689f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_142 N_B1_c_165_n N_Y_c_307_n 6.07813e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B1_M1009_g N_Y_c_290_n 0.0153799f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_144 B1 N_Y_c_290_n 0.0544915f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_145 N_B1_c_165_n N_Y_c_290_n 0.00439029f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_146 N_B1_M1009_g N_Y_c_291_n 8.78222e-19 $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_147 N_B1_M1003_g N_Y_c_296_n 0.00286259f $X=2.235 $Y=2.4 $X2=0 $Y2=0
cc_148 N_B1_M1009_g N_Y_c_293_n 0.00384236f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_149 N_B1_M1009_g N_VGND_c_362_n 0.0113145f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_150 N_B1_M1009_g N_VGND_c_365_n 0.00383152f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B1_M1009_g N_VGND_c_368_n 0.00758569f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_152 N_C1_M1002_g N_VPWR_c_233_n 0.005209f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_153 N_C1_M1002_g N_VPWR_c_226_n 0.00987892f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_154 N_C1_M1002_g N_A_159_368#_c_262_n 0.00206182f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_155 N_C1_M1002_g N_Y_c_307_n 0.0136486f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_156 N_C1_M1004_g N_Y_c_290_n 0.0145657f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_157 N_C1_c_197_n N_Y_c_290_n 0.00680871f $X=2.715 $Y=1.515 $X2=0 $Y2=0
cc_158 N_C1_c_198_n N_Y_c_290_n 0.00121887f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_159 N_C1_c_199_n N_Y_c_290_n 0.0132907f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_160 N_C1_M1004_g N_Y_c_291_n 0.0102372f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_161 N_C1_M1002_g N_Y_c_295_n 0.00190089f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_162 N_C1_c_198_n N_Y_c_295_n 0.00467488f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_163 N_C1_c_199_n N_Y_c_295_n 0.0159673f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_164 N_C1_M1002_g N_Y_c_296_n 0.0176177f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_165 N_C1_M1004_g N_VGND_c_362_n 0.00607661f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_166 N_C1_M1004_g N_VGND_c_367_n 0.00434272f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_167 N_C1_M1004_g N_VGND_c_368_n 0.00825192f $X=2.7 $Y=0.74 $X2=0 $Y2=0
cc_168 N_VPWR_M1008_d N_A_159_368#_c_264_n 0.00787899f $X=1.245 $Y=1.84 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_228_n N_A_159_368#_c_264_n 0.0273365f $X=1.47 $Y=2.76 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_227_n N_A_159_368#_c_261_n 0.0177747f $X=0.48 $Y=2.455 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_228_n N_A_159_368#_c_261_n 0.0139497f $X=1.47 $Y=2.76 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_231_n N_A_159_368#_c_261_n 0.0144776f $X=1.265 $Y=3.33 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_226_n N_A_159_368#_c_261_n 0.0118404f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_228_n N_A_159_368#_c_262_n 0.0139497f $X=1.47 $Y=2.76 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_233_n N_A_159_368#_c_262_n 0.0144588f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_226_n N_A_159_368#_c_262_n 0.0118347f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_VPWR_M1008_d N_Y_c_307_n 0.0135816f $X=1.245 $Y=1.84 $X2=0 $Y2=0
cc_178 N_VPWR_c_233_n N_Y_c_296_n 0.014549f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_226_n N_Y_c_296_n 0.0119743f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_180 N_A_159_368#_M1007_d N_Y_c_307_n 0.00753427f $X=0.795 $Y=1.84 $X2=0 $Y2=0
cc_181 N_A_159_368#_M1000_d N_Y_c_307_n 0.00639613f $X=1.875 $Y=1.84 $X2=0 $Y2=0
cc_182 N_A_159_368#_c_264_n N_Y_c_307_n 0.0446711f $X=1.845 $Y=2.375 $X2=0 $Y2=0
cc_183 N_A_159_368#_c_261_n N_Y_c_307_n 0.0149529f $X=0.93 $Y=2.41 $X2=0 $Y2=0
cc_184 N_A_159_368#_c_262_n N_Y_c_307_n 0.0171646f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_185 N_A_159_368#_c_261_n N_Y_c_302_n 0.00249984f $X=0.93 $Y=2.41 $X2=0 $Y2=0
cc_186 N_A_159_368#_c_262_n N_Y_c_296_n 0.0184946f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_187 A_465_368# N_Y_c_307_n 0.0090141f $X=2.325 $Y=1.84 $X2=2.775 $Y2=2.035
cc_188 N_Y_c_290_n N_VGND_M1009_d 0.00309832f $X=2.75 $Y=1.095 $X2=0 $Y2=0
cc_189 N_Y_c_293_n N_VGND_c_361_n 0.0189403f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_190 N_Y_c_290_n N_VGND_c_362_n 0.024241f $X=2.75 $Y=1.095 $X2=0 $Y2=0
cc_191 N_Y_c_291_n N_VGND_c_362_n 0.0191903f $X=2.915 $Y=0.515 $X2=0 $Y2=0
cc_192 N_Y_c_293_n N_VGND_c_362_n 0.0196004f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_193 N_Y_c_293_n N_VGND_c_365_n 0.0417862f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_194 N_Y_c_291_n N_VGND_c_367_n 0.0145639f $X=2.915 $Y=0.515 $X2=0 $Y2=0
cc_195 N_Y_c_291_n N_VGND_c_368_n 0.0119984f $X=2.915 $Y=0.515 $X2=0 $Y2=0
cc_196 N_Y_c_293_n N_VGND_c_368_n 0.0341885f $X=2.04 $Y=0.765 $X2=0 $Y2=0
cc_197 N_Y_c_292_n A_159_74# 0.00366293f $X=1.085 $Y=0.765 $X2=-0.19 $Y2=-0.245
cc_198 N_Y_c_293_n A_231_74# 0.00122878f $X=2.04 $Y=0.765 $X2=-0.19 $Y2=-0.245

* File: sky130_fd_sc_ms__dlxbn_1.pxi.spice
* Created: Fri Aug 28 17:28:44 2020
* 
x_PM_SKY130_FD_SC_MS__DLXBN_1%D N_D_M1020_g N_D_c_143_n N_D_M1000_g N_D_c_149_n
+ D N_D_c_145_n N_D_c_146_n PM_SKY130_FD_SC_MS__DLXBN_1%D
x_PM_SKY130_FD_SC_MS__DLXBN_1%GATE_N N_GATE_N_M1003_g N_GATE_N_M1001_g GATE_N
+ N_GATE_N_c_183_n N_GATE_N_c_186_n PM_SKY130_FD_SC_MS__DLXBN_1%GATE_N
x_PM_SKY130_FD_SC_MS__DLXBN_1%A_232_82# N_A_232_82#_M1003_d N_A_232_82#_M1001_d
+ N_A_232_82#_c_223_n N_A_232_82#_c_224_n N_A_232_82#_M1008_g
+ N_A_232_82#_M1021_g N_A_232_82#_c_226_n N_A_232_82#_M1012_g
+ N_A_232_82#_c_227_n N_A_232_82#_c_228_n N_A_232_82#_M1006_g
+ N_A_232_82#_c_229_n N_A_232_82#_c_230_n N_A_232_82#_c_239_n
+ N_A_232_82#_c_240_n N_A_232_82#_c_231_n N_A_232_82#_c_241_n
+ N_A_232_82#_c_232_n N_A_232_82#_c_243_n N_A_232_82#_c_233_n
+ N_A_232_82#_c_234_n N_A_232_82#_c_235_n N_A_232_82#_c_236_n
+ PM_SKY130_FD_SC_MS__DLXBN_1%A_232_82#
x_PM_SKY130_FD_SC_MS__DLXBN_1%A_27_120# N_A_27_120#_M1020_s N_A_27_120#_M1000_s
+ N_A_27_120#_M1002_g N_A_27_120#_M1013_g N_A_27_120#_c_358_n
+ N_A_27_120#_c_359_n N_A_27_120#_c_360_n N_A_27_120#_c_361_n
+ N_A_27_120#_c_364_n N_A_27_120#_c_362_n PM_SKY130_FD_SC_MS__DLXBN_1%A_27_120#
x_PM_SKY130_FD_SC_MS__DLXBN_1%A_343_80# N_A_343_80#_M1008_s N_A_343_80#_M1021_s
+ N_A_343_80#_M1014_g N_A_343_80#_M1010_g N_A_343_80#_c_431_n
+ N_A_343_80#_c_432_n N_A_343_80#_c_442_n N_A_343_80#_c_443_n
+ N_A_343_80#_c_433_n N_A_343_80#_c_434_n N_A_343_80#_c_435_n
+ N_A_343_80#_c_436_n N_A_343_80#_c_437_n N_A_343_80#_c_438_n
+ N_A_343_80#_c_439_n PM_SKY130_FD_SC_MS__DLXBN_1%A_343_80#
x_PM_SKY130_FD_SC_MS__DLXBN_1%A_863_294# N_A_863_294#_M1005_d
+ N_A_863_294#_M1015_d N_A_863_294#_M1011_g N_A_863_294#_M1004_g
+ N_A_863_294#_M1019_g N_A_863_294#_c_533_n N_A_863_294#_M1009_g
+ N_A_863_294#_M1016_g N_A_863_294#_c_535_n N_A_863_294#_M1017_g
+ N_A_863_294#_c_536_n N_A_863_294#_c_537_n N_A_863_294#_c_548_n
+ N_A_863_294#_c_538_n N_A_863_294#_c_539_n N_A_863_294#_c_550_n
+ N_A_863_294#_c_540_n N_A_863_294#_c_541_n N_A_863_294#_c_542_n
+ N_A_863_294#_c_543_n PM_SKY130_FD_SC_MS__DLXBN_1%A_863_294#
x_PM_SKY130_FD_SC_MS__DLXBN_1%A_653_79# N_A_653_79#_M1012_d N_A_653_79#_M1014_d
+ N_A_653_79#_M1005_g N_A_653_79#_M1015_g N_A_653_79#_c_650_n
+ N_A_653_79#_c_651_n N_A_653_79#_c_652_n N_A_653_79#_c_669_n
+ N_A_653_79#_c_653_n N_A_653_79#_c_654_n N_A_653_79#_c_655_n
+ PM_SKY130_FD_SC_MS__DLXBN_1%A_653_79#
x_PM_SKY130_FD_SC_MS__DLXBN_1%A_1350_424# N_A_1350_424#_M1017_d
+ N_A_1350_424#_M1016_d N_A_1350_424#_M1018_g N_A_1350_424#_M1007_g
+ N_A_1350_424#_c_727_n N_A_1350_424#_c_728_n N_A_1350_424#_c_729_n
+ N_A_1350_424#_c_730_n N_A_1350_424#_c_731_n N_A_1350_424#_c_732_n
+ PM_SKY130_FD_SC_MS__DLXBN_1%A_1350_424#
x_PM_SKY130_FD_SC_MS__DLXBN_1%VPWR N_VPWR_M1000_d N_VPWR_M1021_d N_VPWR_M1011_d
+ N_VPWR_M1019_d N_VPWR_M1018_s N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n
+ N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n
+ N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n VPWR
+ N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_770_n N_VPWR_c_786_n N_VPWR_c_787_n
+ PM_SKY130_FD_SC_MS__DLXBN_1%VPWR
x_PM_SKY130_FD_SC_MS__DLXBN_1%Q N_Q_M1009_s N_Q_M1019_s N_Q_c_861_n N_Q_c_862_n
+ N_Q_c_858_n Q Q Q PM_SKY130_FD_SC_MS__DLXBN_1%Q
x_PM_SKY130_FD_SC_MS__DLXBN_1%Q_N N_Q_N_M1007_d N_Q_N_M1018_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_MS__DLXBN_1%Q_N
x_PM_SKY130_FD_SC_MS__DLXBN_1%VGND N_VGND_M1020_d N_VGND_M1008_d N_VGND_M1004_d
+ N_VGND_M1009_d N_VGND_M1007_s N_VGND_c_908_n N_VGND_c_909_n N_VGND_c_910_n
+ N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n N_VGND_c_914_n VGND
+ N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n
+ N_VGND_c_920_n N_VGND_c_921_n PM_SKY130_FD_SC_MS__DLXBN_1%VGND
cc_1 VNB N_D_c_143_n 0.0164541f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.758
cc_2 VNB D 0.00437541f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_c_145_n 0.0189654f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_4 VNB N_D_c_146_n 0.0222513f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.26
cc_5 VNB N_GATE_N_M1003_g 0.0420743f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.875
cc_6 VNB N_GATE_N_c_183_n 0.00687508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_232_82#_c_223_n 0.016132f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.54
cc_8 VNB N_A_232_82#_c_224_n 0.0226333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_232_82#_M1021_g 0.0140073f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_10 VNB N_A_232_82#_c_226_n 0.0145234f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.26
cc_11 VNB N_A_232_82#_c_227_n 0.0417178f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_12 VNB N_A_232_82#_c_228_n 0.00604536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_232_82#_c_229_n 0.00640516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_232_82#_c_230_n 0.00486834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_232_82#_c_231_n 0.011184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_232_82#_c_232_n 0.0024711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_232_82#_c_233_n 0.0195475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_82#_c_234_n 0.00141834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_232_82#_c_235_n 0.041699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_232_82#_c_236_n 0.0143228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_120#_M1002_g 0.00456957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_120#_M1013_g 0.0223764f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.425
cc_23 VNB N_A_27_120#_c_358_n 0.00895674f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_24 VNB N_A_27_120#_c_359_n 8.28199e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_120#_c_360_n 0.0336675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_120#_c_361_n 0.0239341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_120#_c_362_n 0.0263096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_343_80#_c_431_n 0.00179992f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_29 VNB N_A_343_80#_c_432_n 0.00400209f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_30 VNB N_A_343_80#_c_433_n 0.00444373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_343_80#_c_434_n 0.00239781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_343_80#_c_435_n 0.0146255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_343_80#_c_436_n 0.0454641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_343_80#_c_437_n 0.00326651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_343_80#_c_438_n 0.0168172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_343_80#_c_439_n 0.0199151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_863_294#_M1004_g 0.0369209f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.425
cc_38 VNB N_A_863_294#_M1019_g 0.00394929f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.595
cc_39 VNB N_A_863_294#_c_533_n 0.0204282f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_40 VNB N_A_863_294#_M1016_g 0.00361627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_863_294#_c_535_n 0.0176098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_863_294#_c_536_n 0.050158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_863_294#_c_537_n 0.0509199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_863_294#_c_538_n 0.00721625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_863_294#_c_539_n 0.013466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_863_294#_c_540_n 0.00419193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_863_294#_c_541_n 0.00171367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_863_294#_c_542_n 0.0170976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_863_294#_c_543_n 0.00173151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_653_79#_M1015_g 0.00172196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_653_79#_c_650_n 0.00590375f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_52 VNB N_A_653_79#_c_651_n 0.0222757f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.26
cc_53 VNB N_A_653_79#_c_652_n 0.00557721f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.595
cc_54 VNB N_A_653_79#_c_653_n 0.00455729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_653_79#_c_654_n 0.0349554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_653_79#_c_655_n 0.0218926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1350_424#_M1018_g 0.00221841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1350_424#_M1007_g 0.0293581f $X=-0.19 $Y=-0.245 $X2=0.592
+ $Y2=1.425
cc_59 VNB N_A_1350_424#_c_727_n 0.0466895f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_60 VNB N_A_1350_424#_c_728_n 0.0173848f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.26
cc_61 VNB N_A_1350_424#_c_729_n 0.0113311f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.595
cc_62 VNB N_A_1350_424#_c_730_n 4.1627e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1350_424#_c_731_n 0.00775186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1350_424#_c_732_n 8.96211e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VPWR_c_770_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_858_n 0.00234071f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_67 VNB Q 0.00788781f $X=-0.19 $Y=-0.245 $X2=0.592 $Y2=1.26
cc_68 VNB Q 0.00173648f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.595
cc_69 VNB Q_N 0.0547907f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.54
cc_70 VNB N_VGND_c_908_n 0.0124753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_909_n 0.020983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_910_n 0.0232086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_911_n 0.0519142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_912_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_913_n 0.0347932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_914_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_915_n 0.0194297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_916_n 0.0530251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_917_n 0.0216681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_918_n 0.0192716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_919_n 0.479662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_920_n 0.0208183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_921_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VPB N_D_c_143_n 0.00701196f $X=-0.19 $Y=1.66 $X2=0.592 $Y2=1.758
cc_85 VPB N_D_M1000_g 0.0291989f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.54
cc_86 VPB N_D_c_149_n 0.0179255f $X=-0.19 $Y=1.66 $X2=0.592 $Y2=1.93
cc_87 VPB D 0.00268093f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_88 VPB N_GATE_N_M1001_g 0.0268663f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.54
cc_89 VPB N_GATE_N_c_183_n 0.0272148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_GATE_N_c_186_n 0.00320413f $X=-0.19 $Y=1.66 $X2=0.592 $Y2=1.425
cc_91 VPB N_A_232_82#_M1021_g 0.0339348f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_92 VPB N_A_232_82#_M1006_g 0.0219566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_232_82#_c_239_n 0.0263583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_232_82#_c_240_n 0.00139443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_232_82#_c_241_n 0.0046072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_232_82#_c_232_n 0.0117398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_232_82#_c_243_n 0.0102963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_232_82#_c_233_n 0.0160842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_232_82#_c_234_n 9.52679e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_120#_M1002_g 0.0289716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_120#_c_364_n 0.0506408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_120#_c_362_n 0.0208812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_343_80#_M1014_g 0.0263092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_343_80#_c_432_n 6.37444e-19 $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.595
cc_105 VPB N_A_343_80#_c_442_n 0.00904665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_343_80#_c_443_n 0.00840821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_343_80#_c_437_n 0.0112652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_343_80#_c_438_n 0.0132182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_863_294#_M1011_g 0.0243265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_863_294#_M1019_g 0.0287662f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.595
cc_111 VPB N_A_863_294#_M1016_g 0.0455433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_863_294#_c_536_n 0.0074202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_863_294#_c_548_n 0.00597164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_863_294#_c_539_n 0.0152468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_863_294#_c_550_n 0.0125238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_863_294#_c_541_n 0.00299376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_863_294#_c_542_n 0.0167711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_653_79#_M1015_g 0.0261286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_653_79#_c_650_n 0.00571365f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_120 VPB N_A_1350_424#_M1018_g 0.0308243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_1350_424#_c_730_n 0.0165242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_771_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_772_n 0.0125441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_773_n 0.0561033f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_774_n 0.0401278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_775_n 0.0111271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_776_n 0.0214822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_777_n 0.0218747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_778_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_779_n 0.0355762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_780_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_781_n 0.0200096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_782_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_783_n 0.03922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_784_n 0.0200671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_770_n 0.126489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_786_n 0.00613689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_787_n 0.0103609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_Q_c_861_n 0.011966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_Q_c_862_n 0.00387358f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_141 VPB N_Q_c_858_n 0.00142931f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_142 VPB Q_N 0.0538045f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.54
cc_143 D N_GATE_N_M1003_g 0.00318577f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_144 N_D_c_145_n N_GATE_N_M1003_g 0.0179436f $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_145 N_D_c_146_n N_GATE_N_M1003_g 0.0215568f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_146 N_D_M1000_g N_GATE_N_M1001_g 0.014197f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_147 N_D_c_143_n N_GATE_N_c_183_n 0.0174584f $X=0.592 $Y=1.758 $X2=0 $Y2=0
cc_148 D N_GATE_N_c_183_n 0.00220012f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_149 N_D_c_143_n N_GATE_N_c_186_n 2.63139e-19 $X=0.592 $Y=1.758 $X2=0 $Y2=0
cc_150 N_D_M1000_g N_GATE_N_c_186_n 0.00354458f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_151 N_D_c_149_n N_GATE_N_c_186_n 2.01987e-19 $X=0.592 $Y=1.93 $X2=0 $Y2=0
cc_152 D N_GATE_N_c_186_n 0.019301f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_153 N_D_c_146_n N_A_232_82#_c_230_n 0.00153265f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_154 D N_A_232_82#_c_231_n 0.0143907f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_155 N_D_c_145_n N_A_232_82#_c_231_n 2.43963e-19 $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_156 D N_A_232_82#_c_232_n 0.00518677f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_157 D N_A_27_120#_c_358_n 0.0120455f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_158 N_D_c_145_n N_A_27_120#_c_358_n 0.00373347f $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_159 N_D_c_146_n N_A_27_120#_c_358_n 0.0102926f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_160 D N_A_27_120#_c_361_n 7.4097e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_161 N_D_c_146_n N_A_27_120#_c_361_n 0.0116922f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_162 N_D_M1000_g N_A_27_120#_c_364_n 0.0181023f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_163 N_D_c_149_n N_A_27_120#_c_364_n 0.00369492f $X=0.592 $Y=1.93 $X2=0 $Y2=0
cc_164 D N_A_27_120#_c_364_n 0.00966208f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_165 N_D_M1000_g N_A_27_120#_c_362_n 0.0035594f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_166 D N_A_27_120#_c_362_n 0.0511223f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_167 N_D_c_146_n N_A_27_120#_c_362_n 0.0195681f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_168 N_D_M1000_g N_VPWR_c_771_n 0.0157718f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_169 D N_VPWR_c_771_n 0.00337254f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_170 N_D_M1000_g N_VPWR_c_777_n 0.00460063f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_171 N_D_M1000_g N_VPWR_c_770_n 0.00912759f $X=0.675 $Y=2.54 $X2=0 $Y2=0
cc_172 N_D_c_146_n N_VGND_c_915_n 0.0032796f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_173 N_D_c_146_n N_VGND_c_919_n 0.00476395f $X=0.592 $Y=1.26 $X2=0 $Y2=0
cc_174 N_GATE_N_c_186_n N_A_232_82#_M1001_d 4.575e-19 $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_175 N_GATE_N_M1003_g N_A_232_82#_c_230_n 0.00956489f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_176 N_GATE_N_M1003_g N_A_232_82#_c_231_n 0.00783859f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_177 N_GATE_N_c_183_n N_A_232_82#_c_231_n 0.00471269f $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_178 N_GATE_N_c_186_n N_A_232_82#_c_231_n 0.0158201f $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_179 N_GATE_N_M1001_g N_A_232_82#_c_241_n 0.00310867f $X=1.175 $Y=2.54 $X2=0
+ $Y2=0
cc_180 N_GATE_N_c_183_n N_A_232_82#_c_241_n 2.30408e-19 $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_181 N_GATE_N_c_186_n N_A_232_82#_c_241_n 0.00338538f $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_182 N_GATE_N_M1003_g N_A_232_82#_c_232_n 0.0014664f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_183 N_GATE_N_M1001_g N_A_232_82#_c_232_n 0.00481811f $X=1.175 $Y=2.54 $X2=0
+ $Y2=0
cc_184 N_GATE_N_c_183_n N_A_232_82#_c_232_n 0.00769376f $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_185 N_GATE_N_c_186_n N_A_232_82#_c_232_n 0.035269f $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_186 N_GATE_N_M1001_g N_A_232_82#_c_243_n 0.00579551f $X=1.175 $Y=2.54 $X2=0
+ $Y2=0
cc_187 N_GATE_N_M1003_g N_A_232_82#_c_235_n 0.00858776f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_188 N_GATE_N_M1003_g N_A_27_120#_c_358_n 0.0178682f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_189 N_GATE_N_M1003_g N_A_27_120#_c_361_n 0.00161607f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_186_n N_A_27_120#_c_364_n 0.00140581f $X=1.17 $Y=1.795 $X2=0
+ $Y2=0
cc_191 N_GATE_N_c_186_n N_VPWR_M1000_d 6.41387e-19 $X=1.17 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_192 N_GATE_N_M1001_g N_VPWR_c_771_n 0.00345319f $X=1.175 $Y=2.54 $X2=0 $Y2=0
cc_193 N_GATE_N_c_183_n N_VPWR_c_771_n 2.16117e-19 $X=1.17 $Y=1.795 $X2=0 $Y2=0
cc_194 N_GATE_N_c_186_n N_VPWR_c_771_n 0.00192769f $X=1.17 $Y=1.795 $X2=0 $Y2=0
cc_195 N_GATE_N_M1001_g N_VPWR_c_783_n 0.005209f $X=1.175 $Y=2.54 $X2=0 $Y2=0
cc_196 N_GATE_N_M1001_g N_VPWR_c_770_n 0.00987293f $X=1.175 $Y=2.54 $X2=0 $Y2=0
cc_197 N_GATE_N_M1003_g N_VGND_c_916_n 0.00414982f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_198 N_GATE_N_M1003_g N_VGND_c_919_n 0.00533081f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_199 N_GATE_N_M1003_g N_VGND_c_920_n 0.00546687f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_200 N_A_232_82#_M1021_g N_A_27_120#_M1002_g 0.0402896f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_201 N_A_232_82#_c_239_n N_A_27_120#_M1002_g 0.0131549f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_202 N_A_232_82#_c_224_n N_A_27_120#_M1013_g 0.0237669f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_203 N_A_232_82#_c_226_n N_A_27_120#_M1013_g 0.0246783f $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_204 N_A_232_82#_M1003_d N_A_27_120#_c_358_n 0.00711247f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_205 N_A_232_82#_c_224_n N_A_27_120#_c_358_n 0.0155711f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_206 N_A_232_82#_c_230_n N_A_27_120#_c_358_n 0.0207561f $X=1.3 $Y=1.005 $X2=0
+ $Y2=0
cc_207 N_A_232_82#_c_231_n N_A_27_120#_c_358_n 0.00794673f $X=1.74 $Y=1.415
+ $X2=0 $Y2=0
cc_208 N_A_232_82#_c_235_n N_A_27_120#_c_358_n 0.00257007f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_209 N_A_232_82#_c_224_n N_A_27_120#_c_359_n 0.00648234f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_210 N_A_232_82#_c_226_n N_A_27_120#_c_359_n 5.46252e-19 $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_211 N_A_232_82#_c_229_n N_A_27_120#_c_359_n 0.00100162f $X=2.235 $Y=1.325
+ $X2=0 $Y2=0
cc_212 N_A_232_82#_c_228_n N_A_27_120#_c_360_n 0.0246783f $X=3.265 $Y=1.185
+ $X2=0 $Y2=0
cc_213 N_A_232_82#_c_229_n N_A_27_120#_c_360_n 0.0209442f $X=2.235 $Y=1.325
+ $X2=0 $Y2=0
cc_214 N_A_232_82#_c_239_n N_A_343_80#_M1021_s 0.00751229f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_215 N_A_232_82#_M1006_g N_A_343_80#_M1014_g 0.0115515f $X=3.95 $Y=2.17 $X2=0
+ $Y2=0
cc_216 N_A_232_82#_c_239_n N_A_343_80#_M1014_g 0.0160248f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_217 N_A_232_82#_c_240_n N_A_343_80#_M1014_g 8.44988e-19 $X=4.06 $Y=2.39 $X2=0
+ $Y2=0
cc_218 N_A_232_82#_c_224_n N_A_343_80#_c_431_n 0.00824133f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_219 N_A_232_82#_c_230_n N_A_343_80#_c_431_n 0.0118197f $X=1.3 $Y=1.005 $X2=0
+ $Y2=0
cc_220 N_A_232_82#_c_231_n N_A_343_80#_c_431_n 0.0152496f $X=1.74 $Y=1.415 $X2=0
+ $Y2=0
cc_221 N_A_232_82#_c_235_n N_A_343_80#_c_431_n 0.0106127f $X=1.74 $Y=1.325 $X2=0
+ $Y2=0
cc_222 N_A_232_82#_c_223_n N_A_343_80#_c_432_n 0.00614272f $X=2.145 $Y=1.325
+ $X2=0 $Y2=0
cc_223 N_A_232_82#_c_224_n N_A_343_80#_c_432_n 0.00532923f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_224 N_A_232_82#_M1021_g N_A_343_80#_c_432_n 0.0095182f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_225 N_A_232_82#_c_229_n N_A_343_80#_c_432_n 0.00278586f $X=2.235 $Y=1.325
+ $X2=0 $Y2=0
cc_226 N_A_232_82#_c_230_n N_A_343_80#_c_432_n 0.00541044f $X=1.3 $Y=1.005 $X2=0
+ $Y2=0
cc_227 N_A_232_82#_c_231_n N_A_343_80#_c_432_n 0.0200983f $X=1.74 $Y=1.415 $X2=0
+ $Y2=0
cc_228 N_A_232_82#_c_232_n N_A_343_80#_c_432_n 0.00766455f $X=1.455 $Y=2.32
+ $X2=0 $Y2=0
cc_229 N_A_232_82#_c_235_n N_A_343_80#_c_432_n 8.70862e-19 $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_230 N_A_232_82#_M1021_g N_A_343_80#_c_442_n 0.0160951f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_231 N_A_232_82#_c_239_n N_A_343_80#_c_442_n 0.0257362f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_232 N_A_232_82#_c_223_n N_A_343_80#_c_443_n 0.00456618f $X=2.145 $Y=1.325
+ $X2=0 $Y2=0
cc_233 N_A_232_82#_M1021_g N_A_343_80#_c_443_n 0.0104277f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_234 N_A_232_82#_c_239_n N_A_343_80#_c_443_n 0.0263523f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_235 N_A_232_82#_c_231_n N_A_343_80#_c_443_n 0.00268721f $X=1.74 $Y=1.415
+ $X2=0 $Y2=0
cc_236 N_A_232_82#_c_232_n N_A_343_80#_c_443_n 0.0366456f $X=1.455 $Y=2.32 $X2=0
+ $Y2=0
cc_237 N_A_232_82#_c_235_n N_A_343_80#_c_443_n 0.00129458f $X=1.74 $Y=1.325
+ $X2=0 $Y2=0
cc_238 N_A_232_82#_c_226_n N_A_343_80#_c_433_n 0.0186865f $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_239 N_A_232_82#_c_228_n N_A_343_80#_c_433_n 0.00556466f $X=3.265 $Y=1.185
+ $X2=0 $Y2=0
cc_240 N_A_232_82#_c_236_n N_A_343_80#_c_433_n 0.001094f $X=3.912 $Y=1.47 $X2=0
+ $Y2=0
cc_241 N_A_232_82#_c_226_n N_A_343_80#_c_434_n 0.00438387f $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_242 N_A_232_82#_c_226_n N_A_343_80#_c_435_n 0.00971484f $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_243 N_A_232_82#_c_227_n N_A_343_80#_c_435_n 0.00318759f $X=3.72 $Y=1.185
+ $X2=0 $Y2=0
cc_244 N_A_232_82#_c_226_n N_A_343_80#_c_436_n 0.0026279f $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_245 N_A_232_82#_c_228_n N_A_343_80#_c_437_n 9.58254e-19 $X=3.265 $Y=1.185
+ $X2=0 $Y2=0
cc_246 N_A_232_82#_c_239_n N_A_343_80#_c_437_n 0.023831f $X=3.975 $Y=2.475 $X2=0
+ $Y2=0
cc_247 N_A_232_82#_c_228_n N_A_343_80#_c_438_n 0.0194401f $X=3.265 $Y=1.185
+ $X2=0 $Y2=0
cc_248 N_A_232_82#_c_233_n N_A_343_80#_c_438_n 0.0116557f $X=3.94 $Y=1.635 $X2=0
+ $Y2=0
cc_249 N_A_232_82#_c_227_n N_A_343_80#_c_439_n 0.00302518f $X=3.72 $Y=1.185
+ $X2=0 $Y2=0
cc_250 N_A_232_82#_c_234_n N_A_343_80#_c_439_n 2.0142e-19 $X=4.06 $Y=1.635 $X2=0
+ $Y2=0
cc_251 N_A_232_82#_M1006_g N_A_863_294#_M1011_g 0.0264604f $X=3.95 $Y=2.17 $X2=0
+ $Y2=0
cc_252 N_A_232_82#_c_239_n N_A_863_294#_M1011_g 0.00106319f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_253 N_A_232_82#_c_240_n N_A_863_294#_M1011_g 0.00614948f $X=4.06 $Y=2.39
+ $X2=0 $Y2=0
cc_254 N_A_232_82#_c_227_n N_A_863_294#_M1004_g 0.00572479f $X=3.72 $Y=1.185
+ $X2=0 $Y2=0
cc_255 N_A_232_82#_M1006_g N_A_863_294#_c_541_n 2.51205e-19 $X=3.95 $Y=2.17
+ $X2=0 $Y2=0
cc_256 N_A_232_82#_c_240_n N_A_863_294#_c_541_n 0.00713378f $X=4.06 $Y=2.39
+ $X2=0 $Y2=0
cc_257 N_A_232_82#_c_233_n N_A_863_294#_c_541_n 3.76643e-19 $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_258 N_A_232_82#_c_234_n N_A_863_294#_c_541_n 0.0258564f $X=4.06 $Y=1.635
+ $X2=0 $Y2=0
cc_259 N_A_232_82#_c_233_n N_A_863_294#_c_542_n 0.0206865f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_260 N_A_232_82#_c_234_n N_A_863_294#_c_542_n 0.00183089f $X=4.06 $Y=1.635
+ $X2=0 $Y2=0
cc_261 N_A_232_82#_c_239_n N_A_653_79#_M1014_d 0.0062843f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_262 N_A_232_82#_M1006_g N_A_653_79#_c_650_n 0.00195167f $X=3.95 $Y=2.17 $X2=0
+ $Y2=0
cc_263 N_A_232_82#_c_240_n N_A_653_79#_c_650_n 0.00941211f $X=4.06 $Y=2.39 $X2=0
+ $Y2=0
cc_264 N_A_232_82#_c_234_n N_A_653_79#_c_650_n 0.02456f $X=4.06 $Y=1.635 $X2=0
+ $Y2=0
cc_265 N_A_232_82#_c_236_n N_A_653_79#_c_650_n 0.00758336f $X=3.912 $Y=1.47
+ $X2=0 $Y2=0
cc_266 N_A_232_82#_c_234_n N_A_653_79#_c_651_n 7.55144e-19 $X=4.06 $Y=1.635
+ $X2=0 $Y2=0
cc_267 N_A_232_82#_c_226_n N_A_653_79#_c_652_n 0.00817513f $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_268 N_A_232_82#_c_227_n N_A_653_79#_c_652_n 0.028451f $X=3.72 $Y=1.185 $X2=0
+ $Y2=0
cc_269 N_A_232_82#_c_233_n N_A_653_79#_c_652_n 0.00610918f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_270 N_A_232_82#_c_234_n N_A_653_79#_c_652_n 0.0237395f $X=4.06 $Y=1.635 $X2=0
+ $Y2=0
cc_271 N_A_232_82#_c_236_n N_A_653_79#_c_652_n 0.00856005f $X=3.912 $Y=1.47
+ $X2=0 $Y2=0
cc_272 N_A_232_82#_c_239_n N_A_653_79#_c_669_n 0.0371845f $X=3.975 $Y=2.475
+ $X2=0 $Y2=0
cc_273 N_A_232_82#_c_233_n N_A_653_79#_c_669_n 0.00319471f $X=3.94 $Y=1.635
+ $X2=0 $Y2=0
cc_274 N_A_232_82#_c_239_n N_VPWR_M1021_d 0.00533673f $X=3.975 $Y=2.475 $X2=0
+ $Y2=0
cc_275 N_A_232_82#_c_241_n N_VPWR_c_771_n 0.0259229f $X=1.4 $Y=2.405 $X2=0 $Y2=0
cc_276 N_A_232_82#_M1021_g N_VPWR_c_772_n 0.00405737f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_277 N_A_232_82#_c_239_n N_VPWR_c_772_n 0.021216f $X=3.975 $Y=2.475 $X2=0
+ $Y2=0
cc_278 N_A_232_82#_M1006_g N_VPWR_c_774_n 4.15871e-19 $X=3.95 $Y=2.17 $X2=0
+ $Y2=0
cc_279 N_A_232_82#_c_239_n N_VPWR_c_774_n 0.00917364f $X=3.975 $Y=2.475 $X2=0
+ $Y2=0
cc_280 N_A_232_82#_c_240_n N_VPWR_c_774_n 0.0150194f $X=4.06 $Y=2.39 $X2=0 $Y2=0
cc_281 N_A_232_82#_M1021_g N_VPWR_c_783_n 0.00562877f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_282 N_A_232_82#_c_243_n N_VPWR_c_783_n 0.0145232f $X=1.455 $Y=2.475 $X2=0
+ $Y2=0
cc_283 N_A_232_82#_M1021_g N_VPWR_c_770_n 0.00595788f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_284 N_A_232_82#_c_239_n N_VPWR_c_770_n 0.0776779f $X=3.975 $Y=2.475 $X2=0
+ $Y2=0
cc_285 N_A_232_82#_c_241_n N_VPWR_c_770_n 0.00457292f $X=1.4 $Y=2.405 $X2=0
+ $Y2=0
cc_286 N_A_232_82#_c_243_n N_VPWR_c_770_n 0.0119642f $X=1.455 $Y=2.475 $X2=0
+ $Y2=0
cc_287 N_A_232_82#_c_239_n A_574_392# 0.00467744f $X=3.975 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_232_82#_c_240_n A_808_392# 0.00476342f $X=4.06 $Y=2.39 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_232_82#_c_226_n N_VGND_c_911_n 9.62964e-19 $X=3.19 $Y=1.11 $X2=0
+ $Y2=0
cc_290 N_A_232_82#_c_224_n N_VGND_c_916_n 0.00806779f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_291 N_A_232_82#_c_224_n N_VGND_c_919_n 0.00536257f $X=2.22 $Y=1.25 $X2=0
+ $Y2=0
cc_292 N_A_27_120#_c_358_n N_A_343_80#_M1008_s 0.0119208f $X=2.535 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_293 N_A_27_120#_M1002_g N_A_343_80#_M1014_g 0.0711814f $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_294 N_A_27_120#_c_358_n N_A_343_80#_c_431_n 0.0362929f $X=2.535 $Y=0.665
+ $X2=0 $Y2=0
cc_295 N_A_27_120#_c_359_n N_A_343_80#_c_431_n 0.00913096f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_296 N_A_27_120#_M1002_g N_A_343_80#_c_432_n 6.74446e-19 $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_297 N_A_27_120#_c_359_n N_A_343_80#_c_432_n 0.0200982f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_298 N_A_27_120#_c_360_n N_A_343_80#_c_432_n 0.0012296f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_299 N_A_27_120#_c_359_n N_A_343_80#_c_442_n 0.00909208f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_300 N_A_27_120#_c_360_n N_A_343_80#_c_442_n 0.00297528f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_301 N_A_27_120#_M1013_g N_A_343_80#_c_433_n 0.00984909f $X=2.8 $Y=0.715 $X2=0
+ $Y2=0
cc_302 N_A_27_120#_c_358_n N_A_343_80#_c_433_n 0.0133618f $X=2.535 $Y=0.665
+ $X2=0 $Y2=0
cc_303 N_A_27_120#_c_359_n N_A_343_80#_c_433_n 0.0536237f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_304 N_A_27_120#_M1013_g N_A_343_80#_c_434_n 0.00392088f $X=2.8 $Y=0.715 $X2=0
+ $Y2=0
cc_305 N_A_27_120#_M1002_g N_A_343_80#_c_437_n 0.0272844f $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_306 N_A_27_120#_c_359_n N_A_343_80#_c_437_n 0.0184951f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_307 N_A_27_120#_c_360_n N_A_343_80#_c_437_n 0.00296483f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_308 N_A_27_120#_M1002_g N_A_343_80#_c_438_n 0.0131756f $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_309 N_A_27_120#_c_360_n N_A_343_80#_c_438_n 0.00688029f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_310 N_A_27_120#_c_364_n N_VPWR_c_771_n 0.0234195f $X=0.38 $Y=2.265 $X2=0
+ $Y2=0
cc_311 N_A_27_120#_M1002_g N_VPWR_c_772_n 0.00973899f $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_312 N_A_27_120#_M1002_g N_VPWR_c_773_n 0.00490827f $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_313 N_A_27_120#_c_364_n N_VPWR_c_777_n 0.0199902f $X=0.38 $Y=2.265 $X2=0
+ $Y2=0
cc_314 N_A_27_120#_M1002_g N_VPWR_c_770_n 0.00472461f $X=2.78 $Y=2.46 $X2=0
+ $Y2=0
cc_315 N_A_27_120#_c_364_n N_VPWR_c_770_n 0.0165461f $X=0.38 $Y=2.265 $X2=0
+ $Y2=0
cc_316 N_A_27_120#_c_358_n N_VGND_M1020_d 0.0117644f $X=2.535 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_317 N_A_27_120#_c_358_n N_VGND_M1008_d 0.0108232f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_318 N_A_27_120#_c_359_n N_VGND_M1008_d 0.00479298f $X=2.7 $Y=1.415 $X2=0
+ $Y2=0
cc_319 N_A_27_120#_M1013_g N_VGND_c_911_n 0.00432157f $X=2.8 $Y=0.715 $X2=0
+ $Y2=0
cc_320 N_A_27_120#_c_358_n N_VGND_c_911_n 0.00342596f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_321 N_A_27_120#_c_358_n N_VGND_c_915_n 0.00346124f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_322 N_A_27_120#_c_361_n N_VGND_c_915_n 0.00779317f $X=0.27 $Y=0.665 $X2=0
+ $Y2=0
cc_323 N_A_27_120#_M1013_g N_VGND_c_916_n 0.00177422f $X=2.8 $Y=0.715 $X2=0
+ $Y2=0
cc_324 N_A_27_120#_c_358_n N_VGND_c_916_n 0.0501284f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_325 N_A_27_120#_M1013_g N_VGND_c_919_n 0.00537853f $X=2.8 $Y=0.715 $X2=0
+ $Y2=0
cc_326 N_A_27_120#_c_358_n N_VGND_c_919_n 0.055622f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_327 N_A_27_120#_c_361_n N_VGND_c_919_n 0.0108955f $X=0.27 $Y=0.665 $X2=0
+ $Y2=0
cc_328 N_A_27_120#_c_358_n N_VGND_c_920_n 0.0245693f $X=2.535 $Y=0.665 $X2=0
+ $Y2=0
cc_329 N_A_343_80#_c_436_n N_A_863_294#_M1004_g 0.0354855f $X=4.095 $Y=0.34
+ $X2=0 $Y2=0
cc_330 N_A_343_80#_c_435_n N_A_653_79#_M1012_d 0.00289102f $X=4.095 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_331 N_A_343_80#_M1014_g N_A_653_79#_c_650_n 0.00238377f $X=3.2 $Y=2.46 $X2=0
+ $Y2=0
cc_332 N_A_343_80#_c_433_n N_A_653_79#_c_650_n 0.00877411f $X=3.12 $Y=1.47 $X2=0
+ $Y2=0
cc_333 N_A_343_80#_c_437_n N_A_653_79#_c_650_n 0.0361324f $X=3.12 $Y=1.845 $X2=0
+ $Y2=0
cc_334 N_A_343_80#_c_438_n N_A_653_79#_c_650_n 0.00249021f $X=3.25 $Y=1.635
+ $X2=0 $Y2=0
cc_335 N_A_343_80#_c_435_n N_A_653_79#_c_651_n 0.00295108f $X=4.095 $Y=0.34
+ $X2=0 $Y2=0
cc_336 N_A_343_80#_c_439_n N_A_653_79#_c_651_n 0.00629255f $X=4.095 $Y=0.505
+ $X2=0 $Y2=0
cc_337 N_A_343_80#_c_433_n N_A_653_79#_c_652_n 0.0383019f $X=3.12 $Y=1.47 $X2=0
+ $Y2=0
cc_338 N_A_343_80#_c_435_n N_A_653_79#_c_652_n 0.0460543f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_339 N_A_343_80#_c_436_n N_A_653_79#_c_652_n 0.00386325f $X=4.095 $Y=0.34
+ $X2=0 $Y2=0
cc_340 N_A_343_80#_c_439_n N_A_653_79#_c_652_n 0.0106624f $X=4.095 $Y=0.505
+ $X2=0 $Y2=0
cc_341 N_A_343_80#_M1014_g N_A_653_79#_c_669_n 0.00646944f $X=3.2 $Y=2.46 $X2=0
+ $Y2=0
cc_342 N_A_343_80#_c_437_n N_A_653_79#_c_669_n 0.0043748f $X=3.12 $Y=1.845 $X2=0
+ $Y2=0
cc_343 N_A_343_80#_c_438_n N_A_653_79#_c_669_n 0.00247985f $X=3.25 $Y=1.635
+ $X2=0 $Y2=0
cc_344 N_A_343_80#_c_442_n N_VPWR_M1021_d 0.00283824f $X=2.655 $Y=1.965 $X2=0
+ $Y2=0
cc_345 N_A_343_80#_M1014_g N_VPWR_c_772_n 0.00171177f $X=3.2 $Y=2.46 $X2=0 $Y2=0
cc_346 N_A_343_80#_M1014_g N_VPWR_c_773_n 0.00553757f $X=3.2 $Y=2.46 $X2=0 $Y2=0
cc_347 N_A_343_80#_M1014_g N_VPWR_c_770_n 0.00540034f $X=3.2 $Y=2.46 $X2=0 $Y2=0
cc_348 N_A_343_80#_c_435_n N_VGND_c_908_n 0.0100907f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_349 N_A_343_80#_c_436_n N_VGND_c_908_n 0.00302969f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_350 N_A_343_80#_c_434_n N_VGND_c_911_n 0.0121867f $X=3.205 $Y=0.38 $X2=0
+ $Y2=0
cc_351 N_A_343_80#_c_435_n N_VGND_c_911_n 0.0687728f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_352 N_A_343_80#_c_436_n N_VGND_c_911_n 0.00659816f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_353 N_A_343_80#_c_434_n N_VGND_c_916_n 0.00770007f $X=3.205 $Y=0.38 $X2=0
+ $Y2=0
cc_354 N_A_343_80#_c_434_n N_VGND_c_919_n 0.00660921f $X=3.205 $Y=0.38 $X2=0
+ $Y2=0
cc_355 N_A_343_80#_c_435_n N_VGND_c_919_n 0.0384913f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_356 N_A_343_80#_c_436_n N_VGND_c_919_n 0.0104196f $X=4.095 $Y=0.34 $X2=0
+ $Y2=0
cc_357 N_A_343_80#_c_433_n A_575_79# 0.00464502f $X=3.12 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_358 N_A_343_80#_c_434_n A_575_79# 0.00147159f $X=3.205 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_359 N_A_863_294#_M1011_g N_A_653_79#_M1015_g 0.0120958f $X=4.435 $Y=2.17
+ $X2=0 $Y2=0
cc_360 N_A_863_294#_c_548_n N_A_653_79#_M1015_g 0.0137308f $X=5.22 $Y=1.805
+ $X2=0 $Y2=0
cc_361 N_A_863_294#_c_539_n N_A_653_79#_M1015_g 0.00272319f $X=5.39 $Y=1.89
+ $X2=0 $Y2=0
cc_362 N_A_863_294#_c_550_n N_A_653_79#_M1015_g 0.0160961f $X=5.385 $Y=1.905
+ $X2=0 $Y2=0
cc_363 N_A_863_294#_c_541_n N_A_653_79#_M1015_g 0.00109658f $X=4.48 $Y=1.635
+ $X2=0 $Y2=0
cc_364 N_A_863_294#_c_542_n N_A_653_79#_M1015_g 0.00746849f $X=4.48 $Y=1.635
+ $X2=0 $Y2=0
cc_365 N_A_863_294#_M1004_g N_A_653_79#_c_651_n 0.0157461f $X=4.575 $Y=0.825
+ $X2=0 $Y2=0
cc_366 N_A_863_294#_c_548_n N_A_653_79#_c_651_n 0.00983898f $X=5.22 $Y=1.805
+ $X2=0 $Y2=0
cc_367 N_A_863_294#_c_541_n N_A_653_79#_c_651_n 0.0246969f $X=4.48 $Y=1.635
+ $X2=0 $Y2=0
cc_368 N_A_863_294#_c_542_n N_A_653_79#_c_651_n 0.00128251f $X=4.48 $Y=1.635
+ $X2=0 $Y2=0
cc_369 N_A_863_294#_M1004_g N_A_653_79#_c_652_n 0.00152312f $X=4.575 $Y=0.825
+ $X2=0 $Y2=0
cc_370 N_A_863_294#_M1004_g N_A_653_79#_c_653_n 0.00154982f $X=4.575 $Y=0.825
+ $X2=0 $Y2=0
cc_371 N_A_863_294#_c_536_n N_A_653_79#_c_653_n 2.85519e-19 $X=6.065 $Y=1.435
+ $X2=0 $Y2=0
cc_372 N_A_863_294#_c_548_n N_A_653_79#_c_653_n 0.0246782f $X=5.22 $Y=1.805
+ $X2=0 $Y2=0
cc_373 N_A_863_294#_c_539_n N_A_653_79#_c_653_n 0.0226111f $X=5.39 $Y=1.89 $X2=0
+ $Y2=0
cc_374 N_A_863_294#_c_540_n N_A_653_79#_c_653_n 0.0104466f $X=5.475 $Y=1.27
+ $X2=0 $Y2=0
cc_375 N_A_863_294#_c_541_n N_A_653_79#_c_653_n 0.00448327f $X=4.48 $Y=1.635
+ $X2=0 $Y2=0
cc_376 N_A_863_294#_c_543_n N_A_653_79#_c_653_n 0.00105254f $X=5.382 $Y=0.96
+ $X2=0 $Y2=0
cc_377 N_A_863_294#_M1004_g N_A_653_79#_c_654_n 0.0181141f $X=4.575 $Y=0.825
+ $X2=0 $Y2=0
cc_378 N_A_863_294#_c_536_n N_A_653_79#_c_654_n 0.0205786f $X=6.065 $Y=1.435
+ $X2=0 $Y2=0
cc_379 N_A_863_294#_c_548_n N_A_653_79#_c_654_n 0.00126186f $X=5.22 $Y=1.805
+ $X2=0 $Y2=0
cc_380 N_A_863_294#_c_539_n N_A_653_79#_c_654_n 0.00730427f $X=5.39 $Y=1.89
+ $X2=0 $Y2=0
cc_381 N_A_863_294#_c_540_n N_A_653_79#_c_654_n 0.00117986f $X=5.475 $Y=1.27
+ $X2=0 $Y2=0
cc_382 N_A_863_294#_c_541_n N_A_653_79#_c_654_n 2.97104e-19 $X=4.48 $Y=1.635
+ $X2=0 $Y2=0
cc_383 N_A_863_294#_M1004_g N_A_653_79#_c_655_n 0.0172907f $X=4.575 $Y=0.825
+ $X2=0 $Y2=0
cc_384 N_A_863_294#_c_538_n N_A_653_79#_c_655_n 0.00473741f $X=5.37 $Y=0.535
+ $X2=0 $Y2=0
cc_385 N_A_863_294#_c_540_n N_A_653_79#_c_655_n 0.0056455f $X=5.475 $Y=1.27
+ $X2=0 $Y2=0
cc_386 N_A_863_294#_c_543_n N_A_653_79#_c_655_n 0.00189095f $X=5.382 $Y=0.96
+ $X2=0 $Y2=0
cc_387 N_A_863_294#_c_537_n N_A_1350_424#_c_727_n 0.00861428f $X=6.66 $Y=1.392
+ $X2=0 $Y2=0
cc_388 N_A_863_294#_c_533_n N_A_1350_424#_c_729_n 3.07525e-19 $X=6.17 $Y=1.185
+ $X2=0 $Y2=0
cc_389 N_A_863_294#_c_535_n N_A_1350_424#_c_729_n 0.013134f $X=6.68 $Y=1.185
+ $X2=0 $Y2=0
cc_390 N_A_863_294#_c_537_n N_A_1350_424#_c_729_n 0.00585128f $X=6.66 $Y=1.392
+ $X2=0 $Y2=0
cc_391 N_A_863_294#_M1019_g N_A_1350_424#_c_730_n 0.00154902f $X=6.155 $Y=2.4
+ $X2=0 $Y2=0
cc_392 N_A_863_294#_M1016_g N_A_1350_424#_c_730_n 0.0331085f $X=6.66 $Y=2.54
+ $X2=0 $Y2=0
cc_393 N_A_863_294#_M1016_g N_A_1350_424#_c_732_n 0.00103708f $X=6.66 $Y=2.54
+ $X2=0 $Y2=0
cc_394 N_A_863_294#_c_537_n N_A_1350_424#_c_732_n 0.0144941f $X=6.66 $Y=1.392
+ $X2=0 $Y2=0
cc_395 N_A_863_294#_c_548_n N_VPWR_M1011_d 0.00263949f $X=5.22 $Y=1.805 $X2=0
+ $Y2=0
cc_396 N_A_863_294#_M1011_g N_VPWR_c_774_n 0.0168802f $X=4.435 $Y=2.17 $X2=0
+ $Y2=0
cc_397 N_A_863_294#_c_548_n N_VPWR_c_774_n 0.0301529f $X=5.22 $Y=1.805 $X2=0
+ $Y2=0
cc_398 N_A_863_294#_c_550_n N_VPWR_c_774_n 0.0285604f $X=5.385 $Y=1.905 $X2=0
+ $Y2=0
cc_399 N_A_863_294#_c_541_n N_VPWR_c_774_n 0.0115733f $X=4.48 $Y=1.635 $X2=0
+ $Y2=0
cc_400 N_A_863_294#_c_542_n N_VPWR_c_774_n 6.26347e-19 $X=4.48 $Y=1.635 $X2=0
+ $Y2=0
cc_401 N_A_863_294#_M1019_g N_VPWR_c_775_n 0.00384612f $X=6.155 $Y=2.4 $X2=0
+ $Y2=0
cc_402 N_A_863_294#_M1016_g N_VPWR_c_775_n 0.0042237f $X=6.66 $Y=2.54 $X2=0
+ $Y2=0
cc_403 N_A_863_294#_c_537_n N_VPWR_c_775_n 0.00467029f $X=6.66 $Y=1.392 $X2=0
+ $Y2=0
cc_404 N_A_863_294#_M1016_g N_VPWR_c_776_n 0.00554988f $X=6.66 $Y=2.54 $X2=0
+ $Y2=0
cc_405 N_A_863_294#_M1019_g N_VPWR_c_779_n 0.00481245f $X=6.155 $Y=2.4 $X2=0
+ $Y2=0
cc_406 N_A_863_294#_c_550_n N_VPWR_c_779_n 0.0113165f $X=5.385 $Y=1.905 $X2=0
+ $Y2=0
cc_407 N_A_863_294#_M1016_g N_VPWR_c_781_n 0.005209f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_408 N_A_863_294#_M1011_g N_VPWR_c_770_n 0.00352022f $X=4.435 $Y=2.17 $X2=0
+ $Y2=0
cc_409 N_A_863_294#_M1019_g N_VPWR_c_770_n 0.00859641f $X=6.155 $Y=2.4 $X2=0
+ $Y2=0
cc_410 N_A_863_294#_M1016_g N_VPWR_c_770_n 0.00987261f $X=6.66 $Y=2.54 $X2=0
+ $Y2=0
cc_411 N_A_863_294#_c_550_n N_VPWR_c_770_n 0.0118362f $X=5.385 $Y=1.905 $X2=0
+ $Y2=0
cc_412 N_A_863_294#_M1019_g N_Q_c_861_n 0.0162171f $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_413 N_A_863_294#_M1019_g N_Q_c_862_n 0.00441429f $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A_863_294#_c_536_n N_Q_c_862_n 0.00734325f $X=6.065 $Y=1.435 $X2=0
+ $Y2=0
cc_415 N_A_863_294#_c_539_n N_Q_c_862_n 0.00714072f $X=5.39 $Y=1.89 $X2=0 $Y2=0
cc_416 N_A_863_294#_c_550_n N_Q_c_862_n 0.0744123f $X=5.385 $Y=1.905 $X2=0 $Y2=0
cc_417 N_A_863_294#_M1019_g N_Q_c_858_n 0.00879467f $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A_863_294#_c_533_n N_Q_c_858_n 0.0028946f $X=6.17 $Y=1.185 $X2=0 $Y2=0
cc_419 N_A_863_294#_M1016_g N_Q_c_858_n 0.00182685f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_420 N_A_863_294#_c_536_n N_Q_c_858_n 0.012774f $X=6.065 $Y=1.435 $X2=0 $Y2=0
cc_421 N_A_863_294#_c_537_n N_Q_c_858_n 0.0156816f $X=6.66 $Y=1.392 $X2=0 $Y2=0
cc_422 N_A_863_294#_c_539_n N_Q_c_858_n 0.0314075f $X=5.39 $Y=1.89 $X2=0 $Y2=0
cc_423 N_A_863_294#_c_540_n N_Q_c_858_n 0.00498203f $X=5.475 $Y=1.27 $X2=0 $Y2=0
cc_424 N_A_863_294#_c_533_n Q 0.00768219f $X=6.17 $Y=1.185 $X2=0 $Y2=0
cc_425 N_A_863_294#_c_535_n Q 3.33005e-19 $X=6.68 $Y=1.185 $X2=0 $Y2=0
cc_426 N_A_863_294#_c_538_n Q 0.0251784f $X=5.37 $Y=0.535 $X2=0 $Y2=0
cc_427 N_A_863_294#_c_533_n Q 0.00185548f $X=6.17 $Y=1.185 $X2=0 $Y2=0
cc_428 N_A_863_294#_c_536_n Q 0.00751058f $X=6.065 $Y=1.435 $X2=0 $Y2=0
cc_429 N_A_863_294#_c_543_n Q 0.0251784f $X=5.382 $Y=0.96 $X2=0 $Y2=0
cc_430 N_A_863_294#_M1004_g N_VGND_c_908_n 0.00548813f $X=4.575 $Y=0.825 $X2=0
+ $Y2=0
cc_431 N_A_863_294#_c_538_n N_VGND_c_908_n 0.0238985f $X=5.37 $Y=0.535 $X2=0
+ $Y2=0
cc_432 N_A_863_294#_c_533_n N_VGND_c_909_n 0.00770657f $X=6.17 $Y=1.185 $X2=0
+ $Y2=0
cc_433 N_A_863_294#_c_535_n N_VGND_c_909_n 0.00410027f $X=6.68 $Y=1.185 $X2=0
+ $Y2=0
cc_434 N_A_863_294#_c_537_n N_VGND_c_909_n 0.00940372f $X=6.66 $Y=1.392 $X2=0
+ $Y2=0
cc_435 N_A_863_294#_c_535_n N_VGND_c_910_n 0.00409144f $X=6.68 $Y=1.185 $X2=0
+ $Y2=0
cc_436 N_A_863_294#_M1004_g N_VGND_c_911_n 0.00420632f $X=4.575 $Y=0.825 $X2=0
+ $Y2=0
cc_437 N_A_863_294#_c_533_n N_VGND_c_913_n 0.00422942f $X=6.17 $Y=1.185 $X2=0
+ $Y2=0
cc_438 N_A_863_294#_c_538_n N_VGND_c_913_n 0.0156453f $X=5.37 $Y=0.535 $X2=0
+ $Y2=0
cc_439 N_A_863_294#_c_535_n N_VGND_c_917_n 0.00426181f $X=6.68 $Y=1.185 $X2=0
+ $Y2=0
cc_440 N_A_863_294#_M1004_g N_VGND_c_919_n 0.00472204f $X=4.575 $Y=0.825 $X2=0
+ $Y2=0
cc_441 N_A_863_294#_c_533_n N_VGND_c_919_n 0.00793595f $X=6.17 $Y=1.185 $X2=0
+ $Y2=0
cc_442 N_A_863_294#_c_535_n N_VGND_c_919_n 0.00487769f $X=6.68 $Y=1.185 $X2=0
+ $Y2=0
cc_443 N_A_863_294#_c_538_n N_VGND_c_919_n 0.012945f $X=5.37 $Y=0.535 $X2=0
+ $Y2=0
cc_444 N_A_653_79#_M1015_g N_VPWR_c_774_n 0.00960411f $X=5.16 $Y=2.32 $X2=0
+ $Y2=0
cc_445 N_A_653_79#_M1015_g N_VPWR_c_779_n 0.00597358f $X=5.16 $Y=2.32 $X2=0
+ $Y2=0
cc_446 N_A_653_79#_M1015_g N_VPWR_c_770_n 0.00624688f $X=5.16 $Y=2.32 $X2=0
+ $Y2=0
cc_447 N_A_653_79#_M1015_g N_Q_c_861_n 0.00213431f $X=5.16 $Y=2.32 $X2=0 $Y2=0
cc_448 N_A_653_79#_M1015_g N_Q_c_862_n 0.00193893f $X=5.16 $Y=2.32 $X2=0 $Y2=0
cc_449 N_A_653_79#_c_655_n Q 0.00104531f $X=5.07 $Y=1.22 $X2=0 $Y2=0
cc_450 N_A_653_79#_c_651_n N_VGND_c_908_n 0.01517f $X=4.89 $Y=1.215 $X2=0 $Y2=0
cc_451 N_A_653_79#_c_653_n N_VGND_c_908_n 0.011731f $X=5.055 $Y=1.215 $X2=0
+ $Y2=0
cc_452 N_A_653_79#_c_654_n N_VGND_c_908_n 8.46342e-19 $X=5.055 $Y=1.385 $X2=0
+ $Y2=0
cc_453 N_A_653_79#_c_655_n N_VGND_c_908_n 0.0103449f $X=5.07 $Y=1.22 $X2=0 $Y2=0
cc_454 N_A_653_79#_c_655_n N_VGND_c_913_n 0.00445602f $X=5.07 $Y=1.22 $X2=0
+ $Y2=0
cc_455 N_A_653_79#_c_655_n N_VGND_c_919_n 0.00866521f $X=5.07 $Y=1.22 $X2=0
+ $Y2=0
cc_456 N_A_1350_424#_c_730_n N_VPWR_c_775_n 0.034761f $X=6.89 $Y=2.265 $X2=0
+ $Y2=0
cc_457 N_A_1350_424#_M1018_g N_VPWR_c_776_n 0.00649215f $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_458 N_A_1350_424#_c_727_n N_VPWR_c_776_n 0.00600559f $X=7.565 $Y=1.465 $X2=0
+ $Y2=0
cc_459 N_A_1350_424#_c_730_n N_VPWR_c_776_n 0.0846938f $X=6.89 $Y=2.265 $X2=0
+ $Y2=0
cc_460 N_A_1350_424#_c_731_n N_VPWR_c_776_n 0.0181512f $X=7.335 $Y=1.465 $X2=0
+ $Y2=0
cc_461 N_A_1350_424#_c_730_n N_VPWR_c_781_n 0.0152183f $X=6.89 $Y=2.265 $X2=0
+ $Y2=0
cc_462 N_A_1350_424#_M1018_g N_VPWR_c_784_n 0.005209f $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_463 N_A_1350_424#_M1018_g N_VPWR_c_770_n 0.00991141f $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_464 N_A_1350_424#_c_730_n N_VPWR_c_770_n 0.0125283f $X=6.89 $Y=2.265 $X2=0
+ $Y2=0
cc_465 N_A_1350_424#_c_729_n N_Q_c_858_n 0.00437285f $X=6.895 $Y=0.835 $X2=0
+ $Y2=0
cc_466 N_A_1350_424#_c_730_n N_Q_c_858_n 0.0125726f $X=6.89 $Y=2.265 $X2=0 $Y2=0
cc_467 N_A_1350_424#_c_732_n N_Q_c_858_n 0.0089399f $X=6.892 $Y=1.465 $X2=0
+ $Y2=0
cc_468 N_A_1350_424#_M1018_g Q_N 0.0247772f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_469 N_A_1350_424#_M1007_g Q_N 0.018165f $X=7.67 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A_1350_424#_c_728_n Q_N 0.0127834f $X=7.655 $Y=1.465 $X2=0 $Y2=0
cc_471 N_A_1350_424#_c_729_n Q_N 0.00481564f $X=6.895 $Y=0.835 $X2=0 $Y2=0
cc_472 N_A_1350_424#_c_730_n Q_N 0.00542516f $X=6.89 $Y=2.265 $X2=0 $Y2=0
cc_473 N_A_1350_424#_c_731_n Q_N 0.0217011f $X=7.335 $Y=1.465 $X2=0 $Y2=0
cc_474 N_A_1350_424#_c_729_n N_VGND_c_909_n 0.0237555f $X=6.895 $Y=0.835 $X2=0
+ $Y2=0
cc_475 N_A_1350_424#_M1007_g N_VGND_c_910_n 0.00647103f $X=7.67 $Y=0.74 $X2=0
+ $Y2=0
cc_476 N_A_1350_424#_c_727_n N_VGND_c_910_n 0.006602f $X=7.565 $Y=1.465 $X2=0
+ $Y2=0
cc_477 N_A_1350_424#_c_729_n N_VGND_c_910_n 0.0390482f $X=6.895 $Y=0.835 $X2=0
+ $Y2=0
cc_478 N_A_1350_424#_c_731_n N_VGND_c_910_n 0.0176257f $X=7.335 $Y=1.465 $X2=0
+ $Y2=0
cc_479 N_A_1350_424#_c_729_n N_VGND_c_917_n 0.00837462f $X=6.895 $Y=0.835 $X2=0
+ $Y2=0
cc_480 N_A_1350_424#_M1007_g N_VGND_c_918_n 0.00428607f $X=7.67 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A_1350_424#_M1007_g N_VGND_c_919_n 0.0081058f $X=7.67 $Y=0.74 $X2=0
+ $Y2=0
cc_482 N_A_1350_424#_c_729_n N_VGND_c_919_n 0.0109536f $X=6.895 $Y=0.835 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_775_n N_Q_c_861_n 0.0342911f $X=6.385 $Y=2.265 $X2=0 $Y2=0
cc_484 N_VPWR_c_779_n N_Q_c_861_n 0.0160061f $X=6.3 $Y=3.33 $X2=0 $Y2=0
cc_485 N_VPWR_c_770_n N_Q_c_861_n 0.0130981f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_486 N_VPWR_c_776_n Q_N 0.0396567f $X=7.43 $Y=1.985 $X2=0 $Y2=0
cc_487 N_VPWR_c_784_n Q_N 0.0147721f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_488 N_VPWR_c_770_n Q_N 0.0121589f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_489 Q N_VGND_c_909_n 0.0309648f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_490 Q N_VGND_c_913_n 0.0149802f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_491 Q N_VGND_c_919_n 0.0123195f $X=5.915 $Y=0.47 $X2=0 $Y2=0
cc_492 Q_N N_VGND_c_910_n 0.0301457f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_493 Q_N N_VGND_c_918_n 0.0147721f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_494 Q_N N_VGND_c_919_n 0.0121589f $X=7.835 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__bufbuf_8.pex.spice
* Created: Wed Sep  2 11:59:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%A 1 3 6 8 12
c34 6 0 8.22433e-20 $X=0.495 $Y=0.835
c35 1 0 1.94207e-19 $X=0.505 $Y=1.77
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.515 $X2=0.405 $Y2=1.515
r37 8 12 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.405 $Y2=1.565
r38 4 11 38.5662 $w=2.97e-07 $l=2.00237e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.417 $Y2=1.515
r39 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.835
r40 1 11 48.8089 $w=2.97e-07 $l=2.95745e-07 $layer=POLY_cond $X=0.505 $Y=1.77
+ $X2=0.417 $Y2=1.515
r41 1 3 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=0.505 $Y=1.77
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%A_27_112# 1 2 9 13 17 19 21 23 25 26 27 28
+ 34
r73 34 37 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.465
+ $X2=0.98 $Y2=1.63
r74 34 36 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.465
+ $X2=0.98 $Y2=1.3
r75 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.465 $X2=0.975 $Y2=1.465
r76 27 33 9.02499 $w=2.87e-07 $l=2.13014e-07 $layer=LI1_cond $X=0.835 $Y=1.63
+ $X2=0.945 $Y2=1.465
r77 27 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.835 $Y=1.63
+ $X2=0.835 $Y2=1.95
r78 25 33 15.7282 $w=2.87e-07 $l=4.5722e-07 $layer=LI1_cond $X=0.75 $Y=1.095
+ $X2=0.945 $Y2=1.465
r79 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.75 $Y=1.095
+ $X2=0.445 $Y2=1.095
r80 24 30 3.51781 $w=2.5e-07 $l=1.33e-07 $layer=LI1_cond $X=0.38 $Y=2.075
+ $X2=0.247 $Y2=2.075
r81 23 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.75 $Y=2.075
+ $X2=0.835 $Y2=1.95
r82 23 24 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=2.075
+ $X2=0.38 $Y2=2.075
r83 19 30 3.30621 $w=2.65e-07 $l=1.25e-07 $layer=LI1_cond $X=0.247 $Y=2.2
+ $X2=0.247 $Y2=2.075
r84 19 21 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=0.247 $Y=2.2
+ $X2=0.247 $Y2=2.535
r85 15 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r86 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.835
r87 13 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.075 $Y=0.74
+ $X2=1.075 $Y2=1.3
r88 9 37 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.03 $Y=2.4 $X2=1.03
+ $Y2=1.63
r89 2 30 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.06
r90 2 21 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.535
r91 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%A_224_368# 1 2 9 13 17 21 25 29 33 37 40 48
+ 52 53 54 55 56 65
c99 54 0 8.22433e-20 $X=1.302 $Y=1.13
c100 52 0 1.94207e-19 $X=1.255 $Y=1.985
c101 25 0 2.25722e-20 $X=2.925 $Y=0.74
r102 64 65 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.925 $Y=1.465
+ $X2=2.94 $Y2=1.465
r103 63 64 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.495 $Y=1.465
+ $X2=2.925 $Y2=1.465
r104 62 63 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.49 $Y=1.465
+ $X2=2.495 $Y2=1.465
r105 59 60 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.04 $Y=1.465
+ $X2=2.065 $Y2=1.465
r106 56 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.95 $Y=1.465
+ $X2=2.04 $Y2=1.465
r107 52 53 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=1.985
+ $X2=1.285 $Y2=1.82
r108 49 62 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.37 $Y=1.465
+ $X2=2.49 $Y2=1.465
r109 49 60 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.37 $Y=1.465
+ $X2=2.065 $Y2=1.465
r110 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.465 $X2=2.37 $Y2=1.465
r111 46 56 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.69 $Y=1.465
+ $X2=1.95 $Y2=1.465
r112 45 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.69 $Y=1.465
+ $X2=2.37 $Y2=1.465
r113 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.465 $X2=1.69 $Y2=1.465
r114 43 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.465
+ $X2=1.395 $Y2=1.465
r115 43 45 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.48 $Y=1.465
+ $X2=1.69 $Y2=1.465
r116 41 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=1.63
+ $X2=1.395 $Y2=1.465
r117 41 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.395 $Y=1.63
+ $X2=1.395 $Y2=1.82
r118 40 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=1.3
+ $X2=1.395 $Y2=1.465
r119 40 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.395 $Y=1.3
+ $X2=1.395 $Y2=1.13
r120 35 54 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=1.302 $Y=0.953
+ $X2=1.302 $Y2=1.13
r121 35 37 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=1.302 $Y=0.953
+ $X2=1.302 $Y2=0.515
r122 31 52 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.285 $Y=2.015
+ $X2=1.285 $Y2=1.985
r123 31 33 23.6399 $w=3.88e-07 $l=8e-07 $layer=LI1_cond $X=1.285 $Y=2.015
+ $X2=1.285 $Y2=2.815
r124 27 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.94 $Y=1.63
+ $X2=2.94 $Y2=1.465
r125 27 29 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.94 $Y=1.63
+ $X2=2.94 $Y2=2.4
r126 23 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.3
+ $X2=2.925 $Y2=1.465
r127 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.925 $Y=1.3
+ $X2=2.925 $Y2=0.74
r128 19 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.3
+ $X2=2.495 $Y2=1.465
r129 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.495 $Y=1.3
+ $X2=2.495 $Y2=0.74
r130 15 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.63
+ $X2=2.49 $Y2=1.465
r131 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.49 $Y=1.63
+ $X2=2.49 $Y2=2.4
r132 11 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.3
+ $X2=2.065 $Y2=1.465
r133 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.065 $Y=1.3
+ $X2=2.065 $Y2=0.74
r134 7 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.63
+ $X2=2.04 $Y2=1.465
r135 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.04 $Y=1.63 $X2=2.04
+ $Y2=2.4
r136 2 52 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.84 $X2=1.255 $Y2=1.985
r137 2 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.84 $X2=1.255 $Y2=2.815
r138 1 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.37 $X2=1.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%A_334_368# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 77 79 81 83 87 91 94 100 108 110 132
c202 110 0 2.25722e-20 $X=2.71 $Y=0.965
r203 131 132 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.635 $Y=1.465
+ $X2=6.645 $Y2=1.465
r204 130 131 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.205 $Y=1.465
+ $X2=6.635 $Y2=1.465
r205 129 130 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.465
+ $X2=6.205 $Y2=1.465
r206 126 127 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=5.705 $Y=1.465
+ $X2=5.745 $Y2=1.465
r207 125 126 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=5.295 $Y=1.465
+ $X2=5.705 $Y2=1.465
r208 124 125 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.215 $Y=1.465
+ $X2=5.295 $Y2=1.465
r209 123 124 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.84 $Y=1.465
+ $X2=5.215 $Y2=1.465
r210 122 123 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.785 $Y=1.465
+ $X2=4.84 $Y2=1.465
r211 121 122 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=4.39 $Y=1.465
+ $X2=4.785 $Y2=1.465
r212 120 121 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.355 $Y=1.465
+ $X2=4.39 $Y2=1.465
r213 119 120 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=3.94 $Y=1.465
+ $X2=4.355 $Y2=1.465
r214 118 119 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=3.855 $Y=1.465
+ $X2=3.94 $Y2=1.465
r215 114 116 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.425 $Y=1.465
+ $X2=3.44 $Y2=1.465
r216 112 113 7.83639 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.897 $Y=1.465
+ $X2=2.897 $Y2=1.63
r217 110 112 13.1437 $w=4.53e-07 $l=5e-07 $layer=LI1_cond $X=2.897 $Y=0.965
+ $X2=2.897 $Y2=1.465
r218 101 129 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=5.895 $Y=1.465
+ $X2=6.195 $Y2=1.465
r219 101 127 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.895 $Y=1.465
+ $X2=5.745 $Y2=1.465
r220 100 101 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=5.895
+ $Y=1.465 $X2=5.895 $Y2=1.465
r221 98 118 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.515 $Y=1.465
+ $X2=3.855 $Y2=1.465
r222 98 116 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.515 $Y=1.465
+ $X2=3.44 $Y2=1.465
r223 97 100 83.1156 $w=3.28e-07 $l=2.38e-06 $layer=LI1_cond $X=3.515 $Y=1.465
+ $X2=5.895 $Y2=1.465
r224 97 98 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=3.515
+ $Y=1.465 $X2=3.515 $Y2=1.465
r225 95 112 2.61955 $w=3.3e-07 $l=2.28e-07 $layer=LI1_cond $X=3.125 $Y=1.465
+ $X2=2.897 $Y2=1.465
r226 95 97 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.125 $Y=1.465
+ $X2=3.515 $Y2=1.465
r227 94 108 3.46198 $w=2.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.775 $Y=1.82
+ $X2=2.715 $Y2=1.905
r228 94 113 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.82
+ $X2=2.775 $Y2=1.63
r229 89 108 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=1.99
+ $X2=2.715 $Y2=1.905
r230 89 91 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=2.715 $Y=1.99
+ $X2=2.715 $Y2=2.815
r231 88 104 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=1.905
+ $X2=1.815 $Y2=1.905
r232 87 108 3.05049 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=1.905
+ $X2=2.715 $Y2=1.905
r233 87 88 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.55 $Y=1.905
+ $X2=1.98 $Y2=1.905
r234 86 106 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.935 $Y=1.005
+ $X2=1.81 $Y2=1.005
r235 86 110 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=1.935 $Y=1.005
+ $X2=2.67 $Y2=1.005
r236 81 106 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=0.88
+ $X2=1.81 $Y2=1.005
r237 81 83 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.81 $Y=0.88
+ $X2=1.81 $Y2=0.515
r238 77 104 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=1.99
+ $X2=1.815 $Y2=1.905
r239 77 79 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=1.99
+ $X2=1.815 $Y2=2.815
r240 73 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.635 $Y=1.3
+ $X2=6.635 $Y2=1.465
r241 73 75 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.635 $Y=1.3
+ $X2=6.635 $Y2=0.74
r242 69 132 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.63
+ $X2=6.645 $Y2=1.465
r243 69 71 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.645 $Y=1.63
+ $X2=6.645 $Y2=2.4
r244 65 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=1.465
r245 65 67 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=0.74
r246 61 129 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=1.465
r247 61 63 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=2.4
r248 57 127 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.745 $Y=1.63
+ $X2=5.745 $Y2=1.465
r249 57 59 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.745 $Y=1.63
+ $X2=5.745 $Y2=2.4
r250 53 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.705 $Y=1.3
+ $X2=5.705 $Y2=1.465
r251 53 55 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.705 $Y=1.3
+ $X2=5.705 $Y2=0.74
r252 49 125 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.295 $Y=1.63
+ $X2=5.295 $Y2=1.465
r253 49 51 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.295 $Y=1.63
+ $X2=5.295 $Y2=2.4
r254 45 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.3
+ $X2=5.215 $Y2=1.465
r255 45 47 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.215 $Y=1.3
+ $X2=5.215 $Y2=0.74
r256 41 123 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.63
+ $X2=4.84 $Y2=1.465
r257 41 43 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.84 $Y=1.63
+ $X2=4.84 $Y2=2.4
r258 37 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=1.465
r259 37 39 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=0.74
r260 33 121 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=1.63
+ $X2=4.39 $Y2=1.465
r261 33 35 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.39 $Y=1.63
+ $X2=4.39 $Y2=2.4
r262 29 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=1.465
r263 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=0.74
r264 25 119 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.63
+ $X2=3.94 $Y2=1.465
r265 25 27 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.94 $Y=1.63
+ $X2=3.94 $Y2=2.4
r266 21 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.3
+ $X2=3.855 $Y2=1.465
r267 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.855 $Y=1.3
+ $X2=3.855 $Y2=0.74
r268 17 116 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.63
+ $X2=3.44 $Y2=1.465
r269 17 19 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.44 $Y=1.63
+ $X2=3.44 $Y2=2.4
r270 13 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.3
+ $X2=3.425 $Y2=1.465
r271 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.425 $Y=1.3
+ $X2=3.425 $Y2=0.74
r272 4 108 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.84 $X2=2.715 $Y2=1.985
r273 4 91 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.84 $X2=2.715 $Y2=2.815
r274 3 104 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.84 $X2=1.815 $Y2=1.985
r275 3 79 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.84 $X2=1.815 $Y2=2.815
r276 2 110 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.965
r277 1 106 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.37 $X2=1.85 $Y2=0.965
r278 1 83 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.37 $X2=1.85 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%VPWR 1 2 3 4 5 6 7 24 28 30 34 38 42 46 50
+ 52 54 58 60 65 70 75 80 86 89 92 95 98 101 105
r108 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r110 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 84 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 84 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r118 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r119 81 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.105 $Y=3.33
+ $X2=5.97 $Y2=3.33
r120 81 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=3.33
+ $X2=6.48 $Y2=3.33
r121 80 104 4.41691 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.967 $Y2=3.33
r122 80 83 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 79 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r124 79 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 76 98 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.067 $Y2=3.33
r127 76 78 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 75 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.97 $Y2=3.33
r129 75 78 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 74 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 74 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r133 71 95 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.162 $Y2=3.33
r134 71 73 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 70 98 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.93 $Y=3.33
+ $X2=5.067 $Y2=3.33
r136 70 73 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.93 $Y=3.33
+ $X2=4.56 $Y2=3.33
r137 69 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 66 86 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=0.742 $Y2=3.33
r141 66 68 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 65 89 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.265 $Y2=3.33
r143 65 68 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 60 86 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.742 $Y2=3.33
r147 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 58 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r149 58 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r150 54 57 26.4495 $w=3.03e-07 $l=7e-07 $layer=LI1_cond $X=6.887 $Y=2.115
+ $X2=6.887 $Y2=2.815
r151 52 104 3.14133 $w=3.05e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.887 $Y=3.245
+ $X2=6.967 $Y2=3.33
r152 52 57 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=6.887 $Y=3.245
+ $X2=6.887 $Y2=2.815
r153 48 101 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=3.245
+ $X2=5.97 $Y2=3.33
r154 48 50 40.1221 $w=2.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.97 $Y=3.245
+ $X2=5.97 $Y2=2.305
r155 44 98 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.067 $Y=3.245
+ $X2=5.067 $Y2=3.33
r156 44 46 39.3926 $w=2.73e-07 $l=9.4e-07 $layer=LI1_cond $X=5.067 $Y=3.245
+ $X2=5.067 $Y2=2.305
r157 40 95 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.162 $Y=3.245
+ $X2=4.162 $Y2=3.33
r158 40 42 42.4822 $w=2.53e-07 $l=9.4e-07 $layer=LI1_cond $X=4.162 $Y=3.245
+ $X2=4.162 $Y2=2.305
r159 39 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=3.33
+ $X2=3.215 $Y2=3.33
r160 38 95 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.162 $Y2=3.33
r161 38 39 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.38 $Y2=3.33
r162 34 37 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.215 $Y=1.985
+ $X2=3.215 $Y2=2.815
r163 32 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=3.33
r164 32 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=2.815
r165 31 89 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.265 $Y2=3.33
r166 30 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=3.215 $Y2=3.33
r167 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=2.38 $Y2=3.33
r168 26 89 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=3.245
+ $X2=2.265 $Y2=3.33
r169 26 28 46.0977 $w=2.28e-07 $l=9.2e-07 $layer=LI1_cond $X=2.265 $Y=3.245
+ $X2=2.265 $Y2=2.325
r170 22 86 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=3.33
r171 22 24 23.0489 $w=3.53e-07 $l=7.1e-07 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=2.535
r172 7 57 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.875 $Y2=2.815
r173 7 54 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.875 $Y2=2.115
r174 6 50 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.835
+ $Y=1.84 $X2=5.97 $Y2=2.305
r175 5 46 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.93
+ $Y=1.84 $X2=5.065 $Y2=2.305
r176 4 42 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.03
+ $Y=1.84 $X2=4.165 $Y2=2.305
r177 3 37 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.84 $X2=3.215 $Y2=2.815
r178 3 34 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.84 $X2=3.215 $Y2=1.985
r179 2 28 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=2.13
+ $Y=1.84 $X2=2.265 $Y2=2.325
r180 1 24 600 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.74 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 41 42 45 49
+ 53 57 61 63 65 69 70 71 75
r113 71 75 7.80543 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.96 $Y=1.665
+ $X2=6.665 $Y2=1.665
r114 65 67 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.42 $Y=1.985
+ $X2=6.42 $Y2=2.815
r115 63 65 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.42 $Y=1.97
+ $X2=6.42 $Y2=1.985
r116 59 61 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=6.42 $Y=0.88
+ $X2=6.42 $Y2=0.515
r117 58 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.655 $Y=1.885
+ $X2=5.52 $Y2=1.885
r118 57 63 5.08453 $w=5.54e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.255 $Y=1.885
+ $X2=6.42 $Y2=1.97
r119 57 75 4.84477 $w=5.54e-07 $l=5.08232e-07 $layer=LI1_cond $X=6.255 $Y=1.885
+ $X2=6.665 $Y2=1.665
r120 57 58 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.255 $Y=1.885
+ $X2=5.655 $Y2=1.885
r121 53 55 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=5.52 $Y=1.985
+ $X2=5.52 $Y2=2.815
r122 51 70 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=1.97
+ $X2=5.52 $Y2=1.885
r123 51 53 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.52 $Y=1.97
+ $X2=5.52 $Y2=1.985
r124 50 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.745 $Y=1.885
+ $X2=4.62 $Y2=1.885
r125 49 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.385 $Y=1.885
+ $X2=5.52 $Y2=1.885
r126 49 50 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.385 $Y=1.885
+ $X2=4.745 $Y2=1.885
r127 45 47 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.62 $Y=1.985
+ $X2=4.62 $Y2=2.815
r128 43 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=1.97
+ $X2=4.62 $Y2=1.885
r129 43 45 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=4.62 $Y=1.97
+ $X2=4.62 $Y2=1.985
r130 41 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=1.885
+ $X2=4.62 $Y2=1.885
r131 41 42 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.495 $Y=1.885
+ $X2=3.83 $Y2=1.885
r132 38 40 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=4.57 $Y=1.005
+ $X2=5.46 $Y2=1.005
r133 36 38 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=3.805 $Y=1.005
+ $X2=4.57 $Y2=1.005
r134 35 75 14.5343 $w=5.54e-07 $l=8.40357e-07 $layer=LI1_cond $X=6.255 $Y=1.005
+ $X2=6.665 $Y2=1.665
r135 35 59 4.73129 $w=5.54e-07 $l=2.18746e-07 $layer=LI1_cond $X=6.255 $Y=1.005
+ $X2=6.42 $Y2=0.88
r136 35 40 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=6.255 $Y=1.005
+ $X2=5.46 $Y2=1.005
r137 31 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=3.697 $Y=1.985
+ $X2=3.697 $Y2=2.815
r138 29 42 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=3.697 $Y=1.97
+ $X2=3.83 $Y2=1.885
r139 29 31 0.652326 $w=2.63e-07 $l=1.5e-08 $layer=LI1_cond $X=3.697 $Y=1.97
+ $X2=3.697 $Y2=1.985
r140 25 36 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.805 $Y2=1.005
r141 25 27 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.64 $Y=0.88
+ $X2=3.64 $Y2=0.515
r142 8 67 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=2.815
r143 8 65 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=1.985
r144 7 55 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.84 $X2=5.52 $Y2=2.815
r145 7 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.84 $X2=5.52 $Y2=1.985
r146 6 47 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.84 $X2=4.615 $Y2=2.815
r147 6 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.84 $X2=4.615 $Y2=1.985
r148 5 33 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.84 $X2=3.715 $Y2=2.815
r149 5 31 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.84 $X2=3.715 $Y2=1.985
r150 4 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.37 $X2=6.42 $Y2=0.515
r151 3 40 182 $w=1.7e-07 $l=6.74667e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.37 $X2=5.46 $Y2=0.965
r152 2 38 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.965
r153 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.37 $X2=3.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_8%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 50 52 57 62 67 72 77 82 88 91 94 97 100 103 107
r101 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r102 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r103 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r104 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r106 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r107 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r108 86 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r109 86 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r110 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r111 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=5.92 $Y2=0
r112 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=0
+ $X2=6.48 $Y2=0
r113 82 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.977 $Y2=0
r114 82 85 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.48 $Y2=0
r115 81 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r116 81 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r117 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r118 78 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r119 78 80 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r120 77 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.92 $Y2=0
r121 77 80 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.52 $Y2=0
r122 76 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r123 76 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r124 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r125 73 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.14
+ $Y2=0
r126 73 75 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=0
+ $X2=4.56 $Y2=0
r127 72 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r128 72 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.56 $Y2=0
r129 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r130 68 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r131 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=4.14
+ $Y2=0
r132 67 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.6
+ $Y2=0
r133 66 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r134 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r135 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r136 63 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.28
+ $Y2=0
r137 63 65 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=0
+ $X2=2.64 $Y2=0
r138 62 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r139 62 65 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r140 61 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r141 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r142 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r143 58 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r144 58 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r145 57 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.28
+ $Y2=0
r146 57 60 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.2
+ $Y2=0
r147 55 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r148 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r149 52 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r150 52 54 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r151 50 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r152 50 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r153 50 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r154 46 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r155 46 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r156 42 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r157 42 44 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.545
r158 38 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r159 38 40 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.545
r160 34 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r161 34 36 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.545
r162 30 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r163 30 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.545
r164 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r165 26 28 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.545
r166 22 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r167 22 24 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.675
r168 7 48 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.71
+ $Y=0.37 $X2=6.92 $Y2=0.515
r169 6 44 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.37 $X2=5.92 $Y2=0.545
r170 5 40 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.545
r171 4 36 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.14 $Y2=0.545
r172 3 32 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.14 $Y2=0.545
r173 2 28 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.37 $X2=2.28 $Y2=0.545
r174 1 24 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.79 $Y2=0.675
.ends


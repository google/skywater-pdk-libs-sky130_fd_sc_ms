* File: sky130_fd_sc_ms__o2111ai_1.pxi.spice
* Created: Fri Aug 28 17:51:57 2020
* 
x_PM_SKY130_FD_SC_MS__O2111AI_1%D1 N_D1_M1008_g N_D1_M1006_g D1 N_D1_c_56_n
+ N_D1_c_57_n PM_SKY130_FD_SC_MS__O2111AI_1%D1
x_PM_SKY130_FD_SC_MS__O2111AI_1%C1 N_C1_M1007_g N_C1_M1009_g C1 C1 C1
+ N_C1_c_85_n N_C1_c_86_n PM_SKY130_FD_SC_MS__O2111AI_1%C1
x_PM_SKY130_FD_SC_MS__O2111AI_1%B1 N_B1_M1000_g N_B1_M1004_g B1 N_B1_c_124_n
+ N_B1_c_125_n N_B1_c_126_n PM_SKY130_FD_SC_MS__O2111AI_1%B1
x_PM_SKY130_FD_SC_MS__O2111AI_1%A2 N_A2_M1002_g N_A2_M1003_g A2 N_A2_c_158_n
+ N_A2_c_159_n PM_SKY130_FD_SC_MS__O2111AI_1%A2
x_PM_SKY130_FD_SC_MS__O2111AI_1%A1 N_A1_M1001_g N_A1_c_191_n N_A1_M1005_g A1
+ N_A1_c_193_n PM_SKY130_FD_SC_MS__O2111AI_1%A1
x_PM_SKY130_FD_SC_MS__O2111AI_1%VPWR N_VPWR_M1008_s N_VPWR_M1009_d
+ N_VPWR_M1001_d N_VPWR_c_217_n N_VPWR_c_218_n N_VPWR_c_219_n N_VPWR_c_220_n
+ N_VPWR_c_221_n N_VPWR_c_222_n VPWR N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_216_n PM_SKY130_FD_SC_MS__O2111AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O2111AI_1%Y N_Y_M1006_s N_Y_M1008_d N_Y_M1004_d
+ N_Y_c_258_n N_Y_c_261_n N_Y_c_262_n N_Y_c_263_n N_Y_c_264_n N_Y_c_259_n
+ N_Y_c_265_n Y Y Y N_Y_c_266_n PM_SKY130_FD_SC_MS__O2111AI_1%Y
x_PM_SKY130_FD_SC_MS__O2111AI_1%A_368_74# N_A_368_74#_M1000_d
+ N_A_368_74#_M1005_d N_A_368_74#_c_321_n N_A_368_74#_c_318_n
+ N_A_368_74#_c_319_n N_A_368_74#_c_320_n
+ PM_SKY130_FD_SC_MS__O2111AI_1%A_368_74#
x_PM_SKY130_FD_SC_MS__O2111AI_1%VGND N_VGND_M1002_d N_VGND_c_346_n VGND
+ N_VGND_c_347_n N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n
+ PM_SKY130_FD_SC_MS__O2111AI_1%VGND
cc_1 VNB N_D1_M1008_g 0.00715433f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.4
cc_2 VNB D1 0.00350742f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_D1_c_56_n 0.0350627f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_4 VNB N_D1_c_57_n 0.0217968f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.22
cc_5 VNB N_C1_M1009_g 0.00688061f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.74
cc_6 VNB C1 0.00553803f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_C1_c_85_n 0.0302626f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.295
cc_8 VNB N_C1_c_86_n 0.0172466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_M1004_g 0.00698513f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.74
cc_10 VNB N_B1_c_124_n 0.0272566f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_11 VNB N_B1_c_125_n 0.0102576f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_12 VNB N_B1_c_126_n 0.0190408f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.22
cc_13 VNB N_A2_M1003_g 0.00632425f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.74
cc_14 VNB A2 0.0144016f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_A2_c_158_n 0.0289335f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_16 VNB N_A2_c_159_n 0.0186396f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.22
cc_17 VNB N_A1_M1001_g 0.0093905f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.4
cc_18 VNB N_A1_c_191_n 0.0247091f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.22
cc_19 VNB A1 0.00922063f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A1_c_193_n 0.0588931f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.55
cc_21 VNB N_VPWR_c_216_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_258_n 0.0309816f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_23 VNB N_Y_c_259_n 0.0331431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_368_74#_c_318_n 0.00289626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_368_74#_c_319_n 0.00716806f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_26 VNB N_A_368_74#_c_320_n 0.021252f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.295
cc_27 VNB N_VGND_c_346_n 0.00739995f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.74
cc_28 VNB N_VGND_c_347_n 0.0659727f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.385
cc_29 VNB N_VGND_c_348_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_349_n 0.219739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_350_n 0.00786346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_D1_M1008_g 0.0248898f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=2.4
cc_33 VPB N_C1_M1009_g 0.0238885f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=0.74
cc_34 VPB N_B1_M1004_g 0.0233499f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=0.74
cc_35 VPB N_A2_M1003_g 0.023181f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=0.74
cc_36 VPB N_A1_M1001_g 0.029635f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=2.4
cc_37 VPB N_VPWR_c_217_n 0.0476286f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.385
cc_38 VPB N_VPWR_c_218_n 0.00666562f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.385
cc_39 VPB N_VPWR_c_219_n 0.0127942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_220_n 0.0555804f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_221_n 0.0142356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_222_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_223_n 0.0212158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_224_n 0.0312467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_225_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_216_n 0.0781978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_258_n 0.00311325f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.385
cc_48 VPB N_Y_c_261_n 0.0157847f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.385
cc_49 VPB N_Y_c_262_n 0.0148348f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.22
cc_50 VPB N_Y_c_263_n 0.0165547f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.55
cc_51 VPB N_Y_c_264_n 0.00253059f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.385
cc_52 VPB N_Y_c_265_n 0.00785442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_Y_c_266_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 N_D1_M1008_g N_C1_M1009_g 0.0231601f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_55 D1 C1 0.028682f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_D1_c_57_n C1 0.0100911f $X=0.745 $Y=1.22 $X2=0 $Y2=0
cc_57 D1 N_C1_c_85_n 3.85374e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_D1_c_56_n N_C1_c_85_n 0.0206451f $X=0.745 $Y=1.385 $X2=0 $Y2=0
cc_59 N_D1_c_57_n N_C1_c_86_n 0.0499419f $X=0.745 $Y=1.22 $X2=0 $Y2=0
cc_60 N_D1_M1008_g N_VPWR_c_217_n 0.00534567f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_61 N_D1_M1008_g N_VPWR_c_223_n 0.005209f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_62 N_D1_M1008_g N_VPWR_c_216_n 0.00986837f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_63 N_D1_M1008_g N_Y_c_258_n 0.00442066f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_64 D1 N_Y_c_258_n 0.0186037f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_D1_c_56_n N_Y_c_258_n 0.00678078f $X=0.745 $Y=1.385 $X2=0 $Y2=0
cc_66 N_D1_c_57_n N_Y_c_258_n 0.00317526f $X=0.745 $Y=1.22 $X2=0 $Y2=0
cc_67 N_D1_M1008_g N_Y_c_261_n 0.0149054f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_68 D1 N_Y_c_261_n 0.0221856f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_D1_c_56_n N_Y_c_261_n 0.00105037f $X=0.745 $Y=1.385 $X2=0 $Y2=0
cc_70 D1 N_Y_c_259_n 0.0150353f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_D1_c_56_n N_Y_c_259_n 0.00110088f $X=0.745 $Y=1.385 $X2=0 $Y2=0
cc_72 N_D1_c_57_n N_Y_c_259_n 0.0105771f $X=0.745 $Y=1.22 $X2=0 $Y2=0
cc_73 N_D1_M1008_g N_Y_c_265_n 0.00224432f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_74 D1 N_Y_c_265_n 0.00234631f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_D1_M1008_g N_Y_c_266_n 0.0195664f $X=0.82 $Y=2.4 $X2=0 $Y2=0
cc_76 N_D1_c_57_n N_VGND_c_347_n 0.00433162f $X=0.745 $Y=1.22 $X2=0 $Y2=0
cc_77 N_D1_c_57_n N_VGND_c_349_n 0.00822327f $X=0.745 $Y=1.22 $X2=0 $Y2=0
cc_78 N_C1_M1009_g N_B1_M1004_g 0.0231672f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_79 C1 N_B1_c_124_n 3.45051e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_80 N_C1_c_85_n N_B1_c_124_n 0.0205652f $X=1.285 $Y=1.385 $X2=0 $Y2=0
cc_81 C1 N_B1_c_125_n 0.0299123f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_82 N_C1_c_85_n N_B1_c_125_n 0.00198614f $X=1.285 $Y=1.385 $X2=0 $Y2=0
cc_83 C1 N_B1_c_126_n 0.00865512f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_84 N_C1_c_86_n N_B1_c_126_n 0.0274744f $X=1.285 $Y=1.22 $X2=0 $Y2=0
cc_85 N_C1_M1009_g N_VPWR_c_218_n 0.0107702f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_86 N_C1_M1009_g N_VPWR_c_223_n 0.00401934f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_87 N_C1_M1009_g N_VPWR_c_216_n 0.00599837f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_88 N_C1_M1009_g N_Y_c_263_n 0.00602435f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_89 C1 N_Y_c_263_n 0.00850845f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_90 N_C1_c_85_n N_Y_c_263_n 0.00142789f $X=1.285 $Y=1.385 $X2=0 $Y2=0
cc_91 N_C1_M1009_g N_Y_c_264_n 6.5456e-19 $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_92 C1 N_Y_c_259_n 0.030281f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_93 N_C1_c_86_n N_Y_c_259_n 9.85906e-19 $X=1.285 $Y=1.22 $X2=0 $Y2=0
cc_94 N_C1_M1009_g N_Y_c_265_n 0.00545707f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_95 C1 N_Y_c_265_n 0.0199629f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_96 N_C1_c_85_n N_Y_c_265_n 4.7205e-19 $X=1.285 $Y=1.385 $X2=0 $Y2=0
cc_97 N_C1_M1009_g N_Y_c_266_n 0.0239293f $X=1.27 $Y=2.4 $X2=0 $Y2=0
cc_98 C1 A_182_74# 0.00751072f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_99 C1 A_260_74# 0.00953457f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_100 C1 N_A_368_74#_c_321_n 0.00723659f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_101 C1 N_A_368_74#_c_318_n 0.0160909f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_102 N_C1_c_86_n N_A_368_74#_c_318_n 7.73661e-19 $X=1.285 $Y=1.22 $X2=0 $Y2=0
cc_103 C1 N_VGND_c_347_n 0.00877891f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_C1_c_86_n N_VGND_c_347_n 0.00303293f $X=1.285 $Y=1.22 $X2=0 $Y2=0
cc_105 C1 N_VGND_c_349_n 0.0110375f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_106 N_C1_c_86_n N_VGND_c_349_n 0.00372419f $X=1.285 $Y=1.22 $X2=0 $Y2=0
cc_107 N_B1_M1004_g N_A2_M1003_g 0.0213919f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_108 N_B1_c_124_n A2 4.1351e-19 $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_109 N_B1_c_125_n A2 0.0249496f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_110 N_B1_c_124_n N_A2_c_158_n 0.0214219f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_111 N_B1_c_125_n N_A2_c_158_n 4.15266e-19 $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_112 N_B1_c_126_n N_A2_c_159_n 0.0193073f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_113 N_B1_M1004_g N_VPWR_c_218_n 0.0163325f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_114 N_B1_M1004_g N_VPWR_c_224_n 0.00532442f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_115 N_B1_M1004_g N_VPWR_c_216_n 0.0104097f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B1_M1004_g N_Y_c_263_n 0.0170372f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_117 N_B1_c_124_n N_Y_c_263_n 0.00383587f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_118 N_B1_c_125_n N_Y_c_263_n 0.0295555f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_119 N_B1_M1004_g N_Y_c_264_n 0.0170474f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_120 N_B1_M1004_g N_Y_c_266_n 5.2051e-19 $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_121 N_B1_c_124_n N_A_368_74#_c_321_n 8.8929e-19 $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_122 N_B1_c_125_n N_A_368_74#_c_321_n 0.011699f $X=1.825 $Y=1.385 $X2=0 $Y2=0
cc_123 N_B1_c_126_n N_A_368_74#_c_321_n 0.0027133f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_124 N_B1_c_126_n N_A_368_74#_c_318_n 0.0082564f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_125 N_B1_c_126_n N_VGND_c_346_n 5.94017e-19 $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_126 N_B1_c_126_n N_VGND_c_347_n 0.00445602f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_127 N_B1_c_126_n N_VGND_c_349_n 0.00859779f $X=1.825 $Y=1.22 $X2=0 $Y2=0
cc_128 N_A2_M1003_g N_A1_M1001_g 0.0688833f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_129 A2 N_A1_c_191_n 3.9318e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_159_n N_A1_c_191_n 0.0198738f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_131 A2 A1 0.0290366f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A2_c_158_n A1 2.10483e-19 $X=2.365 $Y=1.385 $X2=0 $Y2=0
cc_133 A2 N_A1_c_193_n 0.00914335f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A2_c_158_n N_A1_c_193_n 0.0214735f $X=2.365 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A2_M1003_g N_VPWR_c_218_n 7.56227e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A2_M1003_g N_VPWR_c_220_n 0.00394073f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A2_M1003_g N_VPWR_c_224_n 0.005209f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A2_M1003_g N_VPWR_c_216_n 0.00983865f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A2_M1003_g N_Y_c_263_n 0.00532176f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_140 A2 N_Y_c_263_n 0.00963966f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A2_c_158_n N_Y_c_263_n 0.00231539f $X=2.365 $Y=1.385 $X2=0 $Y2=0
cc_142 N_A2_M1003_g N_Y_c_264_n 0.02211f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A2_c_159_n N_A_368_74#_c_318_n 0.00267906f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_144 A2 N_A_368_74#_c_319_n 0.0398068f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A2_c_158_n N_A_368_74#_c_319_n 0.00101161f $X=2.365 $Y=1.385 $X2=0
+ $Y2=0
cc_146 N_A2_c_159_n N_A_368_74#_c_319_n 0.0128517f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_147 N_A2_c_159_n N_A_368_74#_c_320_n 8.66094e-19 $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A2_c_159_n N_VGND_c_346_n 0.00759f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A2_c_159_n N_VGND_c_347_n 0.00383152f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A2_c_159_n N_VGND_c_349_n 0.0038476f $X=2.365 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A1_M1001_g N_VPWR_c_220_n 0.0305651f $X=2.83 $Y=2.4 $X2=0 $Y2=0
cc_152 A1 N_VPWR_c_220_n 0.017696f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A1_c_193_n N_VPWR_c_220_n 0.00245199f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_154 N_A1_M1001_g N_VPWR_c_224_n 0.00460063f $X=2.83 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A1_M1001_g N_VPWR_c_216_n 0.00908712f $X=2.83 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A1_M1001_g N_Y_c_263_n 6.75676e-19 $X=2.83 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A1_M1001_g N_Y_c_264_n 0.00319844f $X=2.83 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A1_c_191_n N_A_368_74#_c_319_n 0.013911f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_159 A1 N_A_368_74#_c_319_n 0.0252927f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A1_c_193_n N_A_368_74#_c_319_n 0.00199248f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_161 N_A1_c_191_n N_A_368_74#_c_320_n 0.00854971f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_162 N_A1_c_191_n N_VGND_c_346_n 0.00499784f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A1_c_191_n N_VGND_c_348_n 0.00434272f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A1_c_191_n N_VGND_c_349_n 0.00449889f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_165 N_VPWR_M1008_s N_Y_c_261_n 0.00330887f $X=0.4 $Y=1.84 $X2=0 $Y2=0
cc_166 N_VPWR_c_217_n N_Y_c_261_n 0.0238156f $X=0.545 $Y=2.145 $X2=0 $Y2=0
cc_167 N_VPWR_M1009_d N_Y_c_263_n 0.00571509f $X=1.36 $Y=1.84 $X2=0 $Y2=0
cc_168 N_VPWR_c_218_n N_Y_c_263_n 0.0219853f $X=1.65 $Y=2.145 $X2=0 $Y2=0
cc_169 N_VPWR_c_220_n N_Y_c_263_n 0.00203965f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_170 N_VPWR_c_218_n N_Y_c_264_n 0.0690412f $X=1.65 $Y=2.145 $X2=0 $Y2=0
cc_171 N_VPWR_c_220_n N_Y_c_264_n 0.029939f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_172 N_VPWR_c_224_n N_Y_c_264_n 0.014537f $X=2.89 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_c_216_n N_Y_c_264_n 0.011955f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_217_n N_Y_c_266_n 0.0368013f $X=0.545 $Y=2.145 $X2=0 $Y2=0
cc_175 N_VPWR_c_218_n N_Y_c_266_n 0.0729356f $X=1.65 $Y=2.145 $X2=0 $Y2=0
cc_176 N_VPWR_c_223_n N_Y_c_266_n 0.0188336f $X=1.485 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_c_216_n N_Y_c_266_n 0.0152059f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_178 N_Y_c_259_n N_VGND_c_347_n 0.0296309f $X=0.62 $Y=0.515 $X2=0 $Y2=0
cc_179 N_Y_c_259_n N_VGND_c_349_n 0.024582f $X=0.62 $Y=0.515 $X2=0 $Y2=0
cc_180 N_A_368_74#_c_319_n N_VGND_M1002_d 0.00792129f $X=2.915 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_181 N_A_368_74#_c_318_n N_VGND_c_346_n 0.0105237f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_182 N_A_368_74#_c_319_n N_VGND_c_346_n 0.0207516f $X=2.915 $Y=0.925 $X2=0
+ $Y2=0
cc_183 N_A_368_74#_c_320_n N_VGND_c_346_n 0.0102004f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_184 N_A_368_74#_c_318_n N_VGND_c_347_n 0.0145621f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_185 N_A_368_74#_c_320_n N_VGND_c_348_n 0.0145323f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0
cc_186 N_A_368_74#_c_318_n N_VGND_c_349_n 0.0120343f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_187 N_A_368_74#_c_319_n N_VGND_c_349_n 0.0115465f $X=2.915 $Y=0.925 $X2=0
+ $Y2=0
cc_188 N_A_368_74#_c_320_n N_VGND_c_349_n 0.0119861f $X=3.08 $Y=0.515 $X2=0
+ $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__and2b_2 A_N B VGND VNB VPB VPWR X
M1000 a_505_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=8.742e+11p ps=5.41e+06u
M1001 a_198_48# a_27_74# a_505_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 VPWR a_198_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.45745e+12p pd=9.24e+06u as=3.024e+11p ps=2.78e+06u
M1003 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1004 VGND a_198_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 a_198_48# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1006 VPWR a_27_74# a_198_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 X a_198_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_198_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__dlymetal6s4s_1.pxi.spice
* Created: Wed Sep  2 12:07:18 2020
* 
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A N_A_M1000_g N_A_M1006_g A N_A_c_96_n
+ N_A_c_97_n PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_28_138# N_A_28_138#_M1006_s
+ N_A_28_138#_M1000_s N_A_28_138#_M1002_g N_A_28_138#_M1003_g
+ N_A_28_138#_c_128_n N_A_28_138#_c_141_n N_A_28_138#_c_129_n
+ N_A_28_138#_c_130_n N_A_28_138#_c_131_n N_A_28_138#_c_135_n
+ N_A_28_138#_c_132_n PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_28_138#
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_209_74# N_A_209_74#_M1002_d
+ N_A_209_74#_M1003_d N_A_209_74#_M1007_g N_A_209_74#_M1004_g
+ N_A_209_74#_c_194_n N_A_209_74#_c_195_n N_A_209_74#_c_196_n
+ N_A_209_74#_c_197_n N_A_209_74#_c_202_n N_A_209_74#_c_198_n
+ N_A_209_74#_c_199_n N_A_209_74#_c_200_n N_A_209_74#_c_204_n
+ PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_209_74#
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_316_138# N_A_316_138#_M1007_s
+ N_A_316_138#_M1004_s N_A_316_138#_M1008_g N_A_316_138#_M1009_g
+ N_A_316_138#_c_264_n N_A_316_138#_c_278_n N_A_316_138#_c_265_n
+ N_A_316_138#_c_266_n N_A_316_138#_c_267_n N_A_316_138#_c_271_n
+ N_A_316_138#_c_268_n PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_316_138#
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%X N_X_M1008_d N_X_M1009_d N_X_M1001_g
+ N_X_M1010_g N_X_c_336_n N_X_c_344_n N_X_c_337_n N_X_c_338_n N_X_c_339_n
+ N_X_c_340_n X N_X_c_341_n N_X_c_346_n N_X_c_342_n N_X_c_352_n N_X_c_348_n
+ PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%X
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_604_138# N_A_604_138#_M1001_s
+ N_A_604_138#_M1010_s N_A_604_138#_M1005_g N_A_604_138#_M1011_g
+ N_A_604_138#_c_436_n N_A_604_138#_c_424_n N_A_604_138#_c_425_n
+ N_A_604_138#_c_426_n N_A_604_138#_c_427_n N_A_604_138#_c_431_n
+ N_A_604_138#_c_428_n PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_604_138#
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%VPWR N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_M1010_d N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n VPWR
+ N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_486_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n VPWR
+ PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%VPWR
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_785_74# N_A_785_74#_M1005_d
+ N_A_785_74#_M1011_d N_A_785_74#_c_535_n N_A_785_74#_c_538_n
+ N_A_785_74#_c_536_n N_A_785_74#_c_539_n N_A_785_74#_c_537_n
+ PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%A_785_74#
x_PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%VGND N_VGND_M1006_d N_VGND_M1007_d
+ N_VGND_M1001_d N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n VGND
+ N_VGND_c_571_n N_VGND_c_572_n N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n
+ N_VGND_c_576_n N_VGND_c_577_n N_VGND_c_578_n VGND
+ PM_SKY130_FD_SC_MS__DLYMETAL6S4S_1%VGND
cc_1 VNB N_A_M1000_g 0.00370597f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.05
cc_2 VNB N_A_M1006_g 0.0286178f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.9
cc_3 VNB N_A_c_96_n 0.0390579f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_4 VNB N_A_c_97_n 0.0129985f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_5 VNB N_A_28_138#_M1002_g 0.0217641f $X=-0.19 $Y=-0.245 $X2=0.16 $Y2=1.58
cc_6 VNB N_A_28_138#_M1003_g 0.00334836f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_7 VNB N_A_28_138#_c_128_n 0.00533825f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.605
cc_8 VNB N_A_28_138#_c_129_n 0.00430876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_138#_c_130_n 7.0366e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_138#_c_131_n 0.0201928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_138#_c_132_n 0.0352396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_209_74#_M1007_g 0.0235592f $X=-0.19 $Y=-0.245 $X2=0.16 $Y2=1.58
cc_13 VNB N_A_209_74#_M1004_g 0.00371635f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_14 VNB N_A_209_74#_c_194_n 0.0137727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_209_74#_c_195_n 0.00523129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_209_74#_c_196_n 0.0159058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_209_74#_c_197_n 0.038581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_209_74#_c_198_n 0.00139382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_209_74#_c_199_n 0.00140045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_209_74#_c_200_n 0.00344243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_316_138#_M1008_g 0.0218556f $X=-0.19 $Y=-0.245 $X2=0.16 $Y2=1.58
cc_22 VNB N_A_316_138#_M1009_g 0.00334941f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_23 VNB N_A_316_138#_c_264_n 0.00420983f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.605
cc_24 VNB N_A_316_138#_c_265_n 0.00578839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_316_138#_c_266_n 9.03105e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_316_138#_c_267_n 0.00632352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_316_138#_c_268_n 0.0350051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_M1001_g 0.0234006f $X=-0.19 $Y=-0.245 $X2=0.16 $Y2=1.58
cc_29 VNB N_X_M1010_g 0.00372339f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_30 VNB N_X_c_336_n 0.0147539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_337_n 0.00530393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_338_n 0.0160421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_339_n 0.00190862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_340_n 0.00344243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_341_n 0.042286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_342_n 0.00141397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_604_138#_M1005_g 0.0223301f $X=-0.19 $Y=-0.245 $X2=0.16 $Y2=1.58
cc_38 VNB N_A_604_138#_M1011_g 0.00335659f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_39 VNB N_A_604_138#_c_424_n 0.0029852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_604_138#_c_425_n 0.00174446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_604_138#_c_426_n 0.00547088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_604_138#_c_427_n 9.14932e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_604_138#_c_428_n 0.0339497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_486_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_785_74#_c_535_n 0.0318665f $X=-0.19 $Y=-0.245 $X2=0.16 $Y2=1.58
cc_46 VNB N_A_785_74#_c_536_n 0.00832176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_785_74#_c_537_n 0.0274113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_568_n 0.0187976f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.44
cc_49 VNB N_VGND_c_569_n 0.0125165f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.44
cc_50 VNB N_VGND_c_570_n 0.012298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_571_n 0.0197723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_572_n 0.0312845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_573_n 0.031135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_574_n 0.0302512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_575_n 0.314614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_576_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_577_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_578_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_A_M1000_g 0.0351987f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=2.05
cc_60 VPB N_A_c_97_n 0.00680159f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_61 VPB N_A_28_138#_M1003_g 0.0264301f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_62 VPB N_A_28_138#_c_130_n 0.002828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_28_138#_c_135_n 0.0138694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_209_74#_M1004_g 0.0274775f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_65 VPB N_A_209_74#_c_202_n 0.00566062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_209_74#_c_198_n 0.00417001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_209_74#_c_204_n 0.0302425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_316_138#_M1009_g 0.0264255f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_69 VPB N_A_316_138#_c_266_n 0.00316663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_316_138#_c_271_n 0.00465887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_X_M1010_g 0.0275239f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_72 VPB N_X_c_344_n 0.0287596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB X 0.036744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_346_n 0.00715823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_X_c_342_n 0.00423493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_X_c_348_n 0.0357173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_604_138#_M1011_g 0.0277434f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_78 VPB N_A_604_138#_c_427_n 0.00324941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_604_138#_c_431_n 0.00357166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_487_n 0.0363175f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_81 VPB N_VPWR_c_488_n 0.0332875f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.44
cc_82 VPB N_VPWR_c_489_n 0.0332856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_490_n 0.0209183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_491_n 0.035526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_492_n 0.0348287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_493_n 0.0284932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_486_n 0.14732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_495_n 0.00564836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_496_n 0.00564503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_497_n 0.00564503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_785_74#_c_538_n 0.0366817f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.44
cc_92 VPB N_A_785_74#_c_539_n 0.0164498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_785_74#_c_537_n 0.00789092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_A_28_138#_M1002_g 0.0165166f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_95 N_A_M1000_g N_A_28_138#_M1003_g 0.0223413f $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_96 N_A_M1006_g N_A_28_138#_c_128_n 0.0142256f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_97 N_A_c_96_n N_A_28_138#_c_128_n 0.00134417f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_98 N_A_c_97_n N_A_28_138#_c_128_n 0.00983824f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_99 N_A_M1000_g N_A_28_138#_c_141_n 0.0140609f $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_100 N_A_M1006_g N_A_28_138#_c_129_n 0.0027595f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_101 N_A_c_96_n N_A_28_138#_c_129_n 0.00339828f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_102 N_A_c_97_n N_A_28_138#_c_129_n 0.0202668f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_103 N_A_M1000_g N_A_28_138#_c_130_n 0.00478677f $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_104 N_A_c_97_n N_A_28_138#_c_130_n 0.0122394f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_105 N_A_M1006_g N_A_28_138#_c_131_n 0.00158922f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_106 N_A_c_96_n N_A_28_138#_c_131_n 0.00417844f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_107 N_A_c_97_n N_A_28_138#_c_131_n 0.0209233f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_108 N_A_M1000_g N_A_28_138#_c_135_n 0.00381879f $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_109 N_A_c_96_n N_A_28_138#_c_135_n 7.69058e-19 $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_110 N_A_c_97_n N_A_28_138#_c_135_n 0.0335151f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_111 N_A_M1006_g N_A_28_138#_c_132_n 7.45276e-19 $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_112 N_A_c_96_n N_A_28_138#_c_132_n 0.0206625f $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_113 N_A_c_97_n N_A_28_138#_c_132_n 2.61364e-19 $X=0.39 $Y=1.44 $X2=0 $Y2=0
cc_114 N_A_M1000_g N_A_209_74#_c_202_n 2.24942e-19 $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_115 N_A_M1000_g N_A_209_74#_c_204_n 7.10715e-19 $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_116 N_A_M1000_g N_VPWR_c_487_n 0.00232657f $X=0.49 $Y=2.05 $X2=0 $Y2=0
cc_117 N_A_M1006_g N_VGND_c_568_n 0.00429157f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_118 N_A_M1006_g N_VGND_c_571_n 0.00382655f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_119 N_A_M1006_g N_VGND_c_575_n 0.00451834f $X=0.48 $Y=0.9 $X2=0 $Y2=0
cc_120 N_A_28_138#_M1002_g N_A_209_74#_c_194_n 0.00268996f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_28_138#_M1002_g N_A_209_74#_c_195_n 0.00332518f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_122 N_A_28_138#_c_129_n N_A_209_74#_c_195_n 0.0122064f $X=0.81 $Y=1.605 $X2=0
+ $Y2=0
cc_123 N_A_28_138#_c_132_n N_A_209_74#_c_195_n 8.26384e-19 $X=0.955 $Y=1.44
+ $X2=0 $Y2=0
cc_124 N_A_28_138#_c_132_n N_A_209_74#_c_197_n 0.00507369f $X=0.955 $Y=1.44
+ $X2=0 $Y2=0
cc_125 N_A_28_138#_M1003_g N_A_209_74#_c_202_n 0.00297266f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_126 N_A_28_138#_c_130_n N_A_209_74#_c_202_n 0.00380645f $X=0.81 $Y=1.935
+ $X2=0 $Y2=0
cc_127 N_A_28_138#_c_132_n N_A_209_74#_c_202_n 0.00104646f $X=0.955 $Y=1.44
+ $X2=0 $Y2=0
cc_128 N_A_28_138#_M1003_g N_A_209_74#_c_198_n 0.00525393f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_129 N_A_28_138#_c_130_n N_A_209_74#_c_198_n 0.0111911f $X=0.81 $Y=1.935 $X2=0
+ $Y2=0
cc_130 N_A_28_138#_c_132_n N_A_209_74#_c_199_n 0.00102685f $X=0.955 $Y=1.44
+ $X2=0 $Y2=0
cc_131 N_A_28_138#_c_129_n N_A_209_74#_c_200_n 0.0244957f $X=0.81 $Y=1.605 $X2=0
+ $Y2=0
cc_132 N_A_28_138#_c_132_n N_A_209_74#_c_200_n 0.00341845f $X=0.955 $Y=1.44
+ $X2=0 $Y2=0
cc_133 N_A_28_138#_M1003_g N_A_209_74#_c_204_n 0.0218733f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_134 N_A_28_138#_c_141_n N_A_209_74#_c_204_n 0.00629937f $X=0.725 $Y=2.037
+ $X2=0 $Y2=0
cc_135 N_A_28_138#_c_129_n N_A_209_74#_c_204_n 0.00274452f $X=0.81 $Y=1.605
+ $X2=0 $Y2=0
cc_136 N_A_28_138#_c_130_n N_A_209_74#_c_204_n 4.40431e-19 $X=0.81 $Y=1.935
+ $X2=0 $Y2=0
cc_137 N_A_28_138#_c_135_n N_A_209_74#_c_204_n 0.00216661f $X=0.43 $Y=2.08 $X2=0
+ $Y2=0
cc_138 N_A_28_138#_M1003_g N_A_316_138#_c_271_n 6.34727e-19 $X=1.005 $Y=2.4
+ $X2=0 $Y2=0
cc_139 N_A_28_138#_M1003_g N_X_c_348_n 0.00653278f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_28_138#_c_141_n N_VPWR_M1000_d 0.00689854f $X=0.725 $Y=2.037
+ $X2=-0.19 $Y2=-0.245
cc_141 N_A_28_138#_c_130_n N_VPWR_M1000_d 0.00158317f $X=0.81 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_28_138#_M1003_g N_VPWR_c_487_n 0.00337637f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_143 N_A_28_138#_c_141_n N_VPWR_c_487_n 0.0213377f $X=0.725 $Y=2.037 $X2=0
+ $Y2=0
cc_144 N_A_28_138#_M1003_g N_VPWR_c_491_n 0.00518311f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_145 N_A_28_138#_M1003_g N_VPWR_c_486_n 0.00991001f $X=1.005 $Y=2.4 $X2=0
+ $Y2=0
cc_146 N_A_28_138#_c_128_n N_VGND_M1006_d 0.00119058f $X=0.725 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_28_138#_c_129_n N_VGND_M1006_d 0.00179209f $X=0.81 $Y=1.605 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_28_138#_M1002_g N_VGND_c_568_n 0.0132572f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_28_138#_c_128_n N_VGND_c_568_n 0.00915704f $X=0.725 $Y=1.06 $X2=0
+ $Y2=0
cc_150 N_A_28_138#_c_129_n N_VGND_c_568_n 0.0110081f $X=0.81 $Y=1.605 $X2=0
+ $Y2=0
cc_151 N_A_28_138#_c_132_n N_VGND_c_568_n 3.45021e-19 $X=0.955 $Y=1.44 $X2=0
+ $Y2=0
cc_152 N_A_28_138#_c_131_n N_VGND_c_571_n 0.00444585f $X=0.265 $Y=0.865 $X2=0
+ $Y2=0
cc_153 N_A_28_138#_M1002_g N_VGND_c_572_n 0.00383152f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_28_138#_M1002_g N_VGND_c_575_n 0.00762539f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_155 N_A_28_138#_c_131_n N_VGND_c_575_n 0.00830526f $X=0.265 $Y=0.865 $X2=0
+ $Y2=0
cc_156 N_A_209_74#_M1007_g N_A_316_138#_M1008_g 0.0165204f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_157 N_A_209_74#_M1004_g N_A_316_138#_M1009_g 0.0229978f $X=1.975 $Y=2.05
+ $X2=0 $Y2=0
cc_158 N_A_209_74#_M1007_g N_A_316_138#_c_264_n 0.0140061f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_159 N_A_209_74#_c_196_n N_A_316_138#_c_264_n 0.0113458f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_160 N_A_209_74#_c_197_n N_A_316_138#_c_264_n 0.00326921f $X=1.83 $Y=1.44
+ $X2=0 $Y2=0
cc_161 N_A_209_74#_M1004_g N_A_316_138#_c_278_n 0.0145588f $X=1.975 $Y=2.05
+ $X2=0 $Y2=0
cc_162 N_A_209_74#_M1007_g N_A_316_138#_c_265_n 0.00276635f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_163 N_A_209_74#_c_196_n N_A_316_138#_c_265_n 0.0244444f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_164 N_A_209_74#_c_197_n N_A_316_138#_c_265_n 0.00302017f $X=1.83 $Y=1.44
+ $X2=0 $Y2=0
cc_165 N_A_209_74#_M1004_g N_A_316_138#_c_266_n 0.00674167f $X=1.975 $Y=2.05
+ $X2=0 $Y2=0
cc_166 N_A_209_74#_M1007_g N_A_316_138#_c_267_n 0.00158921f $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_167 N_A_209_74#_c_194_n N_A_316_138#_c_267_n 0.0359881f $X=1.185 $Y=0.57
+ $X2=0 $Y2=0
cc_168 N_A_209_74#_c_196_n N_A_316_138#_c_267_n 0.0233038f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_169 N_A_209_74#_c_197_n N_A_316_138#_c_267_n 0.00407385f $X=1.83 $Y=1.44
+ $X2=0 $Y2=0
cc_170 N_A_209_74#_c_196_n N_A_316_138#_c_271_n 0.0213641f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_171 N_A_209_74#_c_197_n N_A_316_138#_c_271_n 0.00459063f $X=1.83 $Y=1.44
+ $X2=0 $Y2=0
cc_172 N_A_209_74#_c_202_n N_A_316_138#_c_271_n 0.026595f $X=1.222 $Y=1.992
+ $X2=0 $Y2=0
cc_173 N_A_209_74#_c_204_n N_A_316_138#_c_271_n 0.00174864f $X=1.23 $Y=2 $X2=0
+ $Y2=0
cc_174 N_A_209_74#_M1007_g N_A_316_138#_c_268_n 5.933e-19 $X=1.92 $Y=0.9 $X2=0
+ $Y2=0
cc_175 N_A_209_74#_c_196_n N_A_316_138#_c_268_n 2.57095e-19 $X=1.83 $Y=1.44
+ $X2=0 $Y2=0
cc_176 N_A_209_74#_c_197_n N_A_316_138#_c_268_n 0.0207317f $X=1.83 $Y=1.44 $X2=0
+ $Y2=0
cc_177 N_A_209_74#_M1004_g N_X_c_344_n 0.00115812f $X=1.975 $Y=2.05 $X2=0 $Y2=0
cc_178 N_A_209_74#_M1004_g N_X_c_346_n 3.6476e-19 $X=1.975 $Y=2.05 $X2=0 $Y2=0
cc_179 N_A_209_74#_M1004_g N_X_c_352_n 9.11177e-19 $X=1.975 $Y=2.05 $X2=0 $Y2=0
cc_180 N_A_209_74#_M1004_g N_X_c_348_n 0.00541916f $X=1.975 $Y=2.05 $X2=0 $Y2=0
cc_181 N_A_209_74#_c_204_n N_X_c_348_n 0.0681118f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_182 N_A_209_74#_c_204_n N_VPWR_c_487_n 0.0308555f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_183 N_A_209_74#_M1004_g N_VPWR_c_488_n 0.00189879f $X=1.975 $Y=2.05 $X2=0
+ $Y2=0
cc_184 N_A_209_74#_c_204_n N_VPWR_c_491_n 0.022336f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_185 N_A_209_74#_c_204_n N_VPWR_c_486_n 0.012036f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_186 N_A_209_74#_c_194_n N_VGND_c_568_n 0.0252885f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_187 N_A_209_74#_M1007_g N_VGND_c_569_n 0.00261888f $X=1.92 $Y=0.9 $X2=0 $Y2=0
cc_188 N_A_209_74#_c_194_n N_VGND_c_569_n 0.0141693f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_189 N_A_209_74#_M1007_g N_VGND_c_572_n 0.00382655f $X=1.92 $Y=0.9 $X2=0 $Y2=0
cc_190 N_A_209_74#_c_194_n N_VGND_c_572_n 0.0206458f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_191 N_A_209_74#_M1007_g N_VGND_c_575_n 0.00451834f $X=1.92 $Y=0.9 $X2=0 $Y2=0
cc_192 N_A_209_74#_c_194_n N_VGND_c_575_n 0.0111968f $X=1.185 $Y=0.57 $X2=0
+ $Y2=0
cc_193 N_A_316_138#_M1008_g N_X_c_336_n 0.00270228f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_316_138#_M1009_g N_X_c_344_n 0.0146378f $X=2.49 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_316_138#_M1008_g N_X_c_337_n 0.00322309f $X=2.41 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_316_138#_c_265_n N_X_c_337_n 0.0113527f $X=2.25 $Y=1.605 $X2=0 $Y2=0
cc_197 N_A_316_138#_c_268_n N_X_c_337_n 6.2756e-19 $X=2.44 $Y=1.44 $X2=0 $Y2=0
cc_198 N_A_316_138#_c_268_n N_X_c_339_n 0.00316923f $X=2.44 $Y=1.44 $X2=0 $Y2=0
cc_199 N_A_316_138#_c_265_n N_X_c_340_n 0.0247198f $X=2.25 $Y=1.605 $X2=0 $Y2=0
cc_200 N_A_316_138#_c_268_n N_X_c_340_n 0.00326086f $X=2.44 $Y=1.44 $X2=0 $Y2=0
cc_201 N_A_316_138#_M1009_g X 0.00753496f $X=2.49 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_316_138#_c_265_n N_X_c_341_n 2.02801e-19 $X=2.25 $Y=1.605 $X2=0 $Y2=0
cc_203 N_A_316_138#_c_268_n N_X_c_341_n 0.00588998f $X=2.44 $Y=1.44 $X2=0 $Y2=0
cc_204 N_A_316_138#_M1009_g N_X_c_346_n 0.00827378f $X=2.49 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_316_138#_c_278_n N_X_c_346_n 0.0170367f $X=2.165 $Y=2.017 $X2=0 $Y2=0
cc_206 N_A_316_138#_c_265_n N_X_c_346_n 0.00100347f $X=2.25 $Y=1.605 $X2=0 $Y2=0
cc_207 N_A_316_138#_c_266_n N_X_c_346_n 0.0044306f $X=2.25 $Y=1.895 $X2=0 $Y2=0
cc_208 N_A_316_138#_c_268_n N_X_c_346_n 0.00104646f $X=2.44 $Y=1.44 $X2=0 $Y2=0
cc_209 N_A_316_138#_M1009_g N_X_c_342_n 0.00537231f $X=2.49 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_316_138#_c_266_n N_X_c_342_n 0.0102016f $X=2.25 $Y=1.895 $X2=0 $Y2=0
cc_211 N_A_316_138#_M1009_g N_X_c_352_n 0.00553121f $X=2.49 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_316_138#_c_278_n N_X_c_352_n 0.0067603f $X=2.165 $Y=2.017 $X2=0 $Y2=0
cc_213 N_A_316_138#_c_265_n N_X_c_352_n 0.00419195f $X=2.25 $Y=1.605 $X2=0 $Y2=0
cc_214 N_A_316_138#_c_271_n N_X_c_352_n 0.00259488f $X=1.87 $Y=2.06 $X2=0 $Y2=0
cc_215 N_A_316_138#_c_278_n N_X_c_348_n 0.0114592f $X=2.165 $Y=2.017 $X2=0 $Y2=0
cc_216 N_A_316_138#_c_271_n N_X_c_348_n 0.0170914f $X=1.87 $Y=2.06 $X2=0 $Y2=0
cc_217 N_A_316_138#_M1009_g N_A_604_138#_c_431_n 7.05863e-19 $X=2.49 $Y=2.4
+ $X2=0 $Y2=0
cc_218 N_A_316_138#_c_278_n N_VPWR_M1004_d 0.00674386f $X=2.165 $Y=2.017 $X2=0
+ $Y2=0
cc_219 N_A_316_138#_c_266_n N_VPWR_M1004_d 0.00128457f $X=2.25 $Y=1.895 $X2=0
+ $Y2=0
cc_220 N_A_316_138#_M1009_g N_VPWR_c_488_n 0.00371117f $X=2.49 $Y=2.4 $X2=0
+ $Y2=0
cc_221 N_A_316_138#_c_278_n N_VPWR_c_488_n 0.0181196f $X=2.165 $Y=2.017 $X2=0
+ $Y2=0
cc_222 N_A_316_138#_M1009_g N_VPWR_c_492_n 0.00536645f $X=2.49 $Y=2.4 $X2=0
+ $Y2=0
cc_223 N_A_316_138#_M1009_g N_VPWR_c_486_n 0.0104603f $X=2.49 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A_316_138#_c_264_n N_VGND_M1007_d 0.00119058f $X=2.165 $Y=1.06 $X2=0
+ $Y2=0
cc_225 N_A_316_138#_c_265_n N_VGND_M1007_d 0.00179209f $X=2.25 $Y=1.605 $X2=0
+ $Y2=0
cc_226 N_A_316_138#_M1008_g N_VGND_c_569_n 0.0132572f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_227 N_A_316_138#_c_264_n N_VGND_c_569_n 0.00915704f $X=2.165 $Y=1.06 $X2=0
+ $Y2=0
cc_228 N_A_316_138#_c_265_n N_VGND_c_569_n 0.0110081f $X=2.25 $Y=1.605 $X2=0
+ $Y2=0
cc_229 N_A_316_138#_c_267_n N_VGND_c_572_n 0.00427375f $X=1.705 $Y=0.865 $X2=0
+ $Y2=0
cc_230 N_A_316_138#_M1008_g N_VGND_c_573_n 0.00383152f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_316_138#_M1008_g N_VGND_c_575_n 0.00762539f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_316_138#_c_267_n N_VGND_c_575_n 0.00802181f $X=1.705 $Y=0.865 $X2=0
+ $Y2=0
cc_233 N_X_M1001_g N_A_604_138#_M1005_g 0.0165204f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_234 N_X_M1010_g N_A_604_138#_M1011_g 0.0240139f $X=3.46 $Y=2.05 $X2=0 $Y2=0
cc_235 X N_A_604_138#_M1011_g 0.00791354f $X=0.965 $Y=2.32 $X2=0 $Y2=0
cc_236 N_X_c_336_n N_A_604_138#_c_436_n 0.0196927f $X=2.625 $Y=0.57 $X2=0 $Y2=0
cc_237 N_X_M1001_g N_A_604_138#_c_424_n 0.0144149f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_238 N_X_c_338_n N_A_604_138#_c_424_n 0.0113081f $X=3.27 $Y=1.44 $X2=0 $Y2=0
cc_239 N_X_c_341_n N_A_604_138#_c_424_n 0.00521738f $X=3.46 $Y=1.44 $X2=0 $Y2=0
cc_240 N_X_c_338_n N_A_604_138#_c_425_n 0.0175411f $X=3.27 $Y=1.44 $X2=0 $Y2=0
cc_241 N_X_c_339_n N_A_604_138#_c_425_n 0.013174f $X=2.697 $Y=1.075 $X2=0 $Y2=0
cc_242 N_X_c_341_n N_A_604_138#_c_425_n 0.0040983f $X=3.46 $Y=1.44 $X2=0 $Y2=0
cc_243 N_X_M1001_g N_A_604_138#_c_426_n 0.00277296f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_244 N_X_c_338_n N_A_604_138#_c_426_n 0.0246623f $X=3.27 $Y=1.44 $X2=0 $Y2=0
cc_245 N_X_c_341_n N_A_604_138#_c_426_n 0.00335815f $X=3.46 $Y=1.44 $X2=0 $Y2=0
cc_246 N_X_M1010_g N_A_604_138#_c_427_n 0.00625602f $X=3.46 $Y=2.05 $X2=0 $Y2=0
cc_247 N_X_M1010_g N_A_604_138#_c_431_n 0.0174581f $X=3.46 $Y=2.05 $X2=0 $Y2=0
cc_248 N_X_c_338_n N_A_604_138#_c_431_n 0.017135f $X=3.27 $Y=1.44 $X2=0 $Y2=0
cc_249 X N_A_604_138#_c_431_n 0.0269049f $X=0.965 $Y=2.32 $X2=0 $Y2=0
cc_250 N_X_c_341_n N_A_604_138#_c_431_n 0.00570109f $X=3.46 $Y=1.44 $X2=0 $Y2=0
cc_251 N_X_c_346_n N_A_604_138#_c_431_n 0.0228844f $X=2.715 $Y=2 $X2=0 $Y2=0
cc_252 N_X_c_352_n N_A_604_138#_c_431_n 0.00206411f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_253 N_X_M1001_g N_A_604_138#_c_428_n 4.84716e-19 $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_254 N_X_c_338_n N_A_604_138#_c_428_n 2.23289e-19 $X=3.27 $Y=1.44 $X2=0 $Y2=0
cc_255 N_X_c_341_n N_A_604_138#_c_428_n 0.0208182f $X=3.46 $Y=1.44 $X2=0 $Y2=0
cc_256 X N_VPWR_M1010_d 3.78439e-19 $X=0.965 $Y=2.32 $X2=0 $Y2=0
cc_257 N_X_c_348_n N_VPWR_c_487_n 0.00566053f $X=2.405 $Y=2.405 $X2=0 $Y2=0
cc_258 N_X_c_344_n N_VPWR_c_488_n 0.0352186f $X=2.715 $Y=2.815 $X2=0 $Y2=0
cc_259 N_X_c_352_n N_VPWR_c_488_n 2.96851e-19 $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_260 N_X_c_348_n N_VPWR_c_488_n 0.0341338f $X=2.405 $Y=2.405 $X2=0 $Y2=0
cc_261 N_X_M1010_g N_VPWR_c_489_n 0.00190355f $X=3.46 $Y=2.05 $X2=0 $Y2=0
cc_262 X N_VPWR_c_489_n 0.0333454f $X=0.965 $Y=2.32 $X2=0 $Y2=0
cc_263 N_X_c_344_n N_VPWR_c_492_n 0.0213134f $X=2.715 $Y=2.815 $X2=0 $Y2=0
cc_264 N_X_c_344_n N_VPWR_c_486_n 0.0115215f $X=2.715 $Y=2.815 $X2=0 $Y2=0
cc_265 N_X_M1010_g N_A_785_74#_c_538_n 6.21207e-19 $X=3.46 $Y=2.05 $X2=0 $Y2=0
cc_266 X N_A_785_74#_c_538_n 0.0239695f $X=0.965 $Y=2.32 $X2=0 $Y2=0
cc_267 N_X_M1010_g N_A_785_74#_c_539_n 3.47282e-19 $X=3.46 $Y=2.05 $X2=0 $Y2=0
cc_268 X N_A_785_74#_c_539_n 0.0333096f $X=0.965 $Y=2.32 $X2=0 $Y2=0
cc_269 N_X_c_336_n N_VGND_c_569_n 0.0253911f $X=2.625 $Y=0.57 $X2=0 $Y2=0
cc_270 N_X_M1001_g N_VGND_c_570_n 0.00254928f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_271 N_X_c_336_n N_VGND_c_570_n 0.0151085f $X=2.625 $Y=0.57 $X2=0 $Y2=0
cc_272 N_X_M1001_g N_VGND_c_573_n 0.00382655f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_273 N_X_c_336_n N_VGND_c_573_n 0.0238717f $X=2.625 $Y=0.57 $X2=0 $Y2=0
cc_274 N_X_M1001_g N_VGND_c_575_n 0.00451834f $X=3.36 $Y=0.9 $X2=0 $Y2=0
cc_275 N_X_c_336_n N_VGND_c_575_n 0.0129463f $X=2.625 $Y=0.57 $X2=0 $Y2=0
cc_276 N_A_604_138#_c_427_n N_VPWR_M1010_d 6.4105e-19 $X=3.705 $Y=1.895 $X2=0
+ $Y2=0
cc_277 N_A_604_138#_c_431_n N_VPWR_M1010_d 0.00474659f $X=3.235 $Y=2.06 $X2=0
+ $Y2=0
cc_278 N_A_604_138#_M1011_g N_VPWR_c_489_n 0.00368581f $X=3.98 $Y=2.4 $X2=0
+ $Y2=0
cc_279 N_A_604_138#_c_431_n N_VPWR_c_489_n 0.0172041f $X=3.235 $Y=2.06 $X2=0
+ $Y2=0
cc_280 N_A_604_138#_M1011_g N_VPWR_c_493_n 0.00530534f $X=3.98 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_A_604_138#_M1011_g N_VPWR_c_486_n 0.0102761f $X=3.98 $Y=2.4 $X2=0 $Y2=0
cc_282 N_A_604_138#_M1005_g N_A_785_74#_c_535_n 0.00271338f $X=3.85 $Y=0.74
+ $X2=0 $Y2=0
cc_283 N_A_604_138#_M1011_g N_A_785_74#_c_538_n 0.0147098f $X=3.98 $Y=2.4 $X2=0
+ $Y2=0
cc_284 N_A_604_138#_c_431_n N_A_785_74#_c_538_n 0.00157372f $X=3.235 $Y=2.06
+ $X2=0 $Y2=0
cc_285 N_A_604_138#_c_426_n N_A_785_74#_c_536_n 0.00241382f $X=3.705 $Y=1.605
+ $X2=0 $Y2=0
cc_286 N_A_604_138#_c_428_n N_A_785_74#_c_536_n 0.00475928f $X=3.925 $Y=1.44
+ $X2=0 $Y2=0
cc_287 N_A_604_138#_M1011_g N_A_785_74#_c_539_n 0.0111009f $X=3.98 $Y=2.4 $X2=0
+ $Y2=0
cc_288 N_A_604_138#_c_426_n N_A_785_74#_c_539_n 0.00695851f $X=3.705 $Y=1.605
+ $X2=0 $Y2=0
cc_289 N_A_604_138#_c_427_n N_A_785_74#_c_539_n 0.00449799f $X=3.705 $Y=1.895
+ $X2=0 $Y2=0
cc_290 N_A_604_138#_c_431_n N_A_785_74#_c_539_n 0.0255731f $X=3.235 $Y=2.06
+ $X2=0 $Y2=0
cc_291 N_A_604_138#_c_428_n N_A_785_74#_c_539_n 8.37166e-19 $X=3.925 $Y=1.44
+ $X2=0 $Y2=0
cc_292 N_A_604_138#_M1005_g N_A_785_74#_c_537_n 0.00261251f $X=3.85 $Y=0.74
+ $X2=0 $Y2=0
cc_293 N_A_604_138#_M1011_g N_A_785_74#_c_537_n 0.00426536f $X=3.98 $Y=2.4 $X2=0
+ $Y2=0
cc_294 N_A_604_138#_c_426_n N_A_785_74#_c_537_n 0.0310126f $X=3.705 $Y=1.605
+ $X2=0 $Y2=0
cc_295 N_A_604_138#_c_427_n N_A_785_74#_c_537_n 0.00788655f $X=3.705 $Y=1.895
+ $X2=0 $Y2=0
cc_296 N_A_604_138#_c_428_n N_A_785_74#_c_537_n 0.00854303f $X=3.925 $Y=1.44
+ $X2=0 $Y2=0
cc_297 N_A_604_138#_c_424_n N_VGND_M1001_d 0.00119058f $X=3.605 $Y=1.06 $X2=0
+ $Y2=0
cc_298 N_A_604_138#_c_426_n N_VGND_M1001_d 0.00179209f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_299 N_A_604_138#_M1005_g N_VGND_c_570_n 0.0132572f $X=3.85 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_604_138#_c_424_n N_VGND_c_570_n 0.00915704f $X=3.605 $Y=1.06 $X2=0
+ $Y2=0
cc_301 N_A_604_138#_c_426_n N_VGND_c_570_n 0.0110542f $X=3.705 $Y=1.605 $X2=0
+ $Y2=0
cc_302 N_A_604_138#_c_436_n N_VGND_c_573_n 0.00310575f $X=3.145 $Y=0.865 $X2=0
+ $Y2=0
cc_303 N_A_604_138#_M1005_g N_VGND_c_574_n 0.00383152f $X=3.85 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_604_138#_M1005_g N_VGND_c_575_n 0.00762539f $X=3.85 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_604_138#_c_436_n N_VGND_c_575_n 0.00603761f $X=3.145 $Y=0.865 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_489_n N_A_785_74#_c_538_n 0.035258f $X=3.75 $Y=2.475 $X2=0 $Y2=0
cc_307 N_VPWR_c_493_n N_A_785_74#_c_538_n 0.0212959f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_486_n N_A_785_74#_c_538_n 0.0114986f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_M1010_d N_A_785_74#_c_539_n 0.00279104f $X=3.55 $Y=1.84 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_489_n N_A_785_74#_c_539_n 0.0011495f $X=3.75 $Y=2.475 $X2=0
+ $Y2=0
cc_311 N_A_785_74#_c_535_n N_VGND_c_570_n 0.0254826f $X=4.065 $Y=0.57 $X2=0
+ $Y2=0
cc_312 N_A_785_74#_c_535_n N_VGND_c_574_n 0.0270976f $X=4.065 $Y=0.57 $X2=0
+ $Y2=0
cc_313 N_A_785_74#_c_535_n N_VGND_c_575_n 0.0146958f $X=4.065 $Y=0.57 $X2=0
+ $Y2=0

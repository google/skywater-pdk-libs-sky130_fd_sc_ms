# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__a2bb2oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.471000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.470000 2.275000 1.800000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.471000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.420000 0.455000 1.770000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735000 1.350000 8.515000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.115000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.433600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.270000 0.350000 2.520000 0.790000 ;
        RECT 2.270000 0.790000 6.150000 0.960000 ;
        RECT 3.185000 1.720000 4.255000 1.890000 ;
        RECT 3.185000 1.890000 3.355000 2.735000 ;
        RECT 3.210000 0.350000 3.380000 0.790000 ;
        RECT 3.965000 0.960000 6.150000 1.130000 ;
        RECT 3.965000 1.130000 4.255000 1.720000 ;
        RECT 4.085000 1.890000 4.255000 2.735000 ;
        RECT 4.960000 0.770000 6.150000 0.790000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.105000  1.940000 0.435000 2.905000 ;
      RECT 0.105000  2.905000 1.255000 3.075000 ;
      RECT 0.635000  1.130000 3.585000 1.300000 ;
      RECT 0.635000  1.300000 0.885000 2.735000 ;
      RECT 0.940000  0.085000 1.270000 0.960000 ;
      RECT 1.085000  1.940000 1.255000 1.970000 ;
      RECT 1.085000  1.970000 2.235000 2.140000 ;
      RECT 1.085000  2.140000 1.255000 2.905000 ;
      RECT 1.450000  0.350000 1.620000 1.130000 ;
      RECT 1.455000  2.310000 1.705000 3.245000 ;
      RECT 1.800000  0.085000 2.090000 0.885000 ;
      RECT 1.905000  2.140000 2.235000 2.980000 ;
      RECT 2.575000  1.300000 3.585000 1.550000 ;
      RECT 2.655000  1.820000 2.985000 2.905000 ;
      RECT 2.655000  2.905000 4.785000 3.075000 ;
      RECT 2.700000  0.085000 3.030000 0.620000 ;
      RECT 3.555000  2.060000 3.885000 2.905000 ;
      RECT 3.560000  0.085000 3.890000 0.620000 ;
      RECT 4.455000  1.950000 8.385000 2.120000 ;
      RECT 4.455000  2.120000 4.785000 2.905000 ;
      RECT 4.530000  0.350000 6.500000 0.600000 ;
      RECT 4.985000  2.290000 5.155000 3.245000 ;
      RECT 5.355000  2.120000 5.685000 2.980000 ;
      RECT 5.885000  2.290000 6.135000 3.245000 ;
      RECT 6.330000  0.600000 6.500000 1.010000 ;
      RECT 6.330000  1.010000 8.300000 1.180000 ;
      RECT 6.335000  1.820000 6.505000 1.950000 ;
      RECT 6.335000  2.120000 6.505000 2.980000 ;
      RECT 6.680000  0.085000 6.930000 0.840000 ;
      RECT 6.705000  2.290000 6.955000 3.245000 ;
      RECT 7.110000  0.350000 7.360000 1.010000 ;
      RECT 7.155000  2.120000 7.485000 2.980000 ;
      RECT 7.540000  0.085000 7.790000 0.840000 ;
      RECT 7.685000  2.290000 7.855000 3.245000 ;
      RECT 7.970000  0.350000 8.300000 1.010000 ;
      RECT 8.055000  2.120000 8.385000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ms__a2bb2oi_4
END LIBRARY

* File: sky130_fd_sc_ms__dlrtn_4.spice
* Created: Wed Sep  2 12:05:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrtn_4.pex.spice"
.subckt sky130_fd_sc_ms__dlrtn_4  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_D_M1024_g N_A_27_136#_M1024_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1003 N_A_232_98#_M1003_d N_GATE_N_M1003_g N_VGND_M1024_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2886 AS=0.230174 PD=2.26 PS=1.70946 NRD=8.1 NRS=41.52 M=1
+ R=4.93333 SA=75000.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_232_98#_M1020_g N_A_348_392#_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.421076 AS=0.2109 PD=2.11812 PS=2.05 NRD=83.352 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 A_666_74# N_A_27_136#_M1018_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.364174 PD=0.88 PS=1.83188 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75001.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_642_392#_M1017_d N_A_232_98#_M1017_g A_666_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.0768 PD=1.16528 PS=0.88 NRD=8.436 NRS=12.18 M=1
+ R=4.26667 SA=75001.6 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1006 A_839_74# N_A_348_392#_M1006_g N_A_642_392#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.05775 AS=0.0758774 PD=0.695 PS=0.764717 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_888_406#_M1015_g A_839_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.05775 PD=1.41 PS=0.695 NRD=0 NRS=23.568 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_1035_74#_M1009_d N_A_642_392#_M1009_g N_A_888_406#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1026 N_A_1035_74#_M1026_d N_A_642_392#_M1026_g N_A_888_406#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_A_1035_74#_M1026_d N_RESET_B_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_1035_74#_M1021_d N_RESET_B_M1021_g N_VGND_M1002_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A_888_406#_M1001_g N_Q_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_888_406#_M1004_g N_Q_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1004_d N_A_888_406#_M1011_g N_Q_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_888_406#_M1022_g N_Q_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_D_M1013_g N_A_27_136#_M1013_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1007 N_A_232_98#_M1007_d N_GATE_N_M1007_g N_VPWR_M1013_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1554 PD=2.24 PS=1.21 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1008_d N_A_232_98#_M1008_g N_A_348_392#_M1008_s VPB PSHORT L=0.18
+ W=0.84 AD=0.223193 AS=0.2352 PD=1.50652 PS=2.24 NRD=49.4076 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90003.2 A=0.1512 P=2.04 MULT=1
MM1005 A_564_392# N_A_27_136#_M1005_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1
+ AD=0.105 AS=0.265707 PD=1.21 PS=1.79348 NRD=9.8303 NRS=16.7253 M=1 R=5.55556
+ SA=90000.7 SB=90003 A=0.18 P=2.36 MULT=1
MM1028 N_A_642_392#_M1028_d N_A_348_392#_M1028_g A_564_392# VPB PSHORT L=0.18
+ W=1 AD=0.222394 AS=0.105 PD=1.91549 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556
+ SA=90001.1 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1000 A_750_504# N_A_232_98#_M1000_g N_A_642_392#_M1028_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1449 AS=0.0934056 PD=1.11 PS=0.804507 NRD=136.009 NRS=78.5045 M=1
+ R=2.33333 SA=90001.6 SB=90005.5 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_888_406#_M1010_g A_750_504# VPB PSHORT L=0.18 W=0.42
+ AD=0.1358 AS=0.1449 PD=1.04 PS=1.11 NRD=0 NRS=136.009 M=1 R=2.33333 SA=90002.4
+ SB=90004.6 A=0.0756 P=1.2 MULT=1
MM1012 N_A_888_406#_M1012_d N_A_642_392#_M1012_g N_VPWR_M1010_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.2716 PD=1.11 PS=2.08 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90001.7 SB=90003.7 A=0.1512 P=2.04 MULT=1
MM1016 N_A_888_406#_M1012_d N_A_642_392#_M1016_g N_VPWR_M1016_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.1344 PD=1.11 PS=1.16 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90002.2 SB=90003.3 A=0.1512 P=2.04 MULT=1
MM1014 N_A_888_406#_M1014_d N_RESET_B_M1014_g N_VPWR_M1016_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1428 AS=0.1344 PD=1.18 PS=1.16 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90002.7 SB=90002.8 A=0.1512 P=2.04 MULT=1
MM1029 N_A_888_406#_M1014_d N_RESET_B_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1428 AS=0.176486 PD=1.18 PS=1.30714 NRD=3.5066 NRS=18.7544 M=1
+ R=4.66667 SA=90003.2 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1019 N_VPWR_M1029_s N_A_888_406#_M1019_g N_Q_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.235314 AS=0.1512 PD=1.74286 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90002.9 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1023 N_VPWR_M1023_d N_A_888_406#_M1023_g N_Q_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1025 N_VPWR_M1023_d N_A_888_406#_M1025_g N_Q_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2072 PD=1.44 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.8
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1027 N_VPWR_M1027_d N_A_888_406#_M1027_g N_Q_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2072 PD=2.8 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX30_noxref VNB VPB NWDIODE A=18.5628 P=23.68
*
.include "sky130_fd_sc_ms__dlrtn_4.pxi.spice"
*
.ends
*
*

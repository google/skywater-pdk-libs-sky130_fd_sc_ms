* File: sky130_fd_sc_ms__nor3b_4.pxi.spice
* Created: Wed Sep  2 12:16:30 2020
* 
x_PM_SKY130_FD_SC_MS__NOR3B_4%B N_B_M1010_g N_B_M1001_g N_B_M1006_g N_B_M1015_g
+ N_B_M1007_g N_B_M1025_g N_B_M1011_g N_B_M1026_g B B B B N_B_c_123_n
+ PM_SKY130_FD_SC_MS__NOR3B_4%B
x_PM_SKY130_FD_SC_MS__NOR3B_4%A_468_264# N_A_468_264#_M1014_d
+ N_A_468_264#_M1022_d N_A_468_264#_M1002_g N_A_468_264#_M1000_g
+ N_A_468_264#_M1005_g N_A_468_264#_M1004_g N_A_468_264#_M1009_g
+ N_A_468_264#_M1016_g N_A_468_264#_M1012_g N_A_468_264#_M1019_g
+ N_A_468_264#_c_209_n N_A_468_264#_c_219_n N_A_468_264#_c_220_n
+ N_A_468_264#_c_221_n N_A_468_264#_c_210_n N_A_468_264#_c_211_n
+ N_A_468_264#_c_243_p N_A_468_264#_c_212_n N_A_468_264#_c_213_n
+ PM_SKY130_FD_SC_MS__NOR3B_4%A_468_264#
x_PM_SKY130_FD_SC_MS__NOR3B_4%A N_A_c_352_n N_A_M1008_g N_A_M1003_g N_A_c_354_n
+ N_A_M1018_g N_A_M1013_g N_A_c_356_n N_A_M1021_g N_A_M1017_g N_A_c_358_n
+ N_A_M1024_g N_A_M1020_g A N_A_c_361_n N_A_c_362_n
+ PM_SKY130_FD_SC_MS__NOR3B_4%A
x_PM_SKY130_FD_SC_MS__NOR3B_4%C_N N_C_N_c_444_n N_C_N_M1014_g N_C_N_c_447_n
+ N_C_N_M1022_g N_C_N_c_448_n N_C_N_M1023_g C_N N_C_N_c_446_n
+ PM_SKY130_FD_SC_MS__NOR3B_4%C_N
x_PM_SKY130_FD_SC_MS__NOR3B_4%A_27_368# N_A_27_368#_M1001_d N_A_27_368#_M1006_d
+ N_A_27_368#_M1011_d N_A_27_368#_M1005_s N_A_27_368#_M1012_s
+ N_A_27_368#_c_482_n N_A_27_368#_c_483_n N_A_27_368#_c_484_n
+ N_A_27_368#_c_512_p N_A_27_368#_c_485_n N_A_27_368#_c_497_n
+ N_A_27_368#_c_486_n N_A_27_368#_c_487_n N_A_27_368#_c_501_n
+ N_A_27_368#_c_503_n N_A_27_368#_c_488_n PM_SKY130_FD_SC_MS__NOR3B_4%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR3B_4%A_129_368# N_A_129_368#_M1001_s
+ N_A_129_368#_M1007_s N_A_129_368#_M1003_d N_A_129_368#_M1017_d
+ N_A_129_368#_c_548_n N_A_129_368#_c_545_n N_A_129_368#_c_546_n
+ N_A_129_368#_c_570_n N_A_129_368#_c_571_n N_A_129_368#_c_547_n
+ N_A_129_368#_c_553_n N_A_129_368#_c_558_n N_A_129_368#_c_572_n
+ PM_SKY130_FD_SC_MS__NOR3B_4%A_129_368#
x_PM_SKY130_FD_SC_MS__NOR3B_4%Y N_Y_M1010_s N_Y_M1025_s N_Y_M1000_s N_Y_M1016_s
+ N_Y_M1008_d N_Y_M1021_d N_Y_M1002_d N_Y_M1009_d N_Y_c_611_n N_Y_c_612_n
+ N_Y_c_613_n N_Y_c_614_n N_Y_c_637_n N_Y_c_625_n N_Y_c_615_n N_Y_c_616_n
+ N_Y_c_617_n N_Y_c_671_n N_Y_c_618_n N_Y_c_692_n N_Y_c_619_n N_Y_c_620_n
+ N_Y_c_621_n N_Y_c_622_n N_Y_c_623_n N_Y_c_700_n Y
+ PM_SKY130_FD_SC_MS__NOR3B_4%Y
x_PM_SKY130_FD_SC_MS__NOR3B_4%VPWR N_VPWR_M1003_s N_VPWR_M1013_s N_VPWR_M1020_s
+ N_VPWR_M1023_s N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n
+ N_VPWR_c_753_n VPWR N_VPWR_c_754_n N_VPWR_c_755_n N_VPWR_c_756_n
+ N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n N_VPWR_c_760_n N_VPWR_c_748_n
+ PM_SKY130_FD_SC_MS__NOR3B_4%VPWR
x_PM_SKY130_FD_SC_MS__NOR3B_4%VGND N_VGND_M1010_d N_VGND_M1015_d N_VGND_M1026_d
+ N_VGND_M1004_d N_VGND_M1019_d N_VGND_M1018_s N_VGND_M1024_s N_VGND_c_842_n
+ N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n
+ N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n
+ N_VGND_c_853_n VGND N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ N_VGND_c_862_n N_VGND_c_863_n PM_SKY130_FD_SC_MS__NOR3B_4%VGND
cc_1 VNB N_B_M1010_g 0.030989f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_2 VNB N_B_M1015_g 0.0252957f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_B_M1025_g 0.0248983f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_4 VNB N_B_M1026_g 0.023399f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_5 VNB B 0.018482f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_B_c_123_n 0.0772718f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.515
cc_7 VNB N_A_468_264#_M1002_g 4.92448e-19 $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.68
cc_8 VNB N_A_468_264#_M1000_g 0.0222712f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.35
cc_9 VNB N_A_468_264#_M1005_g 4.78582e-19 $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.68
cc_10 VNB N_A_468_264#_M1004_g 0.0220929f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.35
cc_11 VNB N_A_468_264#_M1009_g 4.78476e-19 $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.68
cc_12 VNB N_A_468_264#_M1016_g 0.0226931f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.35
cc_13 VNB N_A_468_264#_M1012_g 5.19442e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_A_468_264#_M1019_g 0.0241345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_468_264#_c_209_n 0.00717215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_468_264#_c_210_n 0.0289376f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_17 VNB N_A_468_264#_c_211_n 0.031855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_468_264#_c_212_n 0.00697138f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.565
cc_19 VNB N_A_468_264#_c_213_n 0.0892919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_352_n 0.0185806f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_21 VNB N_A_M1003_g 0.00708742f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_22 VNB N_A_c_354_n 0.0191883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_M1013_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.35
cc_24 VNB N_A_c_356_n 0.0198403f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_25 VNB N_A_M1017_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_c_358_n 0.0179355f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_27 VNB N_A_M1020_g 0.00652527f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=2.4
cc_28 VNB A 0.00598605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_c_361_n 0.112873f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_30 VNB N_A_c_362_n 0.00358389f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.515
cc_31 VNB N_C_N_c_444_n 0.0236108f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_32 VNB C_N 0.00374395f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_33 VNB N_C_N_c_446_n 0.0736887f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_34 VNB N_Y_c_611_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=2.4
cc_35 VNB N_Y_c_612_n 0.00273768f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_36 VNB N_Y_c_613_n 0.00239855f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_Y_c_614_n 0.00224624f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_38 VNB N_Y_c_615_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_39 VNB N_Y_c_616_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_40 VNB N_Y_c_617_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.515
cc_41 VNB N_Y_c_618_n 0.00240319f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_42 VNB N_Y_c_619_n 0.0028001f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_43 VNB N_Y_c_620_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_44 VNB N_Y_c_621_n 0.00554939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_622_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_623_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB Y 0.00464838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_748_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_842_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_50 VNB N_VGND_c_843_n 0.0454867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_844_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_845_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_53 VNB N_VGND_c_846_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_54 VNB N_VGND_c_847_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_848_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_849_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_57 VNB N_VGND_c_850_n 0.00967485f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.515
cc_58 VNB N_VGND_c_851_n 0.00586131f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.515
cc_59 VNB N_VGND_c_852_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.515
cc_60 VNB N_VGND_c_853_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_854_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_855_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_856_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_857_n 0.0342743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_858_n 0.412273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_859_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_860_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_861_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_862_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_863_n 0.00884799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VPB N_B_M1001_g 0.0252952f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_72 VPB N_B_M1006_g 0.0196385f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_73 VPB N_B_M1007_g 0.0204814f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_74 VPB N_B_M1011_g 0.0206089f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=2.4
cc_75 VPB B 0.0175303f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_76 VPB N_B_c_123_n 0.0140936f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=1.515
cc_77 VPB N_A_468_264#_M1002_g 0.0221168f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.68
cc_78 VPB N_A_468_264#_M1005_g 0.022344f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.68
cc_79 VPB N_A_468_264#_M1009_g 0.0223661f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.68
cc_80 VPB N_A_468_264#_M1012_g 0.0249367f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_81 VPB N_A_468_264#_c_209_n 0.00416382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_468_264#_c_219_n 0.0202058f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_83 VPB N_A_468_264#_c_220_n 0.00329898f $X=-0.19 $Y=1.66 $X2=1.65 $Y2=1.515
cc_84 VPB N_A_468_264#_c_221_n 0.0121029f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=1.515
cc_85 VPB N_A_468_264#_c_211_n 0.00283905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_M1003_g 0.0254017f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_87 VPB N_A_M1013_g 0.020787f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_88 VPB N_A_M1017_g 0.0207885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_M1020_g 0.0230358f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=2.4
cc_90 VPB N_C_N_c_447_n 0.0171504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_C_N_c_448_n 0.0186777f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_92 VPB N_C_N_c_446_n 0.0140773f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_93 VPB N_A_27_368#_c_482_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_94 VPB N_A_27_368#_c_483_n 0.00240659f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_95 VPB N_A_27_368#_c_484_n 0.0100897f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_96 VPB N_A_27_368#_c_485_n 0.00280532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_368#_c_486_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_98 VPB N_A_27_368#_c_487_n 0.00195487f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_99 VPB N_A_27_368#_c_488_n 0.00327011f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_100 VPB N_A_129_368#_c_545_n 0.0131354f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.68
cc_101 VPB N_A_129_368#_c_546_n 0.0019553f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.35
cc_102 VPB N_A_129_368#_c_547_n 0.00225162f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=2.4
cc_103 VPB N_Y_c_625_n 0.00795728f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_104 VPB Y 0.00150284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_749_n 0.010226f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_106 VPB N_VPWR_c_750_n 0.0026822f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_107 VPB N_VPWR_c_751_n 0.0125833f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_108 VPB N_VPWR_c_752_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=2.4
cc_109 VPB N_VPWR_c_753_n 0.0508884f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=1.35
cc_110 VPB N_VPWR_c_754_n 0.110132f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_111 VPB N_VPWR_c_755_n 0.0164205f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_112 VPB N_VPWR_c_756_n 0.017373f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_113 VPB N_VPWR_c_757_n 0.0195748f $X=-0.19 $Y=1.66 $X2=1.65 $Y2=1.515
cc_114 VPB N_VPWR_c_758_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_115 VPB N_VPWR_c_759_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.565
cc_116 VPB N_VPWR_c_760_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_117 VPB N_VPWR_c_748_n 0.0967963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 N_B_c_123_n N_A_468_264#_M1002_g 0.0325713f $X=1.995 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B_M1026_g N_A_468_264#_M1000_g 0.0264048f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_120 N_B_M1026_g N_A_468_264#_c_209_n 2.25772e-19 $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B_M1026_g N_A_468_264#_c_213_n 0.0325713f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_122 B N_A_27_368#_c_482_n 0.0266008f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_123 N_B_M1001_g N_A_27_368#_c_483_n 0.0150267f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B_M1006_g N_A_27_368#_c_483_n 0.0140221f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B_M1007_g N_A_27_368#_c_485_n 0.0147273f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_126 N_B_M1011_g N_A_27_368#_c_485_n 0.00968688f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B_M1007_g N_A_27_368#_c_487_n 6.66876e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_128 N_B_M1011_g N_A_27_368#_c_487_n 0.00823454f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B_M1006_g N_A_129_368#_c_548_n 0.012931f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_130 N_B_M1007_g N_A_129_368#_c_548_n 0.0136684f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_131 B N_A_129_368#_c_548_n 0.0399165f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_132 N_B_c_123_n N_A_129_368#_c_548_n 4.90767e-19 $X=1.995 $Y=1.515 $X2=0
+ $Y2=0
cc_133 N_B_M1011_g N_A_129_368#_c_545_n 0.0184002f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_134 N_B_M1001_g N_A_129_368#_c_553_n 0.0119008f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_135 N_B_M1006_g N_A_129_368#_c_553_n 0.0116958f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_136 N_B_M1007_g N_A_129_368#_c_553_n 5.74809e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_137 B N_A_129_368#_c_553_n 0.0235495f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_138 N_B_c_123_n N_A_129_368#_c_553_n 5.54777e-19 $X=1.995 $Y=1.515 $X2=0
+ $Y2=0
cc_139 N_B_M1006_g N_A_129_368#_c_558_n 5.68615e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B_M1007_g N_A_129_368#_c_558_n 0.0119056f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_141 B N_A_129_368#_c_558_n 0.0228945f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_142 N_B_c_123_n N_A_129_368#_c_558_n 0.00101037f $X=1.995 $Y=1.515 $X2=0
+ $Y2=0
cc_143 N_B_M1010_g N_Y_c_611_n 4.71232e-19 $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_144 N_B_M1015_g N_Y_c_611_n 0.00959262f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_145 N_B_M1025_g N_Y_c_611_n 6.3028e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_146 N_B_M1010_g N_Y_c_612_n 0.00190113f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_147 N_B_M1015_g N_Y_c_612_n 0.0016171f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_148 B N_Y_c_612_n 0.028235f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B_c_123_n N_Y_c_612_n 0.00305f $X=1.995 $Y=1.515 $X2=0 $Y2=0
cc_150 N_B_M1015_g N_Y_c_613_n 5.35648e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B_M1025_g N_Y_c_613_n 0.00916462f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_152 N_B_M1026_g N_Y_c_613_n 0.00924167f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_153 N_B_M1007_g N_Y_c_637_n 3.37347e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_154 N_B_M1011_g N_Y_c_637_n 0.00732172f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_155 N_B_M1015_g N_Y_c_620_n 0.0118691f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B_M1025_g N_Y_c_620_n 0.0118691f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_157 B N_Y_c_620_n 0.0658285f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_158 N_B_c_123_n N_Y_c_620_n 0.00597192f $X=1.995 $Y=1.515 $X2=0 $Y2=0
cc_159 N_B_M1025_g N_Y_c_621_n 0.00220179f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_160 N_B_M1026_g N_Y_c_621_n 0.0177513f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_161 N_B_c_123_n N_Y_c_621_n 0.00260449f $X=1.995 $Y=1.515 $X2=0 $Y2=0
cc_162 N_B_M1007_g Y 2.57774e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B_M1025_g Y 8.28286e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B_M1011_g Y 0.00314843f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B_M1026_g Y 0.00472643f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_166 B Y 0.0265484f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_167 N_B_c_123_n Y 0.00885602f $X=1.995 $Y=1.515 $X2=0 $Y2=0
cc_168 N_B_M1001_g N_VPWR_c_754_n 0.00333926f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_169 N_B_M1006_g N_VPWR_c_754_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B_M1007_g N_VPWR_c_754_n 0.00333926f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_171 N_B_M1011_g N_VPWR_c_754_n 0.00335119f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_172 N_B_M1001_g N_VPWR_c_748_n 0.00426591f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B_M1006_g N_VPWR_c_748_n 0.00422687f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B_M1007_g N_VPWR_c_748_n 0.00423403f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B_M1011_g N_VPWR_c_748_n 0.00422602f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_176 N_B_M1010_g N_VGND_c_843_n 0.00549949f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_177 B N_VGND_c_843_n 0.0239925f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_178 N_B_M1015_g N_VGND_c_844_n 0.00484409f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B_M1025_g N_VGND_c_844_n 0.00484409f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B_M1025_g N_VGND_c_845_n 0.00434272f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B_M1026_g N_VGND_c_845_n 0.00434272f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B_M1026_g N_VGND_c_846_n 0.00417204f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B_M1010_g N_VGND_c_854_n 0.00461464f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B_M1015_g N_VGND_c_854_n 0.00434272f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_185 N_B_M1010_g N_VGND_c_858_n 0.00911596f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B_M1015_g N_VGND_c_858_n 0.00821539f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B_M1025_g N_VGND_c_858_n 0.00821294f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B_M1026_g N_VGND_c_858_n 0.00820772f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_468_264#_M1019_g N_A_c_352_n 0.0161937f $X=3.855 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_468_264#_c_209_n N_A_M1003_g 0.00488235f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_191 N_A_468_264#_c_219_n N_A_M1003_g 0.0141217f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_192 N_A_468_264#_c_219_n N_A_M1013_g 0.0116635f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_193 N_A_468_264#_c_219_n N_A_M1017_g 0.0116635f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_194 N_A_468_264#_c_219_n N_A_M1020_g 0.016899f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_195 N_A_468_264#_c_220_n N_A_M1020_g 6.47579e-19 $X=6.95 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_468_264#_c_209_n N_A_c_361_n 0.00245232f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_197 N_A_468_264#_c_219_n N_A_c_361_n 0.0161563f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_198 N_A_468_264#_c_213_n N_A_c_361_n 0.0161937f $X=3.855 $Y=1.485 $X2=0 $Y2=0
cc_199 N_A_468_264#_M1019_g N_A_c_362_n 4.72901e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_468_264#_c_209_n N_A_c_362_n 0.014508f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_201 N_A_468_264#_c_219_n N_A_c_362_n 0.160908f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_202 N_A_468_264#_c_212_n N_C_N_c_444_n 0.0094203f $X=7.4 $Y=0.5 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_468_264#_c_219_n N_C_N_c_447_n 0.0103668f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_204 N_A_468_264#_c_220_n N_C_N_c_447_n 0.0134502f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_468_264#_c_243_p N_C_N_c_447_n 0.00126234f $X=6.92 $Y=1.805 $X2=0
+ $Y2=0
cc_206 N_A_468_264#_c_220_n N_C_N_c_448_n 8.71028e-19 $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_468_264#_c_221_n N_C_N_c_448_n 0.0126739f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_208 N_A_468_264#_c_219_n C_N 0.00134249f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_209 N_A_468_264#_c_221_n C_N 0.00279147f $X=7.395 $Y=1.805 $X2=0 $Y2=0
cc_210 N_A_468_264#_c_211_n C_N 0.0183654f $X=7.48 $Y=1.72 $X2=0 $Y2=0
cc_211 N_A_468_264#_c_243_p C_N 0.0218449f $X=6.92 $Y=1.805 $X2=0 $Y2=0
cc_212 N_A_468_264#_c_212_n C_N 0.0286132f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_213 N_A_468_264#_c_219_n N_C_N_c_446_n 0.00874303f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_214 N_A_468_264#_c_221_n N_C_N_c_446_n 0.00909837f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_215 N_A_468_264#_c_211_n N_C_N_c_446_n 0.0162405f $X=7.48 $Y=1.72 $X2=0 $Y2=0
cc_216 N_A_468_264#_c_243_p N_C_N_c_446_n 0.00716382f $X=6.92 $Y=1.805 $X2=0
+ $Y2=0
cc_217 N_A_468_264#_c_212_n N_C_N_c_446_n 0.0145695f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_218 N_A_468_264#_c_209_n N_A_27_368#_M1012_s 0.00408381f $X=3.89 $Y=1.485
+ $X2=0 $Y2=0
cc_219 N_A_468_264#_M1009_g N_A_27_368#_c_497_n 0.00926474f $X=3.33 $Y=2.4 $X2=0
+ $Y2=0
cc_220 N_A_468_264#_M1012_g N_A_27_368#_c_497_n 0.00984351f $X=3.78 $Y=2.4 $X2=0
+ $Y2=0
cc_221 N_A_468_264#_M1002_g N_A_27_368#_c_487_n 0.00924373f $X=2.43 $Y=2.4 $X2=0
+ $Y2=0
cc_222 N_A_468_264#_M1005_g N_A_27_368#_c_487_n 0.00133025f $X=2.88 $Y=2.4 $X2=0
+ $Y2=0
cc_223 N_A_468_264#_M1002_g N_A_27_368#_c_501_n 0.00981134f $X=2.43 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_468_264#_M1005_g N_A_27_368#_c_501_n 0.00926474f $X=2.88 $Y=2.4 $X2=0
+ $Y2=0
cc_225 N_A_468_264#_M1002_g N_A_27_368#_c_503_n 4.65366e-19 $X=2.43 $Y=2.4 $X2=0
+ $Y2=0
cc_226 N_A_468_264#_M1005_g N_A_27_368#_c_503_n 0.00430608f $X=2.88 $Y=2.4 $X2=0
+ $Y2=0
cc_227 N_A_468_264#_M1009_g N_A_27_368#_c_503_n 0.00430608f $X=3.33 $Y=2.4 $X2=0
+ $Y2=0
cc_228 N_A_468_264#_M1012_g N_A_27_368#_c_503_n 4.65366e-19 $X=3.78 $Y=2.4 $X2=0
+ $Y2=0
cc_229 N_A_468_264#_M1009_g N_A_27_368#_c_488_n 5.44851e-19 $X=3.33 $Y=2.4 $X2=0
+ $Y2=0
cc_230 N_A_468_264#_M1012_g N_A_27_368#_c_488_n 0.00476329f $X=3.78 $Y=2.4 $X2=0
+ $Y2=0
cc_231 N_A_468_264#_c_219_n N_A_129_368#_M1003_d 0.00165831f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_232 N_A_468_264#_c_219_n N_A_129_368#_M1017_d 0.00165831f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_233 N_A_468_264#_M1002_g N_A_129_368#_c_545_n 0.0116099f $X=2.43 $Y=2.4 $X2=0
+ $Y2=0
cc_234 N_A_468_264#_M1005_g N_A_129_368#_c_545_n 0.0116635f $X=2.88 $Y=2.4 $X2=0
+ $Y2=0
cc_235 N_A_468_264#_M1009_g N_A_129_368#_c_545_n 0.0116635f $X=3.33 $Y=2.4 $X2=0
+ $Y2=0
cc_236 N_A_468_264#_M1012_g N_A_129_368#_c_545_n 0.0157766f $X=3.78 $Y=2.4 $X2=0
+ $Y2=0
cc_237 N_A_468_264#_c_209_n N_A_129_368#_c_545_n 0.0168146f $X=3.89 $Y=1.485
+ $X2=0 $Y2=0
cc_238 N_A_468_264#_c_219_n N_A_129_368#_c_545_n 0.0234174f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_239 N_A_468_264#_c_219_n N_A_129_368#_c_570_n 0.0356639f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_240 N_A_468_264#_c_219_n N_A_129_368#_c_571_n 0.0149351f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_241 N_A_468_264#_c_219_n N_A_129_368#_c_572_n 0.0187124f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_242 N_A_468_264#_M1000_g N_Y_c_613_n 8.87957e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_468_264#_M1000_g N_Y_c_614_n 0.0152745f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_468_264#_c_209_n N_Y_c_614_n 0.00334513f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_245 N_A_468_264#_c_213_n N_Y_c_614_n 0.00250279f $X=3.855 $Y=1.485 $X2=0
+ $Y2=0
cc_246 N_A_468_264#_M1002_g N_Y_c_625_n 0.0145965f $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_468_264#_M1005_g N_Y_c_625_n 0.0122575f $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_468_264#_M1009_g N_Y_c_625_n 0.0122575f $X=3.33 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_468_264#_M1012_g N_Y_c_625_n 0.0104071f $X=3.78 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_468_264#_c_209_n N_Y_c_625_n 0.0903855f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_251 N_A_468_264#_c_213_n N_Y_c_625_n 0.00673897f $X=3.855 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_468_264#_M1000_g N_Y_c_615_n 3.92313e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_468_264#_M1004_g N_Y_c_615_n 3.92313e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_468_264#_M1004_g N_Y_c_616_n 0.0131239f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_468_264#_M1016_g N_Y_c_616_n 0.0115433f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_468_264#_c_209_n N_Y_c_616_n 0.0500092f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_257 N_A_468_264#_c_213_n N_Y_c_616_n 0.00424488f $X=3.855 $Y=1.485 $X2=0
+ $Y2=0
cc_258 N_A_468_264#_M1004_g N_Y_c_617_n 4.13007e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_468_264#_M1016_g N_Y_c_617_n 0.00721977f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_468_264#_M1019_g N_Y_c_617_n 0.00834185f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_468_264#_M1019_g N_Y_c_671_n 0.0120704f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_468_264#_c_209_n N_Y_c_671_n 0.0202341f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_263 N_A_468_264#_c_219_n N_Y_c_671_n 0.00575327f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_264 N_A_468_264#_M1019_g N_Y_c_618_n 6.03013e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_468_264#_M1000_g N_Y_c_621_n 8.44859e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_468_264#_c_209_n N_Y_c_622_n 0.0143381f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_267 N_A_468_264#_c_213_n N_Y_c_622_n 0.00256622f $X=3.855 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_468_264#_M1004_g N_Y_c_623_n 4.68741e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_468_264#_M1016_g N_Y_c_623_n 0.00330557f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_468_264#_M1019_g N_Y_c_623_n 0.00342047f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_468_264#_c_209_n N_Y_c_623_n 0.0276081f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_272 N_A_468_264#_c_213_n N_Y_c_623_n 0.00268454f $X=3.855 $Y=1.485 $X2=0
+ $Y2=0
cc_273 N_A_468_264#_M1000_g Y 0.00326736f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_468_264#_c_209_n Y 0.0172568f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_275 N_A_468_264#_c_213_n Y 0.00776015f $X=3.855 $Y=1.485 $X2=0 $Y2=0
cc_276 N_A_468_264#_c_219_n N_VPWR_M1003_s 0.0036083f $X=6.785 $Y=1.805
+ $X2=-0.19 $Y2=-0.245
cc_277 N_A_468_264#_c_219_n N_VPWR_M1013_s 0.00166235f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_278 N_A_468_264#_c_219_n N_VPWR_M1020_s 0.00321543f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_279 N_A_468_264#_c_221_n N_VPWR_M1023_s 0.00270206f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_280 N_A_468_264#_M1012_g N_VPWR_c_749_n 0.00425493f $X=3.78 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_A_468_264#_c_219_n N_VPWR_c_751_n 0.0236753f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_282 N_A_468_264#_c_220_n N_VPWR_c_751_n 0.0207405f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_283 N_A_468_264#_c_220_n N_VPWR_c_753_n 0.0236749f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A_468_264#_c_221_n N_VPWR_c_753_n 0.0233742f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_285 N_A_468_264#_M1002_g N_VPWR_c_754_n 0.00376977f $X=2.43 $Y=2.4 $X2=0
+ $Y2=0
cc_286 N_A_468_264#_M1005_g N_VPWR_c_754_n 0.00380305f $X=2.88 $Y=2.4 $X2=0
+ $Y2=0
cc_287 N_A_468_264#_M1009_g N_VPWR_c_754_n 0.00380305f $X=3.33 $Y=2.4 $X2=0
+ $Y2=0
cc_288 N_A_468_264#_M1012_g N_VPWR_c_754_n 0.0038135f $X=3.78 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A_468_264#_c_220_n N_VPWR_c_757_n 0.00541659f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_A_468_264#_M1002_g N_VPWR_c_748_n 0.00469163f $X=2.43 $Y=2.4 $X2=0
+ $Y2=0
cc_291 N_A_468_264#_M1005_g N_VPWR_c_748_n 0.00472981f $X=2.88 $Y=2.4 $X2=0
+ $Y2=0
cc_292 N_A_468_264#_M1009_g N_VPWR_c_748_n 0.00472981f $X=3.33 $Y=2.4 $X2=0
+ $Y2=0
cc_293 N_A_468_264#_M1012_g N_VPWR_c_748_n 0.00477074f $X=3.78 $Y=2.4 $X2=0
+ $Y2=0
cc_294 N_A_468_264#_c_220_n N_VPWR_c_748_n 0.00812781f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A_468_264#_M1000_g N_VGND_c_846_n 0.0100169f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_296 N_A_468_264#_M1004_g N_VGND_c_846_n 4.62684e-19 $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_468_264#_M1000_g N_VGND_c_847_n 4.62684e-19 $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_468_264#_M1004_g N_VGND_c_847_n 0.0100169f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_468_264#_M1016_g N_VGND_c_847_n 0.00417204f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_468_264#_M1019_g N_VGND_c_848_n 0.00405455f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_301 N_A_468_264#_c_212_n N_VGND_c_851_n 0.0284697f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_302 N_A_468_264#_M1000_g N_VGND_c_855_n 0.00383152f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_468_264#_M1004_g N_VGND_c_855_n 0.00383152f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_468_264#_M1016_g N_VGND_c_856_n 0.00434272f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_468_264#_M1019_g N_VGND_c_856_n 0.00434272f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_468_264#_c_210_n N_VGND_c_857_n 0.00758556f $X=7.48 $Y=1.01 $X2=0
+ $Y2=0
cc_307 N_A_468_264#_c_212_n N_VGND_c_857_n 0.0349297f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_308 N_A_468_264#_M1000_g N_VGND_c_858_n 0.0075754f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A_468_264#_M1004_g N_VGND_c_858_n 0.0075754f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_310 N_A_468_264#_M1016_g N_VGND_c_858_n 0.00820718f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_311 N_A_468_264#_M1019_g N_VGND_c_858_n 0.00821312f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_312 N_A_468_264#_c_210_n N_VGND_c_858_n 0.00627867f $X=7.48 $Y=1.01 $X2=0
+ $Y2=0
cc_313 N_A_468_264#_c_212_n N_VGND_c_858_n 0.0289999f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_314 N_A_c_358_n N_C_N_c_444_n 0.0116655f $X=6.055 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_315 A N_C_N_c_444_n 0.00650444f $X=6.395 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_316 N_A_M1020_g N_C_N_c_447_n 0.0136604f $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_317 A C_N 0.030054f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_318 A N_C_N_c_446_n 0.0102326f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_319 N_A_c_361_n N_C_N_c_446_n 0.0258741f $X=6.055 $Y=1.385 $X2=0 $Y2=0
cc_320 N_A_M1003_g N_A_129_368#_c_545_n 0.0117729f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_321 N_A_M1003_g N_A_129_368#_c_546_n 2.23201e-19 $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_322 N_A_M1013_g N_A_129_368#_c_546_n 2.23201e-19 $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_323 N_A_M1013_g N_A_129_368#_c_570_n 0.0142562f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_324 N_A_M1017_g N_A_129_368#_c_570_n 0.0142175f $X=5.69 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A_M1020_g N_A_129_368#_c_571_n 0.00236488f $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_326 N_A_M1017_g N_A_129_368#_c_547_n 2.33902e-19 $X=5.69 $Y=2.4 $X2=0 $Y2=0
cc_327 N_A_M1020_g N_A_129_368#_c_547_n 0.00924834f $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_328 N_A_M1003_g N_A_129_368#_c_572_n 0.0157401f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_329 N_A_c_352_n N_Y_c_617_n 6.03013e-19 $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_330 N_A_c_352_n N_Y_c_671_n 0.0127102f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_331 N_A_c_362_n N_Y_c_671_n 0.00246555f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_332 N_A_c_352_n N_Y_c_618_n 0.00834185f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_333 N_A_c_354_n N_Y_c_618_n 0.00907544f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_334 N_A_c_356_n N_Y_c_618_n 8.95441e-19 $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_335 N_A_c_354_n N_Y_c_692_n 0.0121454f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_336 N_A_c_356_n N_Y_c_692_n 0.0128634f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_337 N_A_c_361_n N_Y_c_692_n 0.0141443f $X=6.055 $Y=1.385 $X2=0 $Y2=0
cc_338 N_A_c_362_n N_Y_c_692_n 0.0783501f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_339 N_A_c_354_n N_Y_c_619_n 8.95441e-19 $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_340 N_A_c_356_n N_Y_c_619_n 0.00908017f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_341 N_A_c_358_n N_Y_c_619_n 0.00282572f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_342 N_A_c_352_n N_Y_c_623_n 4.52963e-19 $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_343 N_A_c_352_n N_Y_c_700_n 7.18016e-19 $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_344 N_A_c_354_n N_Y_c_700_n 7.18016e-19 $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_345 N_A_c_361_n N_Y_c_700_n 0.00232761f $X=6.055 $Y=1.385 $X2=0 $Y2=0
cc_346 N_A_c_362_n N_Y_c_700_n 0.021954f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_347 N_A_M1003_g N_VPWR_c_749_n 0.0107927f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A_M1013_g N_VPWR_c_749_n 4.23447e-19 $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_349 N_A_M1003_g N_VPWR_c_750_n 4.77201e-19 $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_350 N_A_M1013_g N_VPWR_c_750_n 0.0113952f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A_M1017_g N_VPWR_c_750_n 0.0112069f $X=5.69 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A_M1020_g N_VPWR_c_750_n 4.81631e-19 $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_353 N_A_M1020_g N_VPWR_c_751_n 0.00381366f $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_354 N_A_M1003_g N_VPWR_c_755_n 0.00460063f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_355 N_A_M1013_g N_VPWR_c_755_n 0.00460063f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_356 N_A_M1017_g N_VPWR_c_756_n 0.00460063f $X=5.69 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A_M1020_g N_VPWR_c_756_n 0.00520636f $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_358 N_A_M1003_g N_VPWR_c_748_n 0.00908554f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A_M1013_g N_VPWR_c_748_n 0.00908554f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A_M1017_g N_VPWR_c_748_n 0.00908554f $X=5.69 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A_M1020_g N_VPWR_c_748_n 0.00986533f $X=6.14 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A_c_352_n N_VGND_c_848_n 0.00405455f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_363 N_A_c_352_n N_VGND_c_849_n 0.00434272f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_364 N_A_c_354_n N_VGND_c_849_n 0.00434272f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_365 N_A_c_354_n N_VGND_c_850_n 0.00460818f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_366 N_A_c_356_n N_VGND_c_850_n 0.00460818f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_367 N_A_c_356_n N_VGND_c_851_n 5.39035e-19 $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_368 N_A_c_358_n N_VGND_c_851_n 0.011573f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_369 A N_VGND_c_851_n 0.00553831f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_370 N_A_c_361_n N_VGND_c_851_n 3.8009e-19 $X=6.055 $Y=1.385 $X2=0 $Y2=0
cc_371 N_A_c_362_n N_VGND_c_851_n 0.016837f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_372 N_A_c_356_n N_VGND_c_852_n 0.00434272f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_373 N_A_c_358_n N_VGND_c_852_n 0.00383152f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_374 N_A_c_352_n N_VGND_c_858_n 0.00821312f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_375 N_A_c_354_n N_VGND_c_858_n 0.00822177f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_376 N_A_c_356_n N_VGND_c_858_n 0.00822835f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_377 N_A_c_358_n N_VGND_c_858_n 0.00758198f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_378 N_C_N_c_447_n N_VPWR_c_751_n 0.00570014f $X=6.725 $Y=1.76 $X2=0 $Y2=0
cc_379 N_C_N_c_447_n N_VPWR_c_753_n 5.91121e-19 $X=6.725 $Y=1.76 $X2=0 $Y2=0
cc_380 N_C_N_c_448_n N_VPWR_c_753_n 0.0132364f $X=7.175 $Y=1.76 $X2=0 $Y2=0
cc_381 N_C_N_c_447_n N_VPWR_c_757_n 0.00465228f $X=6.725 $Y=1.76 $X2=0 $Y2=0
cc_382 N_C_N_c_448_n N_VPWR_c_757_n 0.00401533f $X=7.175 $Y=1.76 $X2=0 $Y2=0
cc_383 N_C_N_c_447_n N_VPWR_c_748_n 0.00555093f $X=6.725 $Y=1.76 $X2=0 $Y2=0
cc_384 N_C_N_c_448_n N_VPWR_c_748_n 0.00465661f $X=7.175 $Y=1.76 $X2=0 $Y2=0
cc_385 N_C_N_c_444_n N_VGND_c_851_n 0.00661609f $X=6.555 $Y=1.22 $X2=0 $Y2=0
cc_386 N_C_N_c_444_n N_VGND_c_857_n 0.00433162f $X=6.555 $Y=1.22 $X2=0 $Y2=0
cc_387 N_C_N_c_444_n N_VGND_c_858_n 0.00822119f $X=6.555 $Y=1.22 $X2=0 $Y2=0
cc_388 N_A_27_368#_c_483_n N_A_129_368#_M1001_s 0.00165831f $X=1.145 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_389 N_A_27_368#_c_485_n N_A_129_368#_M1007_s 0.00245557f $X=2.04 $Y=2.99
+ $X2=0 $Y2=0
cc_390 N_A_27_368#_M1006_d N_A_129_368#_c_548_n 0.00314376f $X=1.095 $Y=1.84
+ $X2=0 $Y2=0
cc_391 N_A_27_368#_c_512_p N_A_129_368#_c_548_n 0.0126919f $X=1.23 $Y=2.455
+ $X2=0 $Y2=0
cc_392 N_A_27_368#_M1011_d N_A_129_368#_c_545_n 0.00331683f $X=2.07 $Y=1.84
+ $X2=0 $Y2=0
cc_393 N_A_27_368#_M1005_s N_A_129_368#_c_545_n 0.00324035f $X=2.97 $Y=1.84
+ $X2=0 $Y2=0
cc_394 N_A_27_368#_M1012_s N_A_129_368#_c_545_n 0.00658775f $X=3.87 $Y=1.84
+ $X2=0 $Y2=0
cc_395 N_A_27_368#_c_485_n N_A_129_368#_c_545_n 0.00425589f $X=2.04 $Y=2.99
+ $X2=0 $Y2=0
cc_396 N_A_27_368#_c_487_n N_A_129_368#_c_545_n 0.0165925f $X=2.205 $Y=2.665
+ $X2=0 $Y2=0
cc_397 N_A_27_368#_c_501_n N_A_129_368#_c_545_n 0.0793935f $X=2.94 $Y=2.745
+ $X2=0 $Y2=0
cc_398 N_A_27_368#_c_488_n N_A_129_368#_c_545_n 0.0206828f $X=4.005 $Y=2.665
+ $X2=0 $Y2=0
cc_399 N_A_27_368#_c_483_n N_A_129_368#_c_553_n 0.0159318f $X=1.145 $Y=2.99
+ $X2=0 $Y2=0
cc_400 N_A_27_368#_c_485_n N_A_129_368#_c_558_n 0.0189699f $X=2.04 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_27_368#_c_501_n N_Y_M1002_d 0.00420242f $X=2.94 $Y=2.745 $X2=0 $Y2=0
cc_402 N_A_27_368#_c_497_n N_Y_M1009_d 0.00420242f $X=3.84 $Y=2.665 $X2=0 $Y2=0
cc_403 N_A_27_368#_M1011_d N_Y_c_637_n 0.00164183f $X=2.07 $Y=1.84 $X2=0 $Y2=0
cc_404 N_A_27_368#_M1005_s N_Y_c_625_n 0.00168223f $X=2.97 $Y=1.84 $X2=0 $Y2=0
cc_405 N_A_27_368#_c_488_n N_VPWR_c_749_n 0.022248f $X=4.005 $Y=2.665 $X2=0
+ $Y2=0
cc_406 N_A_27_368#_c_483_n N_VPWR_c_754_n 0.0439866f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_407 N_A_27_368#_c_484_n N_VPWR_c_754_n 0.0236566f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_408 N_A_27_368#_c_485_n N_VPWR_c_754_n 0.0457135f $X=2.04 $Y=2.99 $X2=0 $Y2=0
cc_409 N_A_27_368#_c_497_n N_VPWR_c_754_n 0.00996337f $X=3.84 $Y=2.665 $X2=0
+ $Y2=0
cc_410 N_A_27_368#_c_486_n N_VPWR_c_754_n 0.0121867f $X=1.23 $Y=2.99 $X2=0 $Y2=0
cc_411 N_A_27_368#_c_487_n N_VPWR_c_754_n 0.0227642f $X=2.205 $Y=2.665 $X2=0
+ $Y2=0
cc_412 N_A_27_368#_c_501_n N_VPWR_c_754_n 0.00996337f $X=2.94 $Y=2.745 $X2=0
+ $Y2=0
cc_413 N_A_27_368#_c_503_n N_VPWR_c_754_n 0.00884253f $X=3.27 $Y=2.745 $X2=0
+ $Y2=0
cc_414 N_A_27_368#_c_488_n N_VPWR_c_754_n 0.00968772f $X=4.005 $Y=2.665 $X2=0
+ $Y2=0
cc_415 N_A_27_368#_c_483_n N_VPWR_c_748_n 0.0246722f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_416 N_A_27_368#_c_484_n N_VPWR_c_748_n 0.0128296f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_417 N_A_27_368#_c_485_n N_VPWR_c_748_n 0.0257527f $X=2.04 $Y=2.99 $X2=0 $Y2=0
cc_418 N_A_27_368#_c_497_n N_VPWR_c_748_n 0.0154919f $X=3.84 $Y=2.665 $X2=0
+ $Y2=0
cc_419 N_A_27_368#_c_486_n N_VPWR_c_748_n 0.00660921f $X=1.23 $Y=2.99 $X2=0
+ $Y2=0
cc_420 N_A_27_368#_c_487_n N_VPWR_c_748_n 0.0123829f $X=2.205 $Y=2.665 $X2=0
+ $Y2=0
cc_421 N_A_27_368#_c_501_n N_VPWR_c_748_n 0.0154919f $X=2.94 $Y=2.745 $X2=0
+ $Y2=0
cc_422 N_A_27_368#_c_503_n N_VPWR_c_748_n 0.0110299f $X=3.27 $Y=2.745 $X2=0
+ $Y2=0
cc_423 N_A_27_368#_c_488_n N_VPWR_c_748_n 0.0111351f $X=4.005 $Y=2.665 $X2=0
+ $Y2=0
cc_424 N_A_129_368#_c_545_n N_Y_M1002_d 0.00320838f $X=4.795 $Y=2.325 $X2=0
+ $Y2=0
cc_425 N_A_129_368#_c_545_n N_Y_M1009_d 0.00324035f $X=4.795 $Y=2.325 $X2=0
+ $Y2=0
cc_426 N_A_129_368#_c_545_n N_Y_c_637_n 0.0139033f $X=4.795 $Y=2.325 $X2=0 $Y2=0
cc_427 N_A_129_368#_c_545_n N_Y_c_625_n 0.0752334f $X=4.795 $Y=2.325 $X2=0 $Y2=0
cc_428 N_A_129_368#_c_545_n N_VPWR_M1003_s 0.00635246f $X=4.795 $Y=2.325
+ $X2=-0.19 $Y2=1.66
cc_429 N_A_129_368#_c_570_n N_VPWR_M1013_s 0.00321662f $X=5.81 $Y=2.145 $X2=0
+ $Y2=0
cc_430 N_A_129_368#_c_545_n N_VPWR_c_749_n 0.0219147f $X=4.795 $Y=2.325 $X2=0
+ $Y2=0
cc_431 N_A_129_368#_c_546_n N_VPWR_c_749_n 0.0144807f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_432 N_A_129_368#_c_546_n N_VPWR_c_750_n 0.0204109f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_433 N_A_129_368#_c_570_n N_VPWR_c_750_n 0.0170259f $X=5.81 $Y=2.145 $X2=0
+ $Y2=0
cc_434 N_A_129_368#_c_547_n N_VPWR_c_750_n 0.0222705f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_435 N_A_129_368#_c_547_n N_VPWR_c_751_n 0.0288238f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_436 N_A_129_368#_c_546_n N_VPWR_c_755_n 0.00780931f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_437 N_A_129_368#_c_547_n N_VPWR_c_756_n 0.0123696f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_438 N_A_129_368#_c_546_n N_VPWR_c_748_n 0.00624184f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_439 N_A_129_368#_c_547_n N_VPWR_c_748_n 0.00981798f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_440 N_Y_c_620_n N_VGND_M1015_d 0.00358162f $X=1.615 $Y=1.08 $X2=0 $Y2=0
cc_441 N_Y_c_614_n N_VGND_M1026_d 9.24827e-19 $X=2.625 $Y=1.065 $X2=0 $Y2=0
cc_442 N_Y_c_621_n N_VGND_M1026_d 0.00158118f $X=2.275 $Y=1.08 $X2=0 $Y2=0
cc_443 N_Y_c_616_n N_VGND_M1004_d 0.00250873f $X=3.475 $Y=1.065 $X2=0 $Y2=0
cc_444 N_Y_c_671_n N_VGND_M1019_d 0.00859297f $X=4.475 $Y=0.965 $X2=0 $Y2=0
cc_445 N_Y_c_692_n N_VGND_M1018_s 0.0104519f $X=5.605 $Y=0.965 $X2=0 $Y2=0
cc_446 N_Y_c_611_n N_VGND_c_843_n 0.0256697f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_447 N_Y_c_612_n N_VGND_c_843_n 0.00630154f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_448 N_Y_c_611_n N_VGND_c_844_n 0.0191765f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_449 N_Y_c_613_n N_VGND_c_844_n 0.0191765f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_450 N_Y_c_620_n N_VGND_c_844_n 0.0248957f $X=1.615 $Y=1.08 $X2=0 $Y2=0
cc_451 N_Y_c_613_n N_VGND_c_845_n 0.0144124f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_452 N_Y_c_613_n N_VGND_c_846_n 0.0180508f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_453 N_Y_c_615_n N_VGND_c_846_n 0.0171736f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_454 N_Y_c_621_n N_VGND_c_846_n 0.0210834f $X=2.275 $Y=1.08 $X2=0 $Y2=0
cc_455 N_Y_c_615_n N_VGND_c_847_n 0.0171736f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_456 N_Y_c_616_n N_VGND_c_847_n 0.0209867f $X=3.475 $Y=1.065 $X2=0 $Y2=0
cc_457 N_Y_c_617_n N_VGND_c_847_n 0.0180508f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_458 N_Y_c_617_n N_VGND_c_848_n 0.0142986f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_459 N_Y_c_671_n N_VGND_c_848_n 0.0248957f $X=4.475 $Y=0.965 $X2=0 $Y2=0
cc_460 N_Y_c_618_n N_VGND_c_848_n 0.0142986f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_461 N_Y_c_618_n N_VGND_c_849_n 0.0145227f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_462 N_Y_c_618_n N_VGND_c_850_n 0.0132136f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_463 N_Y_c_692_n N_VGND_c_850_n 0.0314257f $X=5.605 $Y=0.965 $X2=0 $Y2=0
cc_464 N_Y_c_619_n N_VGND_c_850_n 0.0132136f $X=5.77 $Y=0.515 $X2=0 $Y2=0
cc_465 N_Y_c_619_n N_VGND_c_851_n 0.0206774f $X=5.77 $Y=0.515 $X2=0 $Y2=0
cc_466 N_Y_c_619_n N_VGND_c_852_n 0.0145947f $X=5.77 $Y=0.515 $X2=0 $Y2=0
cc_467 N_Y_c_611_n N_VGND_c_854_n 0.0145639f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_468 N_Y_c_615_n N_VGND_c_855_n 0.00749631f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_469 N_Y_c_617_n N_VGND_c_856_n 0.0144922f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_470 N_Y_c_611_n N_VGND_c_858_n 0.0119984f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_471 N_Y_c_613_n N_VGND_c_858_n 0.0118513f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_472 N_Y_c_615_n N_VGND_c_858_n 0.0062048f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_473 N_Y_c_617_n N_VGND_c_858_n 0.0118826f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_474 N_Y_c_618_n N_VGND_c_858_n 0.0118946f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_475 N_Y_c_619_n N_VGND_c_858_n 0.0120104f $X=5.77 $Y=0.515 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__dlxtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
M1000 Q a_842_405# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=1.54015e+12p ps=1.207e+07u
M1001 VPWR D a_27_120# VPB pshort w=840000u l=180000u
+  ad=1.89385e+12p pd=1.485e+07u as=2.352e+11p ps=2.24e+06u
M1002 a_672_392# a_232_82# a_658_79# VNB nlowvt w=640000u l=150000u
+  ad=2.803e+11p pd=2.53e+06u as=1.536e+11p ps=1.76e+06u
M1003 a_658_79# a_27_120# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_232_82# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VPWR a_842_405# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.528e+11p ps=2.87e+06u
M1006 VGND a_842_405# a_875_139# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 VPWR a_842_405# a_794_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VGND a_232_82# a_369_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_588_392# a_27_120# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1010 VGND a_842_405# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_842_405# a_672_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_672_392# a_369_392# a_588_392# VPB pshort w=1e+06u l=180000u
+  ad=3.83875e+11p pd=2.86e+06u as=0p ps=0u
M1013 a_875_139# a_369_392# a_672_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_842_405# a_672_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 a_794_503# a_232_82# a_672_392# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND D a_27_120# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 a_232_82# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1018 VPWR a_232_82# a_369_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1019 Q a_842_405# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


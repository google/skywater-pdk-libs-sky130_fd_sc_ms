* File: sky130_fd_sc_ms__a2111o_2.spice
* Created: Fri Aug 28 16:55:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2111o_2.pex.spice"
.subckt sky130_fd_sc_ms__a2111o_2  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_91_244#_M1008_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_91_244#_M1009_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_D1_M1013_g N_A_91_244#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1961 PD=1.06 PS=2.01 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_91_244#_M1003_d N_C1_M1003_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75000.7
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_B1_M1012_g N_A_91_244#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=1.31 PS=1.02 NRD=27.564 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1010 A_771_74# N_A2_M1010_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.2109 PD=0.95 PS=1.31 NRD=8.1 NRS=19.452 M=1 R=4.93333 SA=75001.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_91_244#_M1011_d N_A1_M1011_g A_771_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1004_d N_A_91_244#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1004_d N_A_91_244#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 A_447_368# N_D1_M1001_g N_A_91_244#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1176 AS=0.2912 PD=1.33 PS=2.76 NRD=8.7862 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1006 A_525_368# N_C1_M1006_g A_447_368# VPB PSHORT L=0.18 W=1.12 AD=0.2016
+ AS=0.1176 PD=1.48 PS=1.33 NRD=21.9852 NRS=8.7862 M=1 R=6.22222 SA=90000.6
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1000 N_A_633_368#_M1000_d N_B1_M1000_g A_525_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.2016 PD=1.48 PS=1.48 NRD=2.6201 NRS=21.9852 M=1 R=6.22222
+ SA=90001.1 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_633_368#_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.2016 PD=1.48 PS=1.48 NRD=2.6201 NRS=11.426 M=1 R=6.22222
+ SA=90001.6 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1007 N_A_633_368#_M1007_d N_A1_M1007_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2016 PD=2.76 PS=1.48 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90002.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_85 VPB 0 1.2388e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__a2111o_2.pxi.spice"
*
.ends
*
*

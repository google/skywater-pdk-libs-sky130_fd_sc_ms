* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_837_359# a_699_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.38125e+11p pd=2.8e+06u as=2.1627e+12p ps=1.993e+07u
M1001 VGND RESET_B a_895_138# VNB nlowvt w=420000u l=150000u
+  ad=1.91777e+12p pd=1.512e+07u as=1.008e+11p ps=1.32e+06u
M1002 VPWR a_1271_74# a_1525_212# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.226e+11p ps=1.9e+06u
M1003 a_1271_74# a_493_387# a_837_359# VNB nlowvt w=740000u l=150000u
+  ad=4.58e+11p pd=3.28e+06u as=2.405e+11p ps=2.13e+06u
M1004 a_699_463# a_493_387# a_30_78# VPB pshort w=420000u l=180000u
+  ad=2.31e+11p pd=2.78e+06u as=2.289e+11p ps=2.77e+06u
M1005 VGND a_1525_212# a_1481_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_789_463# a_306_119# a_699_463# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 a_1271_74# a_306_119# a_837_359# VPB pshort w=1e+06u l=180000u
+  ad=4.32625e+11p pd=3.6e+06u as=0p ps=0u
M1008 a_895_138# a_837_359# a_817_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 a_1481_493# a_493_387# a_1271_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1010 a_1924_409# a_1271_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1011 VPWR a_837_359# a_789_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND RESET_B a_117_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_493_387# a_306_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.98825e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_30_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR RESET_B a_30_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND CLK a_306_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_699_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1525_212# a_1481_493# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1525_212# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1924_409# a_1271_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_1663_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 a_1525_212# a_1271_74# a_1663_81# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1023 a_837_359# a_699_463# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_817_138# a_493_387# a_699_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1025 VPWR CLK a_306_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1026 a_699_463# a_306_119# a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1027 a_493_387# a_306_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1028 a_117_78# D a_30_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_1924_409# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1030 VPWR a_1924_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q a_1924_409# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1032 a_1481_81# a_306_119# a_1271_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1924_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

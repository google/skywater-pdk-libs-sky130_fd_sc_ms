* File: sky130_fd_sc_ms__nand2_4.spice
* Created: Fri Aug 28 17:41:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand2_4.pex.spice"
.subckt sky130_fd_sc_ms__nand2_4  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_B_M1004_g N_A_27_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1004_d N_B_M1007_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_B_M1010_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1010_d N_B_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1184 PD=1.05 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75002
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_A_27_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_A_27_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15355 AS=0.1295 PD=1.155 PS=1.09 NRD=14.592 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_A_27_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15355 AS=0.2442 PD=1.155 PS=2.14 NRD=7.296 NRS=7.296 M=1 R=4.93333
+ SA=75003.5 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.6048
+ AS=0.3192 PD=2.2 PS=2.81 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90003.5
+ A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1001_d N_B_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12 AD=0.6048
+ AS=0.1792 PD=2.2 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5 SB=90002.2
+ A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1008_s N_A_M1000_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.1792
+ AS=0.7364 PD=1.44 PS=2.435 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002 SB=90001.7
+ A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.3696
+ AS=0.7364 PD=2.9 PS=2.435 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.4 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__nand2_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor2_4.pex.spice
* Created: Wed Sep  2 12:15:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR2_4%A 3 5 7 10 14 16 18 21 23 24 25 26 41
c71 21 0 9.54685e-20 $X=1.855 $Y=2.4
r72 41 42 6.73602 $w=3.22e-07 $l=4.5e-08 $layer=POLY_cond $X=1.81 $Y=1.385
+ $X2=1.855 $Y2=1.385
r73 39 41 26.9441 $w=3.22e-07 $l=1.8e-07 $layer=POLY_cond $X=1.63 $Y=1.385
+ $X2=1.81 $Y2=1.385
r74 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.385 $X2=1.63 $Y2=1.385
r75 37 39 33.6801 $w=3.22e-07 $l=2.25e-07 $layer=POLY_cond $X=1.405 $Y=1.385
+ $X2=1.63 $Y2=1.385
r76 36 37 67.3602 $w=3.22e-07 $l=4.5e-07 $layer=POLY_cond $X=0.955 $Y=1.385
+ $X2=1.405 $Y2=1.385
r77 34 36 51.6429 $w=3.22e-07 $l=3.45e-07 $layer=POLY_cond $X=0.61 $Y=1.385
+ $X2=0.955 $Y2=1.385
r78 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r79 32 34 13.472 $w=3.22e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.385 $X2=0.61
+ $Y2=1.385
r80 31 32 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.385
+ $X2=0.52 $Y2=1.385
r81 26 40 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.365 $X2=1.63
+ $Y2=1.365
r82 25 40 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=1.63 $Y2=1.365
r83 24 25 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=1.2 $Y2=1.365
r84 24 35 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r85 23 35 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r86 19 42 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.55
+ $X2=1.855 $Y2=1.385
r87 19 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.855 $Y=1.55
+ $X2=1.855 $Y2=2.4
r88 16 41 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.22
+ $X2=1.81 $Y2=1.385
r89 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.81 $Y=1.22 $X2=1.81
+ $Y2=0.74
r90 12 37 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.55
+ $X2=1.405 $Y2=1.385
r91 12 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.405 $Y=1.55
+ $X2=1.405 $Y2=2.4
r92 8 36 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=1.385
r93 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=2.4
r94 5 32 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=1.385
r95 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.22 $X2=0.52
+ $Y2=0.74
r96 1 31 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.385
r97 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_4%B 1 3 6 8 10 13 17 21 23 24 25 40
r66 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.385 $X2=4.01 $Y2=1.385
r67 38 40 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.755 $Y=1.385
+ $X2=4.01 $Y2=1.385
r68 36 38 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=3.33 $Y=1.385
+ $X2=3.755 $Y2=1.385
r69 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.385 $X2=3.33 $Y2=1.385
r70 34 36 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=1.385
+ $X2=3.33 $Y2=1.385
r71 33 34 87.4306 $w=3.3e-07 $l=5e-07 $layer=POLY_cond $X=2.755 $Y=1.385
+ $X2=3.255 $Y2=1.385
r72 32 33 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.74 $Y=1.385
+ $X2=2.755 $Y2=1.385
r73 31 32 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=2.305 $Y=1.385
+ $X2=2.74 $Y2=1.385
r74 29 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.29 $Y=1.385
+ $X2=2.305 $Y2=1.385
r75 25 41 2.1803 $w=3.68e-07 $l=7e-08 $layer=LI1_cond $X=4.08 $Y=1.365 $X2=4.01
+ $Y2=1.365
r76 24 41 12.7703 $w=3.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=4.01 $Y2=1.365
r77 24 37 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=3.33 $Y2=1.365
r78 23 37 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.33 $Y2=1.365
r79 19 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.55
+ $X2=3.755 $Y2=1.385
r80 19 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.755 $Y=1.55
+ $X2=3.755 $Y2=2.4
r81 15 34 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.55
+ $X2=3.255 $Y2=1.385
r82 15 17 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.255 $Y=1.55
+ $X2=3.255 $Y2=2.4
r83 11 33 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.55
+ $X2=2.755 $Y2=1.385
r84 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.755 $Y=1.55
+ $X2=2.755 $Y2=2.4
r85 8 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.22
+ $X2=2.74 $Y2=1.385
r86 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.74 $Y=1.22 $X2=2.74
+ $Y2=0.74
r87 4 31 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.55
+ $X2=2.305 $Y2=1.385
r88 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.305 $Y=1.55
+ $X2=2.305 $Y2=2.4
r89 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.22
+ $X2=2.29 $Y2=1.385
r90 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.29 $Y=1.22 $X2=2.29
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_4%A_27_368# 1 2 3 4 5 18 22 23 26 30 35 38 39
+ 42 46 50 54 55
r73 50 53 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=4.005 $Y=1.985
+ $X2=4.005 $Y2=2.815
r74 48 53 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=4.005 $Y=2.905
+ $X2=4.005 $Y2=2.815
r75 47 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=2.99
+ $X2=3.03 $Y2=2.99
r76 46 48 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.865 $Y=2.99
+ $X2=4.005 $Y2=2.905
r77 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.865 $Y=2.99
+ $X2=3.195 $Y2=2.99
r78 42 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.03 $Y=2.145
+ $X2=3.03 $Y2=2.825
r79 40 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.905
+ $X2=3.03 $Y2=2.99
r80 40 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.03 $Y=2.905 $X2=3.03
+ $Y2=2.825
r81 38 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=3.03 $Y2=2.99
r82 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=2.195 $Y2=2.99
r83 35 37 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.055 $Y=1.985
+ $X2=2.055 $Y2=2.815
r84 33 39 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.195 $Y2=2.99
r85 33 37 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.055 $Y2=2.815
r86 32 35 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.055 $Y=1.89
+ $X2=2.055 $Y2=1.985
r87 31 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=1.805
+ $X2=1.18 $Y2=1.805
r88 30 32 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.915 $Y=1.805
+ $X2=2.055 $Y2=1.89
r89 30 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.915 $Y=1.805
+ $X2=1.345 $Y2=1.805
r90 26 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.18 $Y=1.985
+ $X2=1.18 $Y2=2.815
r91 24 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=1.89 $X2=1.18
+ $Y2=1.805
r92 24 26 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.18 $Y=1.89
+ $X2=1.18 $Y2=1.985
r93 22 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=1.805
+ $X2=1.18 $Y2=1.805
r94 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.015 $Y=1.805
+ $X2=0.445 $Y2=1.805
r95 18 20 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r96 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.445 $Y2=1.805
r97 16 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.28 $Y2=1.985
r98 5 53 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.84 $X2=3.98 $Y2=2.815
r99 5 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.84 $X2=3.98 $Y2=1.985
r100 4 45 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=3.03 $Y2=2.825
r101 4 42 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=3.03 $Y2=2.145
r102 3 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.815
r103 3 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=1.985
r104 2 28 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r105 2 26 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r106 1 20 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r107 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_4%VPWR 1 2 11 15 17 19 26 27 30 33
r48 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.63 $Y2=3.33
r52 24 26 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r57 20 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.63 $Y2=3.33
r59 19 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 17 27 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 17 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r63 13 15 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.225
r64 9 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245 $X2=0.73
+ $Y2=3.33
r65 9 11 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.225
r66 2 15 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.225
r67 1 11 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_4%Y 1 2 3 4 13 17 21 23 24 27 31 35 41 42 43
c59 42 0 9.54685e-20 $X=2.53 $Y=1.805
r60 43 45 12.7875 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.557 $Y=1.295
+ $X2=2.557 $Y2=0.925
r61 40 41 9.36207 $w=6.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.595 $Y=0.675
+ $X2=1.69 $Y2=0.675
r62 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.53 $Y=1.97
+ $X2=3.53 $Y2=2.65
r63 33 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.53 $Y=1.89 $X2=3.53
+ $Y2=1.97
r64 32 42 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=1.805
+ $X2=2.53 $Y2=1.805
r65 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.365 $Y=1.805
+ $X2=3.53 $Y2=1.89
r66 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=1.805
+ $X2=2.695 $Y2=1.805
r67 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=1.97
+ $X2=2.53 $Y2=2.65
r68 25 42 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.89 $X2=2.53
+ $Y2=1.805
r69 25 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.53 $Y=1.89 $X2=2.53
+ $Y2=1.97
r70 24 42 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.72 $X2=2.53
+ $Y2=1.805
r71 23 43 4.04312 $w=3.53e-07 $l=1.27789e-07 $layer=LI1_cond $X=2.53 $Y=1.41
+ $X2=2.557 $Y2=1.295
r72 23 24 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.53 $Y=1.41 $X2=2.53
+ $Y2=1.72
r73 19 45 3.00629 $w=3.53e-07 $l=9.97246e-08 $layer=LI1_cond $X=2.525 $Y=0.84
+ $X2=2.557 $Y2=0.925
r74 19 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.525 $Y=0.84
+ $X2=2.525 $Y2=0.515
r75 17 45 5.025 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.36 $Y=0.925
+ $X2=2.557 $Y2=0.925
r76 17 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.36 $Y=0.925
+ $X2=1.69 $Y2=0.925
r77 13 40 4.28446 $w=6.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.355 $Y=0.675
+ $X2=1.595 $Y2=0.675
r78 13 15 3.65964 $w=6.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0.675
+ $X2=1.15 $Y2=0.675
r79 4 37 400 $w=1.7e-07 $l=8.97747e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.53 $Y2=2.65
r80 4 35 400 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.53 $Y2=1.97
r81 3 29 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.84 $X2=2.53 $Y2=2.65
r82 3 27 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.84 $X2=2.53 $Y2=1.97
r83 2 21 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.37 $X2=2.525 $Y2=0.515
r84 1 40 91 $w=1.7e-07 $l=1.06536e-06 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.37 $X2=1.595 $Y2=0.505
r85 1 15 45.5 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_NDIFF $count=4 $X=0.595
+ $Y=0.37 $X2=1.15 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_4%VGND 1 2 3 10 12 16 19 20 21 30 43 46
r34 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r35 43 45 0.477495 $w=1.022e-06 $l=4e-08 $layer=LI1_cond $X=4.04 $Y=0.462
+ $X2=4.08 $Y2=0.462
r36 41 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r37 40 43 10.9824 $w=1.022e-06 $l=9.2e-07 $layer=LI1_cond $X=3.12 $Y=0.462
+ $X2=4.04 $Y2=0.462
r38 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 38 40 1.96967 $w=1.022e-06 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0.462
+ $X2=3.12 $Y2=0.462
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r42 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 30 38 12.137 $w=1.022e-06 $l=5.07281e-07 $layer=LI1_cond $X=2.86 $Y=0
+ $X2=2.955 $Y2=0.462
r44 30 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.64
+ $Y2=0
r45 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r47 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r48 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r49 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 23 35 4.97422 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.235
+ $Y2=0
r51 23 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r52 21 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r53 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r54 19 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r55 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.025
+ $Y2=0
r56 18 32 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.64
+ $Y2=0
r57 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.025
+ $Y2=0
r58 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r59 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.55
r60 10 35 3.0057 $w=3.55e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.292 $Y=0.085
+ $X2=0.235 $Y2=0
r61 10 12 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=0.292 $Y=0.085
+ $X2=0.292 $Y2=0.515
r62 3 43 60.6667 $w=1.7e-07 $l=1.29074e-06 $layer=licon1_NDIFF $count=3 $X=2.815
+ $Y=0.37 $X2=4.04 $Y2=0.505
r63 3 38 60.6667 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=3 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.505
r64 2 16 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.885 $Y=0.37
+ $X2=2.025 $Y2=0.55
r65 1 12 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.305 $Y2=0.515
.ends


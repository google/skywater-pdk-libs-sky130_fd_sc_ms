* File: sky130_fd_sc_ms__sdlclkp_4.pex.spice
* Created: Fri Aug 28 18:15:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%SCE 3 7 9 12 13
r26 12 15 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.62
+ $X2=0.407 $Y2=1.785
r27 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.62
+ $X2=0.407 $Y2=1.455
r28 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.62 $X2=0.385 $Y2=1.62
r29 9 13 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.62
+ $X2=0.385 $Y2=1.62
r30 7 14 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=0.99
+ $X2=0.52 $Y2=1.455
r31 3 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.505 $Y=2.395
+ $X2=0.505 $Y2=1.785
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%GATE 3 7 9 12
c35 9 0 1.03187e-19 $X=1.2 $Y=1.665
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.62 $X2=1
+ $Y2=1.785
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.62 $X2=1
+ $Y2=1.455
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.62
+ $X2=1 $Y2=1.62
r39 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.62 $X2=1
+ $Y2=1.62
r40 7 14 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.995 $Y=0.99
+ $X2=0.995 $Y2=1.455
r41 3 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=2.395
+ $X2=0.925 $Y2=1.785
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%A_354_105# 1 2 9 11 15 19 21 22 25 27 29
+ 31 39
c78 39 0 1.84961e-19 $X=3.405 $Y=1.57
c79 31 0 8.43768e-20 $X=3.09 $Y=1.57
c80 29 0 3.22822e-20 $X=2.53 $Y=1.65
c81 15 0 1.62426e-20 $X=3.645 $Y=0.58
r82 38 39 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.315 $Y=1.57
+ $X2=3.405 $Y2=1.57
r83 32 38 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.09 $Y=1.57
+ $X2=3.315 $Y2=1.57
r84 31 34 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.09 $Y=1.57 $X2=3.09
+ $Y2=1.65
r85 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.57 $X2=3.09 $Y2=1.57
r86 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=1.65
+ $X2=2.53 $Y2=1.65
r87 27 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=1.65
+ $X2=3.09 $Y2=1.65
r88 27 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.925 $Y=1.65
+ $X2=2.695 $Y2=1.65
r89 23 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.735
+ $X2=2.53 $Y2=1.65
r90 23 25 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.53 $Y=1.735
+ $X2=2.53 $Y2=1.975
r91 21 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=1.65
+ $X2=2.53 $Y2=1.65
r92 21 22 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.365 $Y=1.65
+ $X2=2.075 $Y2=1.65
r93 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.95 $Y=1.565
+ $X2=2.075 $Y2=1.65
r94 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.95 $Y=1.565
+ $X2=1.95 $Y2=1.12
r95 13 15 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.645 $Y=1.405
+ $X2=3.645 $Y2=0.58
r96 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.57 $Y=1.48
+ $X2=3.645 $Y2=1.405
r97 11 39 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.48
+ $X2=3.405 $Y2=1.48
r98 7 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.735
+ $X2=3.315 $Y2=1.57
r99 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.315 $Y=1.735
+ $X2=3.315 $Y2=2.315
r100 2 25 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=2.12 $X2=2.53 $Y2=1.975
r101 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.525 $X2=1.91 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%A_324_79# 1 2 7 9 10 11 15 16 17 18 20 22
+ 25 27 30 31 32 34 35 36 38 39 40 44 47 54 55 57 58
c154 44 0 1.46172e-19 $X=5.67 $Y=0.515
c155 39 0 9.27061e-20 $X=5.445 $Y=0.34
c156 35 0 6.61483e-20 $X=4.605 $Y=0.98
c157 30 0 1.62426e-20 $X=2.89 $Y=1.065
c158 27 0 1.84961e-19 $X=2.805 $Y=1.15
c159 15 0 8.43768e-20 $X=2.22 $Y=2.54
c160 11 0 1.84401e-19 $X=1.77 $Y=1.415
r161 55 57 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.53 $Y=1.82
+ $X2=5.53 $Y2=1.01
r162 54 55 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.607 $Y=1.985
+ $X2=5.607 $Y2=1.82
r163 51 58 13.7476 $w=4.45e-07 $l=1.1e-07 $layer=POLY_cond $X=2.352 $Y=1.23
+ $X2=2.352 $Y2=1.12
r164 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.23 $X2=2.41 $Y2=1.23
r165 47 50 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.41 $Y=1.15 $X2=2.41
+ $Y2=1.23
r166 42 57 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=5.64 $Y=0.815
+ $X2=5.64 $Y2=1.01
r167 42 44 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=5.64 $Y=0.815
+ $X2=5.64 $Y2=0.515
r168 41 44 2.65948 $w=3.88e-07 $l=9e-08 $layer=LI1_cond $X=5.64 $Y=0.425
+ $X2=5.64 $Y2=0.515
r169 39 41 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=5.64 $Y2=0.425
r170 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=4.775 $Y2=0.34
r171 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.69 $Y=0.425
+ $X2=4.775 $Y2=0.34
r172 37 38 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.69 $Y=0.425
+ $X2=4.69 $Y2=0.895
r173 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.605 $Y=0.98
+ $X2=4.69 $Y2=0.895
r174 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.605 $Y=0.98
+ $X2=3.935 $Y2=0.98
r175 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.85 $Y=0.895
+ $X2=3.935 $Y2=0.98
r176 33 34 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.85 $Y=0.44
+ $X2=3.85 $Y2=0.895
r177 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=0.355
+ $X2=3.85 $Y2=0.44
r178 31 32 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.765 $Y=0.355
+ $X2=2.975 $Y2=0.355
r179 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.89 $Y=0.44
+ $X2=2.975 $Y2=0.355
r180 29 30 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.89 $Y=0.44
+ $X2=2.89 $Y2=1.065
r181 28 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=1.15
+ $X2=2.41 $Y2=1.15
r182 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=1.15
+ $X2=2.89 $Y2=1.065
r183 27 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.805 $Y=1.15
+ $X2=2.575 $Y2=1.15
r184 23 25 229.339 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=3.85 $Y=3.075
+ $X2=3.85 $Y2=2.485
r185 20 22 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.095 $Y=1.045
+ $X2=3.095 $Y2=0.645
r186 19 58 28.4889 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.575 $Y=1.12
+ $X2=2.352 $Y2=1.12
r187 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.02 $Y=1.12
+ $X2=3.095 $Y2=1.045
r188 18 19 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.02 $Y=1.12
+ $X2=2.575 $Y2=1.12
r189 16 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.76 $Y=3.15
+ $X2=3.85 $Y2=3.075
r190 16 17 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=3.76 $Y=3.15
+ $X2=2.31 $Y2=3.15
r191 15 62 408.145 $w=1.8e-07 $l=1.05e-06 $layer=POLY_cond $X=2.22 $Y=2.54
+ $X2=2.22 $Y2=1.49
r192 13 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.22 $Y=3.075
+ $X2=2.31 $Y2=3.15
r193 13 15 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=2.22 $Y=3.075
+ $X2=2.22 $Y2=2.54
r194 10 62 29.7069 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=2.352 $Y=1.415
+ $X2=2.352 $Y2=1.49
r195 10 51 23.121 $w=4.45e-07 $l=1.85e-07 $layer=POLY_cond $X=2.352 $Y=1.415
+ $X2=2.352 $Y2=1.23
r196 10 11 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.13 $Y=1.415
+ $X2=1.77 $Y2=1.415
r197 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.695 $Y=1.34
+ $X2=1.77 $Y2=1.415
r198 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.695 $Y=1.34
+ $X2=1.695 $Y2=0.895
r199 2 54 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.84 $X2=5.605 $Y2=1.985
r200 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.525
+ $Y=0.37 $X2=5.67 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%A_792_48# 1 2 9 13 17 21 23 26 29 32 33 36
+ 37 39 43 49 50 52 58 63
c129 63 0 1.06371e-19 $X=7.015 $Y=1.465
c130 23 0 6.61483e-20 $X=4.88 $Y=1.82
c131 9 0 1.23505e-19 $X=4.035 $Y=0.58
r132 52 54 10.9068 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.11 $Y=0.83
+ $X2=5.11 $Y2=1.065
r133 44 58 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.125 $Y=1.74
+ $X2=4.27 $Y2=1.74
r134 44 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.125 $Y=1.74
+ $X2=4.035 $Y2=1.74
r135 43 46 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.125 $Y=1.74
+ $X2=4.125 $Y2=1.82
r136 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.125
+ $Y=1.74 $X2=4.125 $Y2=1.74
r137 40 63 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=6.865 $Y=1.465
+ $X2=7.015 $Y2=1.465
r138 40 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.865 $Y=1.465
+ $X2=6.775 $Y2=1.465
r139 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.865
+ $Y=1.465 $X2=6.865 $Y2=1.465
r140 37 39 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.455 $Y=1.465
+ $X2=6.865 $Y2=1.465
r141 35 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.37 $Y=1.63
+ $X2=6.455 $Y2=1.465
r142 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.37 $Y=1.63
+ $X2=6.37 $Y2=2.24
r143 34 50 4.4465 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.27 $Y=2.325
+ $X2=5.075 $Y2=2.325
r144 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.285 $Y=2.325
+ $X2=6.37 $Y2=2.24
r145 33 34 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=6.285 $Y=2.325
+ $X2=5.27 $Y2=2.325
r146 32 49 3.351 $w=2.8e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.185 $Y=1.735
+ $X2=5.075 $Y2=1.82
r147 32 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.185 $Y=1.735
+ $X2=5.185 $Y2=1.065
r148 27 50 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=2.41
+ $X2=5.075 $Y2=2.325
r149 27 29 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=5.075 $Y=2.41
+ $X2=5.075 $Y2=2.73
r150 26 50 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=2.24
+ $X2=5.075 $Y2=2.325
r151 25 49 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=1.905
+ $X2=5.075 $Y2=1.82
r152 25 26 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=5.075 $Y=1.905
+ $X2=5.075 $Y2=2.24
r153 24 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=1.82
+ $X2=4.125 $Y2=1.82
r154 23 49 3.18746 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.88 $Y=1.82
+ $X2=5.075 $Y2=1.82
r155 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.88 $Y=1.82
+ $X2=4.29 $Y2=1.82
r156 19 63 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.015 $Y=1.63
+ $X2=7.015 $Y2=1.465
r157 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.015 $Y=1.63
+ $X2=7.015 $Y2=2.4
r158 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.775 $Y=1.3
+ $X2=6.775 $Y2=1.465
r159 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.775 $Y=1.3
+ $X2=6.775 $Y2=0.74
r160 11 58 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.905
+ $X2=4.27 $Y2=1.74
r161 11 13 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.27 $Y=1.905
+ $X2=4.27 $Y2=2.485
r162 7 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.035 $Y=1.575
+ $X2=4.035 $Y2=1.74
r163 7 9 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=4.035 $Y=1.575
+ $X2=4.035 $Y2=0.58
r164 2 49 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.755 $X2=5.045 $Y2=1.9
r165 2 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.755 $X2=5.045 $Y2=2.73
r166 1 52 182 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.37 $X2=5.11 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%A_634_74# 1 2 9 13 15 18 22 27 29 30 34 37
c78 27 0 1.23505e-19 $X=3.51 $Y=0.775
r79 34 38 40.9837 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.4
+ $X2=4.785 $Y2=1.565
r80 34 37 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.4
+ $X2=4.785 $Y2=1.235
r81 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.765
+ $Y=1.4 $X2=4.765 $Y2=1.4
r82 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.765 $Y=1.32 $X2=4.765
+ $Y2=1.4
r83 25 27 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.33 $Y=0.775
+ $X2=3.51 $Y2=0.775
r84 23 29 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.705 $Y=1.32
+ $X2=3.565 $Y2=1.32
r85 22 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=1.32
+ $X2=4.765 $Y2=1.32
r86 22 23 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=4.6 $Y=1.32
+ $X2=3.705 $Y2=1.32
r87 18 20 21.4025 $w=2.78e-07 $l=5.2e-07 $layer=LI1_cond $X=3.565 $Y=2.07
+ $X2=3.565 $Y2=2.59
r88 16 29 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=1.405
+ $X2=3.565 $Y2=1.32
r89 16 18 27.3705 $w=2.78e-07 $l=6.65e-07 $layer=LI1_cond $X=3.565 $Y=1.405
+ $X2=3.565 $Y2=2.07
r90 15 29 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=3.51 $Y=1.235
+ $X2=3.565 $Y2=1.32
r91 14 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=0.94
+ $X2=3.51 $Y2=0.775
r92 14 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.51 $Y=0.94
+ $X2=3.51 $Y2=1.235
r93 13 37 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.895 $Y=0.74
+ $X2=4.895 $Y2=1.235
r94 9 38 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.82 $Y=2.315
+ $X2=4.82 $Y2=1.565
r95 2 20 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.895 $X2=3.54 $Y2=2.59
r96 2 18 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.895 $X2=3.54 $Y2=2.07
r97 1 25 182 $w=1.7e-07 $l=4.78357e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.37 $X2=3.33 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%CLK 3 5 7 10 12 14 15 24
c55 15 0 1.06371e-19 $X=6 $Y=1.295
c56 12 0 2.38878e-19 $X=6.385 $Y=1.22
r57 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.37 $Y=1.385
+ $X2=6.385 $Y2=1.385
r58 21 23 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.95 $Y=1.385
+ $X2=6.37 $Y2=1.385
r59 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.385 $X2=5.95 $Y2=1.385
r60 19 21 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=5.885 $Y=1.385
+ $X2=5.95 $Y2=1.385
r61 17 19 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=5.835 $Y=1.385
+ $X2=5.885 $Y2=1.385
r62 15 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.95 $Y=1.295 $X2=5.95
+ $Y2=1.385
r63 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.385 $Y=1.22
+ $X2=6.385 $Y2=1.385
r64 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.385 $Y=1.22
+ $X2=6.385 $Y2=0.74
r65 8 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=1.55
+ $X2=6.37 $Y2=1.385
r66 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.37 $Y=1.55 $X2=6.37
+ $Y2=2.4
r67 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.22
+ $X2=5.885 $Y2=1.385
r68 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.885 $Y=1.22 $X2=5.885
+ $Y2=0.74
r69 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.55
+ $X2=5.835 $Y2=1.385
r70 1 3 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=5.835 $Y=1.55
+ $X2=5.835 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%A_1292_368# 1 2 9 13 17 21 25 29 33 37 41
+ 47 49 50 51 52 54 56 62 65 76
c127 37 0 1.19111e-20 $X=9.105 $Y=0.74
r128 75 76 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.09 $Y=1.465
+ $X2=9.105 $Y2=1.465
r129 74 75 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.675 $Y=1.465
+ $X2=9.09 $Y2=1.465
r130 73 74 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=8.595 $Y=1.465
+ $X2=8.675 $Y2=1.465
r131 70 71 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=8.095 $Y=1.465
+ $X2=8.245 $Y2=1.465
r132 69 70 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=7.765 $Y=1.465
+ $X2=8.095 $Y2=1.465
r133 63 73 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=8.27 $Y=1.465
+ $X2=8.595 $Y2=1.465
r134 63 71 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=8.27 $Y=1.465
+ $X2=8.245 $Y2=1.465
r135 62 63 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.27
+ $Y=1.465 $X2=8.27 $Y2=1.465
r136 60 69 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.59 $Y=1.465
+ $X2=7.765 $Y2=1.465
r137 60 66 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.59 $Y=1.465
+ $X2=7.515 $Y2=1.465
r138 59 62 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.59 $Y=1.465
+ $X2=8.27 $Y2=1.465
r139 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.59
+ $Y=1.465 $X2=7.59 $Y2=1.465
r140 57 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.535 $Y=1.465
+ $X2=7.45 $Y2=1.465
r141 57 59 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=7.535 $Y=1.465
+ $X2=7.59 $Y2=1.465
r142 55 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=1.63
+ $X2=7.45 $Y2=1.465
r143 55 56 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.45 $Y=1.63
+ $X2=7.45 $Y2=1.8
r144 54 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=1.3
+ $X2=7.45 $Y2=1.465
r145 53 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.45 $Y=1.13
+ $X2=7.45 $Y2=1.3
r146 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.045
+ $X2=7.45 $Y2=1.13
r147 51 52 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.365 $Y=1.045
+ $X2=7.155 $Y2=1.045
r148 49 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.885
+ $X2=7.45 $Y2=1.8
r149 49 50 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.365 $Y=1.885
+ $X2=6.955 $Y2=1.885
r150 45 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.99 $Y=0.96
+ $X2=7.155 $Y2=1.045
r151 45 47 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.99 $Y=0.96
+ $X2=6.99 $Y2=0.515
r152 41 43 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.79 $Y=1.985
+ $X2=6.79 $Y2=2.815
r153 39 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.79 $Y=1.97
+ $X2=6.955 $Y2=1.885
r154 39 41 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.79 $Y=1.97
+ $X2=6.79 $Y2=1.985
r155 35 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=9.105 $Y2=1.465
r156 35 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.105 $Y=1.3
+ $X2=9.105 $Y2=0.74
r157 31 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.09 $Y=1.63
+ $X2=9.09 $Y2=1.465
r158 31 33 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=9.09 $Y=1.63
+ $X2=9.09 $Y2=2.4
r159 27 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=1.465
r160 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.675 $Y=1.3
+ $X2=8.675 $Y2=0.74
r161 23 73 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.595 $Y=1.63
+ $X2=8.595 $Y2=1.465
r162 23 25 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.595 $Y=1.63
+ $X2=8.595 $Y2=2.4
r163 19 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=1.465
r164 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.245 $Y=1.3
+ $X2=8.245 $Y2=0.74
r165 15 70 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.63
+ $X2=8.095 $Y2=1.465
r166 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.095 $Y=1.63
+ $X2=8.095 $Y2=2.4
r167 11 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=1.465
r168 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.765 $Y=1.3
+ $X2=7.765 $Y2=0.74
r169 7 66 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.515 $Y=1.63
+ $X2=7.515 $Y2=1.465
r170 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.515 $Y=1.63
+ $X2=7.515 $Y2=2.4
r171 2 43 400 $w=1.7e-07 $l=1.128e-06 $layer=licon1_PDIFF $count=1 $X=6.46
+ $Y=1.84 $X2=6.79 $Y2=2.815
r172 2 41 400 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=1 $X=6.46
+ $Y=1.84 $X2=6.79 $Y2=1.985
r173 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.85
+ $Y=0.37 $X2=6.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%VPWR 1 2 3 4 5 6 7 22 24 28 34 38 42 44 46
+ 51 52 53 55 60 68 77 81 90 97 100 103 107
r105 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r106 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r107 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r108 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r110 85 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r111 85 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r112 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r113 82 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.36 $Y2=3.33
r114 82 84 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 81 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.155 $Y=3.33
+ $X2=9.377 $Y2=3.33
r116 81 84 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.155 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 80 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r118 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r119 77 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.36 $Y2=3.33
r120 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 76 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6 $Y2=3.33
r123 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 73 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.31 $Y=3.33
+ $X2=6.145 $Y2=3.33
r125 73 75 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.31 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 72 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r127 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r128 69 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=4.555 $Y2=3.33
r129 69 71 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=5.04 $Y2=3.33
r130 68 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=6.145 $Y2=3.33
r131 68 71 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 67 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r133 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 64 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 60 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.555 $Y2=3.33
r139 60 66 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r140 59 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r141 59 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r143 56 87 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r144 56 58 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r145 55 63 8.47627 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=1.852 $Y=3.33
+ $X2=2.16 $Y2=3.33
r146 55 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r147 55 90 10.7939 $w=6.13e-07 $l=5.55e-07 $layer=LI1_cond $X=1.852 $Y=3.33
+ $X2=1.852 $Y2=2.775
r148 55 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r149 53 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r150 53 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 51 75 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=3.33
+ $X2=6.96 $Y2=3.33
r152 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=3.33
+ $X2=7.29 $Y2=3.33
r153 50 79 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.92 $Y2=3.33
r154 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.29 $Y2=3.33
r155 46 49 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.32 $Y=1.985
+ $X2=9.32 $Y2=2.815
r156 44 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.32 $Y=3.245
+ $X2=9.377 $Y2=3.33
r157 44 49 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.32 $Y=3.245
+ $X2=9.32 $Y2=2.815
r158 40 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=3.33
r159 40 42 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.305
r160 36 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.29 $Y=3.245
+ $X2=7.29 $Y2=3.33
r161 36 38 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=7.29 $Y=3.245
+ $X2=7.29 $Y2=2.305
r162 32 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.145 $Y=3.245
+ $X2=6.145 $Y2=3.33
r163 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.145 $Y=3.245
+ $X2=6.145 $Y2=2.745
r164 28 31 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=4.555 $Y=2.24
+ $X2=4.555 $Y2=2.73
r165 26 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=3.33
r166 26 31 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=2.73
r167 22 87 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r168 22 24 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.12
r169 7 49 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=9.18
+ $Y=1.84 $X2=9.32 $Y2=2.815
r170 7 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.18
+ $Y=1.84 $X2=9.32 $Y2=1.985
r171 6 42 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=8.185
+ $Y=1.84 $X2=8.32 $Y2=2.305
r172 5 38 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=7.105
+ $Y=1.84 $X2=7.29 $Y2=2.305
r173 4 34 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=5.925
+ $Y=1.84 $X2=6.145 $Y2=2.745
r174 3 31 600 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.275 $X2=4.595 $Y2=2.73
r175 3 28 600 $w=1.7e-07 $l=2.51893e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.275 $X2=4.595 $Y2=2.24
r176 2 90 600 $w=1.7e-07 $l=8.41071e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=2.12 $X2=1.99 $Y2=2.775
r177 1 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.975 $X2=0.28 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%A_119_143# 1 2 3 4 15 17 18 22 25 29 32 35
+ 36 38 39
c95 38 0 3.22822e-20 $X=2.525 $Y=0.62
c96 35 0 8.1214e-20 $X=1.655 $Y=2.217
r97 38 39 11.007 $w=5.43e-07 $l=2.2e-07 $layer=LI1_cond $X=2.525 $Y=0.622
+ $X2=2.305 $Y2=0.622
r98 27 29 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.09 $Y=2.31 $X2=3.09
+ $Y2=2.07
r99 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.925 $Y=2.395
+ $X2=3.09 $Y2=2.31
r100 25 35 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=2.925 $Y=2.395
+ $X2=1.655 $Y2=2.395
r101 24 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.7
+ $X2=1.57 $Y2=0.7
r102 24 39 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.655 $Y=0.7
+ $X2=2.305 $Y2=0.7
r103 22 35 7.85017 $w=5.23e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.217
+ $X2=1.655 $Y2=2.217
r104 22 32 9.56863 $w=5.23e-07 $l=4.2e-07 $layer=LI1_cond $X=1.57 $Y=2.217
+ $X2=1.15 $Y2=2.217
r105 21 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.785
+ $X2=1.57 $Y2=0.7
r106 21 22 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=1.57 $Y=0.785
+ $X2=1.57 $Y2=1.955
r107 17 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=0.7
+ $X2=1.57 $Y2=0.7
r108 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.485 $Y=0.7
+ $X2=0.945 $Y2=0.7
r109 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.785
+ $X2=0.945 $Y2=0.7
r110 13 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.78 $Y=0.785
+ $X2=0.78 $Y2=0.99
r111 4 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=2.945
+ $Y=1.895 $X2=3.09 $Y2=2.07
r112 3 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.015
+ $Y=1.975 $X2=1.15 $Y2=2.12
r113 2 38 182 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.37 $X2=2.525 $Y2=0.62
r114 1 15 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.715 $X2=0.78 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%GCLK 1 2 3 4 15 21 23 24 25 26 29 35 38 39
+ 40 42
c70 25 0 1.19111e-20 $X=8.725 $Y=1.045
r71 40 45 4.56667 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.89 $Y=1.295
+ $X2=8.89 $Y2=1.41
r72 40 42 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.89 $Y=1.295
+ $X2=8.89 $Y2=1.045
r73 38 39 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=8.855 $Y=1.8
+ $X2=8.82 $Y2=1.885
r74 38 45 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=8.855 $Y=1.8
+ $X2=8.855 $Y2=1.41
r75 33 42 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=0.96
+ $X2=8.89 $Y2=1.045
r76 33 35 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.89 $Y=0.96
+ $X2=8.89 $Y2=0.515
r77 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.82 $Y=1.985
+ $X2=8.82 $Y2=2.815
r78 27 39 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=1.97
+ $X2=8.82 $Y2=1.885
r79 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.82 $Y=1.97
+ $X2=8.82 $Y2=1.985
r80 25 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=1.045
+ $X2=8.89 $Y2=1.045
r81 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.725 $Y=1.045
+ $X2=8.115 $Y2=1.045
r82 23 39 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.655 $Y=1.885
+ $X2=8.82 $Y2=1.885
r83 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.655 $Y=1.885
+ $X2=8.035 $Y2=1.885
r84 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.99 $Y=0.96
+ $X2=8.115 $Y2=1.045
r85 19 21 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=7.99 $Y=0.96
+ $X2=7.99 $Y2=0.515
r86 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.87 $Y=1.985
+ $X2=7.87 $Y2=2.815
r87 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.87 $Y=1.97
+ $X2=8.035 $Y2=1.885
r88 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.87 $Y=1.97
+ $X2=7.87 $Y2=1.985
r89 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.685
+ $Y=1.84 $X2=8.82 $Y2=2.815
r90 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.685
+ $Y=1.84 $X2=8.82 $Y2=1.985
r91 3 17 400 $w=1.7e-07 $l=1.09955e-06 $layer=licon1_PDIFF $count=1 $X=7.605
+ $Y=1.84 $X2=7.87 $Y2=2.815
r92 3 15 400 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=7.605
+ $Y=1.84 $X2=7.87 $Y2=1.985
r93 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.515
r94 1 21 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=7.84
+ $Y=0.37 $X2=8.03 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_4%VGND 1 2 3 4 5 6 7 22 24 26 30 34 38 42 44
+ 46 49 50 52 53 54 69 73 78 88 94 97 101
r120 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r121 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r122 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r123 88 91 7.33373 $w=4.38e-07 $l=2.8e-07 $layer=LI1_cond $X=1.345 $Y=0
+ $X2=1.345 $Y2=0.28
r124 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r126 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r128 82 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r129 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r130 79 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=0 $X2=8.42
+ $Y2=0
r131 79 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.545 $Y=0
+ $X2=8.88 $Y2=0
r132 78 100 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.235 $Y=0
+ $X2=9.417 $Y2=0
r133 78 81 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.235 $Y=0
+ $X2=8.88 $Y2=0
r134 77 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r135 77 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r136 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r137 74 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.635 $Y=0 $X2=7.51
+ $Y2=0
r138 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.635 $Y=0
+ $X2=7.92 $Y2=0
r139 73 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=0 $X2=8.42
+ $Y2=0
r140 73 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=7.92 $Y2=0
r141 72 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r142 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r143 69 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.385 $Y=0 $X2=7.51
+ $Y2=0
r144 69 71 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.385 $Y=0
+ $X2=6.48 $Y2=0
r145 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r146 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r147 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r148 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r149 62 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r150 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r151 59 62 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=4.08
+ $Y2=0
r152 59 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r153 58 61 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=4.08
+ $Y2=0
r154 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r155 56 88 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.345
+ $Y2=0
r156 56 58 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=0
+ $X2=1.68 $Y2=0
r157 54 68 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6
+ $Y2=0
r158 54 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r159 52 67 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.005 $Y=0 $X2=6
+ $Y2=0
r160 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.005 $Y=0 $X2=6.17
+ $Y2=0
r161 51 71 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.48 $Y2=0
r162 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.17
+ $Y2=0
r163 49 61 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.08
+ $Y2=0
r164 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.27
+ $Y2=0
r165 48 64 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.56 $Y2=0
r166 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.27
+ $Y2=0
r167 44 100 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.417 $Y2=0
r168 44 46 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.36 $Y2=0.515
r169 40 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r170 40 42 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.57
r171 36 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0
r172 36 38 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0.57
r173 32 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=0.085
+ $X2=6.17 $Y2=0
r174 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.17 $Y=0.085
+ $X2=6.17 $Y2=0.515
r175 28 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r176 28 30 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.535
r177 27 84 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r178 26 88 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.345
+ $Y2=0
r179 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=0
+ $X2=0.445 $Y2=0
r180 22 84 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r181 22 24 31.6049 $w=3.28e-07 $l=9.05e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.99
r182 7 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.18
+ $Y=0.37 $X2=9.32 $Y2=0.515
r183 6 42 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=8.32
+ $Y=0.37 $X2=8.46 $Y2=0.57
r184 5 38 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=7.405
+ $Y=0.37 $X2=7.55 $Y2=0.57
r185 4 34 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.96
+ $Y=0.37 $X2=6.17 $Y2=0.515
r186 3 30 182 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=1 $X=4.11
+ $Y=0.37 $X2=4.27 $Y2=0.535
r187 2 91 182 $w=1.7e-07 $l=5.55743e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.715 $X2=1.345 $Y2=0.28
r188 1 24 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.715 $X2=0.28 $Y2=0.99
.ends


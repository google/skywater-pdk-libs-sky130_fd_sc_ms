* File: sky130_fd_sc_ms__xnor2_2.spice
* Created: Wed Sep  2 12:33:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xnor2_2.pex.spice"
.subckt sky130_fd_sc_ms__xnor2_2  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1014 A_151_74# N_A_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.25 PD=0.98 PS=2.44 NRD=10.536 NRS=21.888 M=1 R=4.93333 SA=75000.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_136_368#_M1013_d N_B_M1013_g A_151_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.206875 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A_136_368#_M1004_g N_A_340_107#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2004 AS=0.197775 PD=1.335 PS=2.05 NRD=17.832 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1004_d N_A_136_368#_M1015_g N_A_340_107#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2004 AS=0.1036 PD=1.335 PS=1.02 NRD=18.648 NRS=0 M=1 R=4.93333
+ SA=75000.8 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_340_107#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1912 AS=0.1036 PD=1.365 PS=1.02 NRD=32.976 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1001 N_A_340_107#_M1001_d N_B_M1001_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1912 PD=1.04 PS=1.365 NRD=0 NRS=32.976 M=1 R=4.93333 SA=75001.9
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1005 N_A_340_107#_M1001_d N_B_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1958 PD=1.04 PS=1.375 NRD=0 NRS=33.984 M=1 R=4.93333 SA=75002.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1005_s N_A_M1007_g N_A_340_107#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1958 AS=0.20355 PD=1.375 PS=2.05 NRD=33.984 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_136_368#_M1011_d N_A_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.1575 AS=0.4027 PD=1.315 PS=2.99 NRD=2.9353 NRS=16.7253 M=1 R=5.55556
+ SA=90000.3 SB=90004.3 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_B_M1012_g N_A_136_368#_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.410684 AS=0.1575 PD=1.80189 PS=1.315 NRD=12.805 NRS=3.9203 M=1 R=5.55556
+ SA=90000.8 SB=90003.8 A=0.18 P=2.36 MULT=1
MM1009 N_Y_M1009_d N_A_136_368#_M1009_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.459966 PD=1.39 PS=2.01811 NRD=0 NRS=4.3931 M=1 R=6.22222
+ SA=90001.6 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1009_d N_A_136_368#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.25945 PD=1.39 PS=1.65 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90002.1 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1010_s N_A_M1002_g N_A_641_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.25945 AS=0.2655 PD=1.65 PS=1.66 NRD=14.9326 NRS=15.8191 M=1 R=6.22222
+ SA=90002.7 SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_A_641_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2655 PD=1.39 PS=1.66 NRD=0 NRS=15.8191 M=1 R=6.22222 SA=90003.3
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1000_d N_B_M1003_g N_A_641_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.8
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_A_641_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1792 PD=2.9 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90004.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ms__xnor2_2.pxi.spice"
*
.ends
*
*

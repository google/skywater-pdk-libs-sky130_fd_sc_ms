* File: sky130_fd_sc_ms__sdfrbp_2.pex.spice
* Created: Wed Sep  2 12:30:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%SCE 2 5 7 9 10 12 16 20 23 25 26 28 29 31
+ 32 33 38 48
r88 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.985 $X2=1.385 $Y2=1.985
r89 38 43 10.6155 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.37 $Y=1.985 $X2=1.46
+ $Y2=1.985
r90 38 40 116.283 $w=3.3e-07 $l=6.65e-07 $layer=POLY_cond $X=1.37 $Y=1.985
+ $X2=0.705 $Y2=1.985
r91 33 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.985
+ $X2=1.625 $Y2=1.985
r92 33 48 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.61 $Y=1.985
+ $X2=1.625 $Y2=1.985
r93 33 44 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=1.985
+ $X2=1.385 $Y2=1.985
r94 32 44 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.385 $Y2=1.985
r95 31 32 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.705 $Y=1.985
+ $X2=1.2 $Y2=1.985
r96 31 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.985 $X2=0.705 $Y2=1.985
r97 29 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.455
+ $X2=2.57 $Y2=1.29
r98 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.455 $X2=2.57 $Y2=1.455
r99 26 28 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=1.795 $Y=1.49
+ $X2=2.57 $Y2=1.49
r100 25 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=1.82
+ $X2=1.71 $Y2=1.985
r101 24 26 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.71 $Y=1.62
+ $X2=1.795 $Y2=1.49
r102 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.71 $Y=1.62 $X2=1.71
+ $Y2=1.82
r103 22 40 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.595 $Y=1.985
+ $X2=0.705 $Y2=1.985
r104 22 23 3.90195 $w=3.3e-07 $l=3.32415e-07 $layer=POLY_cond $X=0.595 $Y=1.985
+ $X2=0.335 $Y2=1.82
r105 18 20 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=0.965
+ $X2=0.495 $Y2=0.965
r106 16 46 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.66 $Y=0.605
+ $X2=2.66 $Y2=1.29
r107 10 43 19.4618 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=2.15
+ $X2=1.46 $Y2=1.985
r108 10 12 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=1.46 $Y=2.15
+ $X2=1.46 $Y2=2.64
r109 7 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.965
r110 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.605
r111 3 23 34.7346 $w=1.65e-07 $l=4.06202e-07 $layer=POLY_cond $X=0.505 $Y=2.15
+ $X2=0.335 $Y2=1.82
r112 3 5 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=0.505 $Y=2.15
+ $X2=0.505 $Y2=2.64
r113 2 23 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.41 $Y=1.82
+ $X2=0.335 $Y2=1.82
r114 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.41 $Y=1.04
+ $X2=0.41 $Y2=0.965
r115 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.41 $Y=1.04 $X2=0.41
+ $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_27_79# 1 2 9 13 15 18 21 24 28 31 35 38
+ 39 44
c85 31 0 1.3564e-19 $X=2.275 $Y=2.405
r86 36 44 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.44 $Y=1.995
+ $X2=2.615 $Y2=1.995
r87 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.995 $X2=2.44 $Y2=1.995
r88 33 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.44 $Y=2.32
+ $X2=2.44 $Y2=1.995
r89 32 39 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.28 $Y2=2.405
r90 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=2.44 $Y2=2.32
r91 31 32 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=0.445 $Y2=2.405
r92 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.415 $X2=1.23 $Y2=1.415
r93 26 38 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.415
+ $X2=0.24 $Y2=1.415
r94 26 28 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.365 $Y=1.415
+ $X2=1.23 $Y2=1.415
r95 22 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.49 $X2=0.28
+ $Y2=2.405
r96 22 24 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.28 $Y=2.49 $X2=0.28
+ $Y2=2.65
r97 21 39 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.32
+ $X2=0.28 $Y2=2.405
r98 20 38 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.58
+ $X2=0.24 $Y2=1.415
r99 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.58 $X2=0.2
+ $Y2=2.32
r100 16 38 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.25
+ $X2=0.24 $Y2=1.415
r101 16 18 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.24 $Y=1.25
+ $X2=0.24 $Y2=0.605
r102 15 29 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.4 $Y=1.415
+ $X2=1.23 $Y2=1.415
r103 11 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=2.16
+ $X2=2.615 $Y2=1.995
r104 11 13 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.615 $Y=2.16
+ $X2=2.615 $Y2=2.735
r105 7 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.475 $Y=1.25
+ $X2=1.4 $Y2=1.415
r106 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=1.475 $Y=1.25
+ $X2=1.475 $Y2=0.605
r107 2 24 600 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.65
r108 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.395 $X2=0.28 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%D 3 6 8 11 12 13
r44 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.09
+ $X2=1.925 $Y2=1.255
r45 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.09
+ $X2=1.925 $Y2=0.925
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.09 $X2=1.925 $Y2=1.09
r47 8 12 7.43022 $w=3.78e-07 $l=2.45e-07 $layer=LI1_cond $X=1.68 $Y=1 $X2=1.925
+ $Y2=1
r48 6 14 538.363 $w=1.8e-07 $l=1.385e-06 $layer=POLY_cond $X=1.88 $Y=2.64
+ $X2=1.88 $Y2=1.255
r49 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.865 $Y=0.605
+ $X2=1.865 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%SCD 3 7 11 12 13 14 18
c45 13 0 1.32376e-19 $X=3.12 $Y=1.665
c46 3 0 2.55706e-19 $X=3.035 $Y=2.735
r47 13 14 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r48 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.605 $X2=3.11 $Y2=1.605
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.945
+ $X2=3.11 $Y2=1.605
r50 11 12 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.945
+ $X2=3.11 $Y2=2.11
r51 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.44
+ $X2=3.11 $Y2=1.605
r52 7 10 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=3.05 $Y=0.605
+ $X2=3.05 $Y2=1.44
r53 3 12 242.944 $w=1.8e-07 $l=6.25e-07 $layer=POLY_cond $X=3.035 $Y=2.735
+ $X2=3.035 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%CLK 1 3 6 10 12 15
c52 10 0 5.22915e-20 $X=4.62 $Y=1.61
r53 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.02
+ $Y=1.105 $X2=4.02 $Y2=1.105
r54 12 16 1.31678 $w=5.43e-07 $l=6e-08 $layer=LI1_cond $X=4.08 $Y=1.277 $X2=4.02
+ $Y2=1.277
r55 10 11 5 $w=2.41e-07 $l=2.5e-08 $layer=POLY_cond $X=4.62 $Y=1.61 $X2=4.645
+ $Y2=1.61
r56 9 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.02 $Y=1.445
+ $X2=4.02 $Y2=1.105
r57 9 10 120 $w=2.41e-07 $l=6e-07 $layer=POLY_cond $X=4.02 $Y=1.61 $X2=4.62
+ $Y2=1.61
r58 4 11 9.67267 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.645 $Y=1.775
+ $X2=4.645 $Y2=1.61
r59 4 6 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.645 $Y=1.775
+ $X2=4.645 $Y2=2.495
r60 1 10 13.8727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.62 $Y=1.445
+ $X2=4.62 $Y2=1.61
r61 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.62 $Y=1.445 $X2=4.62
+ $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_1025_119# 1 2 9 11 15 17 19 20 21 24 29
+ 31 32 33 36 39 42 43 44 46 51 53 56 63 64 67 69 71 81
c204 71 0 6.65228e-20 $X=6.045 $Y=1.575
c205 64 0 3.17494e-19 $X=9.475 $Y=1.07
c206 63 0 2.9567e-20 $X=9.475 $Y=1.07
c207 53 0 3.30675e-20 $X=5.405 $Y=1.665
c208 51 0 1.19518e-19 $X=5.525 $Y=1.132
c209 39 0 1.50504e-19 $X=8.155 $Y=0.665
c210 31 0 1.9224e-20 $X=5.525 $Y=1.5
c211 15 0 6.36741e-20 $X=6.54 $Y=0.805
r212 68 81 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=9.615 $Y=2.03
+ $X2=9.7 $Y2=2.03
r213 67 69 5.06676 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.532 $Y=2.03
+ $X2=9.532 $Y2=1.865
r214 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.615
+ $Y=2.03 $X2=9.615 $Y2=2.03
r215 64 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.475 $Y=1.07
+ $X2=9.475 $Y2=1.16
r216 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.475
+ $Y=1.07 $X2=9.475 $Y2=1.07
r217 60 63 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.185 $Y=1.07
+ $X2=9.475 $Y2=1.07
r218 56 58 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.085 $Y=0.395
+ $X2=7.085 $Y2=0.665
r219 53 55 17.4006 $w=3.12e-07 $l=4.45e-07 $layer=LI1_cond $X=5.405 $Y=1.665
+ $X2=5.405 $Y2=2.11
r220 47 63 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.235
+ $X2=9.475 $Y2=1.07
r221 47 69 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=9.475 $Y=1.235
+ $X2=9.475 $Y2=1.865
r222 46 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=0.905
+ $X2=9.185 $Y2=1.07
r223 45 46 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.185 $Y=0.425
+ $X2=9.185 $Y2=0.905
r224 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.1 $Y=0.34
+ $X2=9.185 $Y2=0.425
r225 43 44 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=9.1 $Y=0.34
+ $X2=8.325 $Y2=0.34
r226 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.325 $Y2=0.34
r227 41 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.24 $Y2=0.58
r228 40 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=0.665
+ $X2=7.085 $Y2=0.665
r229 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.155 $Y=0.665
+ $X2=8.24 $Y2=0.58
r230 39 40 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=8.155 $Y=0.665
+ $X2=7.17 $Y2=0.665
r231 37 74 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.665
+ $X2=6.045 $Y2=1.83
r232 37 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.045 $Y=1.665
+ $X2=6.045 $Y2=1.575
r233 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.045
+ $Y=1.665 $X2=6.045 $Y2=1.665
r234 34 53 0.37154 $w=3.3e-07 $l=2.4e-07 $layer=LI1_cond $X=5.645 $Y=1.665
+ $X2=5.405 $Y2=1.665
r235 34 36 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.645 $Y=1.665
+ $X2=6.045 $Y2=1.665
r236 32 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.395
+ $X2=7.085 $Y2=0.395
r237 32 33 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=7 $Y=0.395
+ $X2=5.43 $Y2=0.395
r238 31 53 7.13281 $w=3.12e-07 $l=2.16852e-07 $layer=LI1_cond $X=5.525 $Y=1.5
+ $X2=5.405 $Y2=1.665
r239 30 51 1.74499 $w=2.4e-07 $l=1.43e-07 $layer=LI1_cond $X=5.525 $Y=1.275
+ $X2=5.525 $Y2=1.132
r240 30 31 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=5.525 $Y=1.275
+ $X2=5.525 $Y2=1.5
r241 27 51 10.5135 $w=2.83e-07 $l=2.6e-07 $layer=LI1_cond $X=5.265 $Y=1.132
+ $X2=5.525 $Y2=1.132
r242 27 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.265 $Y=0.99
+ $X2=5.265 $Y2=0.74
r243 26 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.265 $Y=0.48
+ $X2=5.43 $Y2=0.395
r244 26 29 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.265 $Y=0.48
+ $X2=5.265 $Y2=0.74
r245 22 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.7 $Y=2.195
+ $X2=9.7 $Y2=2.03
r246 22 24 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.7 $Y=2.195
+ $X2=9.7 $Y2=2.565
r247 20 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.31 $Y=1.16
+ $X2=9.475 $Y2=1.16
r248 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.31 $Y=1.16
+ $X2=8.95 $Y2=1.16
r249 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.875 $Y=1.085
+ $X2=8.95 $Y2=1.16
r250 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.875 $Y=1.085
+ $X2=8.875 $Y2=0.69
r251 13 15 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.54 $Y=1.5
+ $X2=6.54 $Y2=0.805
r252 12 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.575
+ $X2=6.045 $Y2=1.575
r253 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.465 $Y=1.575
+ $X2=6.54 $Y2=1.5
r254 11 12 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.465 $Y=1.575
+ $X2=6.21 $Y2=1.575
r255 9 74 258.492 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=6.1 $Y=2.495
+ $X2=6.1 $Y2=1.83
r256 2 55 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.935 $X2=5.32 $Y2=2.11
r257 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.125
+ $Y=0.595 $X2=5.265 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_1370_290# 1 2 9 13 17 18 21 22 24 32 33
+ 35
c89 33 0 1.87473e-19 $X=8.845 $Y=0.842
c90 21 0 6.53341e-20 $X=7.21 $Y=1.005
c91 13 0 1.56765e-19 $X=6.93 $Y=0.805
r92 36 38 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.93 $Y=1.615 $X2=6.94
+ $Y2=1.615
r93 31 33 4.47019 $w=4.93e-07 $l=1.85e-07 $layer=LI1_cond $X=8.66 $Y=0.842
+ $X2=8.845 $Y2=0.842
r94 31 32 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=8.66 $Y=0.842
+ $X2=8.495 $Y2=0.842
r95 28 33 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.845 $Y=1.09
+ $X2=8.845 $Y2=0.842
r96 28 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.845 $Y=1.09
+ $X2=8.845 $Y2=1.745
r97 24 26 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=8.785 $Y=1.91
+ $X2=8.785 $Y2=2.59
r98 22 35 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=8.785 $Y=1.89
+ $X2=8.785 $Y2=1.745
r99 22 24 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=8.785 $Y=1.89
+ $X2=8.785 $Y2=1.91
r100 21 32 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=8.495 $Y2=1.005
r101 18 38 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=1.615
+ $X2=6.94 $Y2=1.615
r102 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.105
+ $Y=1.615 $X2=7.105 $Y2=1.615
r103 15 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.105 $Y=1.09
+ $X2=7.21 $Y2=1.005
r104 15 17 27.7273 $w=2.08e-07 $l=5.25e-07 $layer=LI1_cond $X=7.105 $Y=1.09
+ $X2=7.105 $Y2=1.615
r105 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.93 $Y=1.45
+ $X2=6.93 $Y2=1.615
r106 11 13 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.93 $Y=1.45
+ $X2=6.93 $Y2=0.805
r107 7 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.78
+ $X2=6.94 $Y2=1.615
r108 7 9 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=6.94 $Y=1.78
+ $X2=6.94 $Y2=2.495
r109 2 26 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.59
+ $Y=1.735 $X2=8.725 $Y2=2.59
r110 2 24 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.59
+ $Y=1.735 $X2=8.725 $Y2=1.91
r111 1 31 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.52
+ $Y=0.37 $X2=8.66 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%RESET_B 4 7 9 10 14 15 16 17 19 21 24 30 33
+ 36 38 39 40 41 49 52 53 56 59 61 63 72
c215 72 0 1.25229e-19 $X=10.8 $Y=2.035
c216 33 0 1.32376e-19 $X=3.585 $Y=1.985
c217 9 0 1.66e-21 $X=7.245 $Y=0.18
c218 7 0 1.3005e-19 $X=3.585 $Y=2.735
r219 61 64 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.945 $Y=1.985
+ $X2=10.945 $Y2=2.15
r220 61 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.945 $Y=1.985
+ $X2=10.945 $Y2=1.82
r221 61 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.945
+ $Y=1.985 $X2=10.945 $Y2=1.985
r222 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.825
+ $Y=1.96 $X2=7.825 $Y2=1.96
r223 56 58 15.4929 $w=2.8e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=1.98
+ $X2=7.825 $Y2=1.98
r224 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.985 $X2=3.95 $Y2=1.985
r225 49 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r226 47 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r227 43 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r228 41 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r229 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r230 40 41 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r231 39 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r232 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r233 38 39 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r234 34 36 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=10.715 $Y=1.55
+ $X2=10.855 $Y2=1.55
r235 32 52 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=3.675 $Y=1.985
+ $X2=3.95 $Y2=1.985
r236 32 33 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.675 $Y=1.985
+ $X2=3.585 $Y2=1.985
r237 30 64 161.315 $w=1.8e-07 $l=4.15e-07 $layer=POLY_cond $X=11.005 $Y=2.565
+ $X2=11.005 $Y2=2.15
r238 26 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.855 $Y=1.625
+ $X2=10.855 $Y2=1.55
r239 26 63 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=10.855 $Y=1.625
+ $X2=10.855 $Y2=1.82
r240 22 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.475
+ $X2=10.715 $Y2=1.55
r241 22 24 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=10.715 $Y=1.475
+ $X2=10.715 $Y2=0.58
r242 21 56 17.3521 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=7.735 $Y=1.795
+ $X2=7.735 $Y2=1.98
r243 20 21 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=7.735 $Y=1.24
+ $X2=7.735 $Y2=1.795
r244 17 56 36.15 $w=2.8e-07 $l=2.8801e-07 $layer=POLY_cond $X=7.525 $Y=2.165
+ $X2=7.735 $Y2=1.98
r245 17 19 88.3667 $w=1.8e-07 $l=3.3e-07 $layer=POLY_cond $X=7.525 $Y=2.165
+ $X2=7.525 $Y2=2.495
r246 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.66 $Y=1.165
+ $X2=7.735 $Y2=1.24
r247 15 16 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=7.66 $Y=1.165
+ $X2=7.395 $Y2=1.165
r248 12 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.32 $Y=1.09
+ $X2=7.395 $Y2=1.165
r249 12 14 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.32 $Y=1.09
+ $X2=7.32 $Y2=0.805
r250 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.32 $Y=0.255
+ $X2=7.32 $Y2=0.805
r251 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.245 $Y=0.18
+ $X2=7.32 $Y2=0.255
r252 9 10 1845.96 $w=1.5e-07 $l=3.6e-06 $layer=POLY_cond $X=7.245 $Y=0.18
+ $X2=3.645 $Y2=0.18
r253 5 33 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=2.15
+ $X2=3.585 $Y2=1.985
r254 5 7 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=3.585 $Y=2.15
+ $X2=3.585 $Y2=2.735
r255 2 33 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.57 $Y=1.82
+ $X2=3.585 $Y2=1.985
r256 2 4 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.57 $Y=1.82
+ $X2=3.57 $Y2=0.605
r257 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.57 $Y=0.255
+ $X2=3.645 $Y2=0.18
r258 1 4 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.57 $Y=0.255
+ $X2=3.57 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_1223_119# 1 2 3 12 16 18 23 24 25 27 28
+ 30 31
c102 30 0 1.03439e-19 $X=8.425 $Y=1.41
c103 25 0 1.70204e-19 $X=6.83 $Y=2.425
c104 12 0 2.9567e-20 $X=8.445 $Y=0.69
r105 31 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.425 $Y=1.41
+ $X2=8.425 $Y2=1.575
r106 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.425 $Y=1.41
+ $X2=8.425 $Y2=1.245
r107 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.425
+ $Y=1.41 $X2=8.425 $Y2=1.41
r108 28 30 32.0123 $w=3.13e-07 $l=8.75e-07 $layer=LI1_cond $X=7.55 $Y=1.417
+ $X2=8.425 $Y2=1.417
r109 27 38 10.3482 $w=3.36e-07 $l=3.72552e-07 $layer=LI1_cond $X=7.465 $Y=2.32
+ $X2=7.75 $Y2=2.522
r110 26 28 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.465 $Y=1.575
+ $X2=7.55 $Y2=1.417
r111 26 27 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.465 $Y=1.575
+ $X2=7.465 $Y2=2.32
r112 24 27 6.05874 $w=3.36e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.38 $Y=2.425
+ $X2=7.465 $Y2=2.32
r113 24 25 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.38 $Y=2.425
+ $X2=6.83 $Y2=2.425
r114 23 25 6.00066 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.745 $Y=2.34
+ $X2=6.83 $Y2=2.425
r115 23 34 15.5273 $w=3.3e-07 $l=5.06991e-07 $layer=LI1_cond $X=6.745 $Y=2.34
+ $X2=6.325 $Y2=2.532
r116 22 23 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=6.745 $Y=0.95
+ $X2=6.745 $Y2=2.34
r117 18 22 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.66 $Y=0.8
+ $X2=6.745 $Y2=0.95
r118 18 20 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.66 $Y=0.8
+ $X2=6.325 $Y2=0.8
r119 16 41 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=8.5 $Y=2.235
+ $X2=8.5 $Y2=1.575
r120 12 40 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.445 $Y=0.69
+ $X2=8.445 $Y2=1.245
r121 3 38 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=7.615
+ $Y=2.285 $X2=7.75 $Y2=2.52
r122 2 34 600 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=6.19
+ $Y=2.285 $X2=6.325 $Y2=2.53
r123 1 20 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=6.115
+ $Y=0.595 $X2=6.325 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_852_119# 1 2 9 12 14 17 19 20 21 22 23 24
+ 26 29 31 36 37 38 41 43 44 47 50 52 56 60 61
c173 56 0 6.65228e-20 $X=4.49 $Y=1.717
c174 43 0 5.15375e-20 $X=5.595 $Y=1.52
c175 38 0 1.31172e-19 $X=9.04 $Y=1.55
c176 37 0 1.34905e-19 $X=9.85 $Y=1.55
c177 19 0 1.70204e-19 $X=5.595 $Y=3.075
c178 14 0 1.19518e-19 $X=5.52 $Y=1.52
r179 60 61 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.14 $Y=1.52
+ $X2=5.14 $Y2=1.445
r180 59 63 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.61
+ $X2=5.14 $Y2=1.775
r181 59 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.14 $Y=1.61 $X2=5.14
+ $Y2=1.52
r182 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.61 $X2=5.14 $Y2=1.61
r183 56 58 17.3904 $w=4.56e-07 $l=6.5e-07 $layer=LI1_cond $X=4.49 $Y=1.717
+ $X2=5.14 $Y2=1.717
r184 55 56 0.802632 $w=4.56e-07 $l=3e-08 $layer=LI1_cond $X=4.46 $Y=1.717
+ $X2=4.49 $Y2=1.717
r185 50 56 6.58228 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=4.49 $Y=1.445
+ $X2=4.49 $Y2=1.717
r186 49 52 2.99516 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.49 $Y=0.835
+ $X2=4.405 $Y2=0.71
r187 49 50 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.49 $Y=0.835
+ $X2=4.49 $Y2=1.445
r188 45 55 4.25555 $w=2.5e-07 $l=2.73e-07 $layer=LI1_cond $X=4.46 $Y=1.99
+ $X2=4.46 $Y2=1.717
r189 45 47 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=4.46 $Y=1.99
+ $X2=4.46 $Y2=2.11
r190 39 41 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=9.925 $Y=1.475
+ $X2=9.925 $Y2=0.58
r191 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.85 $Y=1.55
+ $X2=9.925 $Y2=1.475
r192 37 38 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.85 $Y=1.55
+ $X2=9.04 $Y2=1.55
r193 34 36 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=8.95 $Y=3.075
+ $X2=8.95 $Y2=2.235
r194 33 38 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.95 $Y=1.625
+ $X2=9.04 $Y2=1.55
r195 33 36 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=8.95 $Y=1.625
+ $X2=8.95 $Y2=2.235
r196 32 44 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.64 $Y=3.15 $X2=6.55
+ $Y2=3.15
r197 31 34 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.86 $Y=3.15
+ $X2=8.95 $Y2=3.075
r198 31 32 1138.34 $w=1.5e-07 $l=2.22e-06 $layer=POLY_cond $X=8.86 $Y=3.15
+ $X2=6.64 $Y2=3.15
r199 27 44 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.55 $Y=3.075
+ $X2=6.55 $Y2=3.15
r200 27 29 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.55 $Y=3.075
+ $X2=6.55 $Y2=2.495
r201 24 26 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=6.04 $Y=1.11
+ $X2=6.04 $Y2=0.805
r202 22 44 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.46 $Y=3.15 $X2=6.55
+ $Y2=3.15
r203 22 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.46 $Y=3.15
+ $X2=5.67 $Y2=3.15
r204 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.965 $Y=1.185
+ $X2=6.04 $Y2=1.11
r205 20 21 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.965 $Y=1.185
+ $X2=5.67 $Y2=1.185
r206 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.595 $Y=3.075
+ $X2=5.67 $Y2=3.15
r207 18 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.595 $Y=1.595
+ $X2=5.595 $Y2=1.52
r208 18 19 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=5.595 $Y=1.595
+ $X2=5.595 $Y2=3.075
r209 17 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.595 $Y=1.445
+ $X2=5.595 $Y2=1.52
r210 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.595 $Y=1.26
+ $X2=5.67 $Y2=1.185
r211 16 17 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.595 $Y=1.26
+ $X2=5.595 $Y2=1.445
r212 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.52
+ $X2=5.14 $Y2=1.52
r213 14 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.52 $Y=1.52
+ $X2=5.595 $Y2=1.52
r214 14 15 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.52 $Y=1.52
+ $X2=5.305 $Y2=1.52
r215 12 63 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.095 $Y=2.495
+ $X2=5.095 $Y2=1.775
r216 9 61 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.05 $Y=0.965
+ $X2=5.05 $Y2=1.445
r217 2 47 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.935 $X2=4.42 $Y2=2.11
r218 1 52 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.595 $X2=4.405 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_2006_373# 1 2 9 13 18 19 20 21 22 23 26
+ 28 29 31 32
c114 22 0 2.94687e-20 $X=11.065 $Y=2.405
c115 21 0 1.34905e-19 $X=10.545 $Y=1.565
c116 20 0 2.52042e-21 $X=11.69 $Y=1.565
c117 13 0 1.25229e-19 $X=10.285 $Y=0.58
r118 37 39 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.12 $Y=2.03
+ $X2=10.285 $Y2=2.03
r119 32 35 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=11.23 $Y=2.405
+ $X2=11.23 $Y2=2.565
r120 30 31 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=11.775 $Y=0.875
+ $X2=11.775 $Y2=1.48
r121 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.69 $Y=0.79
+ $X2=11.775 $Y2=0.875
r122 28 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.69 $Y=0.79
+ $X2=11.455 $Y2=0.79
r123 24 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.29 $Y=0.705
+ $X2=11.455 $Y2=0.79
r124 24 26 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=11.29 $Y=0.705
+ $X2=11.29 $Y2=0.58
r125 22 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=2.405
+ $X2=11.23 $Y2=2.405
r126 22 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.065 $Y=2.405
+ $X2=10.545 $Y2=2.405
r127 20 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.69 $Y=1.565
+ $X2=11.775 $Y2=1.48
r128 20 21 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=11.69 $Y=1.565
+ $X2=10.545 $Y2=1.565
r129 19 39 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=10.405 $Y=2.03
+ $X2=10.285 $Y2=2.03
r130 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.405
+ $Y=2.03 $X2=10.405 $Y2=2.03
r131 16 23 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.405 $Y=2.32
+ $X2=10.545 $Y2=2.405
r132 16 18 11.936 $w=2.78e-07 $l=2.9e-07 $layer=LI1_cond $X=10.405 $Y=2.32
+ $X2=10.405 $Y2=2.03
r133 15 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.405 $Y=1.65
+ $X2=10.545 $Y2=1.565
r134 15 18 15.6403 $w=2.78e-07 $l=3.8e-07 $layer=LI1_cond $X=10.405 $Y=1.65
+ $X2=10.405 $Y2=2.03
r135 11 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.285 $Y=1.865
+ $X2=10.285 $Y2=2.03
r136 11 13 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=10.285 $Y=1.865
+ $X2=10.285 $Y2=0.58
r137 7 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.12 $Y=2.195
+ $X2=10.12 $Y2=2.03
r138 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=10.12 $Y=2.195
+ $X2=10.12 $Y2=2.565
r139 2 35 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.095
+ $Y=2.355 $X2=11.23 $Y2=2.565
r140 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.15
+ $Y=0.37 $X2=11.29 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_1790_74# 1 2 9 11 13 15 19 23 27 31 33 35
+ 39 47 51 56 58 61 64
c146 58 0 1.02173e-19 $X=10.01 $Y=2.365
c147 56 0 1.57754e-19 $X=10.01 $Y=1.045
c148 27 0 2.52042e-21 $X=12.44 $Y=2.4
c149 19 0 7.64129e-20 $X=11.99 $Y=2.4
c150 13 0 1.05882e-19 $X=11.455 $Y=2.565
r151 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.355
+ $Y=1.175 $X2=11.355 $Y2=1.175
r152 59 64 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.095 $Y=1.177
+ $X2=10.01 $Y2=1.177
r153 59 61 54.7954 $w=2.63e-07 $l=1.26e-06 $layer=LI1_cond $X=10.095 $Y=1.177
+ $X2=11.355 $Y2=1.177
r154 57 64 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.01 $Y=1.31
+ $X2=10.01 $Y2=1.177
r155 57 58 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=10.01 $Y=1.31
+ $X2=10.01 $Y2=2.365
r156 56 64 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=10.01 $Y=1.045
+ $X2=10.01 $Y2=1.177
r157 55 56 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.01 $Y=0.735
+ $X2=10.01 $Y2=1.045
r158 51 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=0.57
+ $X2=10.01 $Y2=0.735
r159 51 53 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.925 $Y=0.57
+ $X2=9.655 $Y2=0.57
r160 47 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.53
+ $X2=10.01 $Y2=2.365
r161 47 49 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=9.925 $Y=2.53
+ $X2=9.37 $Y2=2.53
r162 41 42 13.8758 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=11.99 $Y=1.422
+ $X2=12.085 $Y2=1.422
r163 37 46 21.2229 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=12.99 $Y=1.255
+ $X2=12.99 $Y2=1.422
r164 37 39 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=12.99 $Y=1.255
+ $X2=12.99 $Y2=0.69
r165 33 46 6.57273 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=12.945 $Y=1.422
+ $X2=12.99 $Y2=1.422
r166 33 44 62.8061 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=12.945 $Y=1.422
+ $X2=12.515 $Y2=1.422
r167 33 35 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=12.945 $Y=1.585
+ $X2=12.945 $Y2=2.46
r168 29 44 21.2229 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=12.515 $Y=1.255
+ $X2=12.515 $Y2=1.422
r169 29 31 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.515 $Y=1.255
+ $X2=12.515 $Y2=0.74
r170 25 44 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.44 $Y=1.422
+ $X2=12.515 $Y2=1.422
r171 25 42 51.8515 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=12.44 $Y=1.422
+ $X2=12.085 $Y2=1.422
r172 25 27 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=12.44 $Y=1.585
+ $X2=12.44 $Y2=2.4
r173 21 42 21.2229 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=12.085 $Y=1.255
+ $X2=12.085 $Y2=1.422
r174 21 23 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.085 $Y=1.255
+ $X2=12.085 $Y2=0.74
r175 17 41 16.9318 $w=1.8e-07 $l=1.68e-07 $layer=POLY_cond $X=11.99 $Y=1.59
+ $X2=11.99 $Y2=1.422
r176 17 19 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=11.99 $Y=1.59
+ $X2=11.99 $Y2=2.4
r177 16 62 36.297 $w=3.28e-07 $l=3.76776e-07 $layer=POLY_cond $X=11.545 $Y=1.422
+ $X2=11.272 $Y2=1.175
r178 15 41 12.9493 $w=3.35e-07 $l=9e-08 $layer=POLY_cond $X=11.9 $Y=1.422
+ $X2=11.99 $Y2=1.422
r179 15 16 61.1493 $w=3.35e-07 $l=3.55e-07 $layer=POLY_cond $X=11.9 $Y=1.422
+ $X2=11.545 $Y2=1.422
r180 11 16 34.4294 $w=3.28e-07 $l=2.08192e-07 $layer=POLY_cond $X=11.455 $Y=1.59
+ $X2=11.545 $Y2=1.422
r181 11 13 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=11.455 $Y=1.59
+ $X2=11.455 $Y2=2.565
r182 7 62 38.5876 $w=3.28e-07 $l=2.67047e-07 $layer=POLY_cond $X=11.075 $Y=1.01
+ $X2=11.272 $Y2=1.175
r183 7 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.075 $Y=1.01
+ $X2=11.075 $Y2=0.58
r184 2 49 600 $w=1.7e-07 $l=9.45714e-07 $layer=licon1_PDIFF $count=1 $X=9.04
+ $Y=1.735 $X2=9.37 $Y2=2.53
r185 1 53 182 $w=1.7e-07 $l=7.98765e-07 $layer=licon1_NDIFF $count=1 $X=8.95
+ $Y=0.37 $X2=9.655 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_2607_392# 1 2 9 13 17 21 23 27 31 35 41
+ 44
r50 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.8
+ $Y=1.465 $X2=13.8 $Y2=1.465
r51 39 44 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=13.325 $Y=1.465
+ $X2=13.195 $Y2=1.465
r52 39 41 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=13.325 $Y=1.465
+ $X2=13.8 $Y2=1.465
r53 35 37 31.4706 $w=2.58e-07 $l=7.1e-07 $layer=LI1_cond $X=13.195 $Y=2.105
+ $X2=13.195 $Y2=2.815
r54 33 44 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.63
+ $X2=13.195 $Y2=1.465
r55 33 35 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=13.195 $Y=1.63
+ $X2=13.195 $Y2=2.105
r56 29 44 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.3
+ $X2=13.195 $Y2=1.465
r57 29 31 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=13.195 $Y=1.3
+ $X2=13.195 $Y2=0.515
r58 26 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=14.385 $Y=1.465
+ $X2=14.4 $Y2=1.465
r59 25 26 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=13.97 $Y=1.465
+ $X2=14.385 $Y2=1.465
r60 24 25 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=13.935 $Y=1.465
+ $X2=13.97 $Y2=1.465
r61 23 42 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.8 $Y2=1.465
r62 23 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.935 $Y2=1.465
r63 19 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.4 $Y=1.3
+ $X2=14.4 $Y2=1.465
r64 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.4 $Y=1.3 $X2=14.4
+ $Y2=0.74
r65 15 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.385 $Y=1.63
+ $X2=14.385 $Y2=1.465
r66 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=14.385 $Y=1.63
+ $X2=14.385 $Y2=2.4
r67 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.97 $Y=1.3
+ $X2=13.97 $Y2=1.465
r68 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.97 $Y=1.3
+ $X2=13.97 $Y2=0.74
r69 7 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.935 $Y=1.63
+ $X2=13.935 $Y2=1.465
r70 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.935 $Y=1.63
+ $X2=13.935 $Y2=2.4
r71 2 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=13.035
+ $Y=1.96 $X2=13.17 $Y2=2.815
r72 2 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.035
+ $Y=1.96 $X2=13.17 $Y2=2.105
r73 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.065
+ $Y=0.37 $X2=13.205 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 59 65 69 71 76 77 79 80 81 88 106 110 115 120 125 133 136 138 141 144 151 154
+ 157 161
r181 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r182 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r183 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r184 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r185 142 148 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.32 $Y2=3.33
r186 141 142 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r187 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r188 135 136 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.072
+ $X2=1.4 $Y2=3.072
r189 131 135 0.611135 $w=6.83e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=3.072
+ $X2=1.235 $Y2=3.072
r190 131 133 18.0422 $w=6.83e-07 $l=5.85e-07 $layer=LI1_cond $X=1.2 $Y=3.072
+ $X2=0.615 $Y2=3.072
r191 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r192 129 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r193 129 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r194 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r195 126 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=13.71 $Y2=3.33
r196 126 128 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=14.16 $Y2=3.33
r197 125 160 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.687 $Y2=3.33
r198 125 128 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.16 $Y2=3.33
r199 124 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r200 124 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r201 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r202 121 154 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.83 $Y=3.33
+ $X2=12.685 $Y2=3.33
r203 121 123 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.83 $Y=3.33
+ $X2=13.2 $Y2=3.33
r204 120 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.71 $Y2=3.33
r205 120 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.2 $Y2=3.33
r206 119 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r207 119 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r208 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r209 116 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.85 $Y=3.33
+ $X2=11.725 $Y2=3.33
r210 116 118 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.85 $Y=3.33
+ $X2=12.24 $Y2=3.33
r211 115 154 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.685 $Y2=3.33
r212 115 118 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.24 $Y2=3.33
r213 114 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r214 114 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r215 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r216 111 113 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=11.28 $Y2=3.33
r217 110 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.6 $Y=3.33
+ $X2=11.725 $Y2=3.33
r218 110 113 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.6 $Y=3.33
+ $X2=11.28 $Y2=3.33
r219 109 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r220 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r221 106 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=8.315 $Y2=3.33
r222 106 108 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=7.92 $Y2=3.33
r223 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r224 102 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r225 101 104 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r226 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r227 99 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r228 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r229 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r230 96 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r231 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r232 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r233 93 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.28 $Y2=3.33
r234 93 95 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.6 $Y2=3.33
r235 92 139 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r236 92 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r237 91 136 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.4 $Y2=3.33
r238 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r239 88 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.28 $Y2=3.33
r240 88 91 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=1.68 $Y2=3.33
r241 86 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r242 85 133 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.615 $Y2=3.33
r243 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r244 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r245 81 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r246 79 104 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.07 $Y=3.33
+ $X2=6.96 $Y2=3.33
r247 79 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.07 $Y=3.33
+ $X2=7.195 $Y2=3.33
r248 78 108 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.92 $Y2=3.33
r249 78 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.195 $Y2=3.33
r250 76 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r251 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r252 75 101 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r253 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r254 71 74 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=14.635 $Y=1.985
+ $X2=14.635 $Y2=2.815
r255 69 160 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.687 $Y2=3.33
r256 69 74 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.635 $Y2=2.815
r257 65 68 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.71 $Y=1.985
+ $X2=13.71 $Y2=2.815
r258 63 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=3.33
r259 63 68 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=2.815
r260 59 62 29.0098 $w=2.88e-07 $l=7.3e-07 $layer=LI1_cond $X=12.685 $Y=2.085
+ $X2=12.685 $Y2=2.815
r261 57 154 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.685 $Y=3.245
+ $X2=12.685 $Y2=3.33
r262 57 62 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=12.685 $Y=3.245
+ $X2=12.685 $Y2=2.815
r263 53 56 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.725 $Y=1.985
+ $X2=11.725 $Y2=2.815
r264 51 151 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.725 $Y=3.245
+ $X2=11.725 $Y2=3.33
r265 51 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.725 $Y=3.245
+ $X2=11.725 $Y2=2.815
r266 50 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.44 $Y=3.33
+ $X2=8.315 $Y2=3.33
r267 49 111 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=10.562 $Y=3.33
+ $X2=10.86 $Y2=3.33
r268 49 148 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r269 49 144 10.1516 $w=5.93e-07 $l=5.05e-07 $layer=LI1_cond $X=10.562 $Y=3.33
+ $X2=10.562 $Y2=2.825
r270 49 50 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=10.265 $Y=3.33
+ $X2=8.44 $Y2=3.33
r271 45 48 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.315 $Y=1.91
+ $X2=8.315 $Y2=2.59
r272 43 141 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.315 $Y=3.245
+ $X2=8.315 $Y2=3.33
r273 43 48 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=8.315 $Y=3.245
+ $X2=8.315 $Y2=2.59
r274 39 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=3.245
+ $X2=7.195 $Y2=3.33
r275 39 41 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=7.195 $Y=3.245
+ $X2=7.195 $Y2=2.845
r276 35 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r277 35 37 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.88
r278 31 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=3.33
r279 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=2.78
r280 10 74 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.475
+ $Y=1.84 $X2=14.61 $Y2=2.815
r281 10 71 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.475
+ $Y=1.84 $X2=14.61 $Y2=1.985
r282 9 68 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.84 $X2=13.71 $Y2=2.815
r283 9 65 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.84 $X2=13.71 $Y2=1.985
r284 8 62 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.84 $X2=12.665 $Y2=2.815
r285 8 59 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.84 $X2=12.665 $Y2=2.085
r286 7 56 600 $w=1.7e-07 $l=5.59285e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=2.355 $X2=11.765 $Y2=2.815
r287 7 53 300 $w=1.7e-07 $l=4.67226e-07 $layer=licon1_PDIFF $count=2 $X=11.545
+ $Y=2.355 $X2=11.765 $Y2=1.985
r288 6 144 600 $w=1.7e-07 $l=6.20806e-07 $layer=licon1_PDIFF $count=1 $X=10.21
+ $Y=2.355 $X2=10.56 $Y2=2.825
r289 5 48 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=8.15
+ $Y=1.735 $X2=8.275 $Y2=2.59
r290 5 45 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.15
+ $Y=1.735 $X2=8.275 $Y2=1.91
r291 4 41 600 $w=1.7e-07 $l=6.54523e-07 $layer=licon1_PDIFF $count=1 $X=7.03
+ $Y=2.285 $X2=7.235 $Y2=2.845
r292 3 37 600 $w=1.7e-07 $l=1.01025e-06 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=1.935 $X2=4.87 $Y2=2.88
r293 2 33 600 $w=1.7e-07 $l=4.3566e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=2.415 $X2=3.28 $Y2=2.78
r294 1 135 300 $w=1.7e-07 $l=8.52291e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.32 $X2=1.235 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%A_388_79# 1 2 3 4 5 16 22 24 25 27 28 29 31
+ 32 34 36 39 41 42 43 44 45 47 51
c164 47 0 5.15375e-20 $X=6.405 $Y=2
c165 34 0 1.20066e-19 $X=3.83 $Y=2.88
c166 16 0 1.3005e-19 $X=2.775 $Y=2.785
r167 48 49 2.85743 $w=4.91e-07 $l=1.15e-07 $layer=LI1_cond $X=3.72 $Y=2.42
+ $X2=3.72 $Y2=2.535
r168 46 47 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.405 $Y=1.29
+ $X2=6.405 $Y2=2
r169 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=1.205
+ $X2=6.405 $Y2=1.29
r170 44 45 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.32 $Y=1.205
+ $X2=5.99 $Y2=1.205
r171 42 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=2.085
+ $X2=6.405 $Y2=2
r172 42 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.32 $Y=2.085
+ $X2=5.985 $Y2=2.085
r173 41 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.905 $Y=1.12
+ $X2=5.99 $Y2=1.205
r174 40 51 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.905 $Y=0.82
+ $X2=5.825 $Y2=0.735
r175 40 41 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.905 $Y=0.82
+ $X2=5.905 $Y2=1.12
r176 39 55 3.23633 $w=2.3e-07 $l=1.51063e-07 $layer=LI1_cond $X=5.87 $Y=2.445
+ $X2=5.847 $Y2=2.585
r177 38 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.87 $Y=2.17
+ $X2=5.985 $Y2=2.085
r178 38 39 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.87 $Y=2.17
+ $X2=5.87 $Y2=2.445
r179 37 49 6.68641 $w=1.8e-07 $l=2.75e-07 $layer=LI1_cond $X=3.995 $Y=2.535
+ $X2=3.72 $Y2=2.535
r180 36 55 3.71285 $w=1.8e-07 $l=1.60059e-07 $layer=LI1_cond $X=5.71 $Y=2.535
+ $X2=5.847 $Y2=2.585
r181 36 37 105.672 $w=1.78e-07 $l=1.715e-06 $layer=LI1_cond $X=5.71 $Y=2.535
+ $X2=3.995 $Y2=2.535
r182 32 49 2.89173 $w=4.91e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.805 $Y=2.625
+ $X2=3.72 $Y2=2.535
r183 32 34 7.7335 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=3.805 $Y=2.625
+ $X2=3.805 $Y2=2.88
r184 31 48 8.03646 $w=4.91e-07 $l=2.34734e-07 $layer=LI1_cond $X=3.53 $Y=2.32
+ $X2=3.72 $Y2=2.42
r185 30 31 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=3.53 $Y=1.175
+ $X2=3.53 $Y2=2.32
r186 28 48 6.03726 $w=2e-07 $l=2.75e-07 $layer=LI1_cond $X=3.445 $Y=2.42
+ $X2=3.72 $Y2=2.42
r187 28 29 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=3.445 $Y=2.42
+ $X2=2.945 $Y2=2.42
r188 26 29 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.86 $Y=2.52
+ $X2=2.945 $Y2=2.42
r189 26 27 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.86 $Y=2.52
+ $X2=2.86 $Y2=2.66
r190 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.09
+ $X2=3.53 $Y2=1.175
r191 24 25 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.445 $Y=1.09
+ $X2=2.61 $Y2=1.09
r192 20 25 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=2.435 $Y=1.005
+ $X2=2.61 $Y2=1.09
r193 20 22 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=1.005
+ $X2=2.435 $Y2=0.68
r194 16 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.775 $Y=2.785
+ $X2=2.86 $Y2=2.66
r195 16 18 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=2.775 $Y=2.785
+ $X2=2.245 $Y2=2.785
r196 5 55 600 $w=1.7e-07 $l=2.97993e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=2.285 $X2=5.875 $Y2=2.525
r197 4 34 600 $w=1.7e-07 $l=5.36936e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=2.415 $X2=3.83 $Y2=2.88
r198 3 18 600 $w=1.7e-07 $l=5.45436e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=2.32 $X2=2.245 $Y2=2.745
r199 2 51 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.68
+ $Y=0.595 $X2=5.825 $Y2=0.735
r200 1 22 182 $w=1.7e-07 $l=6.21369e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.395 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%Q_N 1 2 7 8 9 16 30
r28 30 31 0.96397 $w=4.33e-07 $l=1e-08 $layer=LI1_cond $X=12.247 $Y=0.925
+ $X2=12.247 $Y2=0.915
r29 25 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.195 $Y=1.985
+ $X2=12.195 $Y2=2.815
r30 9 25 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=12.195 $Y=1.665
+ $X2=12.195 $Y2=1.985
r31 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.195 $Y=1.295
+ $X2=12.195 $Y2=1.665
r32 8 33 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=12.195 $Y=1.295
+ $X2=12.195 $Y2=1.085
r33 7 33 3.95767 $w=4.33e-07 $l=1.23e-07 $layer=LI1_cond $X=12.247 $Y=0.962
+ $X2=12.247 $Y2=1.085
r34 7 30 0.980239 $w=4.33e-07 $l=3.7e-08 $layer=LI1_cond $X=12.247 $Y=0.962
+ $X2=12.247 $Y2=0.925
r35 7 31 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=12.3 $Y=0.877
+ $X2=12.3 $Y2=0.915
r36 7 16 12.642 $w=3.28e-07 $l=3.62e-07 $layer=LI1_cond $X=12.3 $Y=0.877
+ $X2=12.3 $Y2=0.515
r37 2 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.84 $X2=12.215 $Y2=2.815
r38 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.84 $X2=12.215 $Y2=1.985
r39 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.16
+ $Y=0.37 $X2=12.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%Q 1 2 7 10
r16 7 16 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=2.815
r17 7 10 62.7441 $w=2.68e-07 $l=1.47e-06 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=0.515
r18 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.025
+ $Y=1.84 $X2=14.16 $Y2=2.815
r19 2 7 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.025
+ $Y=1.84 $X2=14.16 $Y2=1.985
r20 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.045
+ $Y=0.37 $X2=14.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 52
+ 56 58 60 63 64 66 67 69 70 71 73 99 103 108 114 118 122 124 127 130 134
c157 134 0 6.26159e-21 $X=14.64 $Y=0
r158 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r159 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r160 128 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r161 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r162 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r163 120 122 7.07024 $w=4.93e-07 $l=6.5e-08 $layer=LI1_cond $X=7.92 $Y=0.162
+ $X2=7.985 $Y2=0.162
r164 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r165 117 120 4.95346 $w=4.93e-07 $l=2.05e-07 $layer=LI1_cond $X=7.715 $Y=0.162
+ $X2=7.92 $Y2=0.162
r166 117 118 11.9029 $w=4.93e-07 $l=2.65e-07 $layer=LI1_cond $X=7.715 $Y=0.162
+ $X2=7.45 $Y2=0.162
r167 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r168 112 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r169 112 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r170 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r171 109 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=13.755 $Y2=0
r172 109 111 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=14.16 $Y2=0
r173 108 133 4.34417 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=14.495 $Y=0
+ $X2=14.687 $Y2=0
r174 108 111 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=0
+ $X2=14.16 $Y2=0
r175 107 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r176 107 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r177 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r178 104 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.895 $Y=0
+ $X2=11.77 $Y2=0
r179 104 106 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.895 $Y=0
+ $X2=12.24 $Y2=0
r180 103 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.765 $Y2=0
r181 103 106 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.24 $Y2=0
r182 102 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r183 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r184 99 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.77 $Y2=0
r185 99 101 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.28 $Y2=0
r186 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r187 98 121 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=7.92 $Y2=0
r188 97 122 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=10.32 $Y=0
+ $X2=7.985 $Y2=0
r189 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r190 93 118 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.45
+ $Y2=0
r191 90 93 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r192 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r193 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r194 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r195 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r196 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r197 81 84 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r198 81 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r199 80 83 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r200 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 78 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r202 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r203 76 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r204 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r205 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r206 73 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r207 71 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r208 71 91 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r209 71 93 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r210 69 97 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.32 $Y2=0
r211 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.5 $Y2=0
r212 68 101 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=11.28 $Y2=0
r213 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=10.5 $Y2=0
r214 66 86 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r215 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.835
+ $Y2=0
r216 65 90 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=5.04
+ $Y2=0
r217 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.835
+ $Y2=0
r218 63 83 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.6
+ $Y2=0
r219 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.805
+ $Y2=0
r220 62 86 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.56
+ $Y2=0
r221 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.805
+ $Y2=0
r222 58 133 3.0545 $w=2.85e-07 $l=1.07121e-07 $layer=LI1_cond $X=14.637 $Y=0.085
+ $X2=14.687 $Y2=0
r223 58 60 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=14.637 $Y=0.085
+ $X2=14.637 $Y2=0.515
r224 54 130 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0
r225 54 56 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0.515
r226 53 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.895 $Y=0
+ $X2=12.765 $Y2=0
r227 52 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=0
+ $X2=13.755 $Y2=0
r228 52 53 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=13.67 $Y=0
+ $X2=12.895 $Y2=0
r229 48 127 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.765 $Y=0.085
+ $X2=12.765 $Y2=0
r230 48 50 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=12.765 $Y=0.085
+ $X2=12.765 $Y2=0.545
r231 44 124 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.77 $Y=0.085
+ $X2=11.77 $Y2=0
r232 44 46 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=11.77 $Y=0.085
+ $X2=11.77 $Y2=0.37
r233 40 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0
r234 40 42 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0.58
r235 36 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=0.085
+ $X2=4.835 $Y2=0
r236 36 38 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.835 $Y=0.085
+ $X2=4.835 $Y2=0.74
r237 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0
r238 32 34 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0.605
r239 28 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r240 28 30 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.605
r241 9 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.475
+ $Y=0.37 $X2=14.615 $Y2=0.515
r242 8 56 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=13.6
+ $Y=0.37 $X2=13.755 $Y2=0.515
r243 7 50 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=12.59
+ $Y=0.37 $X2=12.73 $Y2=0.545
r244 6 46 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=11.685
+ $Y=0.225 $X2=11.81 $Y2=0.37
r245 5 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.36
+ $Y=0.37 $X2=10.5 $Y2=0.58
r246 4 117 182 $w=1.7e-07 $l=4.34511e-07 $layer=licon1_NDIFF $count=1 $X=7.395
+ $Y=0.595 $X2=7.715 $Y2=0.325
r247 3 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.695
+ $Y=0.595 $X2=4.835 $Y2=0.74
r248 2 34 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.395 $X2=3.805 $Y2=0.605
r249 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.395 $X2=0.71 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_2%noxref_25 1 2 9 11 12 15
r35 13 15 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.265 $Y=0.425
+ $X2=3.265 $Y2=0.605
r36 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.1 $Y=0.34
+ $X2=3.265 $Y2=0.425
r37 11 12 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=3.1 $Y=0.34
+ $X2=1.345 $Y2=0.34
r38 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.345 $Y2=0.34
r39 7 9 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.22 $Y=0.425 $X2=1.22
+ $Y2=0.605
r40 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.395 $X2=3.265 $Y2=0.605
r41 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.395 $X2=1.26 $Y2=0.605
.ends


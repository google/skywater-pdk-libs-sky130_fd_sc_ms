* File: sky130_fd_sc_ms__fa_2.spice
* Created: Fri Aug 28 17:35:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fa_2.pex.spice"
.subckt sky130_fd_sc_ms__fa_2  VNB VPB A CIN B VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* B	B
* CIN	CIN
* A	A
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_A_M1023_g N_A_27_79#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.18315 AS=0.2109 PD=1.235 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75008.3 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_79#_M1005_d N_B_M1005_g N_VGND_M1023_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.18315 PD=1.31 PS=1.235 NRD=23.508 NRS=23.508 M=1 R=4.93333
+ SA=75000.9 SB=75007.7 A=0.111 P=1.78 MULT=1
MM1030 N_A_339_347#_M1030_d N_CIN_M1030_g N_A_27_79#_M1005_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=1.31 NRD=11.34 NRS=23.508 M=1 R=4.93333
+ SA=75001.6 SB=75007 A=0.111 P=1.78 MULT=1
MM1028 A_487_79# N_B_M1028_g N_A_339_347#_M1030_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1295 PD=0.98 PS=1.09 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75006.5 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_M1027_g A_487_79# VNB NLOWVT L=0.15 W=0.74 AD=0.1961
+ AS=0.0888 PD=1.27 PS=0.98 NRD=14.592 NRS=10.536 M=1 R=4.93333 SA=75002.5
+ SB=75006.1 A=0.111 P=1.78 MULT=1
MM1031 N_A_701_79#_M1031_d N_CIN_M1031_g N_VGND_M1027_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=1.27 NRD=0 NRS=25.944 M=1 R=4.93333 SA=75003.1
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_B_M1018_g N_A_701_79#_M1031_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.193975 AS=0.1036 PD=1.395 PS=1.02 NRD=33.588 NRS=0 M=1 R=4.93333
+ SA=75003.6 SB=75005 A=0.111 P=1.78 MULT=1
MM1021 N_A_701_79#_M1021_d N_A_M1021_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.193975 PD=1.16 PS=1.395 NRD=1.212 NRS=33.588 M=1 R=4.93333
+ SA=75004.2 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1001 N_A_995_347#_M1001_d N_A_339_347#_M1001_g N_A_701_79#_M1021_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=11.34 NRS=11.34 M=1
+ R=4.93333 SA=75004.7 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1024 A_1119_79# N_CIN_M1024_g N_A_995_347#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75005.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1002 A_1205_79# N_B_M1002_g A_1119_79# VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.1036 PD=0.98 PS=1.02 NRD=10.536 NRS=13.776 M=1 R=4.93333 SA=75005.7
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g A_1205_79# VNB NLOWVT L=0.15 W=0.74
+ AD=0.253662 AS=0.0888 PD=1.52 PS=0.98 NRD=23.508 NRS=10.536 M=1 R=4.93333
+ SA=75006.1 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1004 N_COUT_M1004_d N_A_339_347#_M1004_g N_VGND_M1003_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.253662 PD=1.02 PS=1.52 NRD=0 NRS=46.668 M=1 R=4.93333
+ SA=75006.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1012 N_COUT_M1004_d N_A_339_347#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.251275 PD=1.02 PS=1.515 NRD=0 NRS=46.14 M=1 R=4.93333
+ SA=75007.2 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1006 N_SUM_M1006_d N_A_995_347#_M1006_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.251275 PD=1.02 PS=1.515 NRD=0 NRS=46.14 M=1 R=4.93333
+ SA=75007.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_SUM_M1006_d N_A_995_347#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75008.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_27_378#_M1013_s VPB PSHORT L=0.18 W=1
+ AD=0.248562 AS=0.28 PD=1.625 PS=2.56 NRD=14.7553 NRS=0.3152 M=1 R=5.55556
+ SA=90000.2 SB=90007.1 A=0.18 P=2.36 MULT=1
MM1014 N_A_27_378#_M1014_d N_B_M1014_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.248562 PD=1.27 PS=1.625 NRD=0 NRS=23.6203 M=1 R=5.55556
+ SA=90000.7 SB=90006.8 A=0.18 P=2.36 MULT=1
MM1019 N_A_339_347#_M1019_d N_CIN_M1019_g N_A_27_378#_M1014_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.135 PD=1.56 PS=1.27 NRD=32.4853 NRS=0 M=1 R=5.55556
+ SA=90001.2 SB=90006.4 A=0.18 P=2.36 MULT=1
MM1022 A_487_347# N_B_M1022_g N_A_339_347#_M1019_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=1.56 NRD=12.7853 NRS=22.6353 M=1 R=5.55556 SA=90001.9
+ SB=90005.6 A=0.18 P=2.36 MULT=1
MM1025 N_VPWR_M1025_d N_A_M1025_g A_487_347# VPB PSHORT L=0.18 W=1 AD=0.1975
+ AS=0.12 PD=1.395 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90002.3 SB=90005.2
+ A=0.18 P=2.36 MULT=1
MM1026 N_A_686_347#_M1026_d N_CIN_M1026_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=1
+ AD=0.176062 AS=0.1975 PD=1.48 PS=1.395 NRD=0 NRS=23.6203 M=1 R=5.55556
+ SA=90002.9 SB=90004.6 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_686_347#_M1026_d VPB PSHORT L=0.18 W=1
+ AD=0.218562 AS=0.176062 PD=1.565 PS=1.48 NRD=3.9203 NRS=8.8453 M=1 R=5.55556
+ SA=90003 SB=90004.2 A=0.18 P=2.36 MULT=1
MM1009 N_A_686_347#_M1009_d N_A_M1009_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.218562 PD=1.27 PS=1.565 NRD=0 NRS=22.6353 M=1 R=5.55556
+ SA=90003.5 SB=90004 A=0.18 P=2.36 MULT=1
MM1016 N_A_995_347#_M1016_d N_A_339_347#_M1016_g N_A_686_347#_M1009_d VPB PSHORT
+ L=0.18 W=1 AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=10.8153 NRS=0 M=1 R=5.55556
+ SA=90004 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1020 A_1097_347# N_CIN_M1020_g N_A_995_347#_M1016_d VPB PSHORT L=0.18 W=1
+ AD=0.18735 AS=0.165 PD=1.465 PS=1.33 NRD=26.0631 NRS=0 M=1 R=5.55556
+ SA=90004.5 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1029 A_1205_368# N_B_M1029_g A_1097_347# VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.18735 PD=1.24 PS=1.465 NRD=12.7853 NRS=26.0631 M=1 R=5.55556 SA=90004.8
+ SB=90002.9 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_1205_368# VPB PSHORT L=0.18 W=1 AD=0.199811
+ AS=0.12 PD=1.42453 PS=1.24 NRD=23.64 NRS=12.7853 M=1 R=5.55556 SA=90005.3
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1007 N_COUT_M1007_d N_A_339_347#_M1007_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2044 AS=0.223789 PD=1.485 PS=1.59547 NRD=7.0329 NRS=0 M=1
+ R=6.22222 SA=90005.2 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1010 N_COUT_M1007_d N_A_339_347#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2044 AS=0.2856 PD=1.485 PS=1.63 NRD=7.8997 NRS=15.8191 M=1
+ R=6.22222 SA=90005.8 SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1011 N_SUM_M1011_d N_A_995_347#_M1011_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2856 PD=1.39 PS=1.63 NRD=0 NRS=24.625 M=1 R=6.22222
+ SA=90006.5 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1017 N_SUM_M1011_d N_A_995_347#_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=18.2244 P=22.93
c_86 VNB 0 1.3983e-19 $X=0 $Y=0
c_1247 A_1097_347# 0 1.35287e-19 $X=5.485 $Y=1.735
*
.include "sky130_fd_sc_ms__fa_2.pxi.spice"
*
.ends
*
*

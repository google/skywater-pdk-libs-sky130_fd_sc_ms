* File: sky130_fd_sc_ms__nand2b_4.spice
* Created: Wed Sep  2 12:13:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand2b_4.pex.spice"
.subckt sky130_fd_sc_ms__nand2b_4  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_N_M1010_g N_A_31_74#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_31_74#_M1000_g N_A_243_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1000_d N_A_31_74#_M1006_g N_A_243_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_A_31_74#_M1008_g N_A_243_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.15355 AS=0.1036 PD=1.155 PS=1.02 NRD=12.156 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75003 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1008_d N_A_31_74#_M1013_g N_A_243_74#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.15355 AS=0.1036 PD=1.155 PS=1.02 NRD=9.72 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1001 N_A_243_74#_M1013_s N_B_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_243_74#_M1003_d N_B_M1003_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_A_243_74#_M1003_d N_B_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.27935 PD=1.02 PS=1.495 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_A_243_74#_M1009_d N_B_M1009_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.27935 PD=2.05 PS=1.495 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_31_74#_M1002_d N_A_N_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.525 PD=1.11 PS=2.93 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.5
+ SB=90004.2 A=0.1512 P=2.04 MULT=1
MM1005 N_A_31_74#_M1002_d N_A_N_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1614 PD=1.11 PS=1.26429 NRD=0 NRS=18.7544 M=1 R=4.66667
+ SA=90001 SB=90003.8 A=0.1512 P=2.04 MULT=1
MM1011 N_VPWR_M1005_s N_A_31_74#_M1011_g N_Y_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2152 AS=0.364 PD=1.68571 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.2
+ SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_31_74#_M1014_g N_Y_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.8792 AS=0.364 PD=2.69 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1014_d VPB PSHORT L=0.18 W=1.12 AD=0.1624
+ AS=0.8792 PD=1.41 PS=2.69 NRD=2.6201 NRS=4.3931 M=1 R=6.22222 SA=90003.8
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1004_d N_B_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12 AD=0.1624
+ AS=0.3192 PD=1.41 PS=2.81 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX15_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__nand2b_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfxbp_1.spice
* Created: Fri Aug 28 17:24:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfxbp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfxbp_1  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_27_74#_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2017 AS=0.2109 PD=1.35 PS=2.05 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1017 N_A_208_368#_M1017_d N_A_27_74#_M1017_g N_VGND_M1025_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.3252 AS=0.2017 PD=2.59 PS=1.35 NRD=62.34 NRS=4.452 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1009 N_A_423_503#_M1009_d N_D_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.368725 PD=0.7 PS=2.64 NRD=0 NRS=235.116 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_546_447#_M1002_d N_A_27_74#_M1002_g N_A_423_503#_M1009_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0756875 AS=0.0588 PD=0.83 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1012 A_713_102# N_A_208_368#_M1012_g N_A_546_447#_M1002_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0756875 PD=0.63 PS=0.83 NRD=14.28 NRS=12.852 M=1 R=2.8
+ SA=75001.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_701_463#_M1005_g A_713_102# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125675 AS=0.0441 PD=1.03052 PS=0.63 NRD=69.768 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_701_463#_M1008_d N_A_546_447#_M1008_g N_VGND_M1005_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.11825 AS=0.164575 PD=1.13 PS=1.34948 NRD=34.908 NRS=3.264
+ M=1 R=3.66667 SA=75001.7 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1010 N_A_1005_120#_M1010_d N_A_208_368#_M1010_g N_A_701_463#_M1008_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.147026 AS=0.11825 PD=1.23608 PS=1.13 NRD=27.264
+ NRS=0 M=1 R=3.66667 SA=75001.8 SB=75001 A=0.0825 P=1.4 MULT=1
MM1020 A_1143_146# N_A_27_74#_M1020_g N_A_1005_120#_M1010_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.112274 PD=0.66 PS=0.943918 NRD=18.564 NRS=38.568 M=1
+ R=2.8 SA=75002.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1191_120#_M1013_g A_1143_146# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1005_120#_M1018_g N_A_1191_120#_M1018_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.11874 AS=0.15675 PD=0.989147 PS=1.67 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1006 N_Q_M1006_d N_A_1191_120#_M1006_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.15976 PD=2.05 PS=1.33085 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_1191_120#_M1022_g N_A_1644_112#_M1022_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1027 N_Q_N_M1027_d N_A_1644_112#_M1027_g N_VGND_M1022_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.144644 PD=2.05 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_CLK_M1015_g N_A_27_74#_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_A_208_368#_M1014_d N_A_27_74#_M1014_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1021 N_A_423_503#_M1021_d N_D_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=0.42
+ AD=0.140075 AS=0.2219 PD=1.305 PS=2.07 NRD=130.631 NRS=221.999 M=1 R=2.33333
+ SA=90000.3 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1026 N_A_546_447#_M1026_d N_A_208_368#_M1026_g N_A_423_503#_M1021_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.101237 AS=0.140075 PD=1.08 PS=1.305 NRD=0 NRS=130.631 M=1
+ R=2.33333 SA=90000.5 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1003 A_653_508# N_A_27_74#_M1003_g N_A_546_447#_M1026_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.101237 PD=0.66 PS=1.08 NRD=30.4759 NRS=87.2513 M=1
+ R=2.33333 SA=90000.5 SB=90002.8 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_701_463#_M1019_g A_653_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.14875 AS=0.0504 PD=1.12333 PS=0.66 NRD=53.9386 NRS=30.4759 M=1 R=2.33333
+ SA=90000.9 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1011 N_A_701_463#_M1011_d N_A_546_447#_M1011_g N_VPWR_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2415 AS=0.2975 PD=1.415 PS=2.24667 NRD=1.7533 NRS=70.1517
+ M=1 R=4.66667 SA=90001 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1023 N_A_1005_120#_M1023_d N_A_27_74#_M1023_g N_A_701_463#_M1011_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1752 AS=0.2415 PD=1.59333 PS=1.415 NRD=0 NRS=52.7566 M=1
+ R=4.66667 SA=90001.7 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1016 A_1161_482# N_A_208_368#_M1016_g N_A_1005_120#_M1023_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0876 PD=0.63 PS=0.796667 NRD=23.443 NRS=37.5088 M=1
+ R=2.33333 SA=90002.7 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_A_1191_120#_M1004_g A_1161_482# VPB PSHORT L=0.18 W=0.42
+ AD=0.1134 AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333 SA=90003
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1001 N_VPWR_M1001_d N_A_1005_120#_M1001_g N_A_1191_120#_M1001_s VPB PSHORT
+ L=0.18 W=1 AD=0.167453 AS=0.275 PD=1.36321 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1024 N_Q_M1024_d N_A_1191_120#_M1024_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.187547 PD=2.78 PS=1.52679 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_1191_120#_M1007_g N_A_1644_112#_M1007_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.2268 PD=1.23857 PS=2.22 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1000 N_Q_N_M1000_d N_A_1644_112#_M1000_g N_VPWR_M1007_d VPB PSHORT L=0.18
+ W=1.12 AD=0.308 AS=0.196 PD=2.79 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_206 VPB 0 8.5492e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dfxbp_1.pxi.spice"
*
.ends
*
*

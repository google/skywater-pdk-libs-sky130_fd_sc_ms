# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__or4b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__or4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.350000 2.275000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.470000 2.815000 2.150000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.470000 3.355000 2.520000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.350000 1.405000 1.130000 ;
        RECT 1.060000 1.130000 1.230000 1.820000 ;
        RECT 1.060000 1.820000 1.430000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.640000  0.085000 0.890000 0.840000 ;
        RECT 1.575000  0.085000 1.995000 0.780000 ;
        RECT 2.685000  0.085000 3.205000 0.780000 ;
        RECT 3.875000  0.085000 4.205000 0.930000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.650000 2.660000 0.980000 3.245000 ;
        RECT 1.550000 2.730000 2.125000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 1.950000 0.890000 2.320000 ;
      RECT 0.115000 2.320000 2.465000 2.490000 ;
      RECT 0.115000 2.490000 0.445000 2.700000 ;
      RECT 0.130000 0.540000 0.460000 1.010000 ;
      RECT 0.130000 1.010000 0.890000 1.180000 ;
      RECT 0.720000 1.180000 0.890000 1.950000 ;
      RECT 1.400000 1.300000 1.745000 1.630000 ;
      RECT 1.575000 0.960000 3.705000 1.100000 ;
      RECT 1.575000 1.100000 4.235000 1.130000 ;
      RECT 1.575000 1.130000 1.745000 1.300000 ;
      RECT 2.175000 0.450000 2.505000 0.960000 ;
      RECT 2.295000 2.490000 2.465000 2.690000 ;
      RECT 2.295000 2.690000 3.695000 2.860000 ;
      RECT 3.375000 0.450000 3.705000 0.960000 ;
      RECT 3.375000 1.130000 4.235000 1.270000 ;
      RECT 3.525000 1.440000 3.895000 1.770000 ;
      RECT 3.525000 1.770000 3.695000 2.690000 ;
      RECT 3.865000 1.940000 4.235000 2.980000 ;
      RECT 4.065000 1.270000 4.235000 1.940000 ;
  END
END sky130_fd_sc_ms__or4b_2

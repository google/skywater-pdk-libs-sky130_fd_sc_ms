# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o21a_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o21a_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.835000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.180000 1.385000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.955000 1.550000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.465000 1.720000 3.295000 1.890000 ;
        RECT 2.465000 1.890000 2.795000 2.980000 ;
        RECT 2.965000 0.350000 3.295000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
        RECT 0.750000  0.085000 1.235000 0.600000 ;
        RECT 2.465000  0.085000 2.795000 1.050000 ;
        RECT 3.475000  0.085000 3.725000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.840000 3.415000 ;
        RECT 0.335000 1.820000 0.665000 3.245000 ;
        RECT 1.965000 2.060000 2.295000 3.245000 ;
        RECT 2.965000 2.060000 3.295000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.250000 0.340000 0.580000 0.840000 ;
      RECT 0.250000 0.840000 1.735000 1.010000 ;
      RECT 1.325000 1.720000 2.295000 1.890000 ;
      RECT 1.325000 1.890000 1.655000 2.860000 ;
      RECT 1.405000 0.340000 1.735000 0.840000 ;
      RECT 1.905000 0.340000 2.295000 1.010000 ;
      RECT 2.125000 1.010000 2.295000 1.220000 ;
      RECT 2.125000 1.220000 2.645000 1.550000 ;
      RECT 2.125000 1.550000 2.295000 1.720000 ;
  END
END sky130_fd_sc_ms__o21a_2

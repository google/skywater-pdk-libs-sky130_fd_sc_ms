* File: sky130_fd_sc_ms__a221o_4.pxi.spice
* Created: Fri Aug 28 17:00:58 2020
* 
x_PM_SKY130_FD_SC_MS__A221O_4%A1 N_A1_M1009_g N_A1_c_157_n N_A1_M1016_g
+ N_A1_c_159_n N_A1_c_160_n N_A1_M1011_g N_A1_c_162_n N_A1_M1018_g N_A1_c_164_n
+ N_A1_c_165_n A1 A1 N_A1_c_167_n PM_SKY130_FD_SC_MS__A221O_4%A1
x_PM_SKY130_FD_SC_MS__A221O_4%A2 N_A2_M1001_g N_A2_M1022_g N_A2_M1003_g
+ N_A2_c_226_n N_A2_M1027_g N_A2_c_227_n A2 N_A2_c_229_n
+ PM_SKY130_FD_SC_MS__A221O_4%A2
x_PM_SKY130_FD_SC_MS__A221O_4%A_154_135# N_A_154_135#_M1009_d
+ N_A_154_135#_M1024_d N_A_154_135#_M1012_d N_A_154_135#_M1000_s
+ N_A_154_135#_c_302_n N_A_154_135#_M1006_g N_A_154_135#_c_287_n
+ N_A_154_135#_M1005_g N_A_154_135#_M1008_g N_A_154_135#_c_288_n
+ N_A_154_135#_M1015_g N_A_154_135#_M1010_g N_A_154_135#_c_289_n
+ N_A_154_135#_M1021_g N_A_154_135#_c_290_n N_A_154_135#_M1013_g
+ N_A_154_135#_c_291_n N_A_154_135#_M1023_g N_A_154_135#_c_292_n
+ N_A_154_135#_c_307_n N_A_154_135#_c_293_n N_A_154_135#_c_325_n
+ N_A_154_135#_c_294_n N_A_154_135#_c_295_n N_A_154_135#_c_296_n
+ N_A_154_135#_c_334_p N_A_154_135#_c_297_n N_A_154_135#_c_363_p
+ N_A_154_135#_c_298_n N_A_154_135#_c_299_n N_A_154_135#_c_300_n
+ N_A_154_135#_c_301_n PM_SKY130_FD_SC_MS__A221O_4%A_154_135#
x_PM_SKY130_FD_SC_MS__A221O_4%C1 N_C1_M1024_g N_C1_M1000_g N_C1_M1025_g
+ N_C1_c_497_n N_C1_c_498_n N_C1_c_499_n N_C1_M1026_g C1 C1
+ PM_SKY130_FD_SC_MS__A221O_4%C1
x_PM_SKY130_FD_SC_MS__A221O_4%B2 N_B2_M1017_g N_B2_M1002_g N_B2_c_563_n
+ N_B2_c_564_n N_B2_c_565_n N_B2_M1019_g N_B2_M1004_g N_B2_c_567_n N_B2_c_568_n
+ N_B2_c_569_n N_B2_c_570_n N_B2_c_571_n B2 N_B2_c_572_n N_B2_c_573_n
+ PM_SKY130_FD_SC_MS__A221O_4%B2
x_PM_SKY130_FD_SC_MS__A221O_4%B1 N_B1_M1007_g N_B1_M1012_g N_B1_M1014_g
+ N_B1_M1020_g N_B1_c_658_n B1 B1 N_B1_c_660_n N_B1_c_666_n
+ PM_SKY130_FD_SC_MS__A221O_4%B1
x_PM_SKY130_FD_SC_MS__A221O_4%VPWR N_VPWR_M1016_d N_VPWR_M1018_d N_VPWR_M1003_s
+ N_VPWR_M1008_s N_VPWR_M1013_s N_VPWR_c_708_n N_VPWR_c_709_n N_VPWR_c_710_n
+ N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_713_n N_VPWR_c_714_n N_VPWR_c_715_n
+ N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_718_n N_VPWR_c_719_n VPWR
+ N_VPWR_c_720_n N_VPWR_c_721_n N_VPWR_c_707_n N_VPWR_c_723_n
+ PM_SKY130_FD_SC_MS__A221O_4%VPWR
x_PM_SKY130_FD_SC_MS__A221O_4%A_160_376# N_A_160_376#_M1016_s
+ N_A_160_376#_M1001_d N_A_160_376#_M1002_d N_A_160_376#_M1007_d
+ N_A_160_376#_c_802_n N_A_160_376#_c_796_n N_A_160_376#_c_797_n
+ N_A_160_376#_c_820_n N_A_160_376#_c_798_n N_A_160_376#_c_799_n
+ N_A_160_376#_c_800_n N_A_160_376#_c_838_n N_A_160_376#_c_801_n
+ PM_SKY130_FD_SC_MS__A221O_4%A_160_376#
x_PM_SKY130_FD_SC_MS__A221O_4%X N_X_M1005_d N_X_M1021_d N_X_M1006_d N_X_M1010_d
+ N_X_c_891_n N_X_c_902_n N_X_c_914_n N_X_c_920_n N_X_c_884_n N_X_c_926_n
+ N_X_c_885_n N_X_c_893_n N_X_c_935_n N_X_c_886_n N_X_c_887_n N_X_c_888_n X
+ N_X_c_890_n PM_SKY130_FD_SC_MS__A221O_4%X
x_PM_SKY130_FD_SC_MS__A221O_4%A_1102_392# N_A_1102_392#_M1000_d
+ N_A_1102_392#_M1026_d N_A_1102_392#_M1004_s N_A_1102_392#_M1014_s
+ N_A_1102_392#_c_1004_n N_A_1102_392#_c_1005_n N_A_1102_392#_c_1016_n
+ N_A_1102_392#_c_1006_n N_A_1102_392#_c_1007_n N_A_1102_392#_c_1008_n
+ N_A_1102_392#_c_1009_n PM_SKY130_FD_SC_MS__A221O_4%A_1102_392#
x_PM_SKY130_FD_SC_MS__A221O_4%A_71_135# N_A_71_135#_M1009_s N_A_71_135#_M1011_s
+ N_A_71_135#_M1022_d N_A_71_135#_c_1049_n N_A_71_135#_c_1054_n
+ N_A_71_135#_c_1046_n N_A_71_135#_c_1047_n N_A_71_135#_c_1065_n
+ N_A_71_135#_c_1048_n PM_SKY130_FD_SC_MS__A221O_4%A_71_135#
x_PM_SKY130_FD_SC_MS__A221O_4%VGND N_VGND_M1022_s N_VGND_M1027_s N_VGND_M1015_s
+ N_VGND_M1023_s N_VGND_M1025_s N_VGND_M1019_s N_VGND_c_1099_n N_VGND_c_1100_n
+ N_VGND_c_1101_n N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n
+ N_VGND_c_1105_n N_VGND_c_1106_n N_VGND_c_1107_n N_VGND_c_1108_n
+ N_VGND_c_1109_n N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1162_n VGND N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n
+ N_VGND_c_1116_n N_VGND_c_1117_n N_VGND_c_1118_n N_VGND_c_1119_n
+ N_VGND_c_1120_n PM_SKY130_FD_SC_MS__A221O_4%VGND
x_PM_SKY130_FD_SC_MS__A221O_4%A_1346_123# N_A_1346_123#_M1017_d
+ N_A_1346_123#_M1012_s N_A_1346_123#_M1020_s N_A_1346_123#_c_1258_n
+ N_A_1346_123#_c_1241_n N_A_1346_123#_c_1242_n N_A_1346_123#_c_1243_n
+ N_A_1346_123#_c_1244_n N_A_1346_123#_c_1245_n N_A_1346_123#_c_1246_n
+ PM_SKY130_FD_SC_MS__A221O_4%A_1346_123#
cc_1 VNB N_A1_M1009_g 0.0126596f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.995
cc_2 VNB N_A1_c_157_n 0.00582894f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.48
cc_3 VNB N_A1_M1016_g 0.0105088f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.38
cc_4 VNB N_A1_c_159_n 0.0143467f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.49
cc_5 VNB N_A1_c_160_n 0.0150623f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.49
cc_6 VNB N_A1_M1011_g 0.0108339f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_7 VNB N_A1_c_162_n 0.0202489f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.54
cc_8 VNB N_A1_M1018_g 0.00763938f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_9 VNB N_A1_c_164_n 0.0147864f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.49
cc_10 VNB N_A1_c_165_n 0.0067715f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.49
cc_11 VNB A1 0.0189889f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_12 VNB N_A1_c_167_n 0.0454186f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_13 VNB N_A2_M1001_g 0.0112412f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.995
cc_14 VNB N_A2_M1022_g 0.0102533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1003_g 0.0104206f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.565
cc_16 VNB N_A2_c_226_n 0.014937f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_17 VNB N_A2_c_227_n 0.0415399f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.49
cc_18 VNB A2 0.00844479f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.49
cc_19 VNB N_A2_c_229_n 0.0443821f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.465
cc_20 VNB N_A_154_135#_c_287_n 0.0179122f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_21 VNB N_A_154_135#_c_288_n 0.0160784f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_22 VNB N_A_154_135#_c_289_n 0.0162363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_154_135#_c_290_n 0.077093f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_24 VNB N_A_154_135#_c_291_n 0.0189669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_154_135#_c_292_n 3.931e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_154_135#_c_293_n 3.95392e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_154_135#_c_294_n 0.0194191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_154_135#_c_295_n 0.00345068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_154_135#_c_296_n 0.00212477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_154_135#_c_297_n 0.0123759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_154_135#_c_298_n 0.0118549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_154_135#_c_299_n 0.00492041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_154_135#_c_300_n 0.0061434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_154_135#_c_301_n 0.00193979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C1_M1024_g 0.0238103f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.995
cc_36 VNB N_C1_M1025_g 0.0228799f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.565
cc_37 VNB N_C1_c_497_n 0.00943777f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_38 VNB N_C1_c_498_n 0.0278067f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_39 VNB N_C1_c_499_n 0.0157726f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.54
cc_40 VNB N_B2_c_563_n 0.059418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_B2_c_564_n 0.00510297f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=0.49
cc_42 VNB N_B2_c_565_n 0.00523521f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.565
cc_43 VNB N_B2_M1019_g 0.0282044f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=0.995
cc_44 VNB N_B2_c_567_n 0.00756482f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.39
cc_45 VNB N_B2_c_568_n 0.0604594f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_46 VNB N_B2_c_569_n 0.00422613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_B2_c_570_n 0.0139812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_B2_c_571_n 0.00620432f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_49 VNB N_B2_c_572_n 0.0468869f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.602
cc_50 VNB N_B2_c_573_n 0.0168974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_B1_M1012_g 0.0277209f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.38
cc_52 VNB N_B1_M1020_g 0.0306491f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.54
cc_53 VNB N_B1_c_658_n 0.0346933f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_54 VNB B1 0.035572f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_55 VNB N_B1_c_660_n 0.062292f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_56 VNB N_VPWR_c_707_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_884_n 0.00279061f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.465
cc_58 VNB N_X_c_885_n 0.00252589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_X_c_886_n 0.0161413f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.49
cc_60 VNB N_X_c_887_n 0.0195019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_X_c_888_n 0.0221701f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.925
cc_62 VNB X 0.00470385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_X_c_890_n 0.00409571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_71_135#_c_1046_n 0.0132978f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_65 VNB N_A_71_135#_c_1047_n 8.4331e-19 $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.38
cc_66 VNB N_A_71_135#_c_1048_n 0.0171478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1099_n 0.0138474f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.49
cc_68 VNB N_VGND_c_1100_n 0.0162981f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.465
cc_69 VNB N_VGND_c_1101_n 0.0140948f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.47
cc_70 VNB N_VGND_c_1102_n 0.0259638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1103_n 0.0184531f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=0.4
cc_72 VNB N_VGND_c_1104_n 0.00304657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1105_n 0.0106636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1106_n 0.0562111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1107_n 0.00326288f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.41
cc_76 VNB N_VGND_c_1108_n 0.00840773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1109_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1110_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1111_n 0.0202649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1112_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1113_n 0.022977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1114_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1115_n 0.0218123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1116_n 0.0572372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1117_n 0.55948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1118_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1119_n 0.013849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1120_n 0.00351416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1346_123#_c_1241_n 0.0126797f $X=-0.19 $Y=-0.245 $X2=1.125
+ $Y2=0.995
cc_90 VNB N_A_1346_123#_c_1242_n 0.00246562f $X=-0.19 $Y=-0.245 $X2=1.28
+ $Y2=1.54
cc_91 VNB N_A_1346_123#_c_1243_n 0.00912157f $X=-0.19 $Y=-0.245 $X2=1.435
+ $Y2=0.49
cc_92 VNB N_A_1346_123#_c_1244_n 0.0127125f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.49
cc_93 VNB N_A_1346_123#_c_1245_n 0.00355281f $X=-0.19 $Y=-0.245 $X2=0.71
+ $Y2=1.39
cc_94 VNB N_A_1346_123#_c_1246_n 0.0255734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VPB N_A1_M1016_g 0.0277916f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=2.38
cc_96 VPB N_A1_M1018_g 0.0288755f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_97 VPB N_A2_M1001_g 0.0272841f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=0.995
cc_98 VPB N_A2_M1003_g 0.0250555f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.565
cc_99 VPB N_A_154_135#_c_302_n 0.0173731f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_100 VPB N_A_154_135#_M1008_g 0.0197006f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.39
cc_101 VPB N_A_154_135#_M1010_g 0.0197006f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=0.84
cc_102 VPB N_A_154_135#_c_290_n 0.0196242f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_103 VPB N_A_154_135#_M1013_g 0.0254624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_154_135#_c_307_n 0.00260596f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.41
cc_105 VPB N_A_154_135#_c_293_n 0.00563034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_154_135#_c_297_n 0.0099801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_154_135#_c_298_n 0.0179164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_154_135#_c_299_n 0.00399505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_C1_M1000_g 0.0227256f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=2.38
cc_110 VPB N_C1_c_498_n 0.0260115f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_111 VPB N_C1_c_499_n 0.00246962f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.54
cc_112 VPB N_C1_M1026_g 0.0240917f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_113 VPB C1 0.015703f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.49
cc_114 VPB N_B2_M1002_g 0.0220449f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=2.38
cc_115 VPB N_B2_c_564_n 0.00346162f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=0.49
cc_116 VPB N_B2_c_565_n 0.00369935f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.565
cc_117 VPB N_B2_M1004_g 0.0247393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B2_c_569_n 0.0151793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_B1_M1007_g 0.0279747f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=0.995
cc_120 VPB N_B1_M1014_g 0.0333679f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.565
cc_121 VPB N_B1_c_658_n 0.0113125f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_122 VPB B1 0.019573f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.465
cc_123 VPB N_B1_c_660_n 0.026591f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=0.47
cc_124 VPB N_B1_c_666_n 0.0125041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_708_n 0.0409052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_709_n 0.00877473f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.49
cc_127 VPB N_VPWR_c_710_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_711_n 0.0112086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_712_n 0.0123263f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_130 VPB N_VPWR_c_713_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_131 VPB N_VPWR_c_714_n 0.0225995f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.49
cc_132 VPB N_VPWR_c_715_n 0.00612909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_716_n 0.0177589f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.602
cc_134 VPB N_VPWR_c_717_n 0.00601813f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.925
cc_135 VPB N_VPWR_c_718_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_719_n 0.00611614f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.41
cc_137 VPB N_VPWR_c_720_n 0.0214857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_721_n 0.116897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_707_n 0.134978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_723_n 0.0346226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_160_376#_c_796_n 0.0295027f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=0.49
cc_142 VPB N_A_160_376#_c_797_n 0.00224119f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.39
cc_143 VPB N_A_160_376#_c_798_n 0.00421146f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.465
cc_144 VPB N_A_160_376#_c_799_n 0.00314826f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=0.84
cc_145 VPB N_A_160_376#_c_800_n 0.0026444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_160_376#_c_801_n 0.00250461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_X_c_891_n 0.016621f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=0.995
cc_148 VPB N_X_c_888_n 0.0139957f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=0.925
cc_149 VPB N_A_1102_392#_c_1004_n 0.0117214f $X=-0.19 $Y=1.66 $X2=1.125
+ $Y2=0.995
cc_150 VPB N_A_1102_392#_c_1005_n 0.00280532f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.38
cc_151 VPB N_A_1102_392#_c_1006_n 0.012632f $X=-0.19 $Y=1.66 $X2=1.125 $Y2=1.465
cc_152 VPB N_A_1102_392#_c_1007_n 0.0381637f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=0.47
cc_153 VPB N_A_1102_392#_c_1008_n 0.00113322f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_154 VPB N_A_1102_392#_c_1009_n 0.00325298f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=0.4
cc_155 N_A1_M1018_g N_A2_M1001_g 0.00963031f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_156 N_A1_c_167_n N_A2_M1022_g 7.29007e-19 $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_157 N_A1_c_162_n N_A2_c_227_n 0.00963031f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_158 N_A1_c_167_n N_A2_c_229_n 0.00509489f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_159 N_A1_M1009_g N_A_154_135#_c_292_n 0.00834817f $X=0.695 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A1_c_157_n N_A_154_135#_c_292_n 0.0033001f $X=0.71 $Y=1.48 $X2=0 $Y2=0
cc_161 N_A1_M1016_g N_A_154_135#_c_292_n 0.00299664f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_162 N_A1_M1011_g N_A_154_135#_c_292_n 0.00409333f $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A1_c_162_n N_A_154_135#_c_292_n 0.00830365f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_164 N_A1_M1018_g N_A_154_135#_c_292_n 0.0010381f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_165 N_A1_M1016_g N_A_154_135#_c_307_n 0.00667657f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_166 N_A1_c_162_n N_A_154_135#_c_298_n 0.0042433f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_167 N_A1_M1018_g N_A_154_135#_c_298_n 0.0142546f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_168 N_A1_M1016_g N_VPWR_c_708_n 0.014279f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_169 N_A1_M1018_g N_VPWR_c_708_n 6.94553e-19 $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_170 N_A1_M1016_g N_VPWR_c_720_n 0.00519349f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_171 N_A1_M1018_g N_VPWR_c_720_n 0.00597358f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_172 N_A1_M1016_g N_VPWR_c_707_n 0.00524044f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_173 N_A1_M1018_g N_VPWR_c_707_n 0.00624688f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_174 N_A1_M1018_g N_VPWR_c_723_n 0.00443101f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_175 N_A1_M1018_g N_A_160_376#_c_802_n 0.0142149f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_176 N_A1_M1016_g N_A_160_376#_c_799_n 0.00624529f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_177 N_A1_M1018_g N_A_160_376#_c_799_n 0.0127296f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_178 N_A1_M1016_g N_X_c_893_n 0.0199318f $X=0.71 $Y=2.38 $X2=0 $Y2=0
cc_179 N_A1_c_162_n N_X_c_893_n 2.0859e-19 $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_180 N_A1_M1018_g N_X_c_893_n 0.0138687f $X=1.28 $Y=2.38 $X2=0 $Y2=0
cc_181 N_A1_M1009_g N_X_c_886_n 0.00525441f $X=0.695 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_M1011_g N_X_c_886_n 0.00455416f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A1_c_162_n N_X_c_886_n 0.00166958f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_184 A1 N_X_c_886_n 0.00437127f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_185 N_A1_M1009_g N_X_c_887_n 0.00206546f $X=0.695 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A1_M1009_g N_X_c_888_n 0.0159795f $X=0.695 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_M1009_g N_A_71_135#_c_1049_n 0.0102992f $X=0.695 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A1_c_159_n N_A_71_135#_c_1049_n 0.00238533f $X=1.05 $Y=0.49 $X2=0 $Y2=0
cc_189 N_A1_M1011_g N_A_71_135#_c_1049_n 0.0131077f $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A1_c_164_n N_A_71_135#_c_1049_n 0.00448161f $X=1.435 $Y=0.49 $X2=0
+ $Y2=0
cc_191 A1 N_A_71_135#_c_1049_n 0.0140569f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_192 A1 N_A_71_135#_c_1054_n 0.00994896f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_193 N_A1_c_164_n N_A_71_135#_c_1046_n 0.00234729f $X=1.435 $Y=0.49 $X2=0
+ $Y2=0
cc_194 A1 N_A_71_135#_c_1046_n 0.0131478f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_195 N_A1_c_167_n N_A_71_135#_c_1046_n 3.82631e-19 $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_196 N_A1_M1011_g N_A_71_135#_c_1047_n 0.00288366f $X=1.125 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A1_c_162_n N_A_71_135#_c_1047_n 0.00529894f $X=1.28 $Y=1.54 $X2=0 $Y2=0
cc_198 N_A1_M1009_g N_A_71_135#_c_1048_n 7.91278e-19 $X=0.695 $Y=0.995 $X2=0
+ $Y2=0
cc_199 A1 N_VGND_c_1099_n 0.0315455f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A1_c_167_n N_VGND_c_1099_n 0.00162808f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_201 N_A1_c_160_n N_VGND_c_1106_n 0.0175556f $X=0.77 $Y=0.49 $X2=0 $Y2=0
cc_202 A1 N_VGND_c_1106_n 0.021134f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_203 N_A1_c_167_n N_VGND_c_1106_n 0.0056689f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_204 A1 N_VGND_c_1108_n 0.0294117f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_205 N_A1_c_160_n N_VGND_c_1117_n 0.0244466f $X=0.77 $Y=0.49 $X2=0 $Y2=0
cc_206 A1 N_VGND_c_1117_n 0.011067f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_207 N_A1_c_167_n N_VGND_c_1117_n 0.00759015f $X=1.6 $Y=0.4 $X2=0 $Y2=0
cc_208 N_A2_c_226_n N_A_154_135#_c_287_n 0.0131106f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_209 N_A2_c_229_n N_A_154_135#_c_287_n 0.00102307f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_210 N_A2_M1003_g N_A_154_135#_c_290_n 0.036974f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_211 N_A2_c_227_n N_A_154_135#_c_290_n 0.0131106f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_212 N_A2_c_227_n N_A_154_135#_c_325_n 3.22675e-19 $X=2.89 $Y=1.405 $X2=0
+ $Y2=0
cc_213 N_A2_M1001_g N_A_154_135#_c_298_n 0.0131515f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_214 N_A2_M1003_g N_A_154_135#_c_298_n 0.0124128f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_215 N_A2_c_227_n N_A_154_135#_c_298_n 0.0127287f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_216 N_A2_M1003_g N_VPWR_c_709_n 0.00488167f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_217 N_A2_M1001_g N_VPWR_c_714_n 0.00597358f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_218 N_A2_M1003_g N_VPWR_c_714_n 0.00597358f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_219 N_A2_M1001_g N_VPWR_c_707_n 0.00624688f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_220 N_A2_M1003_g N_VPWR_c_707_n 0.00624688f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_221 N_A2_M1001_g N_VPWR_c_723_n 0.00445916f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_222 N_A2_M1001_g N_A_160_376#_c_802_n 0.0142149f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_223 N_A2_M1003_g N_A_160_376#_c_796_n 0.0109354f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_224 N_A2_M1001_g N_A_160_376#_c_800_n 0.0130222f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_225 N_A2_M1003_g N_A_160_376#_c_800_n 0.0104356f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_226 N_A2_M1003_g N_X_c_902_n 0.00302381f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_227 N_A2_c_226_n N_X_c_884_n 6.23275e-19 $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_228 N_A2_M1001_g N_X_c_893_n 0.0132193f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_229 N_A2_M1003_g N_X_c_893_n 0.0129917f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_230 N_A2_M1022_g N_X_c_886_n 0.00540271f $X=2.46 $Y=0.935 $X2=0 $Y2=0
cc_231 N_A2_c_226_n N_X_c_886_n 0.00725658f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_232 N_A2_c_227_n N_X_c_886_n 0.00189607f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_233 A2 N_X_c_886_n 8.85114e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_234 N_A2_c_226_n X 7.93272e-19 $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_235 N_A2_c_227_n X 8.83029e-19 $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_236 N_A2_c_226_n N_X_c_890_n 0.00276942f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_237 A2 N_A_71_135#_M1022_d 0.00219033f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_238 N_A2_M1022_g N_A_71_135#_c_1046_n 0.0070549f $X=2.46 $Y=0.935 $X2=0 $Y2=0
cc_239 N_A2_c_226_n N_A_71_135#_c_1046_n 6.08595e-19 $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_240 N_A2_c_227_n N_A_71_135#_c_1046_n 0.0232248f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_241 N_A2_M1022_g N_A_71_135#_c_1065_n 0.00996461f $X=2.46 $Y=0.935 $X2=0
+ $Y2=0
cc_242 A2 N_A_71_135#_c_1065_n 0.0145781f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_243 N_A2_c_229_n N_A_71_135#_c_1065_n 2.47224e-19 $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_244 N_A2_M1022_g N_VGND_c_1099_n 0.00270215f $X=2.46 $Y=0.935 $X2=0 $Y2=0
cc_245 A2 N_VGND_c_1099_n 0.0255727f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_246 N_A2_c_229_n N_VGND_c_1099_n 0.00308142f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_247 N_A2_c_226_n N_VGND_c_1100_n 0.00240899f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_248 A2 N_VGND_c_1100_n 0.0246703f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_249 N_A2_c_229_n N_VGND_c_1100_n 0.00262568f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_250 N_A2_c_227_n N_VGND_c_1108_n 0.00144156f $X=2.89 $Y=1.405 $X2=0 $Y2=0
cc_251 A2 N_VGND_c_1108_n 0.0039865f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_252 N_A2_c_229_n N_VGND_c_1108_n 4.08097e-19 $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_253 N_A2_c_226_n N_VGND_c_1113_n 0.00420632f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_254 A2 N_VGND_c_1113_n 0.0315176f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_255 N_A2_c_229_n N_VGND_c_1113_n 0.00659434f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_256 N_A2_c_226_n N_VGND_c_1117_n 0.00472204f $X=2.89 $Y=1.33 $X2=0 $Y2=0
cc_257 A2 N_VGND_c_1117_n 0.0168113f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_258 N_A2_c_229_n N_VGND_c_1117_n 0.0103546f $X=2.44 $Y=0.34 $X2=0 $Y2=0
cc_259 N_A_154_135#_c_294_n N_C1_M1024_g 0.0128795f $X=5.61 $Y=1.215 $X2=0 $Y2=0
cc_260 N_A_154_135#_c_295_n N_C1_M1024_g 0.0119691f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_261 N_A_154_135#_c_296_n N_C1_M1024_g 8.66403e-19 $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_262 N_A_154_135#_c_299_n N_C1_M1024_g 0.00339201f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_263 N_A_154_135#_c_300_n N_C1_M1024_g 0.00142589f $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_264 N_A_154_135#_c_334_p N_C1_M1000_g 0.00824847f $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_265 N_A_154_135#_c_295_n N_C1_M1025_g 0.00714623f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_266 N_A_154_135#_c_296_n N_C1_M1025_g 0.00509715f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_267 N_A_154_135#_c_300_n N_C1_M1025_g 0.0109783f $X=5.85 $Y=1.215 $X2=0 $Y2=0
cc_268 N_A_154_135#_c_296_n N_C1_c_497_n 0.00730338f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_269 N_A_154_135#_c_301_n N_C1_c_497_n 0.00190788f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_270 N_A_154_135#_c_290_n N_C1_c_498_n 8.07662e-19 $X=4.585 $Y=1.69 $X2=0
+ $Y2=0
cc_271 N_A_154_135#_c_294_n N_C1_c_498_n 0.00190609f $X=5.61 $Y=1.215 $X2=0
+ $Y2=0
cc_272 N_A_154_135#_c_296_n N_C1_c_498_n 0.00580359f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_273 N_A_154_135#_c_334_p N_C1_c_498_n 8.41656e-19 $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_274 N_A_154_135#_c_299_n N_C1_c_498_n 0.00556938f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_275 N_A_154_135#_c_300_n N_C1_c_498_n 0.00463795f $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_276 N_A_154_135#_c_301_n N_C1_c_498_n 0.00502274f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_277 N_A_154_135#_c_297_n N_C1_c_499_n 0.00521072f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_278 N_A_154_135#_c_301_n N_C1_c_499_n 0.00224569f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_279 N_A_154_135#_c_334_p N_C1_M1026_g 0.0106082f $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_280 N_A_154_135#_c_297_n N_C1_M1026_g 0.00537582f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_281 N_A_154_135#_c_301_n N_C1_M1026_g 7.77448e-19 $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_282 N_A_154_135#_c_294_n C1 0.015801f $X=5.61 $Y=1.215 $X2=0 $Y2=0
cc_283 N_A_154_135#_c_296_n C1 0.00864364f $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_284 N_A_154_135#_c_334_p C1 0.0205379f $X=6.085 $Y=2.105 $X2=0 $Y2=0
cc_285 N_A_154_135#_c_299_n C1 0.00900014f $X=4.795 $Y=1.215 $X2=0 $Y2=0
cc_286 N_A_154_135#_c_300_n C1 0.0109932f $X=5.85 $Y=1.215 $X2=0 $Y2=0
cc_287 N_A_154_135#_c_301_n C1 0.0126759f $X=6.085 $Y=1.685 $X2=0 $Y2=0
cc_288 N_A_154_135#_c_297_n N_B2_c_564_n 0.00596468f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_289 N_A_154_135#_c_334_p N_B2_c_565_n 0.00153877f $X=6.085 $Y=2.105 $X2=0
+ $Y2=0
cc_290 N_A_154_135#_c_297_n N_B2_c_565_n 0.0104635f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_291 N_A_154_135#_c_297_n N_B2_M1019_g 0.00307374f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_292 N_A_154_135#_c_297_n N_B2_c_567_n 0.00290892f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_293 N_A_154_135#_c_363_p N_B2_c_567_n 5.1726e-19 $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_294 N_A_154_135#_c_363_p N_B2_c_568_n 2.91453e-19 $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_295 N_A_154_135#_c_297_n N_B2_c_569_n 0.0150798f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_296 N_A_154_135#_c_297_n N_B2_c_570_n 0.00279407f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_297 N_A_154_135#_c_363_p N_B2_c_570_n 2.5461e-19 $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_298 N_A_154_135#_c_296_n N_B2_c_573_n 5.938e-19 $X=6.005 $Y=1.6 $X2=0 $Y2=0
cc_299 N_A_154_135#_c_297_n N_B2_c_573_n 0.00433746f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_300 N_A_154_135#_c_300_n N_B2_c_573_n 2.42029e-19 $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_301 N_A_154_135#_c_297_n N_B1_M1007_g 0.00451089f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_302 N_A_154_135#_c_363_p N_B1_M1012_g 0.0136043f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_303 N_A_154_135#_c_297_n N_B1_M1014_g 0.00601804f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_304 N_A_154_135#_c_363_p N_B1_M1020_g 0.0186666f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_305 N_A_154_135#_c_297_n N_B1_c_658_n 0.019752f $X=8.115 $Y=1.685 $X2=0 $Y2=0
cc_306 N_A_154_135#_c_363_p N_B1_c_658_n 0.0180593f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_307 N_A_154_135#_c_363_p B1 0.00257795f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_308 N_A_154_135#_c_297_n N_B1_c_666_n 0.012701f $X=8.115 $Y=1.685 $X2=0 $Y2=0
cc_309 N_A_154_135#_c_363_p N_B1_c_666_n 0.0238299f $X=8.28 $Y=0.76 $X2=0 $Y2=0
cc_310 N_A_154_135#_c_302_n N_VPWR_c_709_n 0.0107275f $X=3.235 $Y=1.78 $X2=0
+ $Y2=0
cc_311 N_A_154_135#_M1008_g N_VPWR_c_709_n 0.00114128f $X=3.685 $Y=2.4 $X2=0
+ $Y2=0
cc_312 N_A_154_135#_c_302_n N_VPWR_c_710_n 0.00114128f $X=3.235 $Y=1.78 $X2=0
+ $Y2=0
cc_313 N_A_154_135#_M1008_g N_VPWR_c_710_n 0.00995427f $X=3.685 $Y=2.4 $X2=0
+ $Y2=0
cc_314 N_A_154_135#_M1010_g N_VPWR_c_710_n 0.00995427f $X=4.135 $Y=2.4 $X2=0
+ $Y2=0
cc_315 N_A_154_135#_M1013_g N_VPWR_c_710_n 0.00114128f $X=4.585 $Y=2.4 $X2=0
+ $Y2=0
cc_316 N_A_154_135#_M1010_g N_VPWR_c_711_n 0.00114128f $X=4.135 $Y=2.4 $X2=0
+ $Y2=0
cc_317 N_A_154_135#_M1013_g N_VPWR_c_711_n 0.0110558f $X=4.585 $Y=2.4 $X2=0
+ $Y2=0
cc_318 N_A_154_135#_c_302_n N_VPWR_c_716_n 0.00460063f $X=3.235 $Y=1.78 $X2=0
+ $Y2=0
cc_319 N_A_154_135#_M1008_g N_VPWR_c_716_n 0.00460063f $X=3.685 $Y=2.4 $X2=0
+ $Y2=0
cc_320 N_A_154_135#_M1010_g N_VPWR_c_718_n 0.00460063f $X=4.135 $Y=2.4 $X2=0
+ $Y2=0
cc_321 N_A_154_135#_M1013_g N_VPWR_c_718_n 0.00460063f $X=4.585 $Y=2.4 $X2=0
+ $Y2=0
cc_322 N_A_154_135#_c_302_n N_VPWR_c_707_n 0.00450805f $X=3.235 $Y=1.78 $X2=0
+ $Y2=0
cc_323 N_A_154_135#_M1008_g N_VPWR_c_707_n 0.00450805f $X=3.685 $Y=2.4 $X2=0
+ $Y2=0
cc_324 N_A_154_135#_M1010_g N_VPWR_c_707_n 0.00450805f $X=4.135 $Y=2.4 $X2=0
+ $Y2=0
cc_325 N_A_154_135#_M1013_g N_VPWR_c_707_n 0.00450805f $X=4.585 $Y=2.4 $X2=0
+ $Y2=0
cc_326 N_A_154_135#_M1000_s N_A_160_376#_c_796_n 0.00329261f $X=5.95 $Y=1.96
+ $X2=0 $Y2=0
cc_327 N_A_154_135#_c_302_n N_A_160_376#_c_796_n 0.0137027f $X=3.235 $Y=1.78
+ $X2=0 $Y2=0
cc_328 N_A_154_135#_M1008_g N_A_160_376#_c_796_n 0.0129434f $X=3.685 $Y=2.4
+ $X2=0 $Y2=0
cc_329 N_A_154_135#_M1010_g N_A_160_376#_c_796_n 0.0129434f $X=4.135 $Y=2.4
+ $X2=0 $Y2=0
cc_330 N_A_154_135#_M1013_g N_A_160_376#_c_796_n 0.0171425f $X=4.585 $Y=2.4
+ $X2=0 $Y2=0
cc_331 N_A_154_135#_c_293_n N_A_160_376#_c_796_n 0.00439276f $X=4.71 $Y=1.55
+ $X2=0 $Y2=0
cc_332 N_A_154_135#_c_334_p N_A_160_376#_c_796_n 0.0169324f $X=6.085 $Y=2.105
+ $X2=0 $Y2=0
cc_333 N_A_154_135#_c_297_n N_A_160_376#_c_796_n 0.0137719f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_334 N_A_154_135#_c_299_n N_A_160_376#_c_796_n 0.00522344f $X=4.795 $Y=1.215
+ $X2=0 $Y2=0
cc_335 N_A_154_135#_c_334_p N_A_160_376#_c_797_n 0.00499291f $X=6.085 $Y=2.105
+ $X2=0 $Y2=0
cc_336 N_A_154_135#_c_297_n N_A_160_376#_c_797_n 0.0262439f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_337 N_A_154_135#_c_334_p N_A_160_376#_c_820_n 0.00220201f $X=6.085 $Y=2.105
+ $X2=0 $Y2=0
cc_338 N_A_154_135#_c_297_n N_A_160_376#_c_798_n 0.0614905f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_339 N_A_154_135#_c_302_n N_A_160_376#_c_800_n 9.64229e-19 $X=3.235 $Y=1.78
+ $X2=0 $Y2=0
cc_340 N_A_154_135#_c_297_n N_A_160_376#_c_801_n 0.0331386f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_341 N_A_154_135#_c_325_n N_X_c_902_n 0.0750761f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_342 N_A_154_135#_c_302_n N_X_c_914_n 0.0135495f $X=3.235 $Y=1.78 $X2=0 $Y2=0
cc_343 N_A_154_135#_M1008_g N_X_c_914_n 0.0126188f $X=3.685 $Y=2.4 $X2=0 $Y2=0
cc_344 N_A_154_135#_M1010_g N_X_c_914_n 0.0126188f $X=4.135 $Y=2.4 $X2=0 $Y2=0
cc_345 N_A_154_135#_c_290_n N_X_c_914_n 0.001658f $X=4.585 $Y=1.69 $X2=0 $Y2=0
cc_346 N_A_154_135#_M1013_g N_X_c_914_n 0.0136432f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_347 N_A_154_135#_c_293_n N_X_c_914_n 0.0750761f $X=4.71 $Y=1.55 $X2=0 $Y2=0
cc_348 N_A_154_135#_c_287_n N_X_c_920_n 0.0110688f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_349 N_A_154_135#_c_290_n N_X_c_920_n 0.0014255f $X=4.585 $Y=1.69 $X2=0 $Y2=0
cc_350 N_A_154_135#_c_298_n N_X_c_920_n 0.00529375f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_351 N_A_154_135#_c_287_n N_X_c_884_n 0.0085362f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_352 N_A_154_135#_c_288_n N_X_c_884_n 0.00805676f $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_353 N_A_154_135#_c_289_n N_X_c_884_n 5.86626e-19 $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_354 N_A_154_135#_c_288_n N_X_c_926_n 0.0109154f $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_355 N_A_154_135#_c_289_n N_X_c_926_n 0.01168f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_356 N_A_154_135#_c_290_n N_X_c_926_n 0.00535808f $X=4.585 $Y=1.69 $X2=0 $Y2=0
cc_357 N_A_154_135#_c_293_n N_X_c_926_n 0.0182043f $X=4.71 $Y=1.55 $X2=0 $Y2=0
cc_358 N_A_154_135#_c_325_n N_X_c_926_n 0.0348755f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_359 N_A_154_135#_c_288_n N_X_c_885_n 5.76374e-19 $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_360 N_A_154_135#_c_289_n N_X_c_885_n 0.00715462f $X=4.24 $Y=1.35 $X2=0 $Y2=0
cc_361 N_A_154_135#_c_307_n N_X_c_893_n 0.0243535f $X=1.075 $Y=1.665 $X2=0 $Y2=0
cc_362 N_A_154_135#_c_298_n N_X_c_893_n 0.0750761f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_363 N_A_154_135#_c_287_n N_X_c_935_n 9.42568e-19 $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_364 N_A_154_135#_c_288_n N_X_c_935_n 7.32094e-19 $X=3.81 $Y=1.35 $X2=0 $Y2=0
cc_365 N_A_154_135#_c_290_n N_X_c_935_n 0.00289909f $X=4.585 $Y=1.69 $X2=0 $Y2=0
cc_366 N_A_154_135#_c_325_n N_X_c_935_n 0.0111425f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_367 N_A_154_135#_c_298_n N_X_c_935_n 0.00527902f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_368 N_A_154_135#_c_292_n N_X_c_886_n 0.0195291f $X=0.91 $Y=1.165 $X2=0 $Y2=0
cc_369 N_A_154_135#_c_298_n N_X_c_886_n 0.0235768f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_370 N_A_154_135#_c_292_n N_X_c_887_n 0.0022879f $X=0.91 $Y=1.165 $X2=0 $Y2=0
cc_371 N_A_154_135#_c_292_n N_X_c_888_n 0.0132312f $X=0.91 $Y=1.165 $X2=0 $Y2=0
cc_372 N_A_154_135#_c_307_n N_X_c_888_n 0.00743502f $X=1.075 $Y=1.665 $X2=0
+ $Y2=0
cc_373 N_A_154_135#_c_287_n X 0.0047024f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_374 N_A_154_135#_c_290_n X 9.39344e-19 $X=4.585 $Y=1.69 $X2=0 $Y2=0
cc_375 N_A_154_135#_c_325_n X 0.00163342f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_376 N_A_154_135#_c_298_n X 0.00413468f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_377 N_A_154_135#_c_287_n N_X_c_890_n 0.00476106f $X=3.38 $Y=1.35 $X2=0 $Y2=0
cc_378 N_A_154_135#_c_290_n N_X_c_890_n 0.00176444f $X=4.585 $Y=1.69 $X2=0 $Y2=0
cc_379 N_A_154_135#_c_325_n N_X_c_890_n 0.00184559f $X=3.795 $Y=1.55 $X2=0 $Y2=0
cc_380 N_A_154_135#_c_298_n N_X_c_890_n 0.015136f $X=3.595 $Y=1.55 $X2=0 $Y2=0
cc_381 N_A_154_135#_M1000_s N_A_1102_392#_c_1004_n 0.00170332f $X=5.95 $Y=1.96
+ $X2=0 $Y2=0
cc_382 N_A_154_135#_M1009_d N_A_71_135#_c_1049_n 0.00430941f $X=0.77 $Y=0.675
+ $X2=0 $Y2=0
cc_383 N_A_154_135#_c_292_n N_A_71_135#_c_1049_n 0.0160844f $X=0.91 $Y=1.165
+ $X2=0 $Y2=0
cc_384 N_A_154_135#_c_298_n N_A_71_135#_c_1049_n 0.00136585f $X=3.595 $Y=1.55
+ $X2=0 $Y2=0
cc_385 N_A_154_135#_c_292_n N_A_71_135#_c_1054_n 0.00606866f $X=0.91 $Y=1.165
+ $X2=0 $Y2=0
cc_386 N_A_154_135#_c_298_n N_A_71_135#_c_1046_n 0.0899913f $X=3.595 $Y=1.55
+ $X2=0 $Y2=0
cc_387 N_A_154_135#_c_292_n N_A_71_135#_c_1047_n 0.0104031f $X=0.91 $Y=1.165
+ $X2=0 $Y2=0
cc_388 N_A_154_135#_c_298_n N_A_71_135#_c_1047_n 0.0123781f $X=3.595 $Y=1.55
+ $X2=0 $Y2=0
cc_389 N_A_154_135#_c_294_n N_VGND_M1023_s 0.00837877f $X=5.61 $Y=1.215 $X2=0
+ $Y2=0
cc_390 N_A_154_135#_c_299_n N_VGND_M1023_s 0.00115102f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_391 N_A_154_135#_c_287_n N_VGND_c_1100_n 0.00278543f $X=3.38 $Y=1.35 $X2=0
+ $Y2=0
cc_392 N_A_154_135#_c_288_n N_VGND_c_1101_n 0.00209581f $X=3.81 $Y=1.35 $X2=0
+ $Y2=0
cc_393 N_A_154_135#_c_289_n N_VGND_c_1101_n 0.00150779f $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_394 N_A_154_135#_c_289_n N_VGND_c_1102_n 4.82085e-19 $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_395 N_A_154_135#_c_291_n N_VGND_c_1102_n 0.0133684f $X=4.67 $Y=1.35 $X2=0
+ $Y2=0
cc_396 N_A_154_135#_c_294_n N_VGND_c_1102_n 0.0445845f $X=5.61 $Y=1.215 $X2=0
+ $Y2=0
cc_397 N_A_154_135#_c_295_n N_VGND_c_1102_n 0.0151478f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_398 N_A_154_135#_c_299_n N_VGND_c_1102_n 0.00887034f $X=4.795 $Y=1.215 $X2=0
+ $Y2=0
cc_399 N_A_154_135#_c_295_n N_VGND_c_1103_n 0.00646413f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_400 N_A_154_135#_c_295_n N_VGND_c_1104_n 0.00765349f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_401 N_A_154_135#_c_297_n N_VGND_c_1104_n 0.0123214f $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_402 N_A_154_135#_c_300_n N_VGND_c_1104_n 0.00721388f $X=5.85 $Y=1.215 $X2=0
+ $Y2=0
cc_403 N_A_154_135#_c_287_n N_VGND_c_1109_n 0.00466874f $X=3.38 $Y=1.35 $X2=0
+ $Y2=0
cc_404 N_A_154_135#_c_288_n N_VGND_c_1109_n 0.00466874f $X=3.81 $Y=1.35 $X2=0
+ $Y2=0
cc_405 N_A_154_135#_c_295_n N_VGND_c_1111_n 0.00739421f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_406 N_A_154_135#_c_295_n N_VGND_c_1162_n 0.020538f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_407 N_A_154_135#_c_297_n N_VGND_c_1162_n 6.72765e-19 $X=8.115 $Y=1.685 $X2=0
+ $Y2=0
cc_408 N_A_154_135#_c_301_n N_VGND_c_1162_n 0.00376194f $X=6.085 $Y=1.685 $X2=0
+ $Y2=0
cc_409 N_A_154_135#_c_289_n N_VGND_c_1114_n 0.00467453f $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_410 N_A_154_135#_c_291_n N_VGND_c_1114_n 0.00405273f $X=4.67 $Y=1.35 $X2=0
+ $Y2=0
cc_411 N_A_154_135#_c_287_n N_VGND_c_1117_n 0.00505379f $X=3.38 $Y=1.35 $X2=0
+ $Y2=0
cc_412 N_A_154_135#_c_288_n N_VGND_c_1117_n 0.00505379f $X=3.81 $Y=1.35 $X2=0
+ $Y2=0
cc_413 N_A_154_135#_c_289_n N_VGND_c_1117_n 0.00505379f $X=4.24 $Y=1.35 $X2=0
+ $Y2=0
cc_414 N_A_154_135#_c_291_n N_VGND_c_1117_n 0.00424518f $X=4.67 $Y=1.35 $X2=0
+ $Y2=0
cc_415 N_A_154_135#_c_295_n N_VGND_c_1117_n 0.0103323f $X=5.775 $Y=0.745 $X2=0
+ $Y2=0
cc_416 N_A_154_135#_c_297_n N_A_1346_123#_c_1241_n 0.0672585f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_417 N_A_154_135#_c_363_p N_A_1346_123#_c_1241_n 0.0136942f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_418 N_A_154_135#_c_296_n N_A_1346_123#_c_1242_n 0.00406848f $X=6.005 $Y=1.6
+ $X2=0 $Y2=0
cc_419 N_A_154_135#_c_297_n N_A_1346_123#_c_1242_n 0.0273383f $X=8.115 $Y=1.685
+ $X2=0 $Y2=0
cc_420 N_A_154_135#_c_300_n N_A_1346_123#_c_1242_n 6.69459e-19 $X=5.85 $Y=1.215
+ $X2=0 $Y2=0
cc_421 N_A_154_135#_c_363_p N_A_1346_123#_c_1243_n 0.0329533f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_422 N_A_154_135#_M1012_d N_A_1346_123#_c_1244_n 0.00176461f $X=8.14 $Y=0.38
+ $X2=0 $Y2=0
cc_423 N_A_154_135#_c_363_p N_A_1346_123#_c_1244_n 0.0159805f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_424 N_A_154_135#_c_363_p N_A_1346_123#_c_1246_n 0.0166977f $X=8.28 $Y=0.76
+ $X2=0 $Y2=0
cc_425 N_C1_M1026_g N_B2_M1002_g 0.0262367f $X=6.31 $Y=2.46 $X2=0 $Y2=0
cc_426 N_C1_c_499_n N_B2_c_565_n 0.0262367f $X=6.31 $Y=1.715 $X2=0 $Y2=0
cc_427 N_C1_c_499_n N_B2_M1019_g 0.00456705f $X=6.31 $Y=1.715 $X2=0 $Y2=0
cc_428 N_C1_M1025_g N_B2_c_572_n 8.38383e-19 $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_429 N_C1_M1025_g N_B2_c_573_n 0.0107847f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_430 N_C1_M1000_g N_VPWR_c_721_n 0.00333926f $X=5.86 $Y=2.46 $X2=0 $Y2=0
cc_431 N_C1_M1026_g N_VPWR_c_721_n 0.00333926f $X=6.31 $Y=2.46 $X2=0 $Y2=0
cc_432 N_C1_M1000_g N_VPWR_c_707_n 0.0042782f $X=5.86 $Y=2.46 $X2=0 $Y2=0
cc_433 N_C1_M1026_g N_VPWR_c_707_n 0.00422798f $X=6.31 $Y=2.46 $X2=0 $Y2=0
cc_434 N_C1_M1000_g N_A_160_376#_c_796_n 0.0183879f $X=5.86 $Y=2.46 $X2=0 $Y2=0
cc_435 N_C1_c_498_n N_A_160_376#_c_796_n 0.00106638f $X=6.065 $Y=1.515 $X2=0
+ $Y2=0
cc_436 N_C1_M1026_g N_A_160_376#_c_796_n 0.0136056f $X=6.31 $Y=2.46 $X2=0 $Y2=0
cc_437 C1 N_A_160_376#_c_796_n 0.0216811f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_438 N_C1_M1026_g N_A_160_376#_c_797_n 4.94927e-19 $X=6.31 $Y=2.46 $X2=0 $Y2=0
cc_439 N_C1_M1026_g N_A_160_376#_c_820_n 0.00103955f $X=6.31 $Y=2.46 $X2=0 $Y2=0
cc_440 C1 N_A_1102_392#_M1000_d 0.00437939f $X=5.435 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_441 N_C1_M1000_g N_A_1102_392#_c_1004_n 0.0163222f $X=5.86 $Y=2.46 $X2=0
+ $Y2=0
cc_442 N_C1_M1026_g N_A_1102_392#_c_1004_n 0.0153296f $X=6.31 $Y=2.46 $X2=0
+ $Y2=0
cc_443 N_C1_M1024_g N_VGND_c_1102_n 0.00563785f $X=5.56 $Y=0.92 $X2=0 $Y2=0
cc_444 N_C1_M1025_g N_VGND_c_1103_n 0.00379263f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_445 N_C1_M1025_g N_VGND_c_1104_n 0.00215221f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_446 N_C1_c_499_n N_VGND_c_1104_n 0.00291685f $X=6.31 $Y=1.715 $X2=0 $Y2=0
cc_447 N_C1_M1024_g N_VGND_c_1111_n 0.00412501f $X=5.56 $Y=0.92 $X2=0 $Y2=0
cc_448 N_C1_M1025_g N_VGND_c_1111_n 0.00412501f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_449 N_C1_M1025_g N_VGND_c_1162_n 0.00298414f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_450 N_C1_c_497_n N_VGND_c_1162_n 0.00318711f $X=6.22 $Y=1.515 $X2=0 $Y2=0
cc_451 N_C1_M1024_g N_VGND_c_1117_n 0.00476395f $X=5.56 $Y=0.92 $X2=0 $Y2=0
cc_452 N_C1_M1025_g N_VGND_c_1117_n 0.00476395f $X=5.99 $Y=0.92 $X2=0 $Y2=0
cc_453 N_C1_M1025_g N_A_1346_123#_c_1242_n 3.77674e-19 $X=5.99 $Y=0.92 $X2=0
+ $Y2=0
cc_454 N_B2_M1004_g N_B1_M1007_g 0.0227826f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_455 N_B2_c_569_n N_B1_M1007_g 0.00425279f $X=7.475 $Y=1.7 $X2=0 $Y2=0
cc_456 N_B2_c_563_n N_B1_M1012_g 0.0131785f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_457 N_B2_c_567_n N_B1_c_658_n 0.00723084f $X=7.475 $Y=1.625 $X2=0 $Y2=0
cc_458 N_B2_c_568_n N_B1_c_658_n 0.0131785f $X=7.575 $Y=1.33 $X2=0 $Y2=0
cc_459 N_B2_M1002_g N_VPWR_c_721_n 0.00333926f $X=6.76 $Y=2.46 $X2=0 $Y2=0
cc_460 N_B2_M1004_g N_VPWR_c_721_n 0.00333926f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_461 N_B2_M1002_g N_VPWR_c_707_n 0.00422798f $X=6.76 $Y=2.46 $X2=0 $Y2=0
cc_462 N_B2_M1004_g N_VPWR_c_707_n 0.00424948f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_463 N_B2_M1002_g N_A_160_376#_c_796_n 0.011188f $X=6.76 $Y=2.46 $X2=0 $Y2=0
cc_464 N_B2_M1002_g N_A_160_376#_c_797_n 0.00391937f $X=6.76 $Y=2.46 $X2=0 $Y2=0
cc_465 N_B2_c_564_n N_A_160_376#_c_797_n 0.00193695f $X=7.01 $Y=1.7 $X2=0 $Y2=0
cc_466 N_B2_M1004_g N_A_160_376#_c_797_n 0.00112087f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_467 N_B2_M1002_g N_A_160_376#_c_820_n 0.00542687f $X=6.76 $Y=2.46 $X2=0 $Y2=0
cc_468 N_B2_M1004_g N_A_160_376#_c_820_n 0.00928993f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_469 N_B2_M1004_g N_A_160_376#_c_798_n 0.0141331f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_470 N_B2_c_569_n N_A_160_376#_c_798_n 0.00630268f $X=7.475 $Y=1.7 $X2=0 $Y2=0
cc_471 N_B2_M1002_g N_A_160_376#_c_838_n 0.00127873f $X=6.76 $Y=2.46 $X2=0 $Y2=0
cc_472 N_B2_M1004_g N_A_160_376#_c_838_n 0.00603356f $X=7.21 $Y=2.46 $X2=0 $Y2=0
cc_473 N_B2_M1002_g N_A_1102_392#_c_1005_n 0.00818857f $X=6.76 $Y=2.46 $X2=0
+ $Y2=0
cc_474 N_B2_M1004_g N_A_1102_392#_c_1005_n 0.0158794f $X=7.21 $Y=2.46 $X2=0
+ $Y2=0
cc_475 N_B2_M1004_g N_A_1102_392#_c_1016_n 0.00981283f $X=7.21 $Y=2.46 $X2=0
+ $Y2=0
cc_476 N_B2_M1002_g N_A_1102_392#_c_1008_n 0.00619966f $X=6.76 $Y=2.46 $X2=0
+ $Y2=0
cc_477 N_B2_M1004_g N_A_1102_392#_c_1008_n 7.38166e-19 $X=7.21 $Y=2.46 $X2=0
+ $Y2=0
cc_478 N_B2_c_571_n N_VGND_c_1103_n 0.0243585f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_479 N_B2_c_572_n N_VGND_c_1103_n 0.00566684f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_480 N_B2_c_573_n N_VGND_c_1103_n 0.00167326f $X=6.635 $Y=0.505 $X2=0 $Y2=0
cc_481 N_B2_c_573_n N_VGND_c_1104_n 2.51918e-19 $X=6.635 $Y=0.505 $X2=0 $Y2=0
cc_482 N_B2_c_563_n N_VGND_c_1105_n 0.0193089f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_483 N_B2_M1019_g N_VGND_c_1105_n 0.00161245f $X=7.085 $Y=0.935 $X2=0 $Y2=0
cc_484 N_B2_c_568_n N_VGND_c_1105_n 0.00832159f $X=7.575 $Y=1.33 $X2=0 $Y2=0
cc_485 N_B2_c_570_n N_VGND_c_1105_n 4.2102e-19 $X=7.575 $Y=1.405 $X2=0 $Y2=0
cc_486 N_B2_c_571_n N_VGND_c_1105_n 0.029476f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_487 N_B2_c_571_n N_VGND_c_1162_n 0.00386879f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_488 N_B2_c_572_n N_VGND_c_1162_n 0.00127982f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_489 N_B2_c_571_n N_VGND_c_1115_n 0.0366677f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_490 N_B2_c_572_n N_VGND_c_1115_n 0.0181591f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_491 N_B2_c_563_n N_VGND_c_1116_n 0.00693208f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_492 N_B2_c_563_n N_VGND_c_1117_n 0.0256169f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_493 N_B2_M1019_g N_VGND_c_1117_n 7.07849e-19 $X=7.085 $Y=0.935 $X2=0 $Y2=0
cc_494 N_B2_c_571_n N_VGND_c_1117_n 0.0191717f $X=6.845 $Y=0.38 $X2=0 $Y2=0
cc_495 N_B2_c_572_n N_VGND_c_1117_n 0.0100038f $X=6.635 $Y=0.2 $X2=0 $Y2=0
cc_496 N_B2_c_571_n N_A_1346_123#_M1017_d 0.00190525f $X=6.845 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_497 N_B2_c_563_n N_A_1346_123#_c_1258_n 3.49074e-19 $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_498 N_B2_M1019_g N_A_1346_123#_c_1258_n 0.00657116f $X=7.085 $Y=0.935 $X2=0
+ $Y2=0
cc_499 N_B2_c_568_n N_A_1346_123#_c_1258_n 5.93148e-19 $X=7.575 $Y=1.33 $X2=0
+ $Y2=0
cc_500 N_B2_c_571_n N_A_1346_123#_c_1258_n 0.0156219f $X=6.845 $Y=0.38 $X2=0
+ $Y2=0
cc_501 N_B2_c_572_n N_A_1346_123#_c_1258_n 0.00127917f $X=6.635 $Y=0.2 $X2=0
+ $Y2=0
cc_502 N_B2_c_573_n N_A_1346_123#_c_1258_n 0.00526654f $X=6.635 $Y=0.505 $X2=0
+ $Y2=0
cc_503 N_B2_M1019_g N_A_1346_123#_c_1241_n 0.0109993f $X=7.085 $Y=0.935 $X2=0
+ $Y2=0
cc_504 N_B2_c_568_n N_A_1346_123#_c_1241_n 0.00932666f $X=7.575 $Y=1.33 $X2=0
+ $Y2=0
cc_505 N_B2_c_569_n N_A_1346_123#_c_1241_n 3.91025e-19 $X=7.475 $Y=1.7 $X2=0
+ $Y2=0
cc_506 N_B2_c_570_n N_A_1346_123#_c_1241_n 0.00873336f $X=7.575 $Y=1.405 $X2=0
+ $Y2=0
cc_507 N_B2_c_571_n N_A_1346_123#_c_1241_n 2.22629e-19 $X=6.845 $Y=0.38 $X2=0
+ $Y2=0
cc_508 N_B2_c_565_n N_A_1346_123#_c_1242_n 0.00210303f $X=6.85 $Y=1.7 $X2=0
+ $Y2=0
cc_509 N_B2_M1019_g N_A_1346_123#_c_1242_n 0.0030905f $X=7.085 $Y=0.935 $X2=0
+ $Y2=0
cc_510 N_B2_c_573_n N_A_1346_123#_c_1242_n 0.00390184f $X=6.635 $Y=0.505 $X2=0
+ $Y2=0
cc_511 N_B2_c_568_n N_A_1346_123#_c_1243_n 0.0086474f $X=7.575 $Y=1.33 $X2=0
+ $Y2=0
cc_512 N_B2_c_563_n N_A_1346_123#_c_1245_n 0.0017897f $X=7.5 $Y=0.2 $X2=0 $Y2=0
cc_513 N_B1_M1007_g N_VPWR_c_721_n 0.00333926f $X=7.95 $Y=2.46 $X2=0 $Y2=0
cc_514 N_B1_M1014_g N_VPWR_c_721_n 0.00333926f $X=8.44 $Y=2.46 $X2=0 $Y2=0
cc_515 N_B1_M1007_g N_VPWR_c_707_n 0.00425342f $X=7.95 $Y=2.46 $X2=0 $Y2=0
cc_516 N_B1_M1014_g N_VPWR_c_707_n 0.00428215f $X=8.44 $Y=2.46 $X2=0 $Y2=0
cc_517 N_B1_M1007_g N_A_160_376#_c_798_n 0.0141331f $X=7.95 $Y=2.46 $X2=0 $Y2=0
cc_518 N_B1_M1007_g N_A_160_376#_c_801_n 0.0170221f $X=7.95 $Y=2.46 $X2=0 $Y2=0
cc_519 N_B1_M1014_g N_A_160_376#_c_801_n 0.012604f $X=8.44 $Y=2.46 $X2=0 $Y2=0
cc_520 N_B1_c_658_n N_A_160_376#_c_801_n 8.91853e-19 $X=8.57 $Y=1.51 $X2=0 $Y2=0
cc_521 N_B1_M1007_g N_A_1102_392#_c_1016_n 0.0100107f $X=7.95 $Y=2.46 $X2=0
+ $Y2=0
cc_522 N_B1_M1007_g N_A_1102_392#_c_1006_n 0.01615f $X=7.95 $Y=2.46 $X2=0 $Y2=0
cc_523 N_B1_M1014_g N_A_1102_392#_c_1006_n 0.0152288f $X=8.44 $Y=2.46 $X2=0
+ $Y2=0
cc_524 N_B1_M1014_g N_A_1102_392#_c_1007_n 4.6887e-19 $X=8.44 $Y=2.46 $X2=0
+ $Y2=0
cc_525 N_B1_c_660_n N_A_1102_392#_c_1007_n 0.00301248f $X=9.115 $Y=1.465 $X2=0
+ $Y2=0
cc_526 N_B1_c_666_n N_A_1102_392#_c_1007_n 0.0178913f $X=9.095 $Y=1.48 $X2=0
+ $Y2=0
cc_527 N_B1_M1012_g N_VGND_c_1116_n 0.00390708f $X=8.065 $Y=0.7 $X2=0 $Y2=0
cc_528 N_B1_M1020_g N_VGND_c_1116_n 0.00390708f $X=8.495 $Y=0.7 $X2=0 $Y2=0
cc_529 N_B1_M1012_g N_VGND_c_1117_n 0.00542671f $X=8.065 $Y=0.7 $X2=0 $Y2=0
cc_530 N_B1_M1020_g N_VGND_c_1117_n 0.00542671f $X=8.495 $Y=0.7 $X2=0 $Y2=0
cc_531 N_B1_M1012_g N_A_1346_123#_c_1241_n 0.00164273f $X=8.065 $Y=0.7 $X2=0
+ $Y2=0
cc_532 N_B1_c_658_n N_A_1346_123#_c_1241_n 0.00211713f $X=8.57 $Y=1.51 $X2=0
+ $Y2=0
cc_533 N_B1_M1012_g N_A_1346_123#_c_1243_n 0.00195727f $X=8.065 $Y=0.7 $X2=0
+ $Y2=0
cc_534 N_B1_M1012_g N_A_1346_123#_c_1244_n 0.0123852f $X=8.065 $Y=0.7 $X2=0
+ $Y2=0
cc_535 N_B1_M1020_g N_A_1346_123#_c_1244_n 0.0135055f $X=8.495 $Y=0.7 $X2=0
+ $Y2=0
cc_536 N_B1_M1020_g N_A_1346_123#_c_1246_n 4.46492e-19 $X=8.495 $Y=0.7 $X2=0
+ $Y2=0
cc_537 N_B1_c_660_n N_A_1346_123#_c_1246_n 0.00691526f $X=9.115 $Y=1.465 $X2=0
+ $Y2=0
cc_538 N_B1_c_666_n N_A_1346_123#_c_1246_n 0.0186971f $X=9.095 $Y=1.48 $X2=0
+ $Y2=0
cc_539 N_VPWR_M1018_d N_A_160_376#_c_802_n 0.0160942f $X=1.37 $Y=1.88 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_723_n N_A_160_376#_c_802_n 0.0488965f $X=1.9 $Y=2.71 $X2=0 $Y2=0
cc_541 N_VPWR_M1003_s N_A_160_376#_c_796_n 0.00817743f $X=2.715 $Y=1.88 $X2=0
+ $Y2=0
cc_542 N_VPWR_M1008_s N_A_160_376#_c_796_n 0.00322506f $X=3.775 $Y=1.84 $X2=0
+ $Y2=0
cc_543 N_VPWR_M1013_s N_A_160_376#_c_796_n 0.00795195f $X=4.675 $Y=1.84 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_709_n N_A_160_376#_c_796_n 0.0213878f $X=3.01 $Y=2.8 $X2=0 $Y2=0
cc_545 N_VPWR_c_710_n N_A_160_376#_c_796_n 0.0166604f $X=3.91 $Y=2.8 $X2=0 $Y2=0
cc_546 N_VPWR_c_711_n N_A_160_376#_c_796_n 0.0215065f $X=4.81 $Y=2.8 $X2=0 $Y2=0
cc_547 N_VPWR_c_707_n N_A_160_376#_c_796_n 0.0691938f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_708_n N_A_160_376#_c_799_n 0.038767f $X=0.485 $Y=2.345 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_720_n N_A_160_376#_c_799_n 0.0109318f $X=1.395 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_707_n N_A_160_376#_c_799_n 0.0114582f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_723_n N_A_160_376#_c_799_n 0.0118598f $X=1.9 $Y=2.71 $X2=0 $Y2=0
cc_552 N_VPWR_c_709_n N_A_160_376#_c_800_n 0.0106231f $X=3.01 $Y=2.8 $X2=0 $Y2=0
cc_553 N_VPWR_c_714_n N_A_160_376#_c_800_n 0.0108548f $X=2.845 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_707_n N_A_160_376#_c_800_n 0.0114305f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_723_n N_A_160_376#_c_800_n 0.0121364f $X=1.9 $Y=2.71 $X2=0 $Y2=0
cc_556 N_VPWR_c_708_n N_X_c_891_n 0.00313887f $X=0.485 $Y=2.345 $X2=0 $Y2=0
cc_557 N_VPWR_M1003_s N_X_c_902_n 0.00730502f $X=2.715 $Y=1.88 $X2=0 $Y2=0
cc_558 N_VPWR_M1008_s N_X_c_914_n 0.00318055f $X=3.775 $Y=1.84 $X2=0 $Y2=0
cc_559 N_VPWR_M1016_d N_X_c_893_n 0.00682304f $X=0.36 $Y=1.88 $X2=0 $Y2=0
cc_560 N_VPWR_M1018_d N_X_c_893_n 0.0160017f $X=1.37 $Y=1.88 $X2=0 $Y2=0
cc_561 N_VPWR_M1003_s N_X_c_893_n 0.00171404f $X=2.715 $Y=1.88 $X2=0 $Y2=0
cc_562 N_VPWR_c_708_n N_X_c_893_n 0.0190672f $X=0.485 $Y=2.345 $X2=0 $Y2=0
cc_563 N_VPWR_c_711_n N_A_1102_392#_c_1004_n 0.0157109f $X=4.81 $Y=2.8 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_721_n N_A_1102_392#_c_1004_n 0.128194f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_707_n N_A_1102_392#_c_1004_n 0.0710407f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_721_n N_A_1102_392#_c_1006_n 0.0699605f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_707_n N_A_1102_392#_c_1006_n 0.0390913f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_721_n N_A_1102_392#_c_1009_n 0.0236566f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_707_n N_A_1102_392#_c_1009_n 0.0128296f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_570 N_A_160_376#_c_796_n N_X_M1006_d 0.00462319f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_571 N_A_160_376#_c_796_n N_X_M1010_d 0.00462319f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_572 N_A_160_376#_c_796_n N_X_c_902_n 0.0930301f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_573 N_A_160_376#_M1016_s N_X_c_893_n 0.00686982f $X=0.8 $Y=1.88 $X2=0 $Y2=0
cc_574 N_A_160_376#_M1001_d N_X_c_893_n 0.00317105f $X=2.265 $Y=1.88 $X2=0 $Y2=0
cc_575 N_A_160_376#_c_802_n N_X_c_893_n 0.0639189f $X=2.235 $Y=2.345 $X2=0 $Y2=0
cc_576 N_A_160_376#_c_796_n N_X_c_893_n 0.0110064f $X=6.82 $Y=2.445 $X2=0 $Y2=0
cc_577 N_A_160_376#_c_799_n N_X_c_893_n 0.0219052f $X=1.055 $Y=2.345 $X2=0 $Y2=0
cc_578 N_A_160_376#_c_800_n N_X_c_893_n 0.0170939f $X=2.4 $Y=2.345 $X2=0 $Y2=0
cc_579 N_A_160_376#_c_796_n N_A_1102_392#_M1000_d 0.00499847f $X=6.82 $Y=2.445
+ $X2=-0.19 $Y2=1.66
cc_580 N_A_160_376#_c_796_n N_A_1102_392#_M1026_d 0.00471229f $X=6.82 $Y=2.445
+ $X2=0 $Y2=0
cc_581 N_A_160_376#_c_798_n N_A_1102_392#_M1004_s 0.0096385f $X=8.01 $Y=2.025
+ $X2=0 $Y2=0
cc_582 N_A_160_376#_c_796_n N_A_1102_392#_c_1004_n 0.0690105f $X=6.82 $Y=2.445
+ $X2=0 $Y2=0
cc_583 N_A_160_376#_M1002_d N_A_1102_392#_c_1005_n 0.00165831f $X=6.85 $Y=1.96
+ $X2=0 $Y2=0
cc_584 N_A_160_376#_c_796_n N_A_1102_392#_c_1005_n 0.00368894f $X=6.82 $Y=2.445
+ $X2=0 $Y2=0
cc_585 N_A_160_376#_c_838_n N_A_1102_392#_c_1005_n 0.0149732f $X=6.985 $Y=2.445
+ $X2=0 $Y2=0
cc_586 N_A_160_376#_c_820_n N_A_1102_392#_c_1016_n 0.00426956f $X=6.985 $Y=2.36
+ $X2=0 $Y2=0
cc_587 N_A_160_376#_c_798_n N_A_1102_392#_c_1016_n 0.0266856f $X=8.01 $Y=2.025
+ $X2=0 $Y2=0
cc_588 N_A_160_376#_c_838_n N_A_1102_392#_c_1016_n 0.0205757f $X=6.985 $Y=2.445
+ $X2=0 $Y2=0
cc_589 N_A_160_376#_c_801_n N_A_1102_392#_c_1016_n 0.0260981f $X=8.195 $Y=2.105
+ $X2=0 $Y2=0
cc_590 N_A_160_376#_M1007_d N_A_1102_392#_c_1006_n 0.00208352f $X=8.04 $Y=1.96
+ $X2=0 $Y2=0
cc_591 N_A_160_376#_c_801_n N_A_1102_392#_c_1006_n 0.0189764f $X=8.195 $Y=2.105
+ $X2=0 $Y2=0
cc_592 N_A_160_376#_c_801_n N_A_1102_392#_c_1007_n 0.00696138f $X=8.195 $Y=2.105
+ $X2=0 $Y2=0
cc_593 N_X_c_886_n N_A_71_135#_M1009_s 0.0019963f $X=2.975 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_594 N_X_c_887_n N_A_71_135#_M1009_s 7.27654e-19 $X=0.385 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_595 N_X_c_886_n N_A_71_135#_M1011_s 0.00206067f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_596 N_X_c_886_n N_A_71_135#_M1022_d 0.00201585f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_597 N_X_c_886_n N_A_71_135#_c_1049_n 0.012018f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_598 N_X_c_886_n N_A_71_135#_c_1054_n 0.00908056f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_599 N_X_c_886_n N_A_71_135#_c_1046_n 0.0443333f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_600 X N_A_71_135#_c_1046_n 0.00129662f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_601 N_X_c_890_n N_A_71_135#_c_1046_n 0.00793711f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_602 N_X_c_886_n N_A_71_135#_c_1047_n 0.00564678f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_603 N_X_c_886_n N_A_71_135#_c_1065_n 0.00591085f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_604 X N_A_71_135#_c_1065_n 0.00128755f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_605 N_X_c_890_n N_A_71_135#_c_1065_n 9.21622e-19 $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_606 N_X_c_886_n N_A_71_135#_c_1048_n 0.00835176f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_607 N_X_c_887_n N_A_71_135#_c_1048_n 0.00187568f $X=0.385 $Y=1.295 $X2=0
+ $Y2=0
cc_608 N_X_c_888_n N_A_71_135#_c_1048_n 0.0027311f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_609 N_X_c_886_n N_VGND_M1022_s 0.00372485f $X=2.975 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_610 N_X_c_920_n N_VGND_M1027_s 6.98766e-19 $X=3.43 $Y=1.095 $X2=0 $Y2=0
cc_611 N_X_c_886_n N_VGND_M1027_s 3.42314e-19 $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_612 X N_VGND_M1027_s 0.00254293f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_613 N_X_c_890_n N_VGND_M1027_s 0.00512514f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_614 N_X_c_926_n N_VGND_M1015_s 0.00330483f $X=4.29 $Y=1.095 $X2=0 $Y2=0
cc_615 N_X_c_920_n N_VGND_c_1100_n 9.87298e-19 $X=3.43 $Y=1.095 $X2=0 $Y2=0
cc_616 N_X_c_884_n N_VGND_c_1100_n 0.0165971f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_617 X N_VGND_c_1100_n 0.00158234f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_618 N_X_c_890_n N_VGND_c_1100_n 0.0172527f $X=3.12 $Y=1.095 $X2=0 $Y2=0
cc_619 N_X_c_884_n N_VGND_c_1101_n 0.0164685f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_620 N_X_c_926_n N_VGND_c_1101_n 0.0135055f $X=4.29 $Y=1.095 $X2=0 $Y2=0
cc_621 N_X_c_885_n N_VGND_c_1101_n 0.013052f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_622 N_X_c_885_n N_VGND_c_1102_n 0.0201101f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_623 N_X_c_886_n N_VGND_c_1108_n 0.0103398f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_624 N_X_c_884_n N_VGND_c_1109_n 0.0105983f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_625 N_X_c_885_n N_VGND_c_1114_n 0.00718756f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_626 N_X_c_884_n N_VGND_c_1117_n 0.0113894f $X=3.595 $Y=0.645 $X2=0 $Y2=0
cc_627 N_X_c_885_n N_VGND_c_1117_n 0.0083989f $X=4.455 $Y=0.645 $X2=0 $Y2=0
cc_628 N_A_71_135#_c_1046_n N_VGND_M1022_s 9.8611e-19 $X=2.51 $Y=1.325 $X2=-0.19
+ $Y2=-0.245
cc_629 N_A_71_135#_c_1049_n N_VGND_c_1106_n 0.0105986f $X=1.255 $Y=0.82 $X2=0
+ $Y2=0
cc_630 N_A_71_135#_c_1048_n N_VGND_c_1106_n 0.00458739f $X=0.48 $Y=0.83 $X2=0
+ $Y2=0
cc_631 N_A_71_135#_c_1054_n N_VGND_c_1108_n 0.00104849f $X=1.34 $Y=1.035 $X2=0
+ $Y2=0
cc_632 N_A_71_135#_c_1046_n N_VGND_c_1108_n 0.0269989f $X=2.51 $Y=1.325 $X2=0
+ $Y2=0
cc_633 N_A_71_135#_c_1049_n N_VGND_c_1117_n 0.0226601f $X=1.255 $Y=0.82 $X2=0
+ $Y2=0
cc_634 N_A_71_135#_c_1065_n N_VGND_c_1117_n 5.77272e-19 $X=2.675 $Y=1.055 $X2=0
+ $Y2=0
cc_635 N_A_71_135#_c_1048_n N_VGND_c_1117_n 0.00719958f $X=0.48 $Y=0.83 $X2=0
+ $Y2=0
cc_636 N_VGND_c_1104_n N_A_1346_123#_c_1258_n 0.0108698f $X=6.44 $Y=1.115 $X2=0
+ $Y2=0
cc_637 N_VGND_c_1117_n N_A_1346_123#_c_1258_n 8.15299e-19 $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_638 N_VGND_c_1105_n N_A_1346_123#_c_1241_n 0.0205307f $X=7.3 $Y=0.925 $X2=0
+ $Y2=0
cc_639 N_VGND_c_1104_n N_A_1346_123#_c_1242_n 0.00157382f $X=6.44 $Y=1.115 $X2=0
+ $Y2=0
cc_640 N_VGND_c_1105_n N_A_1346_123#_c_1243_n 0.0442411f $X=7.3 $Y=0.925 $X2=0
+ $Y2=0
cc_641 N_VGND_c_1116_n N_A_1346_123#_c_1244_n 0.0650231f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_642 N_VGND_c_1117_n N_A_1346_123#_c_1244_n 0.037428f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1105_n N_A_1346_123#_c_1245_n 0.0122034f $X=7.3 $Y=0.925 $X2=0
+ $Y2=0
cc_644 N_VGND_c_1116_n N_A_1346_123#_c_1245_n 0.0179217f $X=9.36 $Y=0 $X2=0
+ $Y2=0
cc_645 N_VGND_c_1117_n N_A_1346_123#_c_1245_n 0.00971942f $X=9.36 $Y=0 $X2=0
+ $Y2=0

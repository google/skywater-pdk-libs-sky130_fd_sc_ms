* File: sky130_fd_sc_ms__and3_1.pex.spice
* Created: Wed Sep  2 11:57:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND3_1%A 5 7 10 12 16 18 22
r42 18 22 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=0.462
+ $X2=1.085 $Y2=0.462
r43 15 22 17.3781 $w=3.13e-07 $l=4.75e-07 $layer=LI1_cond $X=0.61 $Y=0.412
+ $X2=1.085 $Y2=0.412
r44 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=0.405 $X2=0.61 $Y2=0.405
r45 11 12 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.51 $Y=1.395
+ $X2=0.51 $Y2=1.545
r46 10 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.53 $Y=1 $X2=0.53
+ $Y2=1.395
r47 7 16 19.6204 $w=1.5e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.53 $Y=0.57
+ $X2=0.615 $Y2=0.405
r48 7 10 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.53 $Y=0.57 $X2=0.53
+ $Y2=1
r49 5 12 336.234 $w=1.8e-07 $l=8.65e-07 $layer=POLY_cond $X=0.505 $Y=2.41
+ $X2=0.505 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_1%B 3 7 8 9 13 15
c45 3 0 1.67593e-20 $X=1.055 $Y=2.41
r46 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.595
+ $X2=1.01 $Y2=1.76
r47 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.595
+ $X2=1.01 $Y2=1.43
r48 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.595 $X2=1.01 $Y2=1.595
r49 9 14 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=1.08 $Y=1.665 $X2=1.08
+ $Y2=1.595
r50 8 14 7.63454 $w=4.68e-07 $l=3e-07 $layer=LI1_cond $X=1.08 $Y=1.295 $X2=1.08
+ $Y2=1.595
r51 7 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.09 $Y=1 $X2=1.09
+ $Y2=1.43
r52 3 16 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=1.055 $Y=2.41
+ $X2=1.055 $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_1%C 3 7 9 12
c38 9 0 1.67593e-20 $X=1.68 $Y=1.665
r39 12 15 39.9775 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.615
+ $X2=1.615 $Y2=1.78
r40 12 14 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.615
+ $X2=1.615 $Y2=1.45
r41 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.615 $X2=1.65 $Y2=1.615
r42 7 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.565 $Y=0.92
+ $X2=1.565 $Y2=1.45
r43 3 15 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=1.505 $Y=2.41
+ $X2=1.505 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_1%A_27_398# 1 2 3 10 12 15 19 23 25 29 31 34 35
+ 36 38 45
r80 39 45 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.235 $Y=1.515
+ $X2=2.375 $Y2=1.515
r81 39 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.235 $Y=1.515
+ $X2=2.145 $Y2=1.515
r82 38 41 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=1.515
+ $X2=2.235 $Y2=1.68
r83 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.515 $X2=2.235 $Y2=1.515
r84 34 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.155 $Y=1.95
+ $X2=2.155 $Y2=1.68
r85 32 36 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.4 $Y=2.035
+ $X2=1.257 $Y2=2.035
r86 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.07 $Y=2.035
+ $X2=2.155 $Y2=1.95
r87 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=2.035
+ $X2=1.4 $Y2=2.035
r88 27 36 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.257 $Y=2.12
+ $X2=1.257 $Y2=2.035
r89 27 29 0.606549 $w=2.83e-07 $l=1.5e-08 $layer=LI1_cond $X=1.257 $Y=2.12
+ $X2=1.257 $Y2=2.135
r90 26 35 4.00616 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.48 $Y=2.035
+ $X2=0.297 $Y2=2.035
r91 25 36 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.115 $Y=2.035
+ $X2=1.257 $Y2=2.035
r92 25 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.115 $Y=2.035
+ $X2=0.48 $Y2=2.035
r93 21 35 2.75409 $w=3.47e-07 $l=9.31128e-08 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.297 $Y2=2.035
r94 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.135
r95 17 35 2.75409 $w=3.47e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=1.95
+ $X2=0.297 $Y2=2.035
r96 17 19 31.1002 $w=3.63e-07 $l=9.85e-07 $layer=LI1_cond $X=0.297 $Y=1.95
+ $X2=0.297 $Y2=0.965
r97 13 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.68
+ $X2=2.375 $Y2=1.515
r98 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.375 $Y=1.68
+ $X2=2.375 $Y2=2.4
r99 10 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.145 $Y=1.35
+ $X2=2.145 $Y2=1.515
r100 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.145 $Y=1.35
+ $X2=2.145 $Y2=0.87
r101 3 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=1.99 $X2=1.28 $Y2=2.135
r102 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.99 $X2=0.28 $Y2=2.135
r103 1 19 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.68 $X2=0.315 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r39 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 27 36 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=2.31 $Y=3.33 $X2=1.94
+ $Y2=3.33
r44 27 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.31 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r48 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 22 36 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33 $X2=1.94
+ $Y2=3.33
r50 22 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r54 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 11 36 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=3.33
r58 11 13 14.062 $w=7.38e-07 $l=8.7e-07 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=2.375
r59 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r60 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=2.455
r61 2 13 150 $w=1.7e-07 $l=7.17112e-07 $layer=licon1_PDIFF $count=4 $X=1.595
+ $Y=1.99 $X2=2.145 $Y2=2.375
r62 1 9 600 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.99 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_1%X 1 2 9 15 17 18 19 27 36
r21 24 27 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=2.622 $Y=1.992
+ $X2=2.622 $Y2=2.015
r22 18 19 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.622 $Y=2.405
+ $X2=2.622 $Y2=2.775
r23 17 24 0.849169 $w=2.83e-07 $l=2.1e-08 $layer=LI1_cond $X=2.622 $Y=1.971
+ $X2=2.622 $Y2=1.992
r24 17 36 6.75432 $w=2.83e-07 $l=1.21e-07 $layer=LI1_cond $X=2.622 $Y=1.971
+ $X2=2.622 $Y2=1.85
r25 17 18 14.1124 $w=2.83e-07 $l=3.49e-07 $layer=LI1_cond $X=2.622 $Y=2.056
+ $X2=2.622 $Y2=2.405
r26 17 27 1.6579 $w=2.83e-07 $l=4.1e-08 $layer=LI1_cond $X=2.622 $Y=2.056
+ $X2=2.622 $Y2=2.015
r27 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.18
+ $X2=2.68 $Y2=1.095
r28 11 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.68 $Y=1.18
+ $X2=2.68 $Y2=1.85
r29 7 15 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.36 $Y=1.095 $X2=2.68
+ $Y2=1.095
r30 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.36 $Y=1.01 $X2=2.36
+ $Y2=0.645
r31 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=2.815
r32 2 27 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=2.015
r33 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.22 $Y=0.5
+ $X2=2.36 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_1%VGND 1 6 11 12 13 23 24
r23 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r24 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r25 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r26 16 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r27 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 13 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r29 13 17 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.24
+ $Y2=0
r30 11 20 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.68
+ $Y2=0
r31 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.86
+ $Y2=0
r32 10 23 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.64
+ $Y2=0
r33 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.86
+ $Y2=0
r34 6 8 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.86 $Y=0.645 $X2=1.86
+ $Y2=1.065
r35 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=0.085 $X2=1.86
+ $Y2=0
r36 4 6 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.86 $Y=0.085 $X2=1.86
+ $Y2=0.645
r37 1 8 182 $w=1.7e-07 $l=5.6438e-07 $layer=licon1_NDIFF $count=1 $X=1.64 $Y=0.6
+ $X2=1.86 $Y2=1.065
r38 1 6 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.6 $X2=1.86 $Y2=0.645
.ends


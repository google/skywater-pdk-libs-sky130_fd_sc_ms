* File: sky130_fd_sc_ms__a32o_1.pxi.spice
* Created: Fri Aug 28 17:07:50 2020
* 
x_PM_SKY130_FD_SC_MS__A32O_1%A_84_48# N_A_84_48#_M1011_d N_A_84_48#_M1002_d
+ N_A_84_48#_M1010_g N_A_84_48#_M1008_g N_A_84_48#_c_62_n N_A_84_48#_c_138_p
+ N_A_84_48#_c_67_n N_A_84_48#_c_134_p N_A_84_48#_c_63_n N_A_84_48#_c_64_n
+ N_A_84_48#_c_65_n N_A_84_48#_c_77_p PM_SKY130_FD_SC_MS__A32O_1%A_84_48#
x_PM_SKY130_FD_SC_MS__A32O_1%A3 N_A3_M1003_g N_A3_M1006_g A3 N_A3_c_155_n
+ N_A3_c_156_n PM_SKY130_FD_SC_MS__A32O_1%A3
x_PM_SKY130_FD_SC_MS__A32O_1%A2 N_A2_M1004_g N_A2_M1007_g A2 N_A2_c_192_n
+ N_A2_c_193_n PM_SKY130_FD_SC_MS__A32O_1%A2
x_PM_SKY130_FD_SC_MS__A32O_1%A1 N_A1_c_221_n N_A1_M1011_g N_A1_M1001_g A1
+ N_A1_c_224_n PM_SKY130_FD_SC_MS__A32O_1%A1
x_PM_SKY130_FD_SC_MS__A32O_1%B1 N_B1_M1002_g N_B1_M1005_g B1 N_B1_c_255_n
+ N_B1_c_256_n N_B1_c_257_n PM_SKY130_FD_SC_MS__A32O_1%B1
x_PM_SKY130_FD_SC_MS__A32O_1%B2 N_B2_M1009_g N_B2_M1000_g B2 N_B2_c_288_n
+ N_B2_c_289_n PM_SKY130_FD_SC_MS__A32O_1%B2
x_PM_SKY130_FD_SC_MS__A32O_1%X N_X_M1010_s N_X_M1008_s N_X_c_313_n N_X_c_314_n
+ N_X_c_310_n X X X PM_SKY130_FD_SC_MS__A32O_1%X
x_PM_SKY130_FD_SC_MS__A32O_1%VPWR N_VPWR_M1008_d N_VPWR_M1004_d N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n VPWR N_VPWR_c_340_n
+ N_VPWR_c_341_n N_VPWR_c_335_n N_VPWR_c_343_n PM_SKY130_FD_SC_MS__A32O_1%VPWR
x_PM_SKY130_FD_SC_MS__A32O_1%A_247_368# N_A_247_368#_M1003_d
+ N_A_247_368#_M1001_d N_A_247_368#_M1000_d N_A_247_368#_c_385_n
+ N_A_247_368#_c_386_n N_A_247_368#_c_395_n N_A_247_368#_c_379_n
+ N_A_247_368#_c_380_n N_A_247_368#_c_381_n N_A_247_368#_c_382_n
+ PM_SKY130_FD_SC_MS__A32O_1%A_247_368#
x_PM_SKY130_FD_SC_MS__A32O_1%VGND N_VGND_M1010_d N_VGND_M1009_d N_VGND_c_419_n
+ N_VGND_c_420_n N_VGND_c_421_n VGND N_VGND_c_422_n N_VGND_c_423_n
+ N_VGND_c_424_n PM_SKY130_FD_SC_MS__A32O_1%VGND
cc_1 VNB N_A_84_48#_M1010_g 0.029153f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_M1008_g 0.0019151f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_3 VNB N_A_84_48#_c_62_n 0.00309123f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.3
cc_4 VNB N_A_84_48#_c_63_n 0.00575673f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_5 VNB N_A_84_48#_c_64_n 0.033022f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_6 VNB N_A_84_48#_c_65_n 0.00655964f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=0.595
cc_7 VNB N_A3_M1003_g 0.00644414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A3 0.0058955f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_9 VNB N_A3_c_155_n 0.030289f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.63
cc_10 VNB N_A3_c_156_n 0.0183757f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_11 VNB N_A2_M1004_g 0.00722527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A2 0.00343145f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_13 VNB N_A2_c_192_n 0.031857f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.63
cc_14 VNB N_A2_c_193_n 0.0173277f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_15 VNB N_A1_c_221_n 0.0199178f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.47
cc_16 VNB N_A1_M1001_g 0.00722527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.00392553f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_18 VNB N_A1_c_224_n 0.0369284f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.02
cc_19 VNB N_B1_M1002_g 0.00659705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_255_n 0.0283596f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.63
cc_21 VNB N_B1_c_256_n 0.00901079f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_22 VNB N_B1_c_257_n 0.018627f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_23 VNB N_B2_M1000_g 0.00976783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB B2 0.0174691f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_B2_c_288_n 0.0398898f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.63
cc_26 VNB N_B2_c_289_n 0.020822f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_27 VNB N_X_c_310_n 0.0247148f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.02
cc_28 VNB X 0.0265914f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.3
cc_29 VNB X 0.0139041f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=0.935
cc_30 VNB N_VPWR_c_335_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.3
cc_31 VNB N_VGND_c_419_n 0.0134045f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.63
cc_32 VNB N_VGND_c_420_n 0.0130142f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_33 VNB N_VGND_c_421_n 0.0401609f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.02
cc_34 VNB N_VGND_c_422_n 0.0692324f $X=-0.19 $Y=-0.245 $X2=2.895 $Y2=1.805
cc_35 VNB N_VGND_c_423_n 0.0277248f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_36 VNB N_VGND_c_424_n 0.251223f $X=-0.19 $Y=-0.245 $X2=2.715 $Y2=0.595
cc_37 VPB N_A_84_48#_M1008_g 0.0304802f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_38 VPB N_A_84_48#_c_67_n 0.0407691f $X=-0.19 $Y=1.66 $X2=2.895 $Y2=1.805
cc_39 VPB N_A_84_48#_c_63_n 0.00228043f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_40 VPB N_A3_M1003_g 0.0228146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A2_M1004_g 0.0237191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A1_M1001_g 0.0230713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_B1_M1002_g 0.0212067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_B2_M1000_g 0.0294154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_X_c_313_n 0.0419191f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.63
cc_46 VPB N_X_c_314_n 0.0142473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_X_c_310_n 0.0075735f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.02
cc_48 VPB N_VPWR_c_336_n 0.0152168f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_49 VPB N_VPWR_c_337_n 0.016943f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.02
cc_50 VPB N_VPWR_c_338_n 0.0228926f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=0.935
cc_51 VPB N_VPWR_c_339_n 0.00632158f $X=-0.19 $Y=1.66 $X2=2.895 $Y2=1.805
cc_52 VPB N_VPWR_c_340_n 0.0191572f $X=-0.19 $Y=1.66 $X2=3.06 $Y2=1.97
cc_53 VPB N_VPWR_c_341_n 0.044059f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.465
cc_54 VPB N_VPWR_c_335_n 0.0810747f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.3
cc_55 VPB N_VPWR_c_343_n 0.00747566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_247_368#_c_379_n 0.019349f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.3
cc_57 VPB N_A_247_368#_c_380_n 0.00356803f $X=-0.19 $Y=1.66 $X2=2.2 $Y2=0.935
cc_58 VPB N_A_247_368#_c_381_n 0.0443725f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.805
cc_59 VPB N_A_247_368#_c_382_n 0.0028233f $X=-0.19 $Y=1.66 $X2=3.06 $Y2=2.65
cc_60 N_A_84_48#_M1008_g N_A3_M1003_g 0.0229225f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_84_48#_c_67_n N_A3_M1003_g 0.0168583f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_62 N_A_84_48#_c_63_n N_A3_M1003_g 0.00357937f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_63 N_A_84_48#_c_64_n N_A3_M1003_g 0.00305056f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_64 N_A_84_48#_c_62_n A3 0.00839161f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_65 N_A_84_48#_c_67_n A3 0.0258645f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_66 N_A_84_48#_c_63_n A3 0.0201492f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_67 N_A_84_48#_c_64_n A3 2.8743e-19 $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_68 N_A_84_48#_c_77_p A3 0.0236883f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_69 N_A_84_48#_M1010_g N_A3_c_155_n 0.00180795f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A_84_48#_c_62_n N_A3_c_155_n 6.05416e-19 $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_71 N_A_84_48#_c_67_n N_A3_c_155_n 0.00104472f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_72 N_A_84_48#_c_63_n N_A3_c_155_n 0.00142581f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_73 N_A_84_48#_c_64_n N_A3_c_155_n 0.0156273f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_74 N_A_84_48#_c_77_p N_A3_c_155_n 0.00103401f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_75 N_A_84_48#_M1010_g N_A3_c_156_n 0.0131011f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A_84_48#_c_62_n N_A3_c_156_n 0.00325245f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_77 N_A_84_48#_c_77_p N_A3_c_156_n 0.0126218f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_78 N_A_84_48#_c_67_n N_A2_M1004_g 0.0128046f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_79 N_A_84_48#_c_67_n A2 0.0242683f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_80 N_A_84_48#_c_77_p A2 0.0217461f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_81 N_A_84_48#_c_67_n N_A2_c_192_n 0.00105037f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_82 N_A_84_48#_c_77_p N_A2_c_192_n 8.47471e-19 $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_83 N_A_84_48#_c_65_n N_A2_c_193_n 0.00192815f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_84 N_A_84_48#_c_77_p N_A2_c_193_n 0.0120996f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_85 N_A_84_48#_c_65_n N_A1_c_221_n 0.0107943f $X=2.715 $Y=0.595 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_84_48#_c_77_p N_A1_c_221_n 0.00902659f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_84_48#_c_67_n N_A1_M1001_g 0.0142526f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_88 N_A_84_48#_c_67_n A1 0.0244553f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_89 N_A_84_48#_c_77_p A1 0.0225348f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_90 N_A_84_48#_c_67_n N_A1_c_224_n 0.00138872f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_91 N_A_84_48#_c_65_n N_A1_c_224_n 0.00323172f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_92 N_A_84_48#_c_67_n N_B1_M1002_g 0.0157556f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_93 N_A_84_48#_c_67_n N_B1_c_255_n 0.00396981f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_94 N_A_84_48#_c_65_n N_B1_c_255_n 0.00112001f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_95 N_A_84_48#_c_67_n N_B1_c_256_n 0.0356446f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_96 N_A_84_48#_c_65_n N_B1_c_256_n 0.0260766f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_97 N_A_84_48#_c_65_n N_B1_c_257_n 0.0111626f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_98 N_A_84_48#_c_67_n N_B2_M1000_g 0.00365076f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_99 N_A_84_48#_c_65_n N_B2_c_289_n 0.0016581f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_100 N_A_84_48#_M1008_g N_X_c_313_n 0.013446f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_84_48#_M1008_g N_X_c_314_n 0.00416785f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_84_48#_c_63_n N_X_c_314_n 0.00569781f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_103 N_A_84_48#_c_64_n N_X_c_314_n 2.36763e-19 $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_104 N_A_84_48#_M1010_g N_X_c_310_n 0.0100159f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_84_48#_M1008_g N_X_c_310_n 0.00306277f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_84_48#_c_62_n N_X_c_310_n 0.00523589f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_107 N_A_84_48#_c_63_n N_X_c_310_n 0.0315479f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_108 N_A_84_48#_M1010_g X 0.0142066f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_84_48#_M1010_g X 0.00287471f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_84_48#_c_62_n X 0.00468197f $X=0.71 $Y=1.3 $X2=0 $Y2=0
cc_111 N_A_84_48#_c_63_n X 0.00152458f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_112 N_A_84_48#_c_67_n N_VPWR_M1008_d 0.00236156f $X=2.895 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_84_48#_c_63_n N_VPWR_M1008_d 0.00183989f $X=0.59 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_84_48#_c_67_n N_VPWR_M1004_d 0.00529506f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_115 N_A_84_48#_M1008_g N_VPWR_c_336_n 0.00925629f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A_84_48#_c_67_n N_VPWR_c_336_n 0.0164793f $X=2.895 $Y=1.805 $X2=0 $Y2=0
cc_117 N_A_84_48#_c_63_n N_VPWR_c_336_n 0.0119915f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_118 N_A_84_48#_c_64_n N_VPWR_c_336_n 5.07508e-19 $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_119 N_A_84_48#_M1008_g N_VPWR_c_340_n 0.005209f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_84_48#_M1008_g N_VPWR_c_335_n 0.00990503f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_84_48#_c_67_n N_A_247_368#_M1003_d 0.00165831f $X=2.895 $Y=1.805
+ $X2=-0.19 $Y2=-0.245
cc_122 N_A_84_48#_c_67_n N_A_247_368#_M1001_d 0.00165831f $X=2.895 $Y=1.805
+ $X2=0 $Y2=0
cc_123 N_A_84_48#_c_67_n N_A_247_368#_c_385_n 0.0526608f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_124 N_A_84_48#_c_67_n N_A_247_368#_c_386_n 0.0171782f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_125 N_A_84_48#_c_134_p N_A_247_368#_c_379_n 0.0225479f $X=3.06 $Y=1.97 $X2=0
+ $Y2=0
cc_126 N_A_84_48#_c_67_n N_A_247_368#_c_381_n 0.00352479f $X=2.895 $Y=1.805
+ $X2=0 $Y2=0
cc_127 N_A_84_48#_c_67_n N_A_247_368#_c_382_n 0.0171782f $X=2.895 $Y=1.805 $X2=0
+ $Y2=0
cc_128 N_A_84_48#_c_62_n N_VGND_M1010_d 0.00198882f $X=0.71 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_84_48#_c_138_p N_VGND_M1010_d 0.00372868f $X=0.795 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_84_48#_c_77_p N_VGND_M1010_d 0.0125332f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_84_48#_M1010_g N_VGND_c_419_n 0.00811597f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_84_48#_c_138_p N_VGND_c_419_n 0.0126823f $X=0.795 $Y=0.935 $X2=0
+ $Y2=0
cc_133 N_A_84_48#_c_64_n N_VGND_c_419_n 3.34594e-19 $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_134 N_A_84_48#_c_77_p N_VGND_c_419_n 0.0201945f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_135 N_A_84_48#_c_65_n N_VGND_c_421_n 0.0197562f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_136 N_A_84_48#_c_65_n N_VGND_c_422_n 0.0224837f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_137 N_A_84_48#_M1010_g N_VGND_c_423_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_84_48#_M1010_g N_VGND_c_424_n 0.00829501f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_84_48#_c_138_p N_VGND_c_424_n 0.00149237f $X=0.795 $Y=0.935 $X2=0
+ $Y2=0
cc_140 N_A_84_48#_c_65_n N_VGND_c_424_n 0.0236713f $X=2.715 $Y=0.595 $X2=0 $Y2=0
cc_141 N_A_84_48#_c_77_p N_VGND_c_424_n 0.0387864f $X=2.2 $Y=0.725 $X2=0 $Y2=0
cc_142 N_A_84_48#_c_77_p A_259_94# 0.00736231f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_84_48#_c_77_p A_337_94# 0.013672f $X=2.2 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A3_M1003_g N_A2_M1004_g 0.0341796f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_145 A3 A2 0.0264591f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A3_c_155_n A2 3.99347e-19 $X=1.13 $Y=1.385 $X2=0 $Y2=0
cc_147 A3 N_A2_c_192_n 0.00188716f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A3_c_155_n N_A2_c_192_n 0.0206935f $X=1.13 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A3_c_156_n N_A2_c_193_n 0.049285f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A3_M1003_g N_X_c_314_n 9.5102e-19 $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_151 N_A3_M1003_g N_VPWR_c_336_n 0.00889127f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_152 N_A3_M1003_g N_VPWR_c_338_n 0.00567889f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_153 N_A3_M1003_g N_VPWR_c_335_n 0.00610055f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_154 N_A3_M1003_g N_A_247_368#_c_382_n 0.0119778f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_155 N_A3_c_156_n N_VGND_c_419_n 0.010194f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_156 N_A3_c_156_n N_VGND_c_422_n 0.00507111f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A3_c_156_n N_VGND_c_424_n 0.00514438f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A2_c_193_n N_A1_c_221_n 0.0291659f $X=1.67 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_159 N_A2_M1004_g N_A1_M1001_g 0.0265417f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_160 A2 A1 0.0230669f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A2_c_192_n A1 0.00114936f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_162 A2 N_A1_c_224_n 0.00118009f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A2_c_192_n N_A1_c_224_n 0.0203272f $X=1.67 $Y=1.385 $X2=0 $Y2=0
cc_164 N_A2_M1004_g N_VPWR_c_337_n 0.00828775f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_165 N_A2_M1004_g N_VPWR_c_338_n 0.00567889f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_166 N_A2_M1004_g N_VPWR_c_335_n 0.00610055f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_167 N_A2_M1004_g N_A_247_368#_c_385_n 0.0141331f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_168 N_A2_M1004_g N_A_247_368#_c_382_n 0.0168859f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_169 N_A2_c_193_n N_VGND_c_422_n 0.00507111f $X=1.67 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A2_c_193_n N_VGND_c_424_n 0.00514438f $X=1.67 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A1_M1001_g N_B1_M1002_g 0.0338978f $X=2.335 $Y=2.34 $X2=0 $Y2=0
cc_172 A1 N_B1_c_255_n 3.04283e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A1_c_224_n N_B1_c_255_n 0.0165415f $X=2.335 $Y=1.385 $X2=0 $Y2=0
cc_174 A1 N_B1_c_256_n 0.0293561f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A1_c_224_n N_B1_c_256_n 0.002359f $X=2.335 $Y=1.385 $X2=0 $Y2=0
cc_176 N_A1_c_221_n N_B1_c_257_n 0.00495039f $X=2.15 $Y=1.22 $X2=0 $Y2=0
cc_177 N_A1_M1001_g N_VPWR_c_337_n 0.00639768f $X=2.335 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A1_M1001_g N_VPWR_c_341_n 0.00508554f $X=2.335 $Y=2.34 $X2=0 $Y2=0
cc_179 N_A1_M1001_g N_VPWR_c_335_n 0.00508379f $X=2.335 $Y=2.34 $X2=0 $Y2=0
cc_180 N_A1_M1001_g N_A_247_368#_c_385_n 0.0141331f $X=2.335 $Y=2.34 $X2=0 $Y2=0
cc_181 N_A1_M1001_g N_A_247_368#_c_386_n 8.84614e-19 $X=2.335 $Y=2.34 $X2=0
+ $Y2=0
cc_182 N_A1_M1001_g N_A_247_368#_c_395_n 0.0167732f $X=2.335 $Y=2.34 $X2=0 $Y2=0
cc_183 N_A1_M1001_g N_A_247_368#_c_380_n 0.00216107f $X=2.335 $Y=2.34 $X2=0
+ $Y2=0
cc_184 N_A1_c_221_n N_VGND_c_422_n 0.00484285f $X=2.15 $Y=1.22 $X2=0 $Y2=0
cc_185 N_A1_c_221_n N_VGND_c_424_n 0.00514438f $X=2.15 $Y=1.22 $X2=0 $Y2=0
cc_186 N_B1_M1002_g N_B2_M1000_g 0.0141471f $X=2.785 $Y=2.34 $X2=0 $Y2=0
cc_187 N_B1_c_256_n B2 0.017611f $X=2.84 $Y=1.385 $X2=0 $Y2=0
cc_188 N_B1_c_257_n B2 4.01112e-19 $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_189 N_B1_c_255_n N_B2_c_288_n 0.031246f $X=2.84 $Y=1.385 $X2=0 $Y2=0
cc_190 N_B1_c_256_n N_B2_c_289_n 0.00143086f $X=2.84 $Y=1.385 $X2=0 $Y2=0
cc_191 N_B1_c_257_n N_B2_c_289_n 0.031246f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_192 N_B1_M1002_g N_VPWR_c_341_n 8.89343e-19 $X=2.785 $Y=2.34 $X2=0 $Y2=0
cc_193 N_B1_M1002_g N_A_247_368#_c_386_n 0.00235686f $X=2.785 $Y=2.34 $X2=0
+ $Y2=0
cc_194 N_B1_M1002_g N_A_247_368#_c_395_n 0.0114522f $X=2.785 $Y=2.34 $X2=0 $Y2=0
cc_195 N_B1_M1002_g N_A_247_368#_c_379_n 0.0108527f $X=2.785 $Y=2.34 $X2=0 $Y2=0
cc_196 N_B1_M1002_g N_A_247_368#_c_380_n 0.00141162f $X=2.785 $Y=2.34 $X2=0
+ $Y2=0
cc_197 N_B1_M1002_g N_A_247_368#_c_381_n 4.77651e-19 $X=2.785 $Y=2.34 $X2=0
+ $Y2=0
cc_198 N_B1_c_257_n N_VGND_c_421_n 0.0022187f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_199 N_B1_c_257_n N_VGND_c_422_n 0.00484285f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_200 N_B1_c_257_n N_VGND_c_424_n 0.00514438f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_201 N_B2_M1000_g N_VPWR_c_341_n 8.89343e-19 $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_202 N_B2_M1000_g N_A_247_368#_c_395_n 3.82257e-19 $X=3.335 $Y=2.34 $X2=0
+ $Y2=0
cc_203 N_B2_M1000_g N_A_247_368#_c_379_n 0.0128353f $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_204 N_B2_M1000_g N_A_247_368#_c_381_n 0.0161517f $X=3.335 $Y=2.34 $X2=0 $Y2=0
cc_205 B2 N_A_247_368#_c_381_n 0.0193705f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_206 N_B2_c_288_n N_A_247_368#_c_381_n 0.00429583f $X=3.455 $Y=1.385 $X2=0
+ $Y2=0
cc_207 B2 N_VGND_c_421_n 0.0257644f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_208 N_B2_c_288_n N_VGND_c_421_n 0.00156161f $X=3.455 $Y=1.385 $X2=0 $Y2=0
cc_209 N_B2_c_289_n N_VGND_c_421_n 0.0151934f $X=3.432 $Y=1.22 $X2=0 $Y2=0
cc_210 N_B2_c_289_n N_VGND_c_422_n 0.00421418f $X=3.432 $Y=1.22 $X2=0 $Y2=0
cc_211 N_B2_c_289_n N_VGND_c_424_n 0.00432128f $X=3.432 $Y=1.22 $X2=0 $Y2=0
cc_212 N_X_c_313_n N_VPWR_c_336_n 0.0359411f $X=0.29 $Y=2.815 $X2=0 $Y2=0
cc_213 N_X_c_313_n N_VPWR_c_340_n 0.0163338f $X=0.29 $Y=2.815 $X2=0 $Y2=0
cc_214 N_X_c_313_n N_VPWR_c_335_n 0.0134516f $X=0.29 $Y=2.815 $X2=0 $Y2=0
cc_215 X N_VGND_c_419_n 0.0226903f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_216 X N_VGND_c_423_n 0.0159025f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_217 X N_VGND_c_424_n 0.0131064f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_218 N_VPWR_M1004_d N_A_247_368#_c_385_n 0.014331f $X=1.685 $Y=1.84 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_337_n N_A_247_368#_c_385_n 0.0266856f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_337_n N_A_247_368#_c_395_n 0.0279702f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_341_n N_A_247_368#_c_379_n 0.0667586f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_335_n N_A_247_368#_c_379_n 0.0380121f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_337_n N_A_247_368#_c_380_n 0.0107169f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_341_n N_A_247_368#_c_380_n 0.0236566f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_335_n N_A_247_368#_c_380_n 0.0128296f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_226 N_VPWR_c_336_n N_A_247_368#_c_382_n 0.0223391f $X=0.85 $Y=2.225 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_337_n N_A_247_368#_c_382_n 0.0254386f $X=1.965 $Y=2.565 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_338_n N_A_247_368#_c_382_n 0.00967309f $X=1.8 $Y=3.33 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_335_n N_A_247_368#_c_382_n 0.0111395f $X=3.6 $Y=3.33 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__xor3_4.spice
* Created: Wed Sep  2 12:34:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xor3_4.pex.spice"
.subckt sky130_fd_sc_ms__xor3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_74_294#_M1005_g N_A_27_118#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.24225 AS=0.1824 PD=1.57 PS=1.85 NRD=60.648 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1023 N_A_74_294#_M1023_d N_A_M1023_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.2208 AS=0.24225 PD=1.33 PS=1.57 NRD=29.988 NRS=60.648 M=1 R=4.26667
+ SA=75000.9 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1013 N_A_416_118#_M1013_d N_B_M1013_g N_A_74_294#_M1023_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.125283 AS=0.2208 PD=1.19547 PS=1.33 NRD=0 NRS=46.872 M=1 R=4.26667
+ SA=75001.7 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1018 N_A_27_118#_M1018_d N_A_397_320#_M1018_g N_A_416_118#_M1013_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0966792 AS=0.082217 PD=0.863774 PS=0.784528 NRD=0
+ NRS=20.712 M=1 R=2.8 SA=75002.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_326_392#_M1006_d N_B_M1006_g N_A_27_118#_M1018_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.145875 AS=0.147321 PD=1.115 PS=1.31623 NRD=14.988 NRS=31.872 M=1
+ R=4.26667 SA=75001.9 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1027 N_A_74_294#_M1027_d N_A_397_320#_M1027_g N_A_326_392#_M1006_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2848 AS=0.145875 PD=2.17 PS=1.115 NRD=31.872 NRS=14.988 M=1
+ R=4.26667 SA=75002.5 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_B_M1024_g N_A_397_320#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.42 AS=0.2072 PD=2.67 PS=2.04 NRD=41.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1008 N_A_1221_388#_M1008_d N_A_1155_284#_M1008_g N_A_326_392#_M1008_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1696 AS=0.176 PD=1.17 PS=1.83 NRD=46.872 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1016 N_A_416_118#_M1016_d N_C_M1016_g N_A_1221_388#_M1008_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1696 PD=1.85 PS=1.17 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_1155_284#_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.106521 AS=0.2121 PD=0.847241 PS=1.85 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.4 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1001_d N_A_1221_388#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.187679 AS=0.1036 PD=1.49276 PS=1.02 NRD=5.664 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_1221_388#_M1010_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1010_d N_A_1221_388#_M1011_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_1221_388#_M1020_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A_74_294#_M1002_g N_A_27_118#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1025 N_A_74_294#_M1025_d N_A_M1025_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.186413 AS=0.16 PD=1.47283 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90000.7 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1009 N_A_326_392#_M1009_d N_B_M1009_g N_A_74_294#_M1025_d VPB PSHORT L=0.18
+ W=0.84 AD=0.160735 AS=0.156587 PD=1.35649 PS=1.23717 NRD=0 NRS=19.1484 M=1
+ R=4.66667 SA=90001.2 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1019 N_A_27_118#_M1019_d N_A_397_320#_M1019_g N_A_326_392#_M1009_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.140275 AS=0.122465 PD=1.185 PS=1.03351 NRD=0 NRS=25.3933
+ M=1 R=3.55556 SA=90001.8 SB=90001.4 A=0.1152 P=1.64 MULT=1
MM1021 N_A_416_118#_M1021_d N_B_M1021_g N_A_27_118#_M1019_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1224 AS=0.140275 PD=1.03351 PS=1.185 NRD=24.6053 NRS=43.0839 M=1
+ R=3.55556 SA=90001.9 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1014 N_A_74_294#_M1014_d N_A_397_320#_M1014_g N_A_416_118#_M1021_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.5334 AS=0.16065 PD=2.95 PS=1.35649 NRD=71.511 NRS=0 M=1
+ R=4.66667 SA=90001.9 SB=90000.5 A=0.1512 P=2.04 MULT=1
MM1015 N_VPWR_M1015_d N_B_M1015_g N_A_397_320#_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1003 N_A_1221_388#_M1003_d N_A_1155_284#_M1003_g N_A_416_118#_M1003_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.21 AS=0.3696 PD=1.34 PS=2.56 NRD=52.7566 NRS=36.3465
+ M=1 R=4.66667 SA=90000.3 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1007 N_A_326_392#_M1007_d N_C_M1007_g N_A_1221_388#_M1003_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.21 PD=2.24 PS=1.34 NRD=0 NRS=0 M=1 R=4.66667 SA=90001
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_A_1155_284#_M1000_s VPB PSHORT L=0.18 W=0.64
+ AD=0.282182 AS=0.1792 PD=1.34182 PS=1.84 NRD=118.771 NRS=0 M=1 R=3.55556
+ SA=90000.2 SB=90002.5 A=0.1152 P=1.64 MULT=1
MM1012 N_X_M1012_d N_A_1221_388#_M1012_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.493818 PD=1.39 PS=2.34818 NRD=0 NRS=64.1826 M=1 R=6.22222
+ SA=90000.9 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1017 N_X_M1012_d N_A_1221_388#_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196 PD=1.39 PS=1.47 NRD=0 NRS=13.1793 M=1 R=6.22222 SA=90001.3
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1022 N_X_M1022_d N_A_1221_388#_M1022_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196 PD=1.39 PS=1.47 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.8
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1026 N_X_M1022_d N_A_1221_388#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=20.3484 P=25.6
c_208 VPB 0 1.12299e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__xor3_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfrtp_2.pxi.spice
* Created: Fri Aug 28 17:23:02 2020
* 
x_PM_SKY130_FD_SC_MS__DFRTP_2%D N_D_c_242_n N_D_M1014_g N_D_M1028_g D D D
+ N_D_c_244_n N_D_c_245_n N_D_c_249_n PM_SKY130_FD_SC_MS__DFRTP_2%D
x_PM_SKY130_FD_SC_MS__DFRTP_2%CLK N_CLK_M1016_g N_CLK_M1025_g CLK N_CLK_c_274_n
+ N_CLK_c_275_n PM_SKY130_FD_SC_MS__DFRTP_2%CLK
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_493_387# N_A_493_387#_M1013_d
+ N_A_493_387#_M1027_d N_A_493_387#_c_336_n N_A_493_387#_M1004_g
+ N_A_493_387#_c_338_n N_A_493_387#_c_318_n N_A_493_387#_M1024_g
+ N_A_493_387#_c_320_n N_A_493_387#_M1003_g N_A_493_387#_c_321_n
+ N_A_493_387#_c_322_n N_A_493_387#_M1009_g N_A_493_387#_c_323_n
+ N_A_493_387#_c_324_n N_A_493_387#_c_325_n N_A_493_387#_c_326_n
+ N_A_493_387#_c_327_n N_A_493_387#_c_368_p N_A_493_387#_c_328_n
+ N_A_493_387#_c_329_n N_A_493_387#_c_330_n N_A_493_387#_c_331_n
+ N_A_493_387#_c_332_n N_A_493_387#_c_333_n N_A_493_387#_c_334_n
+ N_A_493_387#_c_335_n N_A_493_387#_c_344_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%A_493_387#
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_837_359# N_A_837_359#_M1023_d
+ N_A_837_359#_M1000_d N_A_837_359#_M1011_g N_A_837_359#_M1008_g
+ N_A_837_359#_c_516_n N_A_837_359#_c_523_n N_A_837_359#_c_517_n
+ N_A_837_359#_c_537_n N_A_837_359#_c_539_n N_A_837_359#_c_524_n
+ N_A_837_359#_c_518_n N_A_837_359#_c_519_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%A_837_359#
x_PM_SKY130_FD_SC_MS__DFRTP_2%RESET_B N_RESET_B_M1012_g N_RESET_B_c_601_n
+ N_RESET_B_M1015_g N_RESET_B_c_602_n N_RESET_B_c_603_n N_RESET_B_M1001_g
+ N_RESET_B_c_605_n N_RESET_B_M1017_g N_RESET_B_M1019_g N_RESET_B_M1021_g
+ N_RESET_B_c_607_n N_RESET_B_c_616_n N_RESET_B_c_617_n N_RESET_B_c_618_n
+ N_RESET_B_c_619_n N_RESET_B_c_620_n N_RESET_B_c_621_n RESET_B
+ N_RESET_B_c_608_n N_RESET_B_c_609_n N_RESET_B_c_623_n N_RESET_B_c_624_n
+ N_RESET_B_c_625_n N_RESET_B_c_626_n PM_SKY130_FD_SC_MS__DFRTP_2%RESET_B
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_699_463# N_A_699_463#_M1026_d
+ N_A_699_463#_M1004_d N_A_699_463#_M1017_d N_A_699_463#_M1023_g
+ N_A_699_463#_M1000_g N_A_699_463#_c_811_n N_A_699_463#_c_812_n
+ N_A_699_463#_c_813_n N_A_699_463#_c_821_n N_A_699_463#_c_822_n
+ N_A_699_463#_c_823_n N_A_699_463#_c_814_n N_A_699_463#_c_815_n
+ N_A_699_463#_c_825_n N_A_699_463#_c_816_n N_A_699_463#_c_826_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%A_699_463#
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_306_119# N_A_306_119#_M1016_s
+ N_A_306_119#_M1025_s N_A_306_119#_M1027_g N_A_306_119#_c_930_n
+ N_A_306_119#_M1013_g N_A_306_119#_c_941_n N_A_306_119#_c_942_n
+ N_A_306_119#_c_943_n N_A_306_119#_c_931_n N_A_306_119#_c_932_n
+ N_A_306_119#_c_933_n N_A_306_119#_M1026_g N_A_306_119#_M1006_g
+ N_A_306_119#_c_946_n N_A_306_119#_M1007_g N_A_306_119#_c_934_n
+ N_A_306_119#_c_949_n N_A_306_119#_M1032_g N_A_306_119#_c_950_n
+ N_A_306_119#_c_936_n N_A_306_119#_c_937_n N_A_306_119#_c_965_n
+ N_A_306_119#_c_938_n N_A_306_119#_c_939_n N_A_306_119#_c_953_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%A_306_119#
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_1525_212# N_A_1525_212#_M1022_d
+ N_A_1525_212#_M1019_d N_A_1525_212#_M1005_g N_A_1525_212#_c_1117_n
+ N_A_1525_212#_M1018_g N_A_1525_212#_c_1109_n N_A_1525_212#_c_1110_n
+ N_A_1525_212#_c_1120_n N_A_1525_212#_c_1111_n N_A_1525_212#_c_1121_n
+ N_A_1525_212#_c_1122_n N_A_1525_212#_c_1123_n N_A_1525_212#_c_1112_n
+ N_A_1525_212#_c_1113_n N_A_1525_212#_c_1114_n N_A_1525_212#_c_1115_n
+ N_A_1525_212#_c_1116_n PM_SKY130_FD_SC_MS__DFRTP_2%A_1525_212#
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_1271_74# N_A_1271_74#_M1003_d
+ N_A_1271_74#_M1007_d N_A_1271_74#_M1022_g N_A_1271_74#_M1002_g
+ N_A_1271_74#_c_1223_n N_A_1271_74#_c_1224_n N_A_1271_74#_M1010_g
+ N_A_1271_74#_M1020_g N_A_1271_74#_c_1226_n N_A_1271_74#_c_1244_n
+ N_A_1271_74#_c_1227_n N_A_1271_74#_c_1237_n N_A_1271_74#_c_1228_n
+ N_A_1271_74#_c_1258_n N_A_1271_74#_c_1346_p N_A_1271_74#_c_1238_n
+ N_A_1271_74#_c_1229_n N_A_1271_74#_c_1230_n N_A_1271_74#_c_1231_n
+ N_A_1271_74#_c_1242_n PM_SKY130_FD_SC_MS__DFRTP_2%A_1271_74#
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_1924_409# N_A_1924_409#_M1020_d
+ N_A_1924_409#_M1010_d N_A_1924_409#_c_1362_n N_A_1924_409#_M1029_g
+ N_A_1924_409#_M1031_g N_A_1924_409#_c_1365_n N_A_1924_409#_M1030_g
+ N_A_1924_409#_M1033_g N_A_1924_409#_c_1368_n N_A_1924_409#_c_1369_n
+ N_A_1924_409#_c_1376_n N_A_1924_409#_c_1370_n N_A_1924_409#_c_1371_n
+ N_A_1924_409#_c_1372_n N_A_1924_409#_c_1373_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%A_1924_409#
x_PM_SKY130_FD_SC_MS__DFRTP_2%VPWR N_VPWR_M1014_s N_VPWR_M1015_d N_VPWR_M1025_d
+ N_VPWR_M1011_d N_VPWR_M1000_s N_VPWR_M1018_d N_VPWR_M1002_d N_VPWR_M1029_s
+ N_VPWR_M1030_s N_VPWR_c_1430_n N_VPWR_c_1431_n N_VPWR_c_1432_n N_VPWR_c_1433_n
+ N_VPWR_c_1434_n N_VPWR_c_1435_n N_VPWR_c_1436_n N_VPWR_c_1437_n
+ N_VPWR_c_1438_n N_VPWR_c_1439_n N_VPWR_c_1440_n N_VPWR_c_1441_n
+ N_VPWR_c_1442_n N_VPWR_c_1443_n VPWR N_VPWR_c_1444_n N_VPWR_c_1445_n
+ N_VPWR_c_1446_n N_VPWR_c_1447_n N_VPWR_c_1448_n N_VPWR_c_1449_n
+ N_VPWR_c_1450_n N_VPWR_c_1451_n N_VPWR_c_1452_n N_VPWR_c_1453_n
+ N_VPWR_c_1454_n N_VPWR_c_1455_n N_VPWR_c_1429_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%VPWR
x_PM_SKY130_FD_SC_MS__DFRTP_2%A_30_78# N_A_30_78#_M1028_s N_A_30_78#_M1026_s
+ N_A_30_78#_M1014_d N_A_30_78#_M1004_s N_A_30_78#_c_1581_n N_A_30_78#_c_1587_n
+ N_A_30_78#_c_1582_n N_A_30_78#_c_1589_n N_A_30_78#_c_1583_n
+ N_A_30_78#_c_1590_n N_A_30_78#_c_1591_n N_A_30_78#_c_1584_n
+ N_A_30_78#_c_1585_n N_A_30_78#_c_1593_n N_A_30_78#_c_1594_n
+ N_A_30_78#_c_1595_n N_A_30_78#_c_1586_n PM_SKY130_FD_SC_MS__DFRTP_2%A_30_78#
x_PM_SKY130_FD_SC_MS__DFRTP_2%Q N_Q_M1031_d N_Q_M1029_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__DFRTP_2%Q
x_PM_SKY130_FD_SC_MS__DFRTP_2%VGND N_VGND_M1012_d N_VGND_M1016_d N_VGND_M1001_d
+ N_VGND_M1005_d N_VGND_M1020_s N_VGND_M1031_s N_VGND_M1033_s N_VGND_c_1723_n
+ N_VGND_c_1724_n N_VGND_c_1725_n N_VGND_c_1726_n N_VGND_c_1727_n
+ N_VGND_c_1728_n N_VGND_c_1729_n N_VGND_c_1730_n N_VGND_c_1731_n VGND
+ N_VGND_c_1732_n N_VGND_c_1733_n N_VGND_c_1734_n N_VGND_c_1735_n
+ N_VGND_c_1736_n N_VGND_c_1737_n N_VGND_c_1738_n N_VGND_c_1739_n
+ N_VGND_c_1740_n N_VGND_c_1741_n N_VGND_c_1742_n
+ PM_SKY130_FD_SC_MS__DFRTP_2%VGND
cc_1 VNB N_D_c_242_n 0.040598f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.828
cc_2 VNB N_D_M1028_g 0.0286454f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_3 VNB N_D_c_244_n 0.0216261f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_245_n 0.0279969f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB CLK 0.00300522f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_6 VNB N_CLK_c_274_n 0.0210699f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_CLK_c_275_n 0.0172003f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_8 VNB N_A_493_387#_c_318_n 0.0121631f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_9 VNB N_A_493_387#_M1024_g 0.0232206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_493_387#_c_320_n 0.0178063f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_11 VNB N_A_493_387#_c_321_n 0.0205353f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_12 VNB N_A_493_387#_c_322_n 0.010064f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_13 VNB N_A_493_387#_c_323_n 0.0092862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_493_387#_c_324_n 0.0306116f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_15 VNB N_A_493_387#_c_325_n 4.48828e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_16 VNB N_A_493_387#_c_326_n 7.02729e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_493_387#_c_327_n 0.00324493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_493_387#_c_328_n 0.0145916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_493_387#_c_329_n 0.00228045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_493_387#_c_330_n 0.0036821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_493_387#_c_331_n 0.00197952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_493_387#_c_332_n 0.0149739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_493_387#_c_333_n 0.00719103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_493_387#_c_334_n 0.0318573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_493_387#_c_335_n 0.00728799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_837_359#_M1008_g 0.0283695f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_27 VNB N_A_837_359#_c_516_n 0.00259049f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_28 VNB N_A_837_359#_c_517_n 0.0109483f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_29 VNB N_A_837_359#_c_518_n 0.00239189f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.035
cc_30 VNB N_A_837_359#_c_519_n 0.00880031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_RESET_B_M1012_g 0.0210264f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.845
cc_32 VNB N_RESET_B_c_601_n 0.0249344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_602_n 0.281591f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_RESET_B_c_603_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_RESET_B_M1001_g 0.034622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_RESET_B_c_605_n 0.0106864f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_37 VNB N_RESET_B_M1021_g 0.0519208f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_38 VNB N_RESET_B_c_607_n 0.0158834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_c_608_n 0.0298051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_609_n 0.00416334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_699_463#_M1023_g 0.0236184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_42 VNB N_A_699_463#_c_811_n 0.026897f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_43 VNB N_A_699_463#_c_812_n 0.0170696f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_44 VNB N_A_699_463#_c_813_n 0.00512369f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.845
cc_45 VNB N_A_699_463#_c_814_n 0.00251544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_699_463#_c_815_n 0.00408962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_699_463#_c_816_n 0.00232245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_306_119#_c_930_n 0.0151539f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_49 VNB N_A_306_119#_c_931_n 0.0335538f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_50 VNB N_A_306_119#_c_932_n 0.0609424f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_51 VNB N_A_306_119#_c_933_n 0.0162512f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_52 VNB N_A_306_119#_c_934_n 0.0126064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_306_119#_M1032_g 0.0521291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_306_119#_c_936_n 0.00783205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_306_119#_c_937_n 0.00751406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_306_119#_c_938_n 4.50268e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_306_119#_c_939_n 0.00281154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1525_212#_M1005_g 0.0235036f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_59 VNB N_A_1525_212#_c_1109_n 0.013872f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_60 VNB N_A_1525_212#_c_1110_n 0.0150411f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_61 VNB N_A_1525_212#_c_1111_n 0.0124228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1525_212#_c_1112_n 0.0141072f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=2.035
cc_63 VNB N_A_1525_212#_c_1113_n 0.00326635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1525_212#_c_1114_n 0.00415979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1525_212#_c_1115_n 0.031534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1525_212#_c_1116_n 0.00288865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1271_74#_M1022_g 0.0561848f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_68 VNB N_A_1271_74#_c_1223_n 0.0155616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1271_74#_c_1224_n 0.0127478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1271_74#_M1020_g 0.0397312f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_71 VNB N_A_1271_74#_c_1226_n 0.00460889f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.165
cc_72 VNB N_A_1271_74#_c_1227_n 0.00477322f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.295
cc_73 VNB N_A_1271_74#_c_1228_n 0.00415183f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=2.035
cc_74 VNB N_A_1271_74#_c_1229_n 0.00523477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1271_74#_c_1230_n 0.00751489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1271_74#_c_1231_n 0.00236307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1924_409#_c_1362_n 0.0140421f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1
cc_78 VNB N_A_1924_409#_M1029_g 0.0102109f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_79 VNB N_A_1924_409#_M1031_g 0.0229651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1924_409#_c_1365_n 0.00938445f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_81 VNB N_A_1924_409#_M1030_g 0.0167069f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.845
cc_82 VNB N_A_1924_409#_M1033_g 0.0260342f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.165
cc_83 VNB N_A_1924_409#_c_1368_n 0.00594745f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.295
cc_84 VNB N_A_1924_409#_c_1369_n 0.0111562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1924_409#_c_1370_n 0.0124224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1924_409#_c_1371_n 0.00109385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1924_409#_c_1372_n 0.00157695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1924_409#_c_1373_n 0.0465967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VPWR_c_1429_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_30_78#_c_1581_n 0.00271393f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_91 VNB N_A_30_78#_c_1582_n 0.00538705f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_92 VNB N_A_30_78#_c_1583_n 0.00219226f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.295
cc_93 VNB N_A_30_78#_c_1584_n 0.00309813f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.035
cc_94 VNB N_A_30_78#_c_1585_n 0.0223919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_30_78#_c_1586_n 0.0064063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1
cc_97 VNB N_VGND_c_1723_n 0.0156168f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_98 VNB N_VGND_c_1724_n 0.0160979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1725_n 0.00612754f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.035
cc_100 VNB N_VGND_c_1726_n 0.0164559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1727_n 0.0191664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1728_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1729_n 0.0507342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1730_n 0.0298099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1731_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1732_n 0.0190943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1733_n 0.0794975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1734_n 0.0578377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1735_n 0.0306389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1736_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1737_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1738_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1739_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1740_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1741_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1742_n 0.608208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VPB N_D_c_242_n 0.0142136f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.828
cc_118 VPB N_D_M1014_g 0.0619609f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.845
cc_119 VPB N_D_c_245_n 0.0227717f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_120 VPB N_D_c_249_n 0.0207699f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_121 VPB N_CLK_M1025_g 0.0245882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB CLK 0.00437152f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_123 VPB N_CLK_c_274_n 0.0110909f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_124 VPB N_A_493_387#_c_336_n 0.0297182f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_125 VPB N_A_493_387#_M1004_g 0.0322988f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_126 VPB N_A_493_387#_c_338_n 0.0223645f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_127 VPB N_A_493_387#_c_318_n 0.0141267f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_128 VPB N_A_493_387#_M1009_g 0.0264133f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_129 VPB N_A_493_387#_c_325_n 0.00712057f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_130 VPB N_A_493_387#_c_326_n 0.00133074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_493_387#_c_330_n 0.00603671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_493_387#_c_344_n 0.0415192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_837_359#_M1011_g 0.0217191f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_134 VPB N_A_837_359#_M1008_g 0.0130466f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_135 VPB N_A_837_359#_c_516_n 0.00239255f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_136 VPB N_A_837_359#_c_523_n 0.0389792f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_137 VPB N_A_837_359#_c_524_n 5.83055e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_837_359#_c_519_n 0.00374365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_RESET_B_c_601_n 0.022558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_M1015_g 0.0484082f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_141 VPB N_RESET_B_c_605_n 0.0183715f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_142 VPB N_RESET_B_M1017_g 0.0261582f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_143 VPB N_RESET_B_M1019_g 0.0260486f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.165
cc_144 VPB N_RESET_B_M1021_g 0.0162636f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_145 VPB N_RESET_B_c_616_n 0.0210083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_c_617_n 0.00526925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_618_n 0.020195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_c_619_n 0.00143938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_620_n 0.003966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_621_n 0.0019787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_609_n 0.00148599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_623_n 0.0269084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_624_n 0.0461593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_625_n 0.0310686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_626_n 0.00930396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_699_463#_M1000_g 0.0256462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_699_463#_c_811_n 0.0122975f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_158 VPB N_A_699_463#_c_812_n 0.00327673f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_159 VPB N_A_699_463#_c_813_n 0.00685279f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_160 VPB N_A_699_463#_c_821_n 0.00171693f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_161 VPB N_A_699_463#_c_822_n 0.00630961f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_162 VPB N_A_699_463#_c_823_n 0.0113177f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.165
cc_163 VPB N_A_699_463#_c_815_n 0.00331109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_699_463#_c_825_n 0.00205239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_699_463#_c_826_n 2.03292e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_306_119#_M1027_g 0.0213503f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_167 VPB N_A_306_119#_c_941_n 0.0730305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_306_119#_c_942_n 0.0552875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_306_119#_c_943_n 0.0106267f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_170 VPB N_A_306_119#_c_932_n 0.0143213f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_171 VPB N_A_306_119#_M1006_g 0.0377293f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.165
cc_172 VPB N_A_306_119#_c_946_n 0.188016f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.295
cc_173 VPB N_A_306_119#_M1007_g 0.0292916f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_174 VPB N_A_306_119#_c_934_n 0.0388192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_306_119#_c_949_n 0.00838544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_306_119#_c_950_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_306_119#_c_937_n 0.00550685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_306_119#_c_938_n 0.00111317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_306_119#_c_953_n 0.00486835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1525_212#_c_1117_n 0.00452844f $X=-0.19 $Y=1.66 $X2=0.155
+ $Y2=1.95
cc_181 VPB N_A_1525_212#_M1018_g 0.0321887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1525_212#_c_1109_n 0.0172903f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_183 VPB N_A_1525_212#_c_1120_n 0.0122081f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_184 VPB N_A_1525_212#_c_1121_n 0.00194708f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.665
cc_185 VPB N_A_1525_212#_c_1122_n 0.00467452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1525_212#_c_1123_n 0.00234171f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.845
cc_187 VPB N_A_1525_212#_c_1113_n 0.0058695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1271_74#_M1002_g 0.0492393f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_189 VPB N_A_1271_74#_c_1223_n 0.00814854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1271_74#_c_1224_n 0.0260612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1271_74#_M1010_g 0.0351319f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_192 VPB N_A_1271_74#_c_1226_n 0.00430295f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.165
cc_193 VPB N_A_1271_74#_c_1237_n 0.00135254f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_194 VPB N_A_1271_74#_c_1238_n 0.0126592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1271_74#_c_1229_n 0.0140489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1271_74#_c_1230_n 4.13852e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1271_74#_c_1231_n 4.64263e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1271_74#_c_1242_n 0.00154868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1924_409#_M1029_g 0.0252871f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_200 VPB N_A_1924_409#_M1030_g 0.0274144f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_201 VPB N_A_1924_409#_c_1376_n 0.0113539f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_202 VPB N_A_1924_409#_c_1371_n 0.00700295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1430_n 0.0109398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1431_n 0.0291509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1432_n 0.00655428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1433_n 0.00129922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1434_n 0.0133892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1435_n 0.0221866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1436_n 0.0244305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1437_n 0.0149609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1438_n 0.0163609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1439_n 0.0228504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1440_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1441_n 0.0638732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1442_n 0.0275707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1443_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1444_n 0.0140508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1445_n 0.017333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1446_n 0.056342f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1447_n 0.0531608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1448_n 0.0209549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1449_n 0.0186759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1450_n 0.0053864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1451_n 0.00485379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1452_n 0.00437061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1453_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1454_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1455_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1429_n 0.108605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_30_78#_c_1587_n 0.00131068f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_231 VPB N_A_30_78#_c_1582_n 0.00818028f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_232 VPB N_A_30_78#_c_1589_n 3.98049e-19 $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_233 VPB N_A_30_78#_c_1590_n 0.0055014f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_234 VPB N_A_30_78#_c_1591_n 0.00145207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_30_78#_c_1584_n 0.00577037f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_236 VPB N_A_30_78#_c_1593_n 0.00279651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_30_78#_c_1594_n 0.0163782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_30_78#_c_1595_n 0.00151936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB Q 0.00231613f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_240 N_D_M1028_g N_RESET_B_M1012_g 0.0245996f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_241 N_D_c_245_n N_RESET_B_M1012_g 9.43739e-19 $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_242 N_D_c_242_n N_RESET_B_c_601_n 0.0245996f $X=0.402 $Y=1.828 $X2=0 $Y2=0
cc_243 N_D_M1014_g N_RESET_B_M1015_g 0.0269045f $X=0.495 $Y=2.845 $X2=0 $Y2=0
cc_244 N_D_c_244_n N_RESET_B_c_608_n 0.0245996f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_245 N_D_c_249_n N_RESET_B_c_623_n 0.0245996f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_246 N_D_M1014_g N_VPWR_c_1431_n 0.01511f $X=0.495 $Y=2.845 $X2=0 $Y2=0
cc_247 N_D_c_245_n N_VPWR_c_1431_n 0.0171637f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_248 N_D_c_249_n N_VPWR_c_1431_n 9.92489e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_249 N_D_M1014_g N_VPWR_c_1432_n 4.81981e-19 $X=0.495 $Y=2.845 $X2=0 $Y2=0
cc_250 N_D_M1014_g N_VPWR_c_1444_n 0.00543892f $X=0.495 $Y=2.845 $X2=0 $Y2=0
cc_251 N_D_M1014_g N_VPWR_c_1429_n 0.0097046f $X=0.495 $Y=2.845 $X2=0 $Y2=0
cc_252 N_D_M1028_g N_A_30_78#_c_1581_n 0.0114706f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_253 N_D_c_245_n N_A_30_78#_c_1581_n 0.00258996f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_254 N_D_M1028_g N_A_30_78#_c_1582_n 0.018142f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_255 N_D_c_245_n N_A_30_78#_c_1582_n 0.088088f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_256 N_D_M1028_g N_A_30_78#_c_1585_n 0.00806237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_257 N_D_c_244_n N_A_30_78#_c_1585_n 0.00161806f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_258 N_D_c_245_n N_A_30_78#_c_1585_n 0.0286676f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_259 N_D_M1014_g N_A_30_78#_c_1593_n 0.00323147f $X=0.495 $Y=2.845 $X2=0 $Y2=0
cc_260 N_D_M1028_g N_VGND_c_1723_n 0.00190636f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_261 N_D_M1028_g N_VGND_c_1730_n 0.00429844f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_262 N_D_M1028_g N_VGND_c_1742_n 0.00539454f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_263 N_CLK_M1025_g N_RESET_B_c_601_n 0.00478461f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_264 N_CLK_c_274_n N_RESET_B_c_601_n 0.00647442f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_265 N_CLK_c_275_n N_RESET_B_c_602_n 0.0102966f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_266 N_CLK_M1025_g N_RESET_B_c_616_n 0.00414582f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_267 CLK N_RESET_B_c_616_n 0.0132561f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_268 N_CLK_c_275_n N_RESET_B_c_608_n 0.00394493f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_269 N_CLK_M1025_g N_A_306_119#_M1027_g 0.0514847f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_270 CLK N_A_306_119#_c_930_n 7.58266e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_271 N_CLK_c_275_n N_A_306_119#_c_930_n 0.0230956f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_272 CLK N_A_306_119#_c_932_n 0.00372412f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_273 N_CLK_c_274_n N_A_306_119#_c_932_n 0.0214524f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_274 N_CLK_c_275_n N_A_306_119#_c_932_n 0.00127928f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_275 N_CLK_c_275_n N_A_306_119#_c_936_n 0.00709082f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_276 N_CLK_M1025_g N_A_306_119#_c_937_n 0.00367655f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_277 CLK N_A_306_119#_c_937_n 0.0353887f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_278 N_CLK_c_274_n N_A_306_119#_c_937_n 0.0030261f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_279 N_CLK_c_275_n N_A_306_119#_c_937_n 0.00365637f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_280 CLK N_A_306_119#_c_965_n 0.0291181f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_281 N_CLK_c_274_n N_A_306_119#_c_965_n 4.6511e-19 $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_282 N_CLK_c_275_n N_A_306_119#_c_965_n 0.0115022f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_283 CLK N_A_306_119#_c_938_n 0.0322106f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_284 N_CLK_c_274_n N_A_306_119#_c_938_n 2.23058e-19 $X=1.91 $Y=1.61 $X2=0
+ $Y2=0
cc_285 N_CLK_c_275_n N_A_306_119#_c_938_n 9.57688e-19 $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_286 CLK N_A_306_119#_c_939_n 0.00199038f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_287 N_CLK_c_274_n N_A_306_119#_c_939_n 0.00114873f $X=1.91 $Y=1.61 $X2=0
+ $Y2=0
cc_288 N_CLK_c_275_n N_A_306_119#_c_939_n 7.14557e-19 $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_289 N_CLK_M1025_g N_A_306_119#_c_953_n 0.00685407f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_290 CLK N_A_306_119#_c_953_n 0.00336717f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_291 N_CLK_c_274_n N_A_306_119#_c_953_n 0.00167789f $X=1.91 $Y=1.61 $X2=0
+ $Y2=0
cc_292 N_CLK_M1025_g N_VPWR_c_1432_n 0.00598165f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_293 N_CLK_M1025_g N_VPWR_c_1433_n 0.0106716f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_294 N_CLK_M1025_g N_VPWR_c_1445_n 0.00401239f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_295 N_CLK_M1025_g N_VPWR_c_1429_n 0.00589267f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_296 N_CLK_M1025_g N_A_30_78#_c_1594_n 0.0178578f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_297 CLK N_A_30_78#_c_1594_n 0.00371797f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_298 CLK N_VGND_M1016_d 0.00290034f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_299 N_CLK_c_275_n N_VGND_c_1723_n 0.00274302f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_300 N_CLK_c_275_n N_VGND_c_1724_n 0.00440713f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_301 N_CLK_c_275_n N_VGND_c_1742_n 9.39239e-19 $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_302 N_A_493_387#_c_328_n N_A_837_359#_M1023_d 0.00224297f $X=7.285 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_303 N_A_493_387#_M1004_g N_A_837_359#_M1011_g 0.00211742f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_304 N_A_493_387#_c_318_n N_A_837_359#_M1008_g 0.00674849f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_305 N_A_493_387#_M1024_g N_A_837_359#_M1008_g 0.0529896f $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_306 N_A_493_387#_c_327_n N_A_837_359#_M1008_g 0.00369436f $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_307 N_A_493_387#_c_333_n N_A_837_359#_M1008_g 0.00720138f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_308 N_A_493_387#_c_318_n N_A_837_359#_c_516_n 4.94823e-19 $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_309 N_A_493_387#_M1024_g N_A_837_359#_c_516_n 0.00126199f $X=4.01 $Y=0.9
+ $X2=0 $Y2=0
cc_310 N_A_493_387#_c_336_n N_A_837_359#_c_523_n 0.00211742f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_311 N_A_493_387#_c_327_n N_A_837_359#_c_517_n 0.0769509f $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_312 N_A_493_387#_c_328_n N_A_837_359#_c_517_n 0.00332639f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_313 N_A_493_387#_c_327_n N_A_837_359#_c_537_n 3.80876e-19 $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_314 N_A_493_387#_c_333_n N_A_837_359#_c_537_n 0.00936402f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_315 N_A_493_387#_c_328_n N_A_837_359#_c_539_n 0.0176299f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_316 N_A_493_387#_c_322_n N_A_837_359#_c_524_n 0.00303542f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_317 N_A_493_387#_c_320_n N_A_837_359#_c_518_n 4.62933e-19 $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_318 N_A_493_387#_c_320_n N_A_837_359#_c_519_n 0.00207614f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_319 N_A_493_387#_M1024_g N_RESET_B_c_602_n 0.00526413f $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_320 N_A_493_387#_c_324_n N_RESET_B_c_602_n 0.0232924f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_321 N_A_493_387#_c_327_n N_RESET_B_c_602_n 0.00282315f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_322 N_A_493_387#_c_332_n N_RESET_B_c_602_n 0.0120895f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_323 N_A_493_387#_c_333_n N_RESET_B_c_602_n 0.00229078f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_324 N_A_493_387#_c_327_n N_RESET_B_M1001_g 0.013523f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_325 N_A_493_387#_c_368_p N_RESET_B_M1001_g 0.00355258f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_326 N_A_493_387#_c_333_n N_RESET_B_M1001_g 0.00620923f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_327 N_A_493_387#_M1027_d N_RESET_B_c_616_n 9.76131e-19 $X=2.465 $Y=1.935
+ $X2=0 $Y2=0
cc_328 N_A_493_387#_c_336_n N_RESET_B_c_616_n 0.00392642f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_329 N_A_493_387#_M1004_g N_RESET_B_c_616_n 0.00651345f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_330 N_A_493_387#_c_338_n N_RESET_B_c_616_n 0.00433669f $X=3.825 $Y=1.68 $X2=0
+ $Y2=0
cc_331 N_A_493_387#_c_325_n N_RESET_B_c_616_n 0.0398351f $X=3.08 $Y=1.77 $X2=0
+ $Y2=0
cc_332 N_A_493_387#_c_326_n N_RESET_B_c_616_n 0.010529f $X=3.33 $Y=1.77 $X2=0
+ $Y2=0
cc_333 N_A_493_387#_c_330_n N_RESET_B_c_618_n 0.0218177f $X=7.12 $Y=2.14 $X2=0
+ $Y2=0
cc_334 N_A_493_387#_c_344_n N_RESET_B_c_618_n 0.00330668f $X=7.315 $Y=2.14 $X2=0
+ $Y2=0
cc_335 N_A_493_387#_c_320_n N_A_699_463#_M1023_g 0.0126968f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_336 N_A_493_387#_c_328_n N_A_699_463#_M1023_g 0.0119914f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_337 N_A_493_387#_c_322_n N_A_699_463#_c_812_n 0.0126968f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_338 N_A_493_387#_M1004_g N_A_699_463#_c_813_n 6.55964e-19 $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_339 N_A_493_387#_c_318_n N_A_699_463#_c_813_n 0.0123218f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_340 N_A_493_387#_M1024_g N_A_699_463#_c_813_n 0.00839185f $X=4.01 $Y=0.9
+ $X2=0 $Y2=0
cc_341 N_A_493_387#_M1004_g N_A_699_463#_c_822_n 0.00430041f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_342 N_A_493_387#_c_338_n N_A_699_463#_c_822_n 0.00108491f $X=3.825 $Y=1.68
+ $X2=0 $Y2=0
cc_343 N_A_493_387#_c_338_n N_A_699_463#_c_816_n 0.0016773f $X=3.825 $Y=1.68
+ $X2=0 $Y2=0
cc_344 N_A_493_387#_c_318_n N_A_699_463#_c_816_n 0.00274419f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_345 N_A_493_387#_M1024_g N_A_699_463#_c_816_n 0.0082711f $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_346 N_A_493_387#_c_324_n N_A_699_463#_c_816_n 0.0353714f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_347 N_A_493_387#_c_333_n N_A_699_463#_c_816_n 0.00147443f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_348 N_A_493_387#_c_325_n N_A_306_119#_M1027_g 9.04289e-19 $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_349 N_A_493_387#_c_323_n N_A_306_119#_c_930_n 0.00452109f $X=2.955 $Y=1.605
+ $X2=0 $Y2=0
cc_350 N_A_493_387#_c_332_n N_A_306_119#_c_930_n 0.00693446f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_351 N_A_493_387#_M1004_g N_A_306_119#_c_941_n 0.0237271f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_352 N_A_493_387#_c_325_n N_A_306_119#_c_941_n 0.0219056f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_353 N_A_493_387#_M1004_g N_A_306_119#_c_942_n 0.0122286f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_354 N_A_493_387#_c_336_n N_A_306_119#_c_931_n 0.0224379f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_355 N_A_493_387#_c_324_n N_A_306_119#_c_931_n 0.00408646f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_356 N_A_493_387#_c_325_n N_A_306_119#_c_931_n 0.00142045f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_357 N_A_493_387#_c_326_n N_A_306_119#_c_931_n 0.00381035f $X=3.33 $Y=1.77
+ $X2=0 $Y2=0
cc_358 N_A_493_387#_c_336_n N_A_306_119#_c_932_n 0.0212577f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_359 N_A_493_387#_c_323_n N_A_306_119#_c_932_n 0.0213221f $X=2.955 $Y=1.605
+ $X2=0 $Y2=0
cc_360 N_A_493_387#_c_325_n N_A_306_119#_c_932_n 0.0070493f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_361 N_A_493_387#_c_332_n N_A_306_119#_c_932_n 0.0055573f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_362 N_A_493_387#_M1024_g N_A_306_119#_c_933_n 0.0194425f $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_363 N_A_493_387#_c_324_n N_A_306_119#_c_933_n 0.00349197f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_364 N_A_493_387#_c_332_n N_A_306_119#_c_933_n 0.00456341f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_365 N_A_493_387#_M1004_g N_A_306_119#_M1006_g 0.0167963f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_366 N_A_493_387#_c_338_n N_A_306_119#_M1006_g 0.00609737f $X=3.825 $Y=1.68
+ $X2=0 $Y2=0
cc_367 N_A_493_387#_c_344_n N_A_306_119#_M1007_g 0.00768262f $X=7.315 $Y=2.14
+ $X2=0 $Y2=0
cc_368 N_A_493_387#_c_321_n N_A_306_119#_c_934_n 0.0197541f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_369 N_A_493_387#_c_330_n N_A_306_119#_c_934_n 0.0166975f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_370 N_A_493_387#_c_335_n N_A_306_119#_c_934_n 0.00239794f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_371 N_A_493_387#_c_344_n N_A_306_119#_c_934_n 0.0260258f $X=7.315 $Y=2.14
+ $X2=0 $Y2=0
cc_372 N_A_493_387#_c_322_n N_A_306_119#_c_949_n 0.0197541f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_373 N_A_493_387#_c_328_n N_A_306_119#_M1032_g 0.00912173f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_374 N_A_493_387#_c_330_n N_A_306_119#_M1032_g 0.00885461f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_375 N_A_493_387#_c_331_n N_A_306_119#_M1032_g 0.0230685f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_376 N_A_493_387#_c_334_n N_A_306_119#_M1032_g 0.0213806f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_377 N_A_493_387#_c_335_n N_A_306_119#_M1032_g 0.0123873f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_378 N_A_493_387#_M1013_d N_A_306_119#_c_965_n 0.00308104f $X=2.535 $Y=0.595
+ $X2=0 $Y2=0
cc_379 N_A_493_387#_c_323_n N_A_306_119#_c_965_n 0.0140566f $X=2.955 $Y=1.605
+ $X2=0 $Y2=0
cc_380 N_A_493_387#_c_332_n N_A_306_119#_c_965_n 0.0114269f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_381 N_A_493_387#_M1013_d N_A_306_119#_c_938_n 0.00162539f $X=2.535 $Y=0.595
+ $X2=0 $Y2=0
cc_382 N_A_493_387#_c_323_n N_A_306_119#_c_938_n 0.03259f $X=2.955 $Y=1.605
+ $X2=0 $Y2=0
cc_383 N_A_493_387#_c_325_n N_A_306_119#_c_938_n 0.0265116f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_384 N_A_493_387#_c_325_n N_A_306_119#_c_953_n 0.00357673f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_385 N_A_493_387#_c_328_n N_A_1525_212#_M1005_g 0.00108131f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_386 N_A_493_387#_c_331_n N_A_1525_212#_M1005_g 0.00485618f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_387 N_A_493_387#_c_335_n N_A_1525_212#_M1005_g 0.00116217f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_388 N_A_493_387#_c_344_n N_A_1525_212#_c_1117_n 0.0264655f $X=7.315 $Y=2.14
+ $X2=0 $Y2=0
cc_389 N_A_493_387#_M1009_g N_A_1525_212#_M1018_g 0.0264655f $X=7.315 $Y=2.675
+ $X2=0 $Y2=0
cc_390 N_A_493_387#_c_330_n N_A_1525_212#_c_1109_n 9.8351e-19 $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_391 N_A_493_387#_c_330_n N_A_1525_212#_c_1114_n 0.00193736f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_392 N_A_493_387#_c_335_n N_A_1525_212#_c_1114_n 0.0239506f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_393 N_A_493_387#_c_335_n N_A_1525_212#_c_1115_n 0.00177987f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_394 N_A_493_387#_c_328_n N_A_1271_74#_M1003_d 0.00941894f $X=7.285 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_395 N_A_493_387#_c_328_n N_A_1271_74#_c_1244_n 0.00860077f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_396 N_A_493_387#_c_320_n N_A_1271_74#_c_1227_n 0.0041612f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_397 N_A_493_387#_c_321_n N_A_1271_74#_c_1227_n 0.010955f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_398 N_A_493_387#_c_330_n N_A_1271_74#_c_1227_n 0.00709969f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_399 N_A_493_387#_c_334_n N_A_1271_74#_c_1227_n 0.00131723f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_400 N_A_493_387#_c_335_n N_A_1271_74#_c_1227_n 0.022475f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_401 N_A_493_387#_M1009_g N_A_1271_74#_c_1237_n 0.0038942f $X=7.315 $Y=2.675
+ $X2=0 $Y2=0
cc_402 N_A_493_387#_c_330_n N_A_1271_74#_c_1237_n 0.0315384f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_403 N_A_493_387#_c_344_n N_A_1271_74#_c_1237_n 0.00236717f $X=7.315 $Y=2.14
+ $X2=0 $Y2=0
cc_404 N_A_493_387#_c_321_n N_A_1271_74#_c_1228_n 0.00400734f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_405 N_A_493_387#_c_328_n N_A_1271_74#_c_1228_n 0.0414158f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_406 N_A_493_387#_c_331_n N_A_1271_74#_c_1228_n 0.0196081f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_407 N_A_493_387#_c_334_n N_A_1271_74#_c_1228_n 0.00763158f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_408 N_A_493_387#_c_335_n N_A_1271_74#_c_1228_n 0.0304853f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_409 N_A_493_387#_M1009_g N_A_1271_74#_c_1258_n 0.014245f $X=7.315 $Y=2.675
+ $X2=0 $Y2=0
cc_410 N_A_493_387#_c_330_n N_A_1271_74#_c_1258_n 0.0233706f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_411 N_A_493_387#_c_344_n N_A_1271_74#_c_1258_n 0.00184821f $X=7.315 $Y=2.14
+ $X2=0 $Y2=0
cc_412 N_A_493_387#_c_330_n N_A_1271_74#_c_1238_n 0.0428804f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_413 N_A_493_387#_c_344_n N_A_1271_74#_c_1238_n 0.00609795f $X=7.315 $Y=2.14
+ $X2=0 $Y2=0
cc_414 N_A_493_387#_c_330_n N_A_1271_74#_c_1230_n 0.0142968f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_415 N_A_493_387#_c_321_n N_A_1271_74#_c_1231_n 0.00176995f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_416 N_A_493_387#_c_330_n N_A_1271_74#_c_1231_n 0.00932939f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_417 N_A_493_387#_M1009_g N_VPWR_c_1437_n 0.0012526f $X=7.315 $Y=2.675 $X2=0
+ $Y2=0
cc_418 N_A_493_387#_M1009_g N_VPWR_c_1447_n 0.00469675f $X=7.315 $Y=2.675 $X2=0
+ $Y2=0
cc_419 N_A_493_387#_M1004_g N_VPWR_c_1429_n 0.00112709f $X=3.405 $Y=2.525 $X2=0
+ $Y2=0
cc_420 N_A_493_387#_M1009_g N_VPWR_c_1429_n 0.00626544f $X=7.315 $Y=2.675 $X2=0
+ $Y2=0
cc_421 N_A_493_387#_M1004_g N_A_30_78#_c_1589_n 0.00440524f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_422 N_A_493_387#_M1024_g N_A_30_78#_c_1583_n 2.83252e-19 $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_423 N_A_493_387#_c_324_n N_A_30_78#_c_1583_n 0.0195044f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_424 N_A_493_387#_c_332_n N_A_30_78#_c_1583_n 0.0437866f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_425 N_A_493_387#_M1004_g N_A_30_78#_c_1590_n 0.0104428f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_426 N_A_493_387#_c_338_n N_A_30_78#_c_1590_n 0.00265751f $X=3.825 $Y=1.68
+ $X2=0 $Y2=0
cc_427 N_A_493_387#_c_326_n N_A_30_78#_c_1590_n 0.0024633f $X=3.33 $Y=1.77 $X2=0
+ $Y2=0
cc_428 N_A_493_387#_c_336_n N_A_30_78#_c_1591_n 0.00243404f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_429 N_A_493_387#_M1004_g N_A_30_78#_c_1591_n 0.0027797f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_430 N_A_493_387#_c_325_n N_A_30_78#_c_1591_n 0.015371f $X=3.08 $Y=1.77 $X2=0
+ $Y2=0
cc_431 N_A_493_387#_c_326_n N_A_30_78#_c_1591_n 0.0109437f $X=3.33 $Y=1.77 $X2=0
+ $Y2=0
cc_432 N_A_493_387#_c_336_n N_A_30_78#_c_1584_n 0.00493197f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_433 N_A_493_387#_c_338_n N_A_30_78#_c_1584_n 0.0132261f $X=3.825 $Y=1.68
+ $X2=0 $Y2=0
cc_434 N_A_493_387#_c_318_n N_A_30_78#_c_1584_n 0.00471312f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_435 N_A_493_387#_c_323_n N_A_30_78#_c_1584_n 0.00648483f $X=2.955 $Y=1.605
+ $X2=0 $Y2=0
cc_436 N_A_493_387#_c_325_n N_A_30_78#_c_1584_n 0.00397431f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_437 N_A_493_387#_c_326_n N_A_30_78#_c_1584_n 0.0252428f $X=3.33 $Y=1.77 $X2=0
+ $Y2=0
cc_438 N_A_493_387#_M1027_d N_A_30_78#_c_1594_n 0.00590913f $X=2.465 $Y=1.935
+ $X2=0 $Y2=0
cc_439 N_A_493_387#_c_325_n N_A_30_78#_c_1594_n 0.0378185f $X=3.08 $Y=1.77 $X2=0
+ $Y2=0
cc_440 N_A_493_387#_c_336_n N_A_30_78#_c_1595_n 7.07705e-19 $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_441 N_A_493_387#_M1004_g N_A_30_78#_c_1595_n 0.00472425f $X=3.405 $Y=2.525
+ $X2=0 $Y2=0
cc_442 N_A_493_387#_c_325_n N_A_30_78#_c_1595_n 0.00110215f $X=3.08 $Y=1.77
+ $X2=0 $Y2=0
cc_443 N_A_493_387#_c_326_n N_A_30_78#_c_1595_n 0.00200148f $X=3.33 $Y=1.77
+ $X2=0 $Y2=0
cc_444 N_A_493_387#_c_336_n N_A_30_78#_c_1586_n 0.00476721f $X=3.405 $Y=1.935
+ $X2=0 $Y2=0
cc_445 N_A_493_387#_c_338_n N_A_30_78#_c_1586_n 7.59196e-19 $X=3.825 $Y=1.68
+ $X2=0 $Y2=0
cc_446 N_A_493_387#_M1024_g N_A_30_78#_c_1586_n 8.19151e-19 $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_447 N_A_493_387#_c_323_n N_A_30_78#_c_1586_n 0.0127435f $X=2.955 $Y=1.605
+ $X2=0 $Y2=0
cc_448 N_A_493_387#_c_326_n N_A_30_78#_c_1586_n 0.0133562f $X=3.33 $Y=1.77 $X2=0
+ $Y2=0
cc_449 N_A_493_387#_c_327_n N_VGND_M1001_d 0.0203479f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_450 N_A_493_387#_c_368_p N_VGND_M1001_d 0.00355743f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_451 N_A_493_387#_c_329_n N_VGND_M1001_d 6.7108e-19 $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_452 N_A_493_387#_c_332_n N_VGND_c_1724_n 0.0309435f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_453 N_A_493_387#_c_328_n N_VGND_c_1725_n 0.00865667f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_454 N_A_493_387#_c_324_n N_VGND_c_1733_n 0.0538549f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_455 N_A_493_387#_c_327_n N_VGND_c_1733_n 0.0408719f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_456 N_A_493_387#_c_368_p N_VGND_c_1733_n 0.00152296f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_457 N_A_493_387#_c_329_n N_VGND_c_1733_n 0.0151294f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_458 N_A_493_387#_c_332_n N_VGND_c_1733_n 0.025157f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_459 N_A_493_387#_c_333_n N_VGND_c_1733_n 0.0124175f $X=4.355 $Y=0.415 $X2=0
+ $Y2=0
cc_460 N_A_493_387#_c_320_n N_VGND_c_1734_n 0.00278271f $X=6.28 $Y=1.195 $X2=0
+ $Y2=0
cc_461 N_A_493_387#_c_327_n N_VGND_c_1734_n 0.00309688f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_462 N_A_493_387#_c_328_n N_VGND_c_1734_n 0.114324f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_463 N_A_493_387#_c_329_n N_VGND_c_1734_n 0.0119604f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_464 N_A_493_387#_c_320_n N_VGND_c_1742_n 0.00358928f $X=6.28 $Y=1.195 $X2=0
+ $Y2=0
cc_465 N_A_493_387#_c_324_n N_VGND_c_1742_n 0.0391622f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_466 N_A_493_387#_c_327_n N_VGND_c_1742_n 0.0190163f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_467 N_A_493_387#_c_328_n N_VGND_c_1742_n 0.0653925f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_468 N_A_493_387#_c_329_n N_VGND_c_1742_n 0.00656672f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_469 N_A_493_387#_c_332_n N_VGND_c_1742_n 0.0174682f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_470 N_A_493_387#_c_333_n N_VGND_c_1742_n 0.00552563f $X=4.355 $Y=0.415 $X2=0
+ $Y2=0
cc_471 N_A_493_387#_c_327_n A_895_138# 0.00134267f $X=5.515 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_472 N_A_837_359#_M1008_g N_RESET_B_c_602_n 0.00559335f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_473 N_A_837_359#_M1008_g N_RESET_B_M1001_g 0.0419644f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_474 N_A_837_359#_c_516_n N_RESET_B_M1001_g 0.00106151f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_475 N_A_837_359#_c_517_n N_RESET_B_M1001_g 0.0122236f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_476 N_A_837_359#_M1008_g N_RESET_B_c_605_n 0.0138048f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_477 N_A_837_359#_c_516_n N_RESET_B_c_605_n 4.52393e-19 $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_478 N_A_837_359#_M1011_g N_RESET_B_M1017_g 0.0167346f $X=4.275 $Y=2.525 $X2=0
+ $Y2=0
cc_479 N_A_837_359#_c_517_n N_RESET_B_c_607_n 0.00269956f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_480 N_A_837_359#_c_516_n N_RESET_B_c_616_n 0.0164056f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_481 N_A_837_359#_c_523_n N_RESET_B_c_616_n 0.0101395f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_482 N_A_837_359#_M1000_d N_RESET_B_c_618_n 0.00136926f $X=5.995 $Y=1.735
+ $X2=0 $Y2=0
cc_483 N_A_837_359#_c_524_n N_RESET_B_c_618_n 0.0386667f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_484 N_A_837_359#_c_523_n N_RESET_B_c_624_n 0.0149913f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_485 N_A_837_359#_c_517_n N_A_699_463#_M1023_g 0.0125065f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_486 N_A_837_359#_c_539_n N_A_699_463#_M1023_g 0.0104935f $X=6.02 $Y=0.86
+ $X2=0 $Y2=0
cc_487 N_A_837_359#_c_518_n N_A_699_463#_M1023_g 0.00268294f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_488 N_A_837_359#_c_519_n N_A_699_463#_M1023_g 0.00639735f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_489 N_A_837_359#_c_524_n N_A_699_463#_M1000_g 0.00552021f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_490 N_A_837_359#_c_517_n N_A_699_463#_c_811_n 0.0091182f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_491 N_A_837_359#_c_518_n N_A_699_463#_c_812_n 0.00470883f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_492 N_A_837_359#_c_519_n N_A_699_463#_c_812_n 0.00552021f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_493 N_A_837_359#_M1008_g N_A_699_463#_c_813_n 0.00204111f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_494 N_A_837_359#_c_516_n N_A_699_463#_c_813_n 0.0736089f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_495 N_A_837_359#_c_523_n N_A_699_463#_c_813_n 0.00568157f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_496 N_A_837_359#_c_537_n N_A_699_463#_c_813_n 0.00118204f $X=4.445 $Y=1.04
+ $X2=0 $Y2=0
cc_497 N_A_837_359#_M1011_g N_A_699_463#_c_821_n 0.00882618f $X=4.275 $Y=2.525
+ $X2=0 $Y2=0
cc_498 N_A_837_359#_c_516_n N_A_699_463#_c_821_n 0.0126011f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_499 N_A_837_359#_c_523_n N_A_699_463#_c_821_n 0.00382824f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_500 N_A_837_359#_M1011_g N_A_699_463#_c_822_n 0.0155802f $X=4.275 $Y=2.525
+ $X2=0 $Y2=0
cc_501 N_A_837_359#_M1011_g N_A_699_463#_c_823_n 0.00159495f $X=4.275 $Y=2.525
+ $X2=0 $Y2=0
cc_502 N_A_837_359#_M1008_g N_A_699_463#_c_823_n 0.00140716f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_503 N_A_837_359#_c_516_n N_A_699_463#_c_823_n 0.0386079f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_504 N_A_837_359#_c_523_n N_A_699_463#_c_823_n 0.00219738f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_505 N_A_837_359#_M1008_g N_A_699_463#_c_814_n 0.00201464f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_506 N_A_837_359#_c_516_n N_A_699_463#_c_814_n 0.0226331f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_507 N_A_837_359#_c_517_n N_A_699_463#_c_814_n 0.0137783f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_508 N_A_837_359#_c_517_n N_A_699_463#_c_815_n 0.0680785f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_509 N_A_837_359#_c_519_n N_A_699_463#_c_815_n 0.0134746f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_510 N_A_837_359#_M1011_g N_A_306_119#_M1006_g 0.0381302f $X=4.275 $Y=2.525
+ $X2=0 $Y2=0
cc_511 N_A_837_359#_M1011_g N_A_306_119#_c_946_n 0.0118063f $X=4.275 $Y=2.525
+ $X2=0 $Y2=0
cc_512 N_A_837_359#_c_524_n N_A_306_119#_c_946_n 0.00434706f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_513 N_A_837_359#_c_524_n N_A_306_119#_M1007_g 0.012708f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_514 N_A_837_359#_c_519_n N_A_306_119#_c_949_n 0.00222494f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_515 N_A_837_359#_c_518_n N_A_1271_74#_c_1227_n 0.00157956f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_516 N_A_837_359#_c_519_n N_A_1271_74#_c_1227_n 0.0283811f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_517 N_A_837_359#_c_524_n N_A_1271_74#_c_1237_n 0.0250147f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_518 N_A_837_359#_c_519_n N_A_1271_74#_c_1237_n 0.00658861f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_519 N_A_837_359#_c_519_n N_A_1271_74#_c_1231_n 0.0129728f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_520 N_A_837_359#_M1011_g N_VPWR_c_1434_n 0.00160965f $X=4.275 $Y=2.525 $X2=0
+ $Y2=0
cc_521 N_A_837_359#_c_517_n N_VPWR_c_1436_n 0.00363319f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_522 N_A_837_359#_c_524_n N_VPWR_c_1436_n 0.0405057f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_523 N_A_837_359#_c_524_n N_VPWR_c_1447_n 0.00664291f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_524 N_A_837_359#_M1011_g N_VPWR_c_1429_n 0.00112709f $X=4.275 $Y=2.525 $X2=0
+ $Y2=0
cc_525 N_A_837_359#_c_524_n N_VPWR_c_1429_n 0.00903857f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_526 N_A_837_359#_c_517_n N_VGND_M1001_d 0.0123032f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_527 N_A_837_359#_M1008_g N_VGND_c_1742_n 2.31769e-19 $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_528 N_A_837_359#_c_517_n A_895_138# 0.00134267f $X=5.855 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_529 N_RESET_B_c_618_n N_A_699_463#_M1000_g 0.0119125f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_530 N_RESET_B_c_607_n N_A_699_463#_c_811_n 0.00991362f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_618_n N_A_699_463#_c_811_n 0.00341453f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_616_n N_A_699_463#_c_813_n 0.0190003f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_533 N_RESET_B_c_616_n N_A_699_463#_c_821_n 0.00957379f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_534 N_RESET_B_M1017_g N_A_699_463#_c_822_n 8.24351e-19 $X=4.895 $Y=2.525
+ $X2=0 $Y2=0
cc_535 N_RESET_B_c_616_n N_A_699_463#_c_822_n 0.0145179f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_RESET_B_c_605_n N_A_699_463#_c_823_n 0.0125326f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_616_n N_A_699_463#_c_823_n 0.0170764f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_RESET_B_c_619_n N_A_699_463#_c_823_n 0.00239892f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_620_n N_A_699_463#_c_823_n 0.0245211f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_RESET_B_c_607_n N_A_699_463#_c_814_n 0.00324317f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_605_n N_A_699_463#_c_815_n 0.0123388f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_607_n N_A_699_463#_c_815_n 0.0034188f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_616_n N_A_699_463#_c_815_n 0.00355574f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_544 N_RESET_B_c_618_n N_A_699_463#_c_815_n 0.0096202f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_545 N_RESET_B_c_619_n N_A_699_463#_c_815_n 0.00343479f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_620_n N_A_699_463#_c_815_n 0.019281f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_624_n N_A_699_463#_c_815_n 0.00736996f $X=5.12 $Y=1.96 $X2=0
+ $Y2=0
cc_548 N_RESET_B_M1017_g N_A_699_463#_c_825_n 0.0113125f $X=4.895 $Y=2.525 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_616_n N_A_699_463#_c_825_n 0.00415846f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_550 N_RESET_B_c_618_n N_A_699_463#_c_825_n 6.95302e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_551 N_RESET_B_c_619_n N_A_699_463#_c_825_n 0.00866835f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_620_n N_A_699_463#_c_825_n 0.0206751f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_624_n N_A_699_463#_c_825_n 0.00187572f $X=5.12 $Y=1.96 $X2=0
+ $Y2=0
cc_554 N_RESET_B_M1017_g N_A_699_463#_c_826_n 7.14937e-19 $X=4.895 $Y=2.525
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_616_n N_A_306_119#_M1027_g 0.0100828f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_602_n N_A_306_119#_c_930_n 0.0101603f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_602_n N_A_306_119#_c_933_n 0.00526413f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_616_n N_A_306_119#_M1006_g 0.00279709f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_RESET_B_M1017_g N_A_306_119#_c_946_n 0.0120141f $X=4.895 $Y=2.525 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_618_n N_A_306_119#_M1007_g 0.00927441f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_618_n N_A_306_119#_c_934_n 0.00740552f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_562 N_RESET_B_M1012_g N_A_306_119#_c_936_n 0.00294809f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_602_n N_A_306_119#_c_936_n 0.0073964f $X=4.715 $Y=0.18 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_616_n N_A_306_119#_c_937_n 0.00308596f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_565 N_RESET_B_c_617_n N_A_306_119#_c_937_n 7.65024e-19 $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_566 N_RESET_B_c_608_n N_A_306_119#_c_937_n 0.00735309f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_609_n N_A_306_119#_c_937_n 0.0586003f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_616_n N_A_306_119#_c_938_n 0.00386848f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_569 N_RESET_B_M1012_g N_A_306_119#_c_939_n 0.00123734f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_570 N_RESET_B_c_609_n N_A_306_119#_c_939_n 8.33963e-19 $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_571 N_RESET_B_M1015_g N_A_306_119#_c_953_n 0.00232337f $X=0.945 $Y=2.845
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_616_n N_A_306_119#_c_953_n 0.0252561f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_617_n N_A_306_119#_c_953_n 0.00199927f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_609_n N_A_306_119#_c_953_n 0.0139899f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_623_n N_A_306_119#_c_953_n 0.00154955f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_RESET_B_M1021_g N_A_1525_212#_M1005_g 0.0164487f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_618_n N_A_1525_212#_c_1117_n 4.99514e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_625_n N_A_1525_212#_c_1117_n 0.0164306f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_626_n N_A_1525_212#_c_1117_n 0.00182389f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_580 N_RESET_B_M1019_g N_A_1525_212#_M1018_g 0.0131127f $X=8.235 $Y=2.675
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_618_n N_A_1525_212#_M1018_g 0.00551679f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_RESET_B_c_621_n N_A_1525_212#_M1018_g 0.00136519f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_626_n N_A_1525_212#_M1018_g 0.00440079f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_584 N_RESET_B_M1021_g N_A_1525_212#_c_1109_n 0.0193933f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_618_n N_A_1525_212#_c_1109_n 0.00138661f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_586 N_RESET_B_c_621_n N_A_1525_212#_c_1109_n 8.33981e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_625_n N_A_1525_212#_c_1109_n 0.00147213f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_626_n N_A_1525_212#_c_1109_n 4.18149e-19 $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_589 N_RESET_B_M1021_g N_A_1525_212#_c_1110_n 0.013811f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_590 N_RESET_B_M1019_g N_A_1525_212#_c_1120_n 0.0106582f $X=8.235 $Y=2.675
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_625_n N_A_1525_212#_c_1120_n 0.00159476f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_592 N_RESET_B_c_626_n N_A_1525_212#_c_1120_n 0.00783328f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_593 N_RESET_B_M1021_g N_A_1525_212#_c_1111_n 0.00343438f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_594 N_RESET_B_M1019_g N_A_1525_212#_c_1121_n 0.00299204f $X=8.235 $Y=2.675
+ $X2=0 $Y2=0
cc_595 N_RESET_B_c_625_n N_A_1525_212#_c_1123_n 8.22326e-19 $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_596 N_RESET_B_c_626_n N_A_1525_212#_c_1123_n 0.0092621f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1021_g N_A_1525_212#_c_1114_n 0.00118187f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_598 N_RESET_B_M1021_g N_A_1525_212#_c_1115_n 0.021263f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_599 N_RESET_B_c_618_n N_A_1271_74#_M1007_d 0.00237528f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_RESET_B_M1021_g N_A_1271_74#_M1022_g 0.0755988f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_601 N_RESET_B_M1019_g N_A_1271_74#_M1002_g 0.015592f $X=8.235 $Y=2.675 $X2=0
+ $Y2=0
cc_602 N_RESET_B_M1021_g N_A_1271_74#_M1002_g 0.00125436f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_603 N_RESET_B_c_625_n N_A_1271_74#_M1002_g 0.00729506f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_626_n N_A_1271_74#_M1002_g 0.00157069f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_605 N_RESET_B_M1021_g N_A_1271_74#_c_1224_n 0.0061479f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_618_n N_A_1271_74#_c_1237_n 0.0172254f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_618_n N_A_1271_74#_c_1258_n 0.0183959f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_618_n N_A_1271_74#_c_1238_n 0.0225824f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_609 N_RESET_B_c_621_n N_A_1271_74#_c_1238_n 0.00231685f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_RESET_B_c_626_n N_A_1271_74#_c_1238_n 0.023913f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_611 N_RESET_B_M1021_g N_A_1271_74#_c_1229_n 0.0108634f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_618_n N_A_1271_74#_c_1229_n 0.00539223f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_621_n N_A_1271_74#_c_1229_n 0.00832147f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_614 N_RESET_B_c_625_n N_A_1271_74#_c_1229_n 0.00115858f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_615 N_RESET_B_c_626_n N_A_1271_74#_c_1229_n 0.0386217f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_618_n N_A_1271_74#_c_1231_n 0.00597955f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_617 N_RESET_B_M1021_g N_A_1271_74#_c_1242_n 0.00100578f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_618 N_RESET_B_c_616_n N_VPWR_M1025_d 0.00508462f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_619 N_RESET_B_M1015_g N_VPWR_c_1431_n 6.26155e-19 $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_620 N_RESET_B_M1015_g N_VPWR_c_1432_n 0.00850624f $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_621 N_RESET_B_M1017_g N_VPWR_c_1434_n 0.00404978f $X=4.895 $Y=2.525 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_616_n N_VPWR_c_1434_n 8.49328e-19 $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_605_n N_VPWR_c_1436_n 0.001224f $X=4.88 $Y=1.795 $X2=0 $Y2=0
cc_624 N_RESET_B_M1017_g N_VPWR_c_1436_n 0.011992f $X=4.895 $Y=2.525 $X2=0 $Y2=0
cc_625 N_RESET_B_c_618_n N_VPWR_c_1436_n 0.0327022f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_626 N_RESET_B_c_619_n N_VPWR_c_1436_n 5.54746e-19 $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_620_n N_VPWR_c_1436_n 0.0200056f $X=5.04 $Y=2.035 $X2=0 $Y2=0
cc_628 N_RESET_B_c_624_n N_VPWR_c_1436_n 0.00128826f $X=5.12 $Y=1.96 $X2=0 $Y2=0
cc_629 N_RESET_B_M1019_g N_VPWR_c_1437_n 0.00411051f $X=8.235 $Y=2.675 $X2=0
+ $Y2=0
cc_630 N_RESET_B_c_621_n N_VPWR_c_1437_n 0.00199704f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_625_n N_VPWR_c_1437_n 0.00137444f $X=8.23 $Y=2.11 $X2=0 $Y2=0
cc_632 N_RESET_B_c_626_n N_VPWR_c_1437_n 0.0262861f $X=8.23 $Y=2.11 $X2=0 $Y2=0
cc_633 N_RESET_B_M1019_g N_VPWR_c_1442_n 0.00602856f $X=8.235 $Y=2.675 $X2=0
+ $Y2=0
cc_634 N_RESET_B_M1015_g N_VPWR_c_1444_n 0.00401239f $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_635 N_RESET_B_M1015_g N_VPWR_c_1429_n 0.00488819f $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_636 N_RESET_B_M1017_g N_VPWR_c_1429_n 0.00112709f $X=4.895 $Y=2.525 $X2=0
+ $Y2=0
cc_637 N_RESET_B_M1019_g N_VPWR_c_1429_n 0.00626544f $X=8.235 $Y=2.675 $X2=0
+ $Y2=0
cc_638 N_RESET_B_M1012_g N_A_30_78#_c_1581_n 0.00371558f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_639 N_RESET_B_M1015_g N_A_30_78#_c_1587_n 3.52564e-19 $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_640 N_RESET_B_M1012_g N_A_30_78#_c_1582_n 0.00906084f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_601_n N_A_30_78#_c_1582_n 0.0116166f $X=1.055 $Y=1.92 $X2=0
+ $Y2=0
cc_642 N_RESET_B_M1015_g N_A_30_78#_c_1582_n 0.00592134f $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_617_n N_A_30_78#_c_1582_n 0.00138196f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_608_n N_A_30_78#_c_1582_n 0.0048756f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_645 N_RESET_B_c_609_n N_A_30_78#_c_1582_n 0.0697209f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_646 N_RESET_B_c_623_n N_A_30_78#_c_1582_n 0.0049908f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_616_n N_A_30_78#_c_1590_n 0.0120842f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_616_n N_A_30_78#_c_1591_n 0.00529145f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_616_n N_A_30_78#_c_1584_n 0.0107437f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_650 N_RESET_B_M1012_g N_A_30_78#_c_1585_n 9.29579e-19 $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_651 N_RESET_B_M1015_g N_A_30_78#_c_1594_n 0.0201669f $X=0.945 $Y=2.845 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_616_n N_A_30_78#_c_1594_n 0.0268925f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_653 N_RESET_B_c_617_n N_A_30_78#_c_1594_n 0.0041963f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_609_n N_A_30_78#_c_1594_n 0.0105468f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_623_n N_A_30_78#_c_1594_n 0.00227033f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_616_n N_A_30_78#_c_1595_n 0.00477961f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_616_n N_A_30_78#_c_1586_n 0.00582999f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_658 N_RESET_B_M1012_g N_VGND_c_1723_n 0.00258417f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_659 N_RESET_B_c_602_n N_VGND_c_1723_n 0.0200565f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_660 N_RESET_B_c_608_n N_VGND_c_1723_n 0.00180633f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_661 N_RESET_B_c_609_n N_VGND_c_1723_n 0.0140897f $X=1.12 $Y=1.305 $X2=0 $Y2=0
cc_662 N_RESET_B_c_602_n N_VGND_c_1724_n 0.0257898f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_663 N_RESET_B_M1021_g N_VGND_c_1725_n 0.0104625f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_664 N_RESET_B_c_603_n N_VGND_c_1730_n 0.00785671f $X=0.975 $Y=0.18 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_602_n N_VGND_c_1732_n 0.0213429f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_666 N_RESET_B_c_602_n N_VGND_c_1733_n 0.0704334f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_667 N_RESET_B_M1021_g N_VGND_c_1735_n 0.0045897f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_668 N_RESET_B_c_602_n N_VGND_c_1742_n 0.0943738f $X=4.715 $Y=0.18 $X2=0 $Y2=0
cc_669 N_RESET_B_c_603_n N_VGND_c_1742_n 0.0111572f $X=0.975 $Y=0.18 $X2=0 $Y2=0
cc_670 N_RESET_B_M1021_g N_VGND_c_1742_n 0.0044912f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_671 N_A_699_463#_c_822_n N_A_306_119#_c_942_n 0.0027623f $X=4.25 $Y=2.41
+ $X2=0 $Y2=0
cc_672 N_A_699_463#_c_813_n N_A_306_119#_c_931_n 2.82786e-19 $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_673 N_A_699_463#_c_813_n N_A_306_119#_c_933_n 0.00106324f $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_674 N_A_699_463#_c_816_n N_A_306_119#_c_933_n 0.00211731f $X=4.015 $Y=0.867
+ $X2=0 $Y2=0
cc_675 N_A_699_463#_c_813_n N_A_306_119#_M1006_g 0.00262322f $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_676 N_A_699_463#_c_822_n N_A_306_119#_M1006_g 0.0211941f $X=4.25 $Y=2.41
+ $X2=0 $Y2=0
cc_677 N_A_699_463#_M1000_g N_A_306_119#_c_946_n 0.0123711f $X=5.905 $Y=2.235
+ $X2=0 $Y2=0
cc_678 N_A_699_463#_c_821_n N_A_306_119#_c_946_n 0.00102735f $X=4.615 $Y=2.41
+ $X2=0 $Y2=0
cc_679 N_A_699_463#_c_822_n N_A_306_119#_c_946_n 0.00348581f $X=4.25 $Y=2.41
+ $X2=0 $Y2=0
cc_680 N_A_699_463#_c_825_n N_A_306_119#_c_946_n 0.00698065f $X=5.12 $Y=2.44
+ $X2=0 $Y2=0
cc_681 N_A_699_463#_c_826_n N_A_306_119#_c_946_n 4.87622e-19 $X=4.7 $Y=2.41
+ $X2=0 $Y2=0
cc_682 N_A_699_463#_M1000_g N_A_306_119#_c_949_n 0.0174126f $X=5.905 $Y=2.235
+ $X2=0 $Y2=0
cc_683 N_A_699_463#_c_821_n N_VPWR_M1011_d 0.0026266f $X=4.615 $Y=2.41 $X2=0
+ $Y2=0
cc_684 N_A_699_463#_c_826_n N_VPWR_M1011_d 0.00142227f $X=4.7 $Y=2.41 $X2=0
+ $Y2=0
cc_685 N_A_699_463#_c_821_n N_VPWR_c_1434_n 0.0152182f $X=4.615 $Y=2.41 $X2=0
+ $Y2=0
cc_686 N_A_699_463#_c_822_n N_VPWR_c_1434_n 0.0121695f $X=4.25 $Y=2.41 $X2=0
+ $Y2=0
cc_687 N_A_699_463#_c_826_n N_VPWR_c_1434_n 0.0114153f $X=4.7 $Y=2.41 $X2=0
+ $Y2=0
cc_688 N_A_699_463#_M1000_g N_VPWR_c_1436_n 0.0168944f $X=5.905 $Y=2.235 $X2=0
+ $Y2=0
cc_689 N_A_699_463#_c_811_n N_VPWR_c_1436_n 0.0075672f $X=5.73 $Y=1.41 $X2=0
+ $Y2=0
cc_690 N_A_699_463#_c_815_n N_VPWR_c_1436_n 0.0131953f $X=5.52 $Y=1.41 $X2=0
+ $Y2=0
cc_691 N_A_699_463#_c_825_n N_VPWR_c_1436_n 0.0145224f $X=5.12 $Y=2.44 $X2=0
+ $Y2=0
cc_692 N_A_699_463#_c_822_n N_VPWR_c_1446_n 0.0200693f $X=4.25 $Y=2.41 $X2=0
+ $Y2=0
cc_693 N_A_699_463#_M1000_g N_VPWR_c_1429_n 9.455e-19 $X=5.905 $Y=2.235 $X2=0
+ $Y2=0
cc_694 N_A_699_463#_c_821_n N_VPWR_c_1429_n 0.0058609f $X=4.615 $Y=2.41 $X2=0
+ $Y2=0
cc_695 N_A_699_463#_c_822_n N_VPWR_c_1429_n 0.0206807f $X=4.25 $Y=2.41 $X2=0
+ $Y2=0
cc_696 N_A_699_463#_c_825_n N_VPWR_c_1429_n 0.0155369f $X=5.12 $Y=2.44 $X2=0
+ $Y2=0
cc_697 N_A_699_463#_c_826_n N_VPWR_c_1429_n 0.0018405f $X=4.7 $Y=2.41 $X2=0
+ $Y2=0
cc_698 N_A_699_463#_c_813_n N_A_30_78#_c_1589_n 4.86922e-19 $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_699 N_A_699_463#_c_822_n N_A_30_78#_c_1589_n 0.00430685f $X=4.25 $Y=2.41
+ $X2=0 $Y2=0
cc_700 N_A_699_463#_c_813_n N_A_30_78#_c_1583_n 0.0049664f $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_701 N_A_699_463#_c_816_n N_A_30_78#_c_1583_n 0.014993f $X=4.015 $Y=0.867
+ $X2=0 $Y2=0
cc_702 N_A_699_463#_c_813_n N_A_30_78#_c_1590_n 0.0136648f $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_703 N_A_699_463#_c_822_n N_A_30_78#_c_1590_n 0.0152881f $X=4.25 $Y=2.41 $X2=0
+ $Y2=0
cc_704 N_A_699_463#_c_813_n N_A_30_78#_c_1584_n 0.0501235f $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_705 N_A_699_463#_c_813_n N_A_30_78#_c_1586_n 0.0139397f $X=4.015 $Y=2.295
+ $X2=0 $Y2=0
cc_706 N_A_699_463#_c_816_n N_A_30_78#_c_1586_n 0.00975559f $X=4.015 $Y=0.867
+ $X2=0 $Y2=0
cc_707 N_A_699_463#_M1023_g N_VGND_c_1733_n 0.0012551f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_708 N_A_699_463#_M1023_g N_VGND_c_1734_n 0.00278271f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_709 N_A_699_463#_M1023_g N_VGND_c_1742_n 0.00358928f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_710 N_A_306_119#_M1032_g N_A_1525_212#_M1005_g 0.0390746f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_711 N_A_306_119#_M1032_g N_A_1525_212#_c_1109_n 0.0184343f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_712 N_A_306_119#_M1032_g N_A_1525_212#_c_1114_n 4.84439e-19 $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_713 N_A_306_119#_M1032_g N_A_1525_212#_c_1115_n 0.0192269f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_714 N_A_306_119#_c_949_n N_A_1271_74#_c_1227_n 2.48308e-19 $X=6.5 $Y=1.66
+ $X2=0 $Y2=0
cc_715 N_A_306_119#_M1007_g N_A_1271_74#_c_1237_n 0.0107145f $X=6.41 $Y=2.31
+ $X2=0 $Y2=0
cc_716 N_A_306_119#_c_934_n N_A_1271_74#_c_1237_n 0.00688552f $X=7.255 $Y=1.66
+ $X2=0 $Y2=0
cc_717 N_A_306_119#_M1032_g N_A_1271_74#_c_1228_n 0.00513624f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_718 N_A_306_119#_M1032_g N_A_1271_74#_c_1230_n 0.00152295f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_719 N_A_306_119#_c_934_n N_A_1271_74#_c_1231_n 0.00502126f $X=7.255 $Y=1.66
+ $X2=0 $Y2=0
cc_720 N_A_306_119#_c_949_n N_A_1271_74#_c_1231_n 0.00503723f $X=6.5 $Y=1.66
+ $X2=0 $Y2=0
cc_721 N_A_306_119#_M1032_g N_A_1271_74#_c_1231_n 2.71569e-19 $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_722 N_A_306_119#_M1027_g N_VPWR_c_1433_n 0.0105012f $X=2.375 $Y=2.495 $X2=0
+ $Y2=0
cc_723 N_A_306_119#_c_941_n N_VPWR_c_1433_n 0.00203408f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_724 N_A_306_119#_c_943_n N_VPWR_c_1433_n 7.08583e-19 $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_725 N_A_306_119#_M1006_g N_VPWR_c_1434_n 0.00575867f $X=3.855 $Y=2.525 $X2=0
+ $Y2=0
cc_726 N_A_306_119#_c_946_n N_VPWR_c_1434_n 0.0252266f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_727 N_A_306_119#_c_946_n N_VPWR_c_1435_n 0.026968f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_728 N_A_306_119#_c_946_n N_VPWR_c_1436_n 0.025641f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_729 N_A_306_119#_M1007_g N_VPWR_c_1436_n 0.00644903f $X=6.41 $Y=2.31 $X2=0
+ $Y2=0
cc_730 N_A_306_119#_M1027_g N_VPWR_c_1446_n 0.00401239f $X=2.375 $Y=2.495 $X2=0
+ $Y2=0
cc_731 N_A_306_119#_c_943_n N_VPWR_c_1446_n 0.0443244f $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_732 N_A_306_119#_c_946_n N_VPWR_c_1447_n 0.0203802f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_306_119#_M1027_g N_VPWR_c_1429_n 0.00500024f $X=2.375 $Y=2.495 $X2=0
+ $Y2=0
cc_734 N_A_306_119#_c_942_n N_VPWR_c_1429_n 0.0234871f $X=3.765 $Y=3.15 $X2=0
+ $Y2=0
cc_735 N_A_306_119#_c_943_n N_VPWR_c_1429_n 0.00587633f $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_736 N_A_306_119#_c_946_n N_VPWR_c_1429_n 0.0663876f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_737 N_A_306_119#_c_950_n N_VPWR_c_1429_n 0.00473439f $X=3.855 $Y=3.15 $X2=0
+ $Y2=0
cc_738 N_A_306_119#_c_936_n N_A_30_78#_c_1582_n 0.0042997f $X=1.675 $Y=0.725
+ $X2=0 $Y2=0
cc_739 N_A_306_119#_c_939_n N_A_30_78#_c_1582_n 0.00486522f $X=1.647 $Y=1.065
+ $X2=0 $Y2=0
cc_740 N_A_306_119#_c_953_n N_A_30_78#_c_1582_n 0.00402797f $X=1.7 $Y=2.11 $X2=0
+ $Y2=0
cc_741 N_A_306_119#_c_941_n N_A_30_78#_c_1589_n 0.00329814f $X=2.88 $Y=3.075
+ $X2=0 $Y2=0
cc_742 N_A_306_119#_M1006_g N_A_30_78#_c_1589_n 4.58537e-19 $X=3.855 $Y=2.525
+ $X2=0 $Y2=0
cc_743 N_A_306_119#_c_931_n N_A_30_78#_c_1583_n 0.00836137f $X=3.435 $Y=1.275
+ $X2=0 $Y2=0
cc_744 N_A_306_119#_c_933_n N_A_30_78#_c_1583_n 0.00852665f $X=3.51 $Y=1.185
+ $X2=0 $Y2=0
cc_745 N_A_306_119#_M1006_g N_A_30_78#_c_1590_n 0.00105368f $X=3.855 $Y=2.525
+ $X2=0 $Y2=0
cc_746 N_A_306_119#_c_941_n N_A_30_78#_c_1591_n 5.6937e-19 $X=2.88 $Y=3.075
+ $X2=0 $Y2=0
cc_747 N_A_306_119#_c_932_n N_A_30_78#_c_1584_n 0.00165379f $X=3.04 $Y=1.275
+ $X2=0 $Y2=0
cc_748 N_A_306_119#_M1025_s N_A_30_78#_c_1594_n 0.00684204f $X=1.57 $Y=1.935
+ $X2=0 $Y2=0
cc_749 N_A_306_119#_M1027_g N_A_30_78#_c_1594_n 0.0149926f $X=2.375 $Y=2.495
+ $X2=0 $Y2=0
cc_750 N_A_306_119#_c_941_n N_A_30_78#_c_1594_n 0.0132721f $X=2.88 $Y=3.075
+ $X2=0 $Y2=0
cc_751 N_A_306_119#_c_953_n N_A_30_78#_c_1594_n 0.0256049f $X=1.7 $Y=2.11 $X2=0
+ $Y2=0
cc_752 N_A_306_119#_c_941_n N_A_30_78#_c_1595_n 0.00281908f $X=2.88 $Y=3.075
+ $X2=0 $Y2=0
cc_753 N_A_306_119#_c_942_n N_A_30_78#_c_1595_n 0.00493823f $X=3.765 $Y=3.15
+ $X2=0 $Y2=0
cc_754 N_A_306_119#_c_931_n N_A_30_78#_c_1586_n 0.0150416f $X=3.435 $Y=1.275
+ $X2=0 $Y2=0
cc_755 N_A_306_119#_c_932_n N_A_30_78#_c_1586_n 8.09864e-19 $X=3.04 $Y=1.275
+ $X2=0 $Y2=0
cc_756 N_A_306_119#_c_965_n N_VGND_M1016_d 0.00731677f $X=2.445 $Y=1.065 $X2=0
+ $Y2=0
cc_757 N_A_306_119#_c_936_n N_VGND_c_1723_n 0.0218337f $X=1.675 $Y=0.725 $X2=0
+ $Y2=0
cc_758 N_A_306_119#_c_930_n N_VGND_c_1724_n 0.00252184f $X=2.46 $Y=1.41 $X2=0
+ $Y2=0
cc_759 N_A_306_119#_c_936_n N_VGND_c_1724_n 0.0110191f $X=1.675 $Y=0.725 $X2=0
+ $Y2=0
cc_760 N_A_306_119#_c_965_n N_VGND_c_1724_n 0.0248957f $X=2.445 $Y=1.065 $X2=0
+ $Y2=0
cc_761 N_A_306_119#_M1032_g N_VGND_c_1725_n 4.38128e-19 $X=7.33 $Y=0.615 $X2=0
+ $Y2=0
cc_762 N_A_306_119#_c_936_n N_VGND_c_1732_n 0.00901682f $X=1.675 $Y=0.725 $X2=0
+ $Y2=0
cc_763 N_A_306_119#_M1032_g N_VGND_c_1734_n 9.34015e-19 $X=7.33 $Y=0.615 $X2=0
+ $Y2=0
cc_764 N_A_306_119#_c_930_n N_VGND_c_1742_n 7.88961e-19 $X=2.46 $Y=1.41 $X2=0
+ $Y2=0
cc_765 N_A_306_119#_c_936_n N_VGND_c_1742_n 0.0106863f $X=1.675 $Y=0.725 $X2=0
+ $Y2=0
cc_766 N_A_1525_212#_c_1110_n N_A_1271_74#_M1022_g 0.0108536f $X=8.68 $Y=1.305
+ $X2=0 $Y2=0
cc_767 N_A_1525_212#_c_1111_n N_A_1271_74#_M1022_g 0.0236543f $X=8.845 $Y=0.615
+ $X2=0 $Y2=0
cc_768 N_A_1525_212#_c_1113_n N_A_1271_74#_M1022_g 0.00397247f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_769 N_A_1525_212#_c_1116_n N_A_1271_74#_M1022_g 0.00478437f $X=8.845 $Y=1.305
+ $X2=0 $Y2=0
cc_770 N_A_1525_212#_c_1120_n N_A_1271_74#_M1002_g 0.0105922f $X=8.715 $Y=2.61
+ $X2=0 $Y2=0
cc_771 N_A_1525_212#_c_1121_n N_A_1271_74#_M1002_g 0.00530253f $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_772 N_A_1525_212#_c_1122_n N_A_1271_74#_M1002_g 0.0135181f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_773 N_A_1525_212#_c_1123_n N_A_1271_74#_M1002_g 0.00277746f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_774 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1223_n 0.00213341f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_775 N_A_1525_212#_c_1113_n N_A_1271_74#_c_1223_n 0.0139731f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_776 N_A_1525_212#_c_1123_n N_A_1271_74#_c_1224_n 0.0010617f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_777 N_A_1525_212#_c_1112_n N_A_1271_74#_c_1224_n 0.00714341f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_778 N_A_1525_212#_c_1113_n N_A_1271_74#_c_1224_n 0.0061655f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_779 N_A_1525_212#_c_1116_n N_A_1271_74#_c_1224_n 0.00565398f $X=8.845
+ $Y=1.305 $X2=0 $Y2=0
cc_780 N_A_1525_212#_c_1121_n N_A_1271_74#_M1010_g 7.68645e-19 $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_781 N_A_1525_212#_c_1122_n N_A_1271_74#_M1010_g 0.00178565f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_782 N_A_1525_212#_c_1113_n N_A_1271_74#_M1010_g 0.00400887f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_783 N_A_1525_212#_c_1111_n N_A_1271_74#_M1020_g 0.00350395f $X=8.845 $Y=0.615
+ $X2=0 $Y2=0
cc_784 N_A_1525_212#_c_1112_n N_A_1271_74#_M1020_g 0.00377053f $X=9.205 $Y=1.305
+ $X2=0 $Y2=0
cc_785 N_A_1525_212#_c_1113_n N_A_1271_74#_M1020_g 0.00338537f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_786 N_A_1525_212#_c_1109_n N_A_1271_74#_c_1238_n 0.0152224f $X=7.735 $Y=1.975
+ $X2=0 $Y2=0
cc_787 N_A_1525_212#_c_1117_n N_A_1271_74#_c_1229_n 2.78407e-19 $X=7.735
+ $Y=2.065 $X2=0 $Y2=0
cc_788 N_A_1525_212#_c_1109_n N_A_1271_74#_c_1229_n 0.0105806f $X=7.735 $Y=1.975
+ $X2=0 $Y2=0
cc_789 N_A_1525_212#_c_1110_n N_A_1271_74#_c_1229_n 0.0522284f $X=8.68 $Y=1.305
+ $X2=0 $Y2=0
cc_790 N_A_1525_212#_c_1114_n N_A_1271_74#_c_1229_n 0.023491f $X=7.79 $Y=1.225
+ $X2=0 $Y2=0
cc_791 N_A_1525_212#_c_1115_n N_A_1271_74#_c_1229_n 0.00116263f $X=7.79 $Y=1.225
+ $X2=0 $Y2=0
cc_792 N_A_1525_212#_c_1116_n N_A_1271_74#_c_1229_n 0.00190438f $X=8.845
+ $Y=1.305 $X2=0 $Y2=0
cc_793 N_A_1525_212#_c_1120_n N_A_1271_74#_c_1242_n 2.74753e-19 $X=8.715 $Y=2.61
+ $X2=0 $Y2=0
cc_794 N_A_1525_212#_c_1122_n N_A_1271_74#_c_1242_n 0.00882758f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_795 N_A_1525_212#_c_1123_n N_A_1271_74#_c_1242_n 0.0119175f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_796 N_A_1525_212#_c_1112_n N_A_1271_74#_c_1242_n 0.00177485f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_797 N_A_1525_212#_c_1113_n N_A_1271_74#_c_1242_n 0.0242588f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_798 N_A_1525_212#_c_1116_n N_A_1271_74#_c_1242_n 0.0257641f $X=8.845 $Y=1.305
+ $X2=0 $Y2=0
cc_799 N_A_1525_212#_c_1122_n N_A_1924_409#_c_1376_n 0.0116529f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_800 N_A_1525_212#_c_1113_n N_A_1924_409#_c_1376_n 0.00461164f $X=9.29
+ $Y=2.105 $X2=0 $Y2=0
cc_801 N_A_1525_212#_c_1111_n N_A_1924_409#_c_1370_n 0.00484112f $X=8.845
+ $Y=0.615 $X2=0 $Y2=0
cc_802 N_A_1525_212#_c_1112_n N_A_1924_409#_c_1370_n 0.00459026f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_803 N_A_1525_212#_c_1113_n N_A_1924_409#_c_1371_n 0.0210731f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_804 N_A_1525_212#_c_1112_n N_A_1924_409#_c_1372_n 0.00528833f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_805 N_A_1525_212#_c_1113_n N_A_1924_409#_c_1372_n 0.0123556f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_806 N_A_1525_212#_c_1122_n N_VPWR_M1002_d 0.00762771f $X=9.205 $Y=2.19 $X2=0
+ $Y2=0
cc_807 N_A_1525_212#_c_1113_n N_VPWR_M1002_d 0.00172994f $X=9.29 $Y=2.105 $X2=0
+ $Y2=0
cc_808 N_A_1525_212#_M1018_g N_VPWR_c_1437_n 0.0110188f $X=7.735 $Y=2.675 $X2=0
+ $Y2=0
cc_809 N_A_1525_212#_c_1120_n N_VPWR_c_1437_n 0.0142734f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_810 N_A_1525_212#_c_1120_n N_VPWR_c_1438_n 0.0123985f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_811 N_A_1525_212#_c_1122_n N_VPWR_c_1438_n 0.0245347f $X=9.205 $Y=2.19 $X2=0
+ $Y2=0
cc_812 N_A_1525_212#_c_1120_n N_VPWR_c_1442_n 0.0118789f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_813 N_A_1525_212#_M1018_g N_VPWR_c_1447_n 0.00522765f $X=7.735 $Y=2.675 $X2=0
+ $Y2=0
cc_814 N_A_1525_212#_M1018_g N_VPWR_c_1429_n 0.005256f $X=7.735 $Y=2.675 $X2=0
+ $Y2=0
cc_815 N_A_1525_212#_c_1120_n N_VPWR_c_1429_n 0.0184861f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_816 N_A_1525_212#_M1005_g N_VGND_c_1725_n 0.00870177f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_817 N_A_1525_212#_c_1110_n N_VGND_c_1725_n 0.00751614f $X=8.68 $Y=1.305 $X2=0
+ $Y2=0
cc_818 N_A_1525_212#_c_1111_n N_VGND_c_1725_n 0.0106511f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_819 N_A_1525_212#_c_1114_n N_VGND_c_1725_n 0.00718492f $X=7.79 $Y=1.225 $X2=0
+ $Y2=0
cc_820 N_A_1525_212#_c_1115_n N_VGND_c_1725_n 9.12984e-19 $X=7.79 $Y=1.225 $X2=0
+ $Y2=0
cc_821 N_A_1525_212#_c_1111_n N_VGND_c_1726_n 0.045283f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_822 N_A_1525_212#_c_1112_n N_VGND_c_1726_n 0.0132803f $X=9.205 $Y=1.305 $X2=0
+ $Y2=0
cc_823 N_A_1525_212#_M1005_g N_VGND_c_1734_n 0.0045897f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_824 N_A_1525_212#_c_1111_n N_VGND_c_1735_n 0.0127604f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_825 N_A_1525_212#_M1005_g N_VGND_c_1742_n 0.0044912f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_826 N_A_1525_212#_c_1111_n N_VGND_c_1742_n 0.011834f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_827 N_A_1271_74#_M1002_g N_A_1924_409#_c_1376_n 8.58951e-19 $X=8.945 $Y=2.675
+ $X2=0 $Y2=0
cc_828 N_A_1271_74#_M1010_g N_A_1924_409#_c_1376_n 0.0174933f $X=9.53 $Y=2.465
+ $X2=0 $Y2=0
cc_829 N_A_1271_74#_c_1226_n N_A_1924_409#_c_1376_n 0.0016406f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_830 N_A_1271_74#_M1020_g N_A_1924_409#_c_1370_n 0.0181066f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_831 N_A_1271_74#_M1010_g N_A_1924_409#_c_1371_n 0.00820455f $X=9.53 $Y=2.465
+ $X2=0 $Y2=0
cc_832 N_A_1271_74#_c_1226_n N_A_1924_409#_c_1371_n 0.00365747f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_833 N_A_1271_74#_M1020_g N_A_1924_409#_c_1372_n 0.00613547f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_834 N_A_1271_74#_c_1226_n N_A_1924_409#_c_1372_n 0.00242696f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_835 N_A_1271_74#_M1020_g N_A_1924_409#_c_1373_n 0.0181431f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_836 N_A_1271_74#_c_1238_n N_VPWR_c_1437_n 0.0018405f $X=7.54 $Y=2.475 $X2=0
+ $Y2=0
cc_837 N_A_1271_74#_M1002_g N_VPWR_c_1438_n 0.00645834f $X=8.945 $Y=2.675 $X2=0
+ $Y2=0
cc_838 N_A_1271_74#_M1010_g N_VPWR_c_1438_n 0.00384793f $X=9.53 $Y=2.465 $X2=0
+ $Y2=0
cc_839 N_A_1271_74#_M1010_g N_VPWR_c_1439_n 0.00480399f $X=9.53 $Y=2.465 $X2=0
+ $Y2=0
cc_840 N_A_1271_74#_M1002_g N_VPWR_c_1442_n 0.00602837f $X=8.945 $Y=2.675 $X2=0
+ $Y2=0
cc_841 N_A_1271_74#_c_1258_n N_VPWR_c_1447_n 0.0205727f $X=7.455 $Y=2.64 $X2=0
+ $Y2=0
cc_842 N_A_1271_74#_c_1346_p N_VPWR_c_1447_n 0.00373537f $X=6.685 $Y=2.64 $X2=0
+ $Y2=0
cc_843 N_A_1271_74#_M1010_g N_VPWR_c_1448_n 0.00601158f $X=9.53 $Y=2.465 $X2=0
+ $Y2=0
cc_844 N_A_1271_74#_M1002_g N_VPWR_c_1429_n 0.00626544f $X=8.945 $Y=2.675 $X2=0
+ $Y2=0
cc_845 N_A_1271_74#_M1010_g N_VPWR_c_1429_n 0.00626544f $X=9.53 $Y=2.465 $X2=0
+ $Y2=0
cc_846 N_A_1271_74#_c_1258_n N_VPWR_c_1429_n 0.0299068f $X=7.455 $Y=2.64 $X2=0
+ $Y2=0
cc_847 N_A_1271_74#_c_1346_p N_VPWR_c_1429_n 0.00557315f $X=6.685 $Y=2.64 $X2=0
+ $Y2=0
cc_848 N_A_1271_74#_c_1258_n A_1481_493# 0.00204811f $X=7.455 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_849 N_A_1271_74#_M1022_g N_VGND_c_1725_n 0.00147575f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_850 N_A_1271_74#_M1022_g N_VGND_c_1726_n 0.00438924f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_851 N_A_1271_74#_c_1223_n N_VGND_c_1726_n 0.00294706f $X=9.44 $Y=1.63 $X2=0
+ $Y2=0
cc_852 N_A_1271_74#_M1020_g N_VGND_c_1726_n 0.00488092f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_853 N_A_1271_74#_M1020_g N_VGND_c_1727_n 0.00412165f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_854 N_A_1271_74#_M1022_g N_VGND_c_1735_n 0.00527282f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_855 N_A_1271_74#_M1020_g N_VGND_c_1736_n 0.00434272f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_856 N_A_1271_74#_M1022_g N_VGND_c_1742_n 0.00534666f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_857 N_A_1271_74#_M1020_g N_VGND_c_1742_n 0.00830282f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_858 N_A_1924_409#_c_1376_n N_VPWR_c_1438_n 0.0180508f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_859 N_A_1924_409#_c_1362_n N_VPWR_c_1439_n 0.00728605f $X=10.475 $Y=1.375
+ $X2=0 $Y2=0
cc_860 N_A_1924_409#_M1029_g N_VPWR_c_1439_n 0.0218803f $X=10.565 $Y=2.4 $X2=0
+ $Y2=0
cc_861 N_A_1924_409#_M1030_g N_VPWR_c_1439_n 6.51046e-19 $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_862 N_A_1924_409#_c_1371_n N_VPWR_c_1439_n 0.072832f $X=9.755 $Y=2.03 $X2=0
+ $Y2=0
cc_863 N_A_1924_409#_c_1372_n N_VPWR_c_1439_n 0.00302521f $X=10.09 $Y=1.465
+ $X2=0 $Y2=0
cc_864 N_A_1924_409#_c_1373_n N_VPWR_c_1439_n 0.00372647f $X=10.09 $Y=1.375
+ $X2=0 $Y2=0
cc_865 N_A_1924_409#_M1030_g N_VPWR_c_1441_n 0.00518749f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_866 N_A_1924_409#_c_1376_n N_VPWR_c_1448_n 0.0111522f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_867 N_A_1924_409#_M1029_g N_VPWR_c_1449_n 0.00532442f $X=10.565 $Y=2.4 $X2=0
+ $Y2=0
cc_868 N_A_1924_409#_M1030_g N_VPWR_c_1449_n 0.00492575f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_869 N_A_1924_409#_M1029_g N_VPWR_c_1429_n 0.0104063f $X=10.565 $Y=2.4 $X2=0
+ $Y2=0
cc_870 N_A_1924_409#_M1030_g N_VPWR_c_1429_n 0.0089429f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_871 N_A_1924_409#_c_1376_n N_VPWR_c_1429_n 0.0115238f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_872 N_A_1924_409#_M1029_g Q 0.0327276f $X=10.565 $Y=2.4 $X2=0 $Y2=0
cc_873 N_A_1924_409#_M1031_g Q 0.0157053f $X=10.6 $Y=0.74 $X2=0 $Y2=0
cc_874 N_A_1924_409#_c_1365_n Q 0.00813241f $X=10.925 $Y=1.375 $X2=0 $Y2=0
cc_875 N_A_1924_409#_M1030_g Q 0.0386825f $X=11.015 $Y=2.4 $X2=0 $Y2=0
cc_876 N_A_1924_409#_M1033_g Q 0.0192861f $X=11.03 $Y=0.74 $X2=0 $Y2=0
cc_877 N_A_1924_409#_c_1368_n Q 0.00396751f $X=10.575 $Y=1.375 $X2=0 $Y2=0
cc_878 N_A_1924_409#_c_1369_n Q 0.00693891f $X=11.015 $Y=1.375 $X2=0 $Y2=0
cc_879 N_A_1924_409#_c_1370_n Q 0.00478422f $X=9.825 $Y=0.515 $X2=0 $Y2=0
cc_880 N_A_1924_409#_c_1372_n Q 0.0113958f $X=10.09 $Y=1.465 $X2=0 $Y2=0
cc_881 N_A_1924_409#_c_1373_n Q 5.0889e-19 $X=10.09 $Y=1.375 $X2=0 $Y2=0
cc_882 N_A_1924_409#_c_1370_n N_VGND_c_1726_n 0.0258169f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_883 N_A_1924_409#_M1031_g N_VGND_c_1727_n 0.00647412f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_884 N_A_1924_409#_c_1370_n N_VGND_c_1727_n 0.051504f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_885 N_A_1924_409#_c_1373_n N_VGND_c_1727_n 0.0102912f $X=10.09 $Y=1.375 $X2=0
+ $Y2=0
cc_886 N_A_1924_409#_M1033_g N_VGND_c_1729_n 0.00647412f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_887 N_A_1924_409#_c_1370_n N_VGND_c_1736_n 0.0145639f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_888 N_A_1924_409#_M1031_g N_VGND_c_1737_n 0.00434272f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_889 N_A_1924_409#_M1033_g N_VGND_c_1737_n 0.00434272f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_890 N_A_1924_409#_M1031_g N_VGND_c_1742_n 0.00825283f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_891 N_A_1924_409#_M1033_g N_VGND_c_1742_n 0.00823925f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_892 N_A_1924_409#_c_1370_n N_VGND_c_1742_n 0.0119984f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1431_n N_A_30_78#_c_1587_n 0.0144417f $X=0.27 $Y=2.845 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1444_n N_A_30_78#_c_1587_n 0.0110259f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1429_n N_A_30_78#_c_1587_n 0.00761614f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1431_n N_A_30_78#_c_1593_n 0.00783618f $X=0.27 $Y=2.845 $X2=0
+ $Y2=0
cc_897 N_VPWR_M1025_d N_A_30_78#_c_1594_n 0.00446117f $X=2.015 $Y=1.935 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1432_n N_A_30_78#_c_1594_n 0.0233375f $X=1.17 $Y=2.88 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1433_n N_A_30_78#_c_1594_n 0.016342f $X=2.15 $Y=2.88 $X2=0 $Y2=0
cc_900 N_VPWR_c_1444_n N_A_30_78#_c_1594_n 0.00240209f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1445_n N_A_30_78#_c_1594_n 0.00942193f $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1446_n N_A_30_78#_c_1594_n 0.00993548f $X=4.42 $Y=3.33 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_1429_n N_A_30_78#_c_1594_n 0.0406792f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1446_n N_A_30_78#_c_1595_n 0.00639259f $X=4.42 $Y=3.33 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1429_n N_A_30_78#_c_1595_n 0.0092373f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1439_n Q 0.0870519f $X=10.315 $Y=1.985 $X2=0 $Y2=0
cc_907 N_VPWR_c_1441_n Q 0.0440104f $X=11.24 $Y=1.985 $X2=0 $Y2=0
cc_908 N_VPWR_c_1449_n Q 0.0144623f $X=11.155 $Y=3.33 $X2=0 $Y2=0
cc_909 N_VPWR_c_1429_n Q 0.0118344f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_910 N_A_30_78#_c_1581_n A_117_78# 0.00232882f $X=0.665 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_911 N_A_30_78#_c_1581_n N_VGND_c_1723_n 0.00655394f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_912 N_A_30_78#_c_1585_n N_VGND_c_1723_n 0.00436551f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_913 N_A_30_78#_c_1581_n N_VGND_c_1730_n 0.00539861f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_914 N_A_30_78#_c_1585_n N_VGND_c_1730_n 0.0131067f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_915 N_A_30_78#_c_1581_n N_VGND_c_1742_n 0.0106165f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_916 N_A_30_78#_c_1585_n N_VGND_c_1742_n 0.0117869f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_917 Q N_VGND_c_1727_n 0.0294122f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_918 Q N_VGND_c_1729_n 0.0294122f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_919 Q N_VGND_c_1737_n 0.0144922f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_920 Q N_VGND_c_1742_n 0.0118826f $X=10.715 $Y=0.47 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.495000 2.170000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.650000 0.350000 10.980000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.415800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.140000 1.285000 2.150000 ;
        RECT 4.955000 1.795000 5.285000 2.150000 ;
        RECT 7.805000 1.920000 8.395000 2.275000 ;
      LAYER mcon ;
        RECT 1.115000 1.950000 1.285000 2.120000 ;
        RECT 4.955000 1.950000 5.125000 2.120000 ;
        RECT 7.835000 1.950000 8.005000 2.120000 ;
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 8.065000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 4.895000 1.920000 5.185000 1.965000 ;
        RECT 4.895000 2.105000 5.185000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.320000 2.275000 1.775000 ;
        RECT 2.045000 1.775000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.520000 0.085000 ;
        RECT  1.030000  0.085000  1.280000 0.830000 ;
        RECT  2.010000  0.085000  2.340000 0.810000 ;
        RECT  4.920000  0.085000  5.345000 0.445000 ;
        RECT  7.770000  0.085000  8.190000 0.715000 ;
        RECT  9.230000  0.085000  9.480000 1.050000 ;
        RECT 10.220000  0.085000 10.470000 1.130000 ;
        RECT 11.160000  0.085000 11.410000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.520000 3.415000 ;
        RECT  0.105000 2.520000  0.435000 3.245000 ;
        RECT  1.005000 2.795000  1.335000 3.245000 ;
        RECT  1.985000 2.795000  2.315000 3.245000 ;
        RECT  4.420000 2.695000  4.750000 3.245000 ;
        RECT  5.515000 1.745000  5.845000 3.245000 ;
        RECT  7.795000 2.445000  8.125000 3.245000 ;
        RECT  9.090000 2.445000  9.420000 3.245000 ;
        RECT 10.150000 1.820000 10.480000 3.245000 ;
        RECT 11.155000 1.820000 11.405000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.130000 0.370000  0.460000 0.660000 ;
      RECT 0.130000 0.660000  0.835000 0.830000 ;
      RECT 0.635000 2.520000  3.375000 2.625000 ;
      RECT 0.635000 2.625000  0.835000 3.055000 ;
      RECT 0.665000 0.830000  0.835000 2.445000 ;
      RECT 0.665000 2.445000  3.375000 2.520000 ;
      RECT 1.455000 0.560000  1.840000 0.980000 ;
      RECT 1.455000 0.980000  2.700000 1.150000 ;
      RECT 1.455000 1.150000  1.625000 1.945000 ;
      RECT 1.455000 1.945000  1.865000 2.275000 ;
      RECT 2.445000 1.150000  2.700000 1.550000 ;
      RECT 2.510000 0.330000  4.440000 0.500000 ;
      RECT 2.510000 0.500000  3.040000 0.810000 ;
      RECT 2.515000 1.550000  2.700000 1.775000 ;
      RECT 2.515000 1.945000  3.080000 1.985000 ;
      RECT 2.515000 1.985000  3.055000 2.025000 ;
      RECT 2.515000 2.025000  3.035000 2.275000 ;
      RECT 2.825000 1.895000  3.420000 1.935000 ;
      RECT 2.825000 1.935000  3.080000 1.945000 ;
      RECT 2.850000 1.855000  3.420000 1.895000 ;
      RECT 2.870000 0.810000  3.040000 1.605000 ;
      RECT 2.870000 1.605000  3.420000 1.855000 ;
      RECT 3.015000 2.625000  3.375000 2.725000 ;
      RECT 3.205000 2.105000  3.760000 2.275000 ;
      RECT 3.205000 2.275000  3.375000 2.445000 ;
      RECT 3.210000 0.670000  3.460000 1.235000 ;
      RECT 3.210000 1.235000  3.760000 1.405000 ;
      RECT 3.545000 2.445000  5.285000 2.525000 ;
      RECT 3.545000 2.525000  4.250000 2.860000 ;
      RECT 3.590000 1.405000  3.760000 2.105000 ;
      RECT 3.630000 0.670000  4.100000 1.065000 ;
      RECT 3.930000 1.065000  4.100000 2.295000 ;
      RECT 3.930000 2.295000  4.785000 2.320000 ;
      RECT 3.930000 2.320000  5.285000 2.445000 ;
      RECT 4.270000 0.500000  4.440000 0.615000 ;
      RECT 4.270000 0.615000  5.685000 0.785000 ;
      RECT 4.270000 0.955000  6.185000 1.125000 ;
      RECT 4.270000 1.125000  4.445000 2.125000 ;
      RECT 4.615000 1.295000  5.685000 1.575000 ;
      RECT 4.615000 1.575000  4.785000 2.295000 ;
      RECT 5.515000 0.255000  7.455000 0.425000 ;
      RECT 5.515000 0.425000  5.685000 0.615000 ;
      RECT 5.855000 0.595000  6.185000 0.955000 ;
      RECT 5.855000 1.125000  6.185000 1.130000 ;
      RECT 6.015000 1.130000  6.185000 1.855000 ;
      RECT 6.015000 1.855000  6.345000 2.755000 ;
      RECT 6.355000 0.595000  7.115000 0.845000 ;
      RECT 6.355000 0.845000  6.525000 1.515000 ;
      RECT 6.355000 1.515000  6.685000 1.685000 ;
      RECT 6.515000 1.685000  6.685000 2.475000 ;
      RECT 6.515000 2.475000  7.625000 2.805000 ;
      RECT 6.725000 1.015000  7.455000 1.345000 ;
      RECT 6.955000 1.345000  7.285000 2.305000 ;
      RECT 7.285000 0.425000  7.455000 1.015000 ;
      RECT 7.455000 1.560000  9.035000 1.730000 ;
      RECT 7.455000 1.730000  7.625000 2.475000 ;
      RECT 7.625000 1.060000  7.955000 1.220000 ;
      RECT 7.625000 1.220000  9.375000 1.390000 ;
      RECT 8.295000 2.445000  8.885000 2.775000 ;
      RECT 8.680000 0.385000  9.010000 1.220000 ;
      RECT 8.705000 1.730000  9.035000 1.890000 ;
      RECT 8.715000 2.105000  9.375000 2.275000 ;
      RECT 8.715000 2.275000  8.885000 2.445000 ;
      RECT 9.205000 1.390000  9.375000 2.105000 ;
      RECT 9.590000 2.030000  9.920000 2.905000 ;
      RECT 9.660000 0.350000  9.990000 1.300000 ;
      RECT 9.660000 1.300000 10.190000 1.630000 ;
      RECT 9.660000 1.630000  9.920000 2.030000 ;
  END
END sky130_fd_sc_ms__dfrtp_2

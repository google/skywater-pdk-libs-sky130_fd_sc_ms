* NGSPICE file created from sky130_fd_sc_ms__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=6.722e+11p ps=3.36e+06u
M1001 a_165_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=7.616e+11p ps=5.84e+06u
M1002 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.32e+11p ps=3.19e+06u
M1003 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1004 Y A2 a_165_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


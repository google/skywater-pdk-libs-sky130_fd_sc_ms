* File: sky130_fd_sc_ms__nor4b_1.pex.spice
* Created: Wed Sep  2 12:16:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR4B_1%D_N 3 7 9 12
c37 12 0 1.706e-19 $X=0.61 $Y=1.275
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.275
+ $X2=0.61 $Y2=1.44
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.275
+ $X2=0.61 $Y2=1.11
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.275 $X2=0.61 $Y2=1.275
r41 9 13 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.275
+ $X2=0.61 $Y2=1.275
r42 7 14 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.67 $Y=0.645
+ $X2=0.67 $Y2=1.11
r43 3 15 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=0.655 $Y=2.26
+ $X2=0.655 $Y2=1.44
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%A 3 7 9 12 13
c37 13 0 2.22943e-19 $X=1.15 $Y=1.515
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.515
+ $X2=1.15 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.515
+ $X2=1.15 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.515 $X2=1.15 $Y2=1.515
r41 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.515
r42 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.24 $Y=0.74 $X2=1.24
+ $Y2=1.35
r43 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.225 $Y=2.4
+ $X2=1.225 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%B 3 7 9 12 13
c38 3 0 1.20528e-19 $X=1.645 $Y=2.4
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.69 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.515
+ $X2=1.69 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.515 $X2=1.69 $Y2=1.515
r42 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=1.515
r43 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.67 $Y=0.74 $X2=1.67
+ $Y2=1.35
r44 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.645 $Y=2.4
+ $X2=1.645 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%C 3 7 9 12 13
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.515
+ $X2=2.23 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.515
+ $X2=2.23 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.515 $X2=2.23 $Y2=1.515
r42 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.22 $Y2=1.515
r43 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.25 $Y=0.74 $X2=2.25
+ $Y2=1.35
r44 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.155 $Y=2.4
+ $X2=2.155 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%A_57_368# 1 2 9 13 19 22 26 29 30 31 35 36
r77 36 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.515
+ $X2=2.77 $Y2=1.68
r78 36 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.515
+ $X2=2.77 $Y2=1.35
r79 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.515 $X2=2.77 $Y2=1.515
r80 32 35 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.65 $Y=1.515
+ $X2=2.77 $Y2=1.515
r81 29 31 1.22049 $w=4.88e-07 $l=5e-08 $layer=LI1_cond $X=0.35 $Y=1.985 $X2=0.35
+ $Y2=2.035
r82 29 30 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.35 $Y=1.985
+ $X2=0.35 $Y2=1.82
r83 23 26 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=0.19 $Y=0.645
+ $X2=0.455 $Y2=0.645
r84 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=1.68
+ $X2=2.65 $Y2=1.515
r85 21 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.65 $Y=1.68 $X2=2.65
+ $Y2=1.95
r86 20 31 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.595 $Y=2.035
+ $X2=0.35 $Y2=2.035
r87 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=2.65 $Y2=1.95
r88 19 20 128.524 $w=1.68e-07 $l=1.97e-06 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=0.595 $Y2=2.035
r89 15 23 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.19 $Y=0.94
+ $X2=0.19 $Y2=0.645
r90 15 30 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.19 $Y=0.94
+ $X2=0.19 $Y2=1.82
r91 13 40 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.725 $Y=2.4
+ $X2=2.725 $Y2=1.68
r92 9 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.68 $Y=0.74 $X2=2.68
+ $Y2=1.35
r93 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=1.84 $X2=0.43 $Y2=1.985
r94 1 26 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.37 $X2=0.455 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%VPWR 1 6 9 10 11 21 22
r26 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r27 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r28 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r29 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r30 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 11 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 9 14 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33 $X2=1
+ $Y2=3.33
r35 8 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=3.33 $X2=1
+ $Y2=3.33
r37 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=3.33
r38 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1 $Y=3.245 $X2=1
+ $Y2=2.455
r39 1 6 300 $w=1.7e-07 $l=7.31471e-07 $layer=licon1_PDIFF $count=2 $X=0.745
+ $Y=1.84 $X2=1 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%Y 1 2 3 12 14 15 18 20 24 25 26 27 43
c61 15 0 6.81849e-20 $X=1.62 $Y=1.095
r62 26 27 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=2.405
+ $X2=3.09 $Y2=2.775
r63 25 43 7.82243 $w=3.68e-07 $l=1.42e-07 $layer=LI1_cond $X=3.09 $Y=1.992
+ $X2=3.09 $Y2=1.85
r64 25 26 10.2163 $w=3.68e-07 $l=3.28e-07 $layer=LI1_cond $X=3.09 $Y=2.077
+ $X2=3.09 $Y2=2.405
r65 22 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=1.18
+ $X2=3.19 $Y2=1.85
r66 21 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.095
+ $X2=2.465 $Y2=1.095
r67 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=1.095
+ $X2=3.19 $Y2=1.18
r68 20 21 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.105 $Y=1.095
+ $X2=2.63 $Y2=1.095
r69 16 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.01
+ $X2=2.465 $Y2=1.095
r70 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.465 $Y=1.01
+ $X2=2.465 $Y2=0.515
r71 14 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=1.095
+ $X2=2.465 $Y2=1.095
r72 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.3 $Y=1.095
+ $X2=1.62 $Y2=1.095
r73 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.455 $Y=1.01
+ $X2=1.62 $Y2=1.095
r74 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.455 $Y=1.01
+ $X2=1.455 $Y2=0.515
r75 3 25 400 $w=1.7e-07 $l=3.31134e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.84 $X2=3.07 $Y2=2.015
r76 3 27 400 $w=1.7e-07 $l=1.0951e-06 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.84 $X2=3.07 $Y2=2.815
r77 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.37 $X2=2.465 $Y2=0.515
r78 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.315
+ $Y=0.37 $X2=1.455 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4B_1%VGND 1 2 3 12 16 18 20 23 24 26 27 28 37 43
r43 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 40 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r45 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 37 42 4.53027 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.08
+ $Y2=0
r47 37 39 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r48 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 28 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 28 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r51 28 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 26 35 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=1.68
+ $Y2=0
r53 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=1.955
+ $Y2=0
r54 25 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.64
+ $Y2=0
r55 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=1.955
+ $Y2=0
r56 23 31 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.72
+ $Y2=0
r57 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.955
+ $Y2=0
r58 22 35 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.68
+ $Y2=0
r59 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.955
+ $Y2=0
r60 18 42 3.23591 $w=3.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=3.08 $Y2=0
r61 18 20 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=2.965 $Y2=0.595
r62 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0
r63 14 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0.595
r64 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=0.085
+ $X2=0.955 $Y2=0
r65 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.955 $Y=0.085
+ $X2=0.955 $Y2=0.645
r66 3 20 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.37 $X2=2.965 $Y2=0.595
r67 2 16 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.37 $X2=1.955 $Y2=0.595
r68 1 12 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=0.745
+ $Y=0.37 $X2=0.955 $Y2=0.645
.ends


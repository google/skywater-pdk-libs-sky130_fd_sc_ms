* File: sky130_fd_sc_ms__or2_4.spice
* Created: Fri Aug 28 18:06:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or2_4.pex.spice"
.subckt sky130_fd_sc_ms__or2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1008 N_X_M1008_d N_A_83_260#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1008_d N_A_83_260#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_83_260#_M1012_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13505 AS=0.1036 PD=1.105 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1012_d N_A_83_260#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13505 AS=0.1295 PD=1.105 PS=1.09 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_83_260#_M1004_d N_A_M1004_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12395 AS=0.1295 PD=1.075 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g N_A_83_260#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.9287 AS=0.12395 PD=3.99 PS=1.075 NRD=0 NRS=8.916 M=1 R=4.93333 SA=75002.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_83_260#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1002 N_X_M1001_d N_A_83_260#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1003 N_X_M1003_d N_A_83_260#_M1003_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1003_d N_A_83_260#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.205298 PD=1.39 PS=1.55849 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1005 N_A_496_388#_M1005_d N_A_M1005_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.183302 PD=1.27 PS=1.39151 NRD=0 NRS=15.7403 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_83_260#_M1007_d N_B_M1007_g N_A_496_388#_M1005_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.5
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1010 N_A_83_260#_M1007_d N_B_M1010_g N_A_496_388#_M1010_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90003
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_A_496_388#_M1010_s N_A_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.305 PD=1.32 PS=2.61 NRD=0 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__or2_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o31a_2.spice
* Created: Wed Sep  2 12:25:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o31a_2.pex.spice"
.subckt sky130_fd_sc_ms__o31a_2  VNB VPB A1 A2 A3 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_55_264#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_55_264#_M1006_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_328_74#_M1010_d N_A1_M1010_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.12765 AS=0.1554 PD=1.085 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.3
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_328_74#_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.12765 PD=1.16 PS=1.085 NRD=5.664 NRS=10.536 M=1 R=4.93333
+ SA=75001.8 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1008 N_A_328_74#_M1008_d N_A3_M1008_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.18315 AS=0.1554 PD=1.235 PS=1.16 NRD=17.016 NRS=17.016 M=1 R=4.93333
+ SA=75002.3 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1003 N_A_55_264#_M1003_d N_B1_M1003_g N_A_328_74#_M1008_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.18315 PD=2.19 PS=1.235 NRD=11.34 NRS=17.832 M=1
+ R=4.93333 SA=75003 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1004_d N_A_55_264#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.182 AS=0.3136 PD=1.445 PS=2.8 NRD=3.5066 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1004_d N_A_55_264#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.182 AS=0.261509 PD=1.445 PS=1.67472 NRD=4.3931 NRS=15.8191 M=1 R=6.22222
+ SA=90000.7 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1007 A_349_392# N_A1_M1007_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.233491 PD=1.24 PS=1.49528 NRD=12.7853 NRS=18.715 M=1 R=5.55556 SA=90001.3
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1009 A_433_392# N_A2_M1009_g A_349_392# VPB PSHORT L=0.18 W=1 AD=0.195 AS=0.12
+ PD=1.39 PS=1.24 NRD=27.5603 NRS=12.7853 M=1 R=5.55556 SA=90001.8 SB=90001.4
+ A=0.18 P=2.36 MULT=1
MM1000 N_A_55_264#_M1000_d N_A3_M1000_g A_433_392# VPB PSHORT L=0.18 W=1 AD=0.18
+ AS=0.195 PD=1.36 PS=1.39 NRD=10.8153 NRS=27.5603 M=1 R=5.55556 SA=90002.3
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_55_264#_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.43 AS=0.18 PD=2.86 PS=1.36 NRD=28.5453 NRS=4.9053 M=1 R=5.55556
+ SA=90002.9 SB=90000.3 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o31a_2.pxi.spice"
*
.ends
*
*

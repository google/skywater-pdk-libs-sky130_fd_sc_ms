* File: sky130_fd_sc_ms__dfrbp_1.spice
* Created: Wed Sep  2 12:02:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfrbp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfrbp_1  VNB VPB D CLK RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1010 A_125_78# N_D_M1010_g N_A_38_78#_M1010_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_RESET_B_M1029_g A_125_78# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1281 AS=0.0504 PD=1.45 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_CLK_M1011_g N_A_307_387#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13745 AS=0.245475 PD=1.115 PS=2.15 NRD=7.296 NRS=7.296 M=1
+ R=4.93333 SA=75000.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1012 N_A_501_387#_M1012_d N_A_307_387#_M1012_g N_VGND_M1011_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2262 AS=0.13745 PD=2.14 PS=1.115 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_709_463#_M1018_d N_A_307_387#_M1018_g N_A_38_78#_M1018_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1017 A_832_119# N_A_501_387#_M1017_g N_A_709_463#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1001 A_910_119# N_A_841_401#_M1001_g A_832_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_RESET_B_M1019_g A_910_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.127288 AS=0.0504 PD=1.01038 PS=0.66 NRD=70.872 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1002 N_A_841_401#_M1002_d N_A_709_463#_M1002_g N_VGND_M1019_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1611 AS=0.193962 PD=1.22 PS=1.53962 NRD=15.936 NRS=15.936
+ M=1 R=4.26667 SA=75001.5 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_1224_74#_M1003_d N_A_501_387#_M1003_g N_A_841_401#_M1002_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.261434 AS=0.1611 PD=1.85962 PS=1.22 NRD=81.552 NRS=15.936
+ M=1 R=4.26667 SA=75002 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1000 A_1434_74# N_A_307_387#_M1000_g N_A_1224_74#_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.171566 PD=0.66 PS=1.22038 NRD=18.564 NRS=52.848 M=1
+ R=2.8 SA=75002.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1482_48#_M1022_g A_1434_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0861 AS=0.0504 PD=0.83 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1026 A_1624_74# N_RESET_B_M1026_g N_VGND_M1022_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0861 PD=0.66 PS=0.83 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_A_1482_48#_M1027_d N_A_1224_74#_M1027_g A_1624_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_Q_N_M1015_d N_A_1224_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_1224_74#_M1013_g N_A_2026_424#_M1013_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.104351 AS=0.15675 PD=0.929457 PS=1.67 NRD=13.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1004 N_Q_M1004_d N_A_2026_424#_M1004_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.140399 PD=2.05 PS=1.25054 NRD=0 NRS=1.62 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_38_78#_M1023_d N_D_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_RESET_B_M1024_g N_A_38_78#_M1023_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0567 PD=1.4 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.6
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_307_387#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3361 PD=1.39 PS=2.92 NRD=0 NRS=13.1793 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_A_501_387#_M1014_d N_A_307_387#_M1014_g N_VPWR_M1006_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1005 N_A_709_463#_M1005_d N_A_501_387#_M1005_g N_A_38_78#_M1005_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1009 A_799_463# N_A_307_387#_M1009_g N_A_709_463#_M1005_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1028 N_VPWR_M1028_d N_A_841_401#_M1028_g A_799_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.133675 AS=0.0441 PD=1.125 PS=0.63 NRD=123.48 NRS=23.443 M=1 R=2.33333
+ SA=90001 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1031 N_A_709_463#_M1031_d N_RESET_B_M1031_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.133675 PD=1.37 PS=1.125 NRD=0 NRS=123.48 M=1 R=2.33333
+ SA=90001.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1016 N_A_841_401#_M1016_d N_A_709_463#_M1016_g N_VPWR_M1016_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1020 N_A_1224_74#_M1020_d N_A_307_387#_M1020_g N_A_841_401#_M1016_d VPB PSHORT
+ L=0.18 W=1 AD=0.258028 AS=0.135 PD=2.21127 PS=1.27 NRD=23.6203 NRS=0 M=1
+ R=5.55556 SA=90000.6 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1033 A_1468_471# N_A_501_387#_M1033_g N_A_1224_74#_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.108372 PD=0.66 PS=0.928732 NRD=30.4759 NRS=60.9715 M=1
+ R=2.33333 SA=90001.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_1482_48#_M1007_g A_1468_471# VPB PSHORT L=0.18 W=0.42
+ AD=0.0693 AS=0.0504 PD=0.75 PS=0.66 NRD=9.3772 NRS=30.4759 M=1 R=2.33333
+ SA=90001.7 SB=90002 A=0.0756 P=1.2 MULT=1
MM1021 N_A_1482_48#_M1021_d N_RESET_B_M1021_g N_VPWR_M1007_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.0693 PD=0.69 PS=0.75 NRD=0 NRS=14.0658 M=1 R=2.33333
+ SA=90002.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1025 N_VPWR_M1025_d N_A_1224_74#_M1025_g N_A_1482_48#_M1021_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.0880091 AS=0.0567 PD=0.793636 PS=0.69 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90002.6 SB=90001 A=0.0756 P=1.2 MULT=1
MM1008 N_Q_N_M1008_d N_A_1224_74#_M1008_g N_VPWR_M1025_d VPB PSHORT L=0.18
+ W=1.12 AD=0.672 AS=0.234691 PD=3.44 PS=2.11636 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.3 SB=90000.5 A=0.2016 P=2.6 MULT=1
MM1030 N_VPWR_M1030_d N_A_1224_74#_M1030_g N_A_2026_424#_M1030_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1518 AS=0.2352 PD=1.24714 PS=2.24 NRD=7.0329 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1032 N_Q_M1032_d N_A_2026_424#_M1032_g N_VPWR_M1030_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2024 PD=2.8 PS=1.66286 NRD=0 NRS=2.6201 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=22.2347 P=27.92
c_121 VNB 0 1.61434e-19 $X=0 $Y=0
c_235 VPB 0 1.13494e-19 $X=0 $Y=3.085
c_1726 A_1468_471# 0 1.03385e-19 $X=7.34 $Y=2.355
*
.include "sky130_fd_sc_ms__dfrbp_1.pxi.spice"
*
.ends
*
*

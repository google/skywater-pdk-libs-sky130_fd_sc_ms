* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_8 A VGND VNB VPB VPWR X
X0 X a_128_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 X a_128_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VGND a_128_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 X a_128_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 X a_128_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 X a_128_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VPWR A a_128_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 X a_128_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 VGND A a_128_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 X a_128_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 VGND a_128_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 VPWR a_128_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 VGND a_128_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 VPWR a_128_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_128_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 VGND a_128_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 VPWR a_128_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 X a_128_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_128_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 VPWR a_128_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__and3b_4.pex.spice
* Created: Fri Aug 28 17:13:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND3B_4%A_N 3 7 9 13
c33 9 0 1.93105e-19 $X=0.72 $Y=1.295
r34 13 15 27.563 $w=3.41e-07 $l=1.95e-07 $layer=POLY_cond $X=0.67 $Y=1.39
+ $X2=0.865 $Y2=1.39
r35 11 13 24.7361 $w=3.41e-07 $l=1.75e-07 $layer=POLY_cond $X=0.495 $Y=1.39
+ $X2=0.67 $Y2=1.39
r36 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.345 $X2=0.67 $Y2=1.345
r37 5 15 17.6972 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.865 $Y=1.6
+ $X2=0.865 $Y2=1.39
r38 5 7 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=0.865 $Y=1.6 $X2=0.865
+ $Y2=2.34
r39 1 11 22.0049 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=1.39
r40 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%A_27_74# 1 2 9 13 17 21 25 28 29 30 33 37 39
+ 40 42 48
c88 48 0 1.93105e-19 $X=1.865 $Y=1.485
c89 21 0 4.59863e-20 $X=1.985 $Y=0.81
r90 47 48 48.513 $w=3.08e-07 $l=3.1e-07 $layer=POLY_cond $X=1.555 $Y=1.485
+ $X2=1.865 $Y2=1.485
r91 46 47 21.9091 $w=3.08e-07 $l=1.4e-07 $layer=POLY_cond $X=1.415 $Y=1.485
+ $X2=1.555 $Y2=1.485
r92 43 46 8.60714 $w=3.08e-07 $l=5.5e-08 $layer=POLY_cond $X=1.36 $Y=1.485
+ $X2=1.415 $Y2=1.485
r93 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.36
+ $Y=1.485 $X2=1.36 $Y2=1.485
r94 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.765
+ $X2=0.64 $Y2=1.765
r95 37 42 11.1634 $w=3.06e-07 $l=3.64692e-07 $layer=LI1_cond $X=1.135 $Y=1.765
+ $X2=1.33 $Y2=1.485
r96 37 38 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.135 $Y=1.765
+ $X2=0.805 $Y2=1.765
r97 33 35 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.64 $Y=1.985
+ $X2=0.64 $Y2=2.695
r98 31 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=1.85 $X2=0.64
+ $Y2=1.765
r99 31 33 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.64 $Y=1.85
+ $X2=0.64 $Y2=1.985
r100 29 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=1.765
+ $X2=0.64 $Y2=1.765
r101 29 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.475 $Y=1.765
+ $X2=0.285 $Y2=1.765
r102 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.68
+ $X2=0.285 $Y2=1.765
r103 28 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.2 $Y=1.68 $X2=0.2
+ $Y2=1.01
r104 23 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.845
+ $X2=0.28 $Y2=1.01
r105 23 25 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=0.845
+ $X2=0.28 $Y2=0.495
r106 19 48 18.7792 $w=3.08e-07 $l=2.16852e-07 $layer=POLY_cond $X=1.985 $Y=1.32
+ $X2=1.865 $Y2=1.485
r107 19 21 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.985 $Y=1.32
+ $X2=1.985 $Y2=0.81
r108 15 48 15.3289 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.65
+ $X2=1.865 $Y2=1.485
r109 15 17 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.865 $Y=1.65
+ $X2=1.865 $Y2=2.34
r110 11 47 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.555 $Y=1.32
+ $X2=1.555 $Y2=1.485
r111 11 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.555 $Y=1.32
+ $X2=1.555 $Y2=0.81
r112 7 46 15.3289 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.65
+ $X2=1.415 $Y2=1.485
r113 7 9 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.415 $Y=1.65
+ $X2=1.415 $Y2=2.34
r114 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.495
+ $Y=1.84 $X2=0.64 $Y2=2.695
r115 2 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.495
+ $Y=1.84 $X2=0.64 $Y2=1.985
r116 1 25 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%B 3 7 11 15 17 18 25
c56 15 0 7.05897e-20 $X=2.915 $Y=0.81
c57 7 0 1.67143e-19 $X=2.415 $Y=0.81
c58 3 0 8.49494e-20 $X=2.415 $Y=2.34
r59 25 26 7.53125 $w=3.2e-07 $l=5e-08 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=2.915 $Y2=1.515
r60 23 25 56.4844 $w=3.2e-07 $l=3.75e-07 $layer=POLY_cond $X=2.49 $Y=1.515
+ $X2=2.865 $Y2=1.515
r61 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.515 $X2=2.49 $Y2=1.515
r62 21 23 11.2969 $w=3.2e-07 $l=7.5e-08 $layer=POLY_cond $X=2.415 $Y=1.515
+ $X2=2.49 $Y2=1.515
r63 18 24 4.02015 $w=4.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.49 $Y2=1.565
r64 17 24 8.84433 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.49 $Y2=1.565
r65 13 26 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=1.515
r66 13 15 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=0.81
r67 9 25 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.68
+ $X2=2.865 $Y2=1.515
r68 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.865 $Y=1.68
+ $X2=2.865 $Y2=2.34
r69 5 21 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.515
r70 5 7 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=0.81
r71 1 21 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.68
+ $X2=2.415 $Y2=1.515
r72 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.415 $Y=1.68
+ $X2=2.415 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%C 3 5 7 10 12 14 16 17 21 26
c58 10 0 9.02718e-20 $X=3.925 $Y=2.34
c59 5 0 1.44963e-19 $X=3.905 $Y=1.205
r60 25 26 38.8612 $w=4.75e-07 $l=9e-08 $layer=POLY_cond $X=3.925 $Y=1.442
+ $X2=4.015 $Y2=1.442
r61 20 23 9.3668 $w=4.75e-07 $l=8e-08 $layer=POLY_cond $X=3.395 $Y=1.442
+ $X2=3.475 $Y2=1.442
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.395
+ $Y=1.515 $X2=3.395 $Y2=1.515
r63 17 21 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.395 $Y2=1.565
r64 14 16 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.335 $Y=1.205
+ $X2=4.335 $Y2=0.79
r65 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.26 $Y=1.28
+ $X2=4.335 $Y2=1.205
r66 12 26 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=4.26 $Y=1.28
+ $X2=4.015 $Y2=1.28
r67 8 25 25.6061 $w=1.8e-07 $l=2.38e-07 $layer=POLY_cond $X=3.925 $Y=1.68
+ $X2=3.925 $Y2=1.442
r68 8 10 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.925 $Y=1.68
+ $X2=3.925 $Y2=2.34
r69 5 25 2.3417 $w=4.75e-07 $l=2e-08 $layer=POLY_cond $X=3.905 $Y=1.442
+ $X2=3.925 $Y2=1.442
r70 5 23 50.3466 $w=4.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.905 $Y=1.442
+ $X2=3.475 $Y2=1.442
r71 5 7 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=3.905 $Y=1.205
+ $X2=3.905 $Y2=0.79
r72 1 23 25.6061 $w=1.8e-07 $l=2.38e-07 $layer=POLY_cond $X=3.475 $Y=1.68
+ $X2=3.475 $Y2=1.442
r73 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.475 $Y=1.68
+ $X2=3.475 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%A_301_368# 1 2 3 4 13 15 16 17 20 22 24 27
+ 29 31 34 36 38 41 45 49 53 57 59 63 66 68 71 74 78 79 82 84 86 87 95
c175 79 0 1.28172e-19 $X=1.67 $Y=1.82
c176 78 0 8.49494e-20 $X=1.64 $Y=1.985
c177 41 0 1.61033e-19 $X=6.225 $Y=0.74
c178 20 0 1.64454e-19 $X=4.845 $Y=0.74
r179 94 95 20.0327 $w=3.97e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.522
+ $X2=5.96 $Y2=1.522
r180 91 92 20.0327 $w=3.97e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.522
+ $X2=5.51 $Y2=1.522
r181 90 91 46.7431 $w=3.97e-07 $l=3.85e-07 $layer=POLY_cond $X=4.96 $Y=1.522
+ $X2=5.345 $Y2=1.522
r182 80 81 2.81784 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.035
+ $X2=1.67 $Y2=2.12
r183 79 82 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.78 $Y=1.82
+ $X2=1.78 $Y2=1.15
r184 78 80 1.47749 $w=3.88e-07 $l=5e-08 $layer=LI1_cond $X=1.67 $Y=1.985
+ $X2=1.67 $Y2=2.035
r185 78 79 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=1.985
+ $X2=1.67 $Y2=1.82
r186 75 94 23.6751 $w=3.97e-07 $l=1.95e-07 $layer=POLY_cond $X=5.6 $Y=1.522
+ $X2=5.795 $Y2=1.522
r187 75 92 10.927 $w=3.97e-07 $l=9e-08 $layer=POLY_cond $X=5.6 $Y=1.522 $X2=5.51
+ $Y2=1.522
r188 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=1.465 $X2=5.6 $Y2=1.465
r189 72 90 4.85642 $w=3.97e-07 $l=4e-08 $layer=POLY_cond $X=4.92 $Y=1.522
+ $X2=4.96 $Y2=1.522
r190 72 88 9.10579 $w=3.97e-07 $l=7.5e-08 $layer=POLY_cond $X=4.92 $Y=1.522
+ $X2=4.845 $Y2=1.522
r191 71 87 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=1.465
+ $X2=4.755 $Y2=1.465
r192 71 74 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.92 $Y=1.465
+ $X2=5.6 $Y2=1.465
r193 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.92
+ $Y=1.465 $X2=4.92 $Y2=1.465
r194 68 87 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.9 $Y=1.545
+ $X2=4.755 $Y2=1.545
r195 66 86 3.49088 $w=2.67e-07 $l=1.33918e-07 $layer=LI1_cond $X=3.815 $Y=1.95
+ $X2=3.717 $Y2=2.035
r196 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=1.63
+ $X2=3.9 $Y2=1.545
r197 65 66 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.815 $Y=1.63
+ $X2=3.815 $Y2=1.95
r198 61 86 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=3.717 $Y=2.12
+ $X2=3.717 $Y2=2.035
r199 61 63 18.7864 $w=3.63e-07 $l=5.95e-07 $layer=LI1_cond $X=3.717 $Y=2.12
+ $X2=3.717 $Y2=2.715
r200 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.035
+ $X2=2.64 $Y2=2.035
r201 59 86 3.01551 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.535 $Y=2.035
+ $X2=3.717 $Y2=2.035
r202 59 60 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.535 $Y=2.035
+ $X2=2.805 $Y2=2.035
r203 55 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=2.12
+ $X2=2.64 $Y2=2.035
r204 55 57 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.64 $Y=2.12
+ $X2=2.64 $Y2=2.715
r205 54 80 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.865 $Y=2.035
+ $X2=1.67 $Y2=2.035
r206 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=2.035
+ $X2=2.64 $Y2=2.035
r207 53 54 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.475 $Y=2.035
+ $X2=1.865 $Y2=2.035
r208 47 82 5.59224 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=1.775 $Y=1.06
+ $X2=1.775 $Y2=1.15
r209 47 49 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=1.775 $Y=1.06
+ $X2=1.775 $Y2=0.87
r210 45 81 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.64 $Y=2.695
+ $X2=1.64 $Y2=2.12
r211 39 95 32.1738 $w=3.97e-07 $l=3.59242e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=5.96 $Y2=1.522
r212 39 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=6.225 $Y2=0.74
r213 36 95 21.283 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=5.96 $Y=1.745
+ $X2=5.96 $Y2=1.522
r214 36 38 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=5.96 $Y=1.745
+ $X2=5.96 $Y2=2.4
r215 32 94 25.678 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.795 $Y=1.3
+ $X2=5.795 $Y2=1.522
r216 32 34 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.795 $Y=1.3
+ $X2=5.795 $Y2=0.74
r217 29 92 21.283 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=5.51 $Y=1.745
+ $X2=5.51 $Y2=1.522
r218 29 31 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=5.51 $Y=1.745
+ $X2=5.51 $Y2=2.4
r219 25 91 25.678 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.345 $Y=1.3
+ $X2=5.345 $Y2=1.522
r220 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.345 $Y=1.3
+ $X2=5.345 $Y2=0.74
r221 22 90 21.283 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=4.96 $Y=1.745
+ $X2=4.96 $Y2=1.522
r222 22 24 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=4.96 $Y=1.745
+ $X2=4.96 $Y2=2.4
r223 18 88 25.678 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.845 $Y=1.3
+ $X2=4.845 $Y2=1.522
r224 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.845 $Y=1.3
+ $X2=4.845 $Y2=0.74
r225 16 88 30.4212 $w=3.97e-07 $l=1.87681e-07 $layer=POLY_cond $X=4.755 $Y=1.67
+ $X2=4.845 $Y2=1.522
r226 16 17 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.755 $Y=1.67
+ $X2=4.6 $Y2=1.67
r227 13 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.51 $Y=1.745
+ $X2=4.6 $Y2=1.67
r228 13 15 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=4.51 $Y=1.745
+ $X2=4.51 $Y2=2.4
r229 4 86 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.84 $X2=3.7 $Y2=2.035
r230 4 63 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.84 $X2=3.7 $Y2=2.715
r231 3 84 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.84 $X2=2.64 $Y2=2.035
r232 3 57 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.84 $X2=2.64 $Y2=2.715
r233 2 78 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.84 $X2=1.64 $Y2=1.985
r234 2 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.84 $X2=1.64 $Y2=2.695
r235 1 49 182 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.49 $X2=1.77 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 41 45 48 49
+ 51 52 53 55 60 65 78 79 82 85 88 91
r96 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r100 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r102 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r104 73 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 70 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.235 $Y2=3.33
r107 70 72 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.4 $Y=3.33 $X2=5.04
+ $Y2=3.33
r108 69 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 66 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.14 $Y2=3.33
r112 66 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 65 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=3.14 $Y2=3.33
r114 65 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 64 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 61 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.14 $Y2=3.33
r119 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 60 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=2.14 $Y2=3.33
r121 60 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 58 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 55 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.14 $Y2=3.33
r125 55 57 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 53 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 53 89 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 51 75 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.07 $Y=3.33 $X2=6
+ $Y2=3.33
r129 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=6.235 $Y2=3.33
r130 50 78 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.4 $Y=3.33 $X2=6.48
+ $Y2=3.33
r131 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.4 $Y=3.33
+ $X2=6.235 $Y2=3.33
r132 48 72 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.07 $Y=3.33 $X2=5.04
+ $Y2=3.33
r133 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=3.33
+ $X2=5.235 $Y2=3.33
r134 47 75 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.4 $Y=3.33 $X2=6
+ $Y2=3.33
r135 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.4 $Y=3.33
+ $X2=5.235 $Y2=3.33
r136 43 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=3.245
+ $X2=6.235 $Y2=3.33
r137 43 45 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=6.235 $Y=3.245
+ $X2=6.235 $Y2=2.25
r138 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=3.245
+ $X2=5.235 $Y2=3.33
r139 39 41 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=5.235 $Y=3.245
+ $X2=5.235 $Y2=2.25
r140 35 38 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.235 $Y=1.985
+ $X2=4.235 $Y2=2.815
r141 33 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.235 $Y=3.245
+ $X2=4.235 $Y2=3.33
r142 33 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.235 $Y=3.245
+ $X2=4.235 $Y2=2.815
r143 32 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.14 $Y2=3.33
r144 31 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=4.235 $Y2=3.33
r145 31 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=3.305 $Y2=3.33
r146 27 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=3.33
r147 27 29 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=2.375
r148 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=3.245
+ $X2=2.14 $Y2=3.33
r149 23 25 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.14 $Y=3.245
+ $X2=2.14 $Y2=2.375
r150 19 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r151 19 21 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.15
r152 6 45 300 $w=1.7e-07 $l=4.93913e-07 $layer=licon1_PDIFF $count=2 $X=6.05
+ $Y=1.84 $X2=6.235 $Y2=2.25
r153 5 41 300 $w=1.7e-07 $l=4.93913e-07 $layer=licon1_PDIFF $count=2 $X=5.05
+ $Y=1.84 $X2=5.235 $Y2=2.25
r154 4 38 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.84 $X2=4.235 $Y2=2.815
r155 4 35 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=4.015
+ $Y=1.84 $X2=4.235 $Y2=1.985
r156 3 29 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.84 $X2=3.14 $Y2=2.375
r157 2 25 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=1.955
+ $Y=1.84 $X2=2.14 $Y2=2.375
r158 1 21 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=0.955
+ $Y=1.84 $X2=1.14 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%X 1 2 3 4 15 19 20 23 25 26 29 35 38 39 41
+ 42 43
c82 42 0 1.61033e-19 $X=6.015 $Y=1.045
c83 20 0 9.02718e-20 $X=4.9 $Y=1.885
r84 43 48 11.0234 $w=2.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.885
r85 40 41 4.30018 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=6.105 $Y=1.885
+ $X2=5.837 $Y2=1.885
r86 39 48 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.365 $Y=1.885
+ $X2=6.48 $Y2=1.885
r87 39 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.365 $Y=1.885
+ $X2=6.105 $Y2=1.885
r88 38 41 1.96316 $w=1.7e-07 $l=2.21459e-07 $layer=LI1_cond $X=6.02 $Y=1.8
+ $X2=5.837 $Y2=1.885
r89 37 42 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.02 $Y=1.13
+ $X2=6.015 $Y2=1.045
r90 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.02 $Y=1.13
+ $X2=6.02 $Y2=1.8
r91 33 42 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=0.96
+ $X2=6.015 $Y2=1.045
r92 33 35 27.4192 $w=1.78e-07 $l=4.45e-07 $layer=LI1_cond $X=6.015 $Y=0.96
+ $X2=6.015 $Y2=0.515
r93 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.735 $Y=1.985
+ $X2=5.735 $Y2=2.815
r94 27 41 1.96316 $w=3.3e-07 $l=1.38109e-07 $layer=LI1_cond $X=5.735 $Y=1.97
+ $X2=5.837 $Y2=1.885
r95 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.735 $Y=1.97
+ $X2=5.735 $Y2=1.985
r96 25 42 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.925 $Y=1.045
+ $X2=6.015 $Y2=1.045
r97 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.925 $Y=1.045
+ $X2=5.215 $Y2=1.045
r98 21 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.09 $Y=0.96
+ $X2=5.215 $Y2=1.045
r99 21 23 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.09 $Y=0.96
+ $X2=5.09 $Y2=0.515
r100 19 41 4.30018 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=5.57 $Y=1.885
+ $X2=5.837 $Y2=1.885
r101 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.57 $Y=1.885
+ $X2=4.9 $Y2=1.885
r102 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.735 $Y=1.985
+ $X2=4.735 $Y2=2.815
r103 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.735 $Y=1.97
+ $X2=4.9 $Y2=1.885
r104 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.735 $Y=1.97
+ $X2=4.735 $Y2=1.985
r105 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.6
+ $Y=1.84 $X2=5.735 $Y2=2.815
r106 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.6
+ $Y=1.84 $X2=5.735 $Y2=1.985
r107 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.84 $X2=4.735 $Y2=2.815
r108 3 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.84 $X2=4.735 $Y2=1.985
r109 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.87
+ $Y=0.37 $X2=6.01 $Y2=0.515
r110 1 23 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.92
+ $Y=0.37 $X2=5.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%VGND 1 2 3 4 5 18 22 26 32 34 36 38 40 45 50
+ 55 60 66 69 72 75 79
c92 79 0 3.3892e-20 $X=6.48 $Y=0
r93 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r97 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r98 64 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r99 64 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r100 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r101 61 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=5.56
+ $Y2=0
r102 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=6
+ $Y2=0
r103 60 78 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.497 $Y2=0
r104 60 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6
+ $Y2=0
r105 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r106 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r107 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r108 56 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.63
+ $Y2=0
r109 56 58 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=5.04
+ $Y2=0
r110 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.56
+ $Y2=0
r111 55 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.04 $Y2=0
r112 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r113 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r114 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r115 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.69
+ $Y2=0
r116 51 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=4.08 $Y2=0
r117 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.63
+ $Y2=0
r118 50 53 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.08 $Y2=0
r119 49 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 46 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.745
+ $Y2=0
r122 46 48 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r123 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.69
+ $Y2=0
r124 45 48 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=3.525 $Y=0
+ $X2=1.2 $Y2=0
r125 43 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r126 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 40 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.745
+ $Y2=0
r128 40 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r129 38 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r130 38 49 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=1.2
+ $Y2=0
r131 34 78 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.497 $Y2=0
r132 34 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.515
r133 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=0.085
+ $X2=5.56 $Y2=0
r134 30 32 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.56 $Y=0.085
+ $X2=5.56 $Y2=0.625
r135 26 28 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.63 $Y=0.515
+ $X2=4.63 $Y2=0.965
r136 24 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0
r137 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0.515
r138 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=0.085
+ $X2=3.69 $Y2=0
r139 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.69 $Y=0.085
+ $X2=3.69 $Y2=0.675
r140 16 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r141 16 18 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.495
r142 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.37 $X2=6.44 $Y2=0.515
r143 4 32 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.42
+ $Y=0.37 $X2=5.56 $Y2=0.625
r144 3 28 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.47 $X2=4.63 $Y2=0.965
r145 3 26 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.47 $X2=4.63 $Y2=0.515
r146 2 22 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.47 $X2=3.69 $Y2=0.675
r147 1 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%A_239_98# 1 2 3 12 14 15 20 22 26
c45 26 0 7.05897e-20 $X=2.2 $Y=0.635
c46 20 0 1.20944e-20 $X=3.13 $Y=0.635
c47 14 0 3.89712e-20 $X=2.035 $Y=0.34
r48 24 26 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.2 $Y=0.595 $X2=2.2
+ $Y2=0.635
r49 22 24 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.2 $Y=0.34 $X2=2.2
+ $Y2=0.595
r50 18 24 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0.595
+ $X2=2.2 $Y2=0.595
r51 18 20 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=2.365 $Y=0.595
+ $X2=3.13 $Y2=0.595
r52 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=2.2 $Y2=0.34
r53 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=1.505 $Y2=0.34
r54 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.505 $Y2=0.34
r55 10 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.34 $Y2=0.635
r56 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.49 $X2=3.13 $Y2=0.635
r57 2 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.49 $X2=2.2 $Y2=0.635
r58 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.195
+ $Y=0.49 $X2=1.34 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_4%A_498_98# 1 2 7 11 14
c30 11 0 3.09417e-19 $X=4.12 $Y=0.615
r31 14 16 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.7 $Y=0.98 $X2=2.7
+ $Y2=1.095
r32 9 11 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=4.16 $Y=1.01
+ $X2=4.16 $Y2=0.615
r33 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=1.095
+ $X2=2.7 $Y2=1.095
r34 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.035 $Y=1.095
+ $X2=4.16 $Y2=1.01
r35 7 8 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.035 $Y=1.095
+ $X2=2.865 $Y2=1.095
r36 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.98
+ $Y=0.47 $X2=4.12 $Y2=0.615
r37 1 14 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.49 $X2=2.7 $Y2=0.98
.ends


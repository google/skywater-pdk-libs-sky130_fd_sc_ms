* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__bufinv_16 A VGND VNB VPB VPWR Y
X0 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X25 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X33 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X34 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X38 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X40 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X41 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X42 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X43 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X44 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X45 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X46 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X47 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X48 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X49 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__a2111oi_4.pex.spice
* Created: Fri Aug 28 16:56:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2111OI_4%D1 3 7 11 13 15 16 18 21 23 24 25 40 41
r69 41 42 2.21779 $w=3.26e-07 $l=1.5e-08 $layer=POLY_cond $X=1.83 $Y=1.385
+ $X2=1.845 $Y2=1.385
r70 39 41 13.3067 $w=3.26e-07 $l=9e-08 $layer=POLY_cond $X=1.74 $Y=1.385
+ $X2=1.83 $Y2=1.385
r71 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.385 $X2=1.74 $Y2=1.385
r72 36 39 50.2699 $w=3.26e-07 $l=3.4e-07 $layer=POLY_cond $X=1.4 $Y=1.385
+ $X2=1.74 $Y2=1.385
r73 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=1.385 $X2=1.4 $Y2=1.385
r74 34 36 0.739264 $w=3.26e-07 $l=5e-09 $layer=POLY_cond $X=1.395 $Y=1.385
+ $X2=1.4 $Y2=1.385
r75 33 34 66.5337 $w=3.26e-07 $l=4.5e-07 $layer=POLY_cond $X=0.945 $Y=1.385
+ $X2=1.395 $Y2=1.385
r76 31 33 33.2669 $w=3.26e-07 $l=2.25e-07 $layer=POLY_cond $X=0.72 $Y=1.385
+ $X2=0.945 $Y2=1.385
r77 29 31 33.2669 $w=3.26e-07 $l=2.25e-07 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.72 $Y2=1.385
r78 25 40 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=1.68 $Y=1.365 $X2=1.74
+ $Y2=1.365
r79 25 37 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.4 $Y2=1.365
r80 24 37 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.365 $X2=1.4
+ $Y2=1.365
r81 23 24 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=1.2 $Y2=1.365
r82 23 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.385 $X2=0.72 $Y2=1.385
r83 19 42 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.55
+ $X2=1.845 $Y2=1.385
r84 19 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.845 $Y=1.55
+ $X2=1.845 $Y2=2.4
r85 16 41 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.22
+ $X2=1.83 $Y2=1.385
r86 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.22 $X2=1.83
+ $Y2=0.74
r87 13 36 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.22 $X2=1.4
+ $Y2=1.385
r88 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.4 $Y=1.22 $X2=1.4
+ $Y2=0.74
r89 9 34 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.55
+ $X2=1.395 $Y2=1.385
r90 9 11 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.395 $Y=1.55
+ $X2=1.395 $Y2=2.4
r91 5 33 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.55
+ $X2=0.945 $Y2=1.385
r92 5 7 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.945 $Y=1.55
+ $X2=0.945 $Y2=2.4
r93 1 29 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=1.385
r94 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%C1 3 5 7 10 14 18 22 24 25 37 38
c77 37 0 2.2789e-19 $X=3.42 $Y=1.515
c78 14 0 1.008e-19 $X=2.745 $Y=2.4
r79 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.42
+ $Y=1.515 $X2=3.42 $Y2=1.515
r80 31 33 37.2747 $w=3.75e-07 $l=2.9e-07 $layer=POLY_cond $X=2.4 $Y=1.545
+ $X2=2.69 $Y2=1.545
r81 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.4
+ $Y=1.515 $X2=2.4 $Y2=1.515
r82 29 31 13.496 $w=3.75e-07 $l=1.05e-07 $layer=POLY_cond $X=2.295 $Y=1.545
+ $X2=2.4 $Y2=1.545
r83 28 29 4.49867 $w=3.75e-07 $l=3.5e-08 $layer=POLY_cond $X=2.26 $Y=1.545
+ $X2=2.295 $Y2=1.545
r84 25 38 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.42
+ $Y2=1.565
r85 24 25 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r86 24 32 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.4 $Y2=1.565
r87 20 37 28.92 $w=3.75e-07 $l=2.25e-07 $layer=POLY_cond $X=3.645 $Y=1.545
+ $X2=3.42 $Y2=1.545
r88 20 22 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=3.645 $Y=1.71
+ $X2=3.645 $Y2=2.4
r89 16 37 28.92 $w=3.75e-07 $l=2.25e-07 $layer=POLY_cond $X=3.195 $Y=1.545
+ $X2=3.42 $Y2=1.545
r90 16 18 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=3.195 $Y=1.71
+ $X2=3.195 $Y2=2.4
r91 12 16 57.84 $w=3.75e-07 $l=4.5e-07 $layer=POLY_cond $X=2.745 $Y=1.545
+ $X2=3.195 $Y2=1.545
r92 12 33 7.06933 $w=3.75e-07 $l=5.5e-08 $layer=POLY_cond $X=2.745 $Y=1.545
+ $X2=2.69 $Y2=1.545
r93 12 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.745 $Y=1.68
+ $X2=2.745 $Y2=2.4
r94 8 33 24.2915 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.69 $Y=1.32
+ $X2=2.69 $Y2=1.545
r95 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.69 $Y=1.32 $X2=2.69
+ $Y2=0.74
r96 5 29 19.9308 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=2.295 $Y=1.77
+ $X2=2.295 $Y2=1.545
r97 5 7 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.295 $Y=1.77 $X2=2.295
+ $Y2=2.4
r98 1 28 24.2915 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.26 $Y=1.32
+ $X2=2.26 $Y2=1.545
r99 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.26 $Y=1.32 $X2=2.26
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%B1 3 7 11 15 19 23 25 26 27 40 41
c70 23 0 1.68901e-19 $X=5.985 $Y=2.4
r71 40 42 11.3323 $w=3.19e-07 $l=7.5e-08 $layer=POLY_cond $X=5.91 $Y=1.515
+ $X2=5.985 $Y2=1.515
r72 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.91
+ $Y=1.515 $X2=5.91 $Y2=1.515
r73 38 40 56.6614 $w=3.19e-07 $l=3.75e-07 $layer=POLY_cond $X=5.535 $Y=1.515
+ $X2=5.91 $Y2=1.515
r74 37 38 67.9937 $w=3.19e-07 $l=4.5e-07 $layer=POLY_cond $X=5.085 $Y=1.515
+ $X2=5.535 $Y2=1.515
r75 36 37 67.9937 $w=3.19e-07 $l=4.5e-07 $layer=POLY_cond $X=4.635 $Y=1.515
+ $X2=5.085 $Y2=1.515
r76 35 36 27.953 $w=3.19e-07 $l=1.85e-07 $layer=POLY_cond $X=4.45 $Y=1.515
+ $X2=4.635 $Y2=1.515
r77 33 35 1.51097 $w=3.19e-07 $l=1e-08 $layer=POLY_cond $X=4.44 $Y=1.515
+ $X2=4.45 $Y2=1.515
r78 33 34 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.44
+ $Y=1.515 $X2=4.44 $Y2=1.515
r79 27 41 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.91 $Y2=1.565
r80 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r81 25 26 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r82 25 34 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.44 $Y2=1.565
r83 21 42 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=1.68
+ $X2=5.985 $Y2=1.515
r84 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.985 $Y=1.68
+ $X2=5.985 $Y2=2.4
r85 17 38 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.68
+ $X2=5.535 $Y2=1.515
r86 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.535 $Y=1.68
+ $X2=5.535 $Y2=2.4
r87 13 37 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.085 $Y=1.68
+ $X2=5.085 $Y2=1.515
r88 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.085 $Y=1.68
+ $X2=5.085 $Y2=2.4
r89 9 36 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.68
+ $X2=4.635 $Y2=1.515
r90 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.635 $Y=1.68
+ $X2=4.635 $Y2=2.4
r91 5 35 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.45 $Y=1.35 $X2=4.45
+ $Y2=1.515
r92 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.45 $Y=1.35 $X2=4.45
+ $Y2=0.74
r93 1 33 63.4608 $w=3.19e-07 $l=4.95681e-07 $layer=POLY_cond $X=4.02 $Y=1.35
+ $X2=4.44 $Y2=1.515
r94 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.02 $Y=1.35 $X2=4.02
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%A1 3 7 11 15 19 23 27 31 33 34 35 53
c81 31 0 1.20142e-20 $X=7.79 $Y=0.74
c82 27 0 1.69181e-19 $X=7.785 $Y=2.4
c83 19 0 1.69181e-19 $X=7.335 $Y=2.4
c84 11 0 1.69181e-19 $X=6.885 $Y=2.4
c85 3 0 1.69181e-19 $X=6.435 $Y=2.4
r86 52 53 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.785 $Y=1.515
+ $X2=7.79 $Y2=1.515
r87 50 52 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.71 $Y=1.515
+ $X2=7.785 $Y2=1.515
r88 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.71
+ $Y=1.515 $X2=7.71 $Y2=1.515
r89 48 50 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=7.36 $Y=1.515
+ $X2=7.71 $Y2=1.515
r90 47 48 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.335 $Y=1.515
+ $X2=7.36 $Y2=1.515
r91 46 47 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=6.93 $Y=1.515
+ $X2=7.335 $Y2=1.515
r92 45 46 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.885 $Y=1.515
+ $X2=6.93 $Y2=1.515
r93 43 45 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.69 $Y=1.515
+ $X2=6.885 $Y2=1.515
r94 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.69
+ $Y=1.515 $X2=6.69 $Y2=1.515
r95 41 43 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=6.5 $Y=1.515
+ $X2=6.69 $Y2=1.515
r96 39 41 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=6.435 $Y=1.515
+ $X2=6.5 $Y2=1.515
r97 35 51 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=7.71 $Y2=1.565
r98 34 51 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.71 $Y2=1.565
r99 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r100 33 44 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.69 $Y2=1.565
r101 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.35
+ $X2=7.79 $Y2=1.515
r102 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.79 $Y=1.35
+ $X2=7.79 $Y2=0.74
r103 25 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.785 $Y=1.68
+ $X2=7.785 $Y2=1.515
r104 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.785 $Y=1.68
+ $X2=7.785 $Y2=2.4
r105 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.36 $Y=1.35
+ $X2=7.36 $Y2=1.515
r106 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.36 $Y=1.35
+ $X2=7.36 $Y2=0.74
r107 17 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.335 $Y=1.68
+ $X2=7.335 $Y2=1.515
r108 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.335 $Y=1.68
+ $X2=7.335 $Y2=2.4
r109 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.93 $Y=1.35
+ $X2=6.93 $Y2=1.515
r110 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.93 $Y=1.35
+ $X2=6.93 $Y2=0.74
r111 9 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.885 $Y=1.68
+ $X2=6.885 $Y2=1.515
r112 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.885 $Y=1.68
+ $X2=6.885 $Y2=2.4
r113 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.5 $Y=1.35 $X2=6.5
+ $Y2=1.515
r114 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.5 $Y=1.35 $X2=6.5
+ $Y2=0.74
r115 1 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.435 $Y=1.68
+ $X2=6.435 $Y2=1.515
r116 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.435 $Y=1.68
+ $X2=6.435 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%A2 3 7 11 15 19 23 27 31 33 34 35 51 53
c75 7 0 1.69181e-19 $X=8.235 $Y=2.4
c76 3 0 2.06049e-19 $X=8.22 $Y=0.74
r77 52 53 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.51 $Y=1.515
+ $X2=9.585 $Y2=1.515
r78 50 52 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=9.39 $Y=1.515
+ $X2=9.51 $Y2=1.515
r79 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.39
+ $Y=1.515 $X2=9.39 $Y2=1.515
r80 48 50 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=9.135 $Y=1.515
+ $X2=9.39 $Y2=1.515
r81 47 48 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=9.08 $Y=1.515
+ $X2=9.135 $Y2=1.515
r82 46 47 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=8.685 $Y=1.515
+ $X2=9.08 $Y2=1.515
r83 45 46 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.65 $Y=1.515
+ $X2=8.685 $Y2=1.515
r84 43 45 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=8.37 $Y=1.515
+ $X2=8.65 $Y2=1.515
r85 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.37
+ $Y=1.515 $X2=8.37 $Y2=1.515
r86 41 43 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.235 $Y=1.515
+ $X2=8.37 $Y2=1.515
r87 39 41 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.22 $Y=1.515
+ $X2=8.235 $Y2=1.515
r88 35 51 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.39
+ $Y2=1.565
r89 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r90 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r91 33 44 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=8.4 $Y=1.565 $X2=8.37
+ $Y2=1.565
r92 29 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.585 $Y=1.68
+ $X2=9.585 $Y2=1.515
r93 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.585 $Y=1.68
+ $X2=9.585 $Y2=2.4
r94 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.51 $Y=1.35
+ $X2=9.51 $Y2=1.515
r95 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.51 $Y=1.35
+ $X2=9.51 $Y2=0.74
r96 21 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.135 $Y=1.68
+ $X2=9.135 $Y2=1.515
r97 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.135 $Y=1.68
+ $X2=9.135 $Y2=2.4
r98 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.08 $Y=1.35
+ $X2=9.08 $Y2=1.515
r99 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.08 $Y=1.35
+ $X2=9.08 $Y2=0.74
r100 13 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.685 $Y=1.68
+ $X2=8.685 $Y2=1.515
r101 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.685 $Y=1.68
+ $X2=8.685 $Y2=2.4
r102 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.65 $Y=1.35
+ $X2=8.65 $Y2=1.515
r103 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.65 $Y=1.35
+ $X2=8.65 $Y2=0.74
r104 5 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=1.68
+ $X2=8.235 $Y2=1.515
r105 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.235 $Y=1.68
+ $X2=8.235 $Y2=2.4
r106 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.22 $Y=1.35
+ $X2=8.22 $Y2=1.515
r107 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.22 $Y=1.35 $X2=8.22
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%A_29_368# 1 2 3 4 5 18 20 21 24 26 28 31
+ 32 36 38 42 46 48
c59 28 0 1.29691e-19 $X=2.07 $Y=2.12
c60 26 0 1.008e-19 $X=1.905 $Y=2.99
r61 39 46 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=2.97 $Y2=2.035
r62 38 48 4.17978 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.705 $Y=2.035
+ $X2=3.87 $Y2=1.97
r63 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.705 $Y=2.035
+ $X2=3.085 $Y2=2.035
r64 34 46 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.12
+ $X2=2.97 $Y2=2.035
r65 34 36 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.97 $Y=2.12
+ $X2=2.97 $Y2=2.57
r66 33 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.035
+ $X2=2.07 $Y2=2.035
r67 32 46 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.855 $Y=2.035
+ $X2=2.97 $Y2=2.035
r68 32 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.855 $Y=2.035
+ $X2=2.235 $Y2=2.035
r69 29 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=2.905 $X2=2.07
+ $Y2=2.815
r70 28 44 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.12 $X2=2.07
+ $Y2=2.035
r71 28 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.07 $Y=2.12
+ $X2=2.07 $Y2=2.815
r72 27 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=2.99
+ $X2=1.17 $Y2=2.99
r73 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=2.07 $Y2=2.905
r74 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=1.255 $Y2=2.99
r75 22 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.99
r76 22 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.225
r77 20 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.17 $Y2=2.99
r78 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.355 $Y2=2.99
r79 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.355 $Y2=2.99
r80 16 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.23 $Y2=2.225
r81 5 48 300 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=2 $X=3.735
+ $Y=1.84 $X2=3.87 $Y2=2.05
r82 4 46 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.835
+ $Y=1.84 $X2=2.97 $Y2=2.035
r83 4 36 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=2.835
+ $Y=1.84 $X2=2.97 $Y2=2.57
r84 3 44 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.035
r85 3 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.815
r86 2 24 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=2.225
r87 1 18 300 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%Y 1 2 3 4 5 6 7 22 23 24 28 30 34 38 40 44
+ 46 50 54 57 59 61 64 67 68 70 74 75 79 84
c125 70 0 4.44094e-20 $X=7.575 $Y=0.95
c126 54 0 1.20142e-20 $X=7.41 $Y=1.022
c127 40 0 9.81988e-20 $X=2.39 $Y=0.925
r128 79 84 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.24 $Y=1.72
+ $X2=0.24 $Y2=1.665
r129 75 79 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.805
+ $X2=0.24 $Y2=1.72
r130 75 84 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=1.65
+ $X2=0.24 $Y2=1.665
r131 74 75 17.7877 $w=2.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.65
r132 70 72 2.51442 $w=3.28e-07 $l=7.2e-08 $layer=LI1_cond $X=7.575 $Y=0.95
+ $X2=7.575 $Y2=1.022
r133 66 68 7.23236 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0.975
+ $X2=6.88 $Y2=0.975
r134 66 67 7.51706 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0.975
+ $X2=6.55 $Y2=0.975
r135 61 62 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.515 $Y=0.925
+ $X2=2.515 $Y2=1.095
r136 56 74 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=1.295
r137 54 72 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=1.022
+ $X2=7.575 $Y2=1.022
r138 54 68 28.4091 $w=2.13e-07 $l=5.3e-07 $layer=LI1_cond $X=7.41 $Y=1.022
+ $X2=6.88 $Y2=1.022
r139 53 64 6.51676 $w=1.87e-07 $l=1.25e-07 $layer=LI1_cond $X=4.32 $Y=1.077
+ $X2=4.195 $Y2=1.077
r140 53 67 120.647 $w=2.03e-07 $l=2.23e-06 $layer=LI1_cond $X=4.32 $Y=1.077
+ $X2=6.55 $Y2=1.077
r141 48 64 0.330231 $w=2.5e-07 $l=1.02e-07 $layer=LI1_cond $X=4.195 $Y=0.975
+ $X2=4.195 $Y2=1.077
r142 48 50 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.195 $Y=0.975
+ $X2=4.195 $Y2=0.515
r143 47 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.095
+ $X2=2.515 $Y2=1.095
r144 46 64 6.51676 $w=1.87e-07 $l=1.33697e-07 $layer=LI1_cond $X=4.07 $Y=1.095
+ $X2=4.195 $Y2=1.077
r145 46 47 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=4.07 $Y=1.095
+ $X2=2.64 $Y2=1.095
r146 42 61 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.84
+ $X2=2.515 $Y2=0.925
r147 42 44 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.515 $Y=0.84
+ $X2=2.515 $Y2=0.515
r148 41 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.925
+ $X2=1.615 $Y2=0.925
r149 40 61 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.39 $Y=0.925
+ $X2=2.515 $Y2=0.925
r150 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.39 $Y=0.925
+ $X2=1.7 $Y2=0.925
r151 36 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.84
+ $X2=1.615 $Y2=0.925
r152 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.615 $Y=0.84
+ $X2=1.615 $Y2=0.495
r153 32 34 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.58 $Y=1.89
+ $X2=1.58 $Y2=1.985
r154 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=1.805
+ $X2=0.72 $Y2=1.805
r155 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.455 $Y=1.805
+ $X2=1.58 $Y2=1.89
r156 30 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.455 $Y=1.805
+ $X2=0.885 $Y2=1.805
r157 26 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.89
+ $X2=0.72 $Y2=1.805
r158 26 28 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.89
+ $X2=0.72 $Y2=1.985
r159 25 75 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.805
+ $X2=0.24 $Y2=1.805
r160 24 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=1.805
+ $X2=0.72 $Y2=1.805
r161 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.555 $Y=1.805
+ $X2=0.355 $Y2=1.805
r162 23 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=0.925
+ $X2=0.24 $Y2=1.01
r163 22 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=0.925
+ $X2=1.615 $Y2=0.925
r164 22 23 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.53 $Y=0.925
+ $X2=0.355 $Y2=0.925
r165 7 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=1.985
r166 6 28 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
r167 5 70 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.435
+ $Y=0.37 $X2=7.575 $Y2=0.95
r168 4 66 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.575
+ $Y=0.37 $X2=6.715 $Y2=0.95
r169 3 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.095
+ $Y=0.37 $X2=4.235 $Y2=0.515
r170 2 61 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.37 $X2=2.475 $Y2=0.965
r171 2 44 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.37 $X2=2.475 $Y2=0.515
r172 1 59 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.925
r173 1 38 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%A_477_368# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
r62 31 33 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=5.76 $Y=2.905 $X2=5.76
+ $Y2=2.405
r63 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=2.99
+ $X2=4.86 $Y2=2.99
r64 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.595 $Y=2.99
+ $X2=5.76 $Y2=2.905
r65 29 30 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.595 $Y=2.99
+ $X2=5.025 $Y2=2.99
r66 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.86 $Y=2.905
+ $X2=4.86 $Y2=2.99
r67 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.86 $Y=2.905 $X2=4.86
+ $Y2=2.405
r68 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=2.99
+ $X2=3.42 $Y2=2.99
r69 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=4.86 $Y2=2.99
r70 23 24 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=3.585 $Y2=2.99
r71 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.905
+ $X2=3.42 $Y2=2.99
r72 19 21 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.42 $Y=2.905
+ $X2=3.42 $Y2=2.42
r73 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.99
+ $X2=3.42 $Y2=2.99
r74 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.255 $Y=2.99
+ $X2=2.685 $Y2=2.99
r75 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.685 $Y2=2.99
r76 13 15 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.56 $Y2=2.455
r77 4 33 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=5.625
+ $Y=1.84 $X2=5.76 $Y2=2.405
r78 3 27 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=4.725
+ $Y=1.84 $X2=4.86 $Y2=2.405
r79 2 21 300 $w=1.7e-07 $l=6.43972e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.84 $X2=3.42 $Y2=2.42
r80 1 15 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.385
+ $Y=1.84 $X2=2.52 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%A_853_368# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 48 50 54 56 58 60 65 69 71 73
c87 48 0 3.38362e-19 $X=8.01 $Y=2.43
c88 42 0 3.38362e-19 $X=7.11 $Y=2.43
c89 36 0 3.38082e-19 $X=6.21 $Y=2.43
r90 58 75 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=9.85 $Y=2.12 $X2=9.85
+ $Y2=1.97
r91 58 60 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=9.85 $Y=2.12
+ $X2=9.85 $Y2=2.4
r92 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=2.035
+ $X2=8.91 $Y2=2.035
r93 56 75 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=9.725 $Y=2.035
+ $X2=9.85 $Y2=1.97
r94 56 57 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.725 $Y=2.035
+ $X2=9.075 $Y2=2.035
r95 52 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=2.12 $X2=8.91
+ $Y2=2.035
r96 52 54 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.91 $Y=2.12
+ $X2=8.91 $Y2=2.815
r97 51 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.095 $Y=2.035
+ $X2=8.01 $Y2=2.035
r98 50 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.91 $Y2=2.035
r99 50 51 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.095 $Y2=2.035
r100 46 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.01 $Y=2.12
+ $X2=8.01 $Y2=2.035
r101 46 48 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.01 $Y=2.12
+ $X2=8.01 $Y2=2.43
r102 45 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=2.035
+ $X2=7.11 $Y2=2.035
r103 44 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.925 $Y=2.035
+ $X2=8.01 $Y2=2.035
r104 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.925 $Y=2.035
+ $X2=7.195 $Y2=2.035
r105 40 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.11 $Y=2.12
+ $X2=7.11 $Y2=2.035
r106 40 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.11 $Y=2.12
+ $X2=7.11 $Y2=2.43
r107 39 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.035
+ $X2=6.21 $Y2=2.035
r108 38 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=2.035
+ $X2=7.11 $Y2=2.035
r109 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.025 $Y=2.035
+ $X2=6.295 $Y2=2.035
r110 34 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=2.12
+ $X2=6.21 $Y2=2.035
r111 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.21 $Y=2.12
+ $X2=6.21 $Y2=2.43
r112 33 65 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.425 $Y=2.035
+ $X2=5.31 $Y2=2.035
r113 32 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=2.035
+ $X2=6.21 $Y2=2.035
r114 32 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.125 $Y=2.035
+ $X2=5.425 $Y2=2.035
r115 28 65 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=2.12
+ $X2=5.31 $Y2=2.035
r116 28 30 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.31 $Y=2.12
+ $X2=5.31 $Y2=2.57
r117 27 63 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.525 $Y=2.035
+ $X2=4.385 $Y2=2.035
r118 26 65 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.195 $Y=2.035
+ $X2=5.31 $Y2=2.035
r119 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.195 $Y=2.035
+ $X2=4.525 $Y2=2.035
r120 22 63 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.385 $Y=2.12
+ $X2=4.385 $Y2=2.035
r121 22 24 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=4.385 $Y=2.12
+ $X2=4.385 $Y2=2.57
r122 7 75 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.675
+ $Y=1.84 $X2=9.81 $Y2=1.985
r123 7 60 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=9.675
+ $Y=1.84 $X2=9.81 $Y2=2.4
r124 6 73 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=8.775
+ $Y=1.84 $X2=8.91 $Y2=2.035
r125 6 54 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.775
+ $Y=1.84 $X2=8.91 $Y2=2.815
r126 5 71 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.84 $X2=8.01 $Y2=2.035
r127 5 48 300 $w=1.7e-07 $l=6.54026e-07 $layer=licon1_PDIFF $count=2 $X=7.875
+ $Y=1.84 $X2=8.01 $Y2=2.43
r128 4 69 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=6.975
+ $Y=1.84 $X2=7.11 $Y2=2.035
r129 4 42 300 $w=1.7e-07 $l=6.54026e-07 $layer=licon1_PDIFF $count=2 $X=6.975
+ $Y=1.84 $X2=7.11 $Y2=2.43
r130 3 67 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=6.075
+ $Y=1.84 $X2=6.21 $Y2=2.035
r131 3 36 300 $w=1.7e-07 $l=6.54026e-07 $layer=licon1_PDIFF $count=2 $X=6.075
+ $Y=1.84 $X2=6.21 $Y2=2.43
r132 2 65 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=5.175
+ $Y=1.84 $X2=5.31 $Y2=2.035
r133 2 30 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=5.175
+ $Y=1.84 $X2=5.31 $Y2=2.57
r134 1 63 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.84 $X2=4.41 $Y2=2.035
r135 1 24 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.84 $X2=4.41 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%VPWR 1 2 3 4 15 17 21 25 29 31 32 33 42 47
+ 54 55 58 61 64
r115 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r117 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 55 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r119 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r120 52 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.525 $Y=3.33
+ $X2=9.4 $Y2=3.33
r121 52 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.525 $Y=3.33
+ $X2=9.84 $Y2=3.33
r122 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r123 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r124 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r125 48 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=3.33
+ $X2=8.42 $Y2=3.33
r126 48 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.545 $Y=3.33
+ $X2=8.88 $Y2=3.33
r127 47 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=9.4 $Y2=3.33
r128 47 50 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=8.88 $Y2=3.33
r129 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r130 46 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r131 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r132 43 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.56 $Y2=3.33
r133 43 45 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 42 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.42 $Y2=3.33
r135 42 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=7.92 $Y2=3.33
r136 41 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r137 40 41 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r138 36 40 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 36 37 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 33 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r141 33 37 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 31 40 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.48 $Y2=3.33
r143 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.66 $Y2=3.33
r144 27 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.4 $Y=3.245
+ $X2=9.4 $Y2=3.33
r145 27 29 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=9.4 $Y=3.245
+ $X2=9.4 $Y2=2.455
r146 23 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=3.33
r147 23 25 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=2.455
r148 19 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=3.245
+ $X2=7.56 $Y2=3.33
r149 19 21 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.56 $Y=3.245
+ $X2=7.56 $Y2=2.375
r150 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.66 $Y2=3.33
r151 17 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=7.56 $Y2=3.33
r152 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=6.825 $Y2=3.33
r153 13 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=3.245
+ $X2=6.66 $Y2=3.33
r154 13 15 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.66 $Y=3.245
+ $X2=6.66 $Y2=2.375
r155 4 29 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=9.225
+ $Y=1.84 $X2=9.36 $Y2=2.455
r156 3 25 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=1.84 $X2=8.46 $Y2=2.455
r157 2 21 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=7.425
+ $Y=1.84 $X2=7.56 $Y2=2.375
r158 1 15 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=1.84 $X2=6.66 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%VGND 1 2 3 4 5 6 21 25 27 31 35 39 42 43
+ 44 46 59 67 74 75 78 82 88 90 93 96
r103 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r104 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r105 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r106 87 88 11.4973 $w=9.23e-07 $l=9.5e-08 $layer=LI1_cond $X=3.805 $Y=0.377
+ $X2=3.9 $Y2=0.377
r107 85 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r108 84 87 2.70378 $w=9.23e-07 $l=2.05e-07 $layer=LI1_cond $X=3.6 $Y=0.377
+ $X2=3.805 $Y2=0.377
r109 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r110 81 84 9.16649 $w=9.23e-07 $l=6.95e-07 $layer=LI1_cond $X=2.905 $Y=0.377
+ $X2=3.6 $Y2=0.377
r111 81 82 11.4973 $w=9.23e-07 $l=9.5e-08 $layer=LI1_cond $X=2.905 $Y=0.377
+ $X2=2.81 $Y2=0.377
r112 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r114 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r115 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.46 $Y=0 $X2=9.295
+ $Y2=0
r116 72 74 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.46 $Y=0 $X2=9.84
+ $Y2=0
r117 71 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r118 71 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r119 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r120 68 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.6 $Y=0 $X2=8.435
+ $Y2=0
r121 68 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.6 $Y=0 $X2=8.88
+ $Y2=0
r122 67 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.13 $Y=0 $X2=9.295
+ $Y2=0
r123 67 70 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=9.13 $Y=0 $X2=8.88
+ $Y2=0
r124 66 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r125 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r126 62 65 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.92
+ $Y2=0
r127 60 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.665
+ $Y2=0
r128 60 62 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.04
+ $Y2=0
r129 59 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.27 $Y=0 $X2=8.435
+ $Y2=0
r130 59 65 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.27 $Y=0 $X2=7.92
+ $Y2=0
r131 58 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r132 57 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.81
+ $Y2=0
r133 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r134 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r135 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r136 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r137 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.185
+ $Y2=0
r138 51 53 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.68
+ $Y2=0
r139 49 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r140 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r141 46 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.185
+ $Y2=0
r142 46 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.72
+ $Y2=0
r143 44 66 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=7.92 $Y2=0
r144 44 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r145 44 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r146 42 53 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.68
+ $Y2=0
r147 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.045
+ $Y2=0
r148 41 57 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.64
+ $Y2=0
r149 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.045
+ $Y2=0
r150 37 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=0.085
+ $X2=9.295 $Y2=0
r151 37 39 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.295 $Y=0.085
+ $X2=9.295 $Y2=0.675
r152 33 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.435 $Y=0.085
+ $X2=8.435 $Y2=0
r153 33 35 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.435 $Y=0.085
+ $X2=8.435 $Y2=0.675
r154 29 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0
r155 29 31 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0.64
r156 27 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.665
+ $Y2=0
r157 27 88 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=3.9
+ $Y2=0
r158 23 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r159 23 25 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.55
r160 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r161 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.55
r162 6 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.37 $X2=9.295 $Y2=0.675
r163 5 35 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.37 $X2=8.435 $Y2=0.675
r164 4 31 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.37 $X2=4.665 $Y2=0.64
r165 3 87 121.333 $w=1.7e-07 $l=1.18271e-06 $layer=licon1_NDIFF $count=1
+ $X=2.765 $Y=0.37 $X2=3.805 $Y2=0.675
r166 3 81 121.333 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1
+ $X=2.765 $Y=0.37 $X2=2.905 $Y2=0.675
r167 2 25 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.37 $X2=2.045 $Y2=0.55
r168 1 21 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.37 $X2=1.185 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__A2111OI_4%A_1228_74# 1 2 3 4 5 18 20 24 25 28 30 34
+ 39 42 43 46
c59 20 0 1.6164e-19 $X=8.005 $Y=0.6
r60 41 43 4.37153 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.145 $Y=0.515
+ $X2=7.25 $Y2=0.515
r61 41 42 4.37153 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.145 $Y=0.515
+ $X2=7.04 $Y2=0.515
r62 39 42 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=6.38 $Y=0.475
+ $X2=7.04 $Y2=0.475
r63 37 39 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.285 $Y=0.515
+ $X2=6.38 $Y2=0.515
r64 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.765 $Y=1.01
+ $X2=9.765 $Y2=0.515
r65 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.95 $Y=1.095
+ $X2=8.865 $Y2=1.095
r66 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.64 $Y=1.095
+ $X2=9.765 $Y2=1.01
r67 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.64 $Y=1.095
+ $X2=8.95 $Y2=1.095
r68 26 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=1.01
+ $X2=8.865 $Y2=1.095
r69 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.865 $Y=1.01
+ $X2=8.865 $Y2=0.515
r70 24 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.78 $Y=1.095
+ $X2=8.865 $Y2=1.095
r71 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.78 $Y=1.095
+ $X2=8.09 $Y2=1.095
r72 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.005 $Y=1.01
+ $X2=8.09 $Y2=1.095
r73 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.005 $Y=1.01
+ $X2=8.005 $Y2=0.965
r74 20 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.005 $Y=0.6
+ $X2=8.005 $Y2=0.475
r75 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.005 $Y=0.6
+ $X2=8.005 $Y2=0.965
r76 18 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=0.475
+ $X2=8.005 $Y2=0.475
r77 18 43 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.92 $Y=0.475
+ $X2=7.25 $Y2=0.475
r78 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.585
+ $Y=0.37 $X2=9.725 $Y2=0.515
r79 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.725
+ $Y=0.37 $X2=8.865 $Y2=0.515
r80 3 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.865
+ $Y=0.37 $X2=8.005 $Y2=0.515
r81 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.865
+ $Y=0.37 $X2=8.005 $Y2=0.965
r82 2 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.005
+ $Y=0.37 $X2=7.145 $Y2=0.515
r83 1 37 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.14
+ $Y=0.37 $X2=6.285 $Y2=0.515
.ends


/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_MS__UDP_DLATCH_P_TB_V
`define SKY130_FD_SC_MS__UDP_DLATCH_P_TB_V

/**
 * udp_dlatch$P: D-latch, gated standard drive / active high
 *               (Q output UDP)
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_ms__udp_dlatch_p.v"

module top();

    // Inputs are registered
    reg D;

    // Outputs are wires
    wire Q;

    initial
    begin
        // Initial state is x for all inputs.
        D = 1'bX;

        #20   D = 1'b0;
        #40   D = 1'b1;
        #60   D = 1'b0;
        #80   D = 1'b1;
        #100  D = 1'bx;
    end

    // Create a clock
    reg GATE;
    initial
    begin
        GATE = 1'b0;
    end

    always
    begin
        #5 GATE = ~GATE;
    end

    sky130_fd_sc_ms__udp_dlatch$P dut (.D(D), .Q(Q), .GATE(GATE));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_MS__UDP_DLATCH_P_TB_V

* File: sky130_fd_sc_ms__dfsbp_1.pxi.spice
* Created: Wed Sep  2 12:03:23 2020
* 
x_PM_SKY130_FD_SC_MS__DFSBP_1%D N_D_c_270_n N_D_M1023_g N_D_M1003_g D D
+ N_D_c_272_n N_D_c_273_n N_D_c_277_n PM_SKY130_FD_SC_MS__DFSBP_1%D
x_PM_SKY130_FD_SC_MS__DFSBP_1%CLK N_CLK_M1032_g N_CLK_M1012_g CLK N_CLK_c_304_n
+ N_CLK_c_305_n PM_SKY130_FD_SC_MS__DFSBP_1%CLK
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_398_74# N_A_398_74#_M1013_d N_A_398_74#_M1019_d
+ N_A_398_74#_c_340_n N_A_398_74#_c_359_n N_A_398_74#_M1009_g
+ N_A_398_74#_M1022_g N_A_398_74#_M1018_g N_A_398_74#_M1005_g
+ N_A_398_74#_c_362_n N_A_398_74#_c_342_n N_A_398_74#_c_363_n
+ N_A_398_74#_c_343_n N_A_398_74#_c_344_n N_A_398_74#_c_364_n
+ N_A_398_74#_c_365_n N_A_398_74#_c_345_n N_A_398_74#_c_346_n
+ N_A_398_74#_c_347_n N_A_398_74#_c_369_n N_A_398_74#_c_370_n
+ N_A_398_74#_c_371_n N_A_398_74#_c_372_n N_A_398_74#_c_373_n
+ N_A_398_74#_c_374_n N_A_398_74#_c_375_n N_A_398_74#_c_376_n
+ N_A_398_74#_c_399_p N_A_398_74#_c_377_n N_A_398_74#_c_378_n
+ N_A_398_74#_c_348_n N_A_398_74#_c_349_n N_A_398_74#_c_350_n
+ N_A_398_74#_c_351_n N_A_398_74#_c_352_n N_A_398_74#_c_380_n
+ N_A_398_74#_c_353_n N_A_398_74#_c_354_n N_A_398_74#_c_381_n
+ N_A_398_74#_c_382_n N_A_398_74#_c_355_n N_A_398_74#_c_356_n
+ N_A_398_74#_c_357_n PM_SKY130_FD_SC_MS__DFSBP_1%A_398_74#
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_779_380# N_A_779_380#_M1015_s
+ N_A_779_380#_M1029_d N_A_779_380#_M1020_g N_A_779_380#_c_631_n
+ N_A_779_380#_M1006_g N_A_779_380#_c_638_n N_A_779_380#_c_639_n
+ N_A_779_380#_c_632_n N_A_779_380#_c_633_n N_A_779_380#_c_640_n
+ N_A_779_380#_c_641_n N_A_779_380#_c_642_n N_A_779_380#_c_634_n
+ N_A_779_380#_c_635_n N_A_779_380#_c_636_n
+ PM_SKY130_FD_SC_MS__DFSBP_1%A_779_380#
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_596_81# N_A_596_81#_M1004_d N_A_596_81#_M1009_d
+ N_A_596_81#_M1029_g N_A_596_81#_c_718_n N_A_596_81#_M1015_g
+ N_A_596_81#_M1001_g N_A_596_81#_M1000_g N_A_596_81#_c_721_n
+ N_A_596_81#_c_722_n N_A_596_81#_c_723_n N_A_596_81#_c_724_n
+ N_A_596_81#_c_725_n N_A_596_81#_c_726_n N_A_596_81#_c_727_n
+ N_A_596_81#_c_728_n N_A_596_81#_c_729_n N_A_596_81#_c_739_n
+ N_A_596_81#_c_730_n N_A_596_81#_c_731_n N_A_596_81#_c_732_n
+ N_A_596_81#_c_733_n N_A_596_81#_c_734_n N_A_596_81#_c_735_n
+ PM_SKY130_FD_SC_MS__DFSBP_1%A_596_81#
x_PM_SKY130_FD_SC_MS__DFSBP_1%SET_B N_SET_B_M1016_g N_SET_B_M1026_g
+ N_SET_B_M1024_g N_SET_B_c_878_n N_SET_B_c_879_n N_SET_B_M1014_g
+ N_SET_B_c_880_n N_SET_B_c_891_n N_SET_B_c_881_n N_SET_B_c_882_n
+ N_SET_B_c_883_n SET_B N_SET_B_c_896_n N_SET_B_c_885_n N_SET_B_c_886_n
+ PM_SKY130_FD_SC_MS__DFSBP_1%SET_B
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_225_74# N_A_225_74#_M1032_s N_A_225_74#_M1012_s
+ N_A_225_74#_M1013_g N_A_225_74#_M1019_g N_A_225_74#_c_1035_n
+ N_A_225_74#_c_1023_n N_A_225_74#_c_1036_n N_A_225_74#_c_1037_n
+ N_A_225_74#_M1004_g N_A_225_74#_M1007_g N_A_225_74#_c_1039_n
+ N_A_225_74#_M1002_g N_A_225_74#_c_1025_n N_A_225_74#_c_1026_n
+ N_A_225_74#_M1031_g N_A_225_74#_c_1028_n N_A_225_74#_c_1029_n
+ N_A_225_74#_c_1030_n N_A_225_74#_c_1046_n N_A_225_74#_c_1031_n
+ N_A_225_74#_c_1048_n N_A_225_74#_c_1049_n N_A_225_74#_c_1050_n
+ N_A_225_74#_c_1032_n N_A_225_74#_c_1033_n N_A_225_74#_c_1052_n
+ PM_SKY130_FD_SC_MS__DFSBP_1%A_225_74#
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_1510_48# N_A_1510_48#_M1011_d
+ N_A_1510_48#_M1017_s N_A_1510_48#_M1028_g N_A_1510_48#_M1010_g
+ N_A_1510_48#_c_1194_n N_A_1510_48#_c_1195_n N_A_1510_48#_c_1196_n
+ N_A_1510_48#_c_1197_n N_A_1510_48#_c_1203_n N_A_1510_48#_c_1198_n
+ N_A_1510_48#_c_1204_n N_A_1510_48#_c_1205_n N_A_1510_48#_c_1199_n
+ N_A_1510_48#_c_1200_n N_A_1510_48#_c_1201_n
+ PM_SKY130_FD_SC_MS__DFSBP_1%A_1510_48#
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_1358_377# N_A_1358_377#_M1018_d
+ N_A_1358_377#_M1002_d N_A_1358_377#_M1014_d N_A_1358_377#_c_1309_n
+ N_A_1358_377#_M1011_g N_A_1358_377#_c_1310_n N_A_1358_377#_c_1311_n
+ N_A_1358_377#_c_1324_n N_A_1358_377#_M1017_g N_A_1358_377#_c_1312_n
+ N_A_1358_377#_M1008_g N_A_1358_377#_M1030_g N_A_1358_377#_c_1314_n
+ N_A_1358_377#_c_1315_n N_A_1358_377#_M1025_g N_A_1358_377#_M1033_g
+ N_A_1358_377#_c_1317_n N_A_1358_377#_c_1318_n N_A_1358_377#_c_1319_n
+ N_A_1358_377#_c_1328_n N_A_1358_377#_c_1341_n N_A_1358_377#_c_1329_n
+ N_A_1358_377#_c_1330_n N_A_1358_377#_c_1320_n N_A_1358_377#_c_1331_n
+ N_A_1358_377#_c_1332_n N_A_1358_377#_c_1333_n N_A_1358_377#_c_1334_n
+ N_A_1358_377#_c_1321_n N_A_1358_377#_c_1335_n N_A_1358_377#_c_1322_n
+ N_A_1358_377#_c_1336_n N_A_1358_377#_c_1337_n N_A_1358_377#_c_1338_n
+ N_A_1358_377#_c_1339_n PM_SKY130_FD_SC_MS__DFSBP_1%A_1358_377#
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_2113_74# N_A_2113_74#_M1025_s
+ N_A_2113_74#_M1033_s N_A_2113_74#_M1027_g N_A_2113_74#_M1021_g
+ N_A_2113_74#_c_1507_n N_A_2113_74#_c_1508_n N_A_2113_74#_c_1509_n
+ N_A_2113_74#_c_1510_n N_A_2113_74#_c_1511_n N_A_2113_74#_c_1512_n
+ N_A_2113_74#_c_1531_n N_A_2113_74#_c_1513_n
+ PM_SKY130_FD_SC_MS__DFSBP_1%A_2113_74#
x_PM_SKY130_FD_SC_MS__DFSBP_1%A_27_80# N_A_27_80#_M1003_s N_A_27_80#_M1004_s
+ N_A_27_80#_M1023_s N_A_27_80#_M1009_s N_A_27_80#_c_1562_n N_A_27_80#_c_1563_n
+ N_A_27_80#_c_1568_n N_A_27_80#_c_1569_n N_A_27_80#_c_1570_n
+ N_A_27_80#_c_1564_n N_A_27_80#_c_1565_n N_A_27_80#_c_1572_n
+ N_A_27_80#_c_1613_n N_A_27_80#_c_1566_n PM_SKY130_FD_SC_MS__DFSBP_1%A_27_80#
x_PM_SKY130_FD_SC_MS__DFSBP_1%VPWR N_VPWR_M1023_d N_VPWR_M1012_d N_VPWR_M1020_d
+ N_VPWR_M1016_d N_VPWR_M1010_d N_VPWR_M1017_d N_VPWR_M1033_d N_VPWR_c_1630_n
+ N_VPWR_c_1631_n N_VPWR_c_1632_n N_VPWR_c_1633_n N_VPWR_c_1634_n
+ N_VPWR_c_1635_n N_VPWR_c_1636_n N_VPWR_c_1637_n N_VPWR_c_1638_n VPWR
+ N_VPWR_c_1639_n N_VPWR_c_1640_n N_VPWR_c_1641_n N_VPWR_c_1642_n
+ N_VPWR_c_1643_n N_VPWR_c_1644_n N_VPWR_c_1645_n N_VPWR_c_1629_n
+ N_VPWR_c_1647_n N_VPWR_c_1648_n N_VPWR_c_1649_n N_VPWR_c_1650_n
+ N_VPWR_c_1651_n N_VPWR_c_1652_n PM_SKY130_FD_SC_MS__DFSBP_1%VPWR
x_PM_SKY130_FD_SC_MS__DFSBP_1%Q_N N_Q_N_M1008_d N_Q_N_M1030_d N_Q_N_c_1769_n Q_N
+ Q_N Q_N Q_N Q_N N_Q_N_c_1771_n Q_N PM_SKY130_FD_SC_MS__DFSBP_1%Q_N
x_PM_SKY130_FD_SC_MS__DFSBP_1%Q N_Q_M1021_d N_Q_M1027_d N_Q_c_1798_n
+ N_Q_c_1799_n Q Q Q Q N_Q_c_1800_n PM_SKY130_FD_SC_MS__DFSBP_1%Q
x_PM_SKY130_FD_SC_MS__DFSBP_1%VGND N_VGND_M1003_d N_VGND_M1032_d N_VGND_M1006_d
+ N_VGND_M1026_d N_VGND_M1024_d N_VGND_M1008_s N_VGND_M1025_d N_VGND_c_1817_n
+ N_VGND_c_1818_n N_VGND_c_1819_n N_VGND_c_1820_n N_VGND_c_1821_n
+ N_VGND_c_1822_n N_VGND_c_1823_n N_VGND_c_1824_n N_VGND_c_1825_n
+ N_VGND_c_1826_n N_VGND_c_1827_n VGND N_VGND_c_1828_n N_VGND_c_1829_n
+ N_VGND_c_1830_n N_VGND_c_1831_n N_VGND_c_1832_n N_VGND_c_1833_n
+ N_VGND_c_1834_n N_VGND_c_1835_n N_VGND_c_1836_n N_VGND_c_1837_n
+ N_VGND_c_1838_n PM_SKY130_FD_SC_MS__DFSBP_1%VGND
cc_1 VNB N_D_c_270_n 0.0419528f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_2 VNB N_D_M1003_g 0.0274789f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_3 VNB N_D_c_272_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_4 VNB N_D_c_273_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_5 VNB N_CLK_M1012_g 0.00393768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB CLK 0.00902946f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_7 VNB N_CLK_c_304_n 0.0323766f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_CLK_c_305_n 0.0199636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_398_74#_c_340_n 0.0171808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.01
cc_10 VNB N_A_398_74#_M1022_g 0.0446757f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_11 VNB N_A_398_74#_c_342_n 0.00892931f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_12 VNB N_A_398_74#_c_343_n 0.0169218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_398_74#_c_344_n 0.00361019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_345_n 0.00319375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_346_n 0.00240575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_347_n 0.0254493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_348_n 0.00221741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_349_n 0.0018239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_350_n 0.00460376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_351_n 0.00217282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_352_n 0.0117768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_353_n 0.004676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_354_n 0.0311252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_355_n 0.00489304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_356_n 0.0220283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_398_74#_c_357_n 0.0177899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_779_380#_c_631_n 0.0184541f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_A_779_380#_c_632_n 0.0192733f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_29 VNB N_A_779_380#_c_633_n 0.011878f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_30 VNB N_A_779_380#_c_634_n 0.0257785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_779_380#_c_635_n 0.0198399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_779_380#_c_636_n 0.0363032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_596_81#_c_718_n 0.00979214f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_A_596_81#_M1015_g 0.031127f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_35 VNB N_A_596_81#_M1001_g 0.0048429f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.855
cc_36 VNB N_A_596_81#_c_721_n 0.00681179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_596_81#_c_722_n 0.00270325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_596_81#_c_723_n 0.0121552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_596_81#_c_724_n 0.00622085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_596_81#_c_725_n 0.0124404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_596_81#_c_726_n 0.00316404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_596_81#_c_727_n 0.00348619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_596_81#_c_728_n 5.61828e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_596_81#_c_729_n 0.0192499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_596_81#_c_730_n 0.00641571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_596_81#_c_731_n 0.00220131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_596_81#_c_732_n 0.00333015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_596_81#_c_733_n 0.0357243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_596_81#_c_734_n 0.0357028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_596_81#_c_735_n 0.0189964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SET_B_M1026_g 0.0548813f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.01
cc_52 VNB N_SET_B_M1024_g 0.0362239f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_53 VNB N_SET_B_c_878_n 0.0174323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_879_n 0.00564647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_880_n 0.00545817f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_56 VNB N_SET_B_c_881_n 0.011778f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_57 VNB N_SET_B_c_882_n 0.00183892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_883_n 9.3748e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_59 VNB SET_B 6.75578e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_60 VNB N_SET_B_c_885_n 0.0380623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_886_n 0.00714345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_225_74#_M1013_g 0.0224618f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_63 VNB N_A_225_74#_c_1023_n 0.0320241f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_64 VNB N_A_225_74#_M1004_g 0.0273819f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_65 VNB N_A_225_74#_c_1025_n 0.00983536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_225_74#_c_1026_n 8.10579e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_225_74#_M1031_g 0.0551903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_225_74#_c_1028_n 0.0129807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_225_74#_c_1029_n 0.0266488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_225_74#_c_1030_n 0.0184718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_225_74#_c_1031_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_225_74#_c_1032_n 0.0030415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_225_74#_c_1033_n 0.0131011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1510_48#_M1028_g 0.0488917f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_75 VNB N_A_1510_48#_c_1194_n 0.0116397f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.175
cc_76 VNB N_A_1510_48#_c_1195_n 0.0163178f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_77 VNB N_A_1510_48#_c_1196_n 0.00463124f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.855
cc_78 VNB N_A_1510_48#_c_1197_n 0.00509151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1510_48#_c_1198_n 0.00694629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1510_48#_c_1199_n 0.00256065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1510_48#_c_1200_n 3.86133e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1510_48#_c_1201_n 0.015955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1358_377#_c_1309_n 0.0201771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1358_377#_c_1310_n 0.0170735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1358_377#_c_1311_n 0.00484113f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.175
cc_86 VNB N_A_1358_377#_c_1312_n 0.022227f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_87 VNB N_A_1358_377#_M1030_g 0.00297705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1358_377#_c_1314_n 0.0770337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1358_377#_c_1315_n 0.072408f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_90 VNB N_A_1358_377#_M1025_g 0.0357041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1358_377#_c_1317_n 0.0350006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1358_377#_c_1318_n 0.0121211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1358_377#_c_1319_n 0.00297161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1358_377#_c_1320_n 0.00561225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1358_377#_c_1321_n 8.84857e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1358_377#_c_1322_n 2.14136e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2113_74#_M1027_g 0.00708251f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_98 VNB N_A_2113_74#_c_1507_n 0.00643367f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.175
cc_99 VNB N_A_2113_74#_c_1508_n 0.00270135f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.855
cc_100 VNB N_A_2113_74#_c_1509_n 8.76539e-19 $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=2.02
cc_101 VNB N_A_2113_74#_c_1510_n 0.00756196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2113_74#_c_1511_n 0.0343004f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.665
cc_103 VNB N_A_2113_74#_c_1512_n 0.00315728f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.855
cc_104 VNB N_A_2113_74#_c_1513_n 0.0226346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_27_80#_c_1562_n 0.0147808f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.175
cc_106 VNB N_A_27_80#_c_1563_n 0.0387846f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.01
cc_107 VNB N_A_27_80#_c_1564_n 0.00707322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_27_80#_c_1565_n 0.00791533f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.855
cc_109 VNB N_A_27_80#_c_1566_n 0.00383527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VPWR_c_1629_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_Q_N_c_1769_n 0.00815532f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_112 VNB Q_N 7.79382e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_113 VNB N_Q_N_c_1771_n 0.0117591f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.02
cc_114 VNB N_Q_c_1798_n 0.0229628f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_115 VNB N_Q_c_1799_n 0.00626527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_Q_c_1800_n 0.0284292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1817_n 0.00901699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1818_n 0.0221343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1819_n 0.00564229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1820_n 0.0168622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1821_n 0.00853376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1822_n 0.0134931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1823_n 0.0101134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1824_n 0.0584454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1825_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1826_n 0.0209428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1827_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1828_n 0.0176596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1829_n 0.0413222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1830_n 0.048518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1831_n 0.034271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1832_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1833_n 0.676277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1834_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1835_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1836_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1837_n 0.0235452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1838_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VPB N_D_c_270_n 0.015511f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_140 VPB N_D_M1023_g 0.0617714f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_141 VPB N_D_c_273_n 0.00196261f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_142 VPB N_D_c_277_n 0.0244074f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_143 VPB N_CLK_M1012_g 0.0238795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_398_74#_c_340_n 0.00445887f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.01
cc_145 VPB N_A_398_74#_c_359_n 0.0199469f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_146 VPB N_A_398_74#_M1009_g 0.0246013f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_147 VPB N_A_398_74#_M1005_g 0.0263939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_398_74#_c_362_n 0.0183712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_398_74#_c_363_n 0.00385362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_398_74#_c_364_n 0.0217985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_398_74#_c_365_n 0.00371777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_398_74#_c_345_n 0.00209213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_398_74#_c_346_n 0.00544086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_398_74#_c_347_n 0.0166802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_398_74#_c_369_n 0.00281843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_398_74#_c_370_n 0.0089583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_398_74#_c_371_n 0.00388407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_398_74#_c_372_n 0.0155543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_398_74#_c_373_n 0.00260538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_398_74#_c_374_n 0.00215642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_398_74#_c_375_n 0.0113219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_398_74#_c_376_n 2.69913e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_398_74#_c_377_n 0.00637994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_398_74#_c_378_n 0.001186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_398_74#_c_349_n 0.00188182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_398_74#_c_380_n 9.12633e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_398_74#_c_381_n 0.00136728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_398_74#_c_382_n 0.039862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_398_74#_c_355_n 0.00507103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_398_74#_c_356_n 0.0145112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_779_380#_M1020_g 0.031113f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_172 VPB N_A_779_380#_c_638_n 0.0103536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_779_380#_c_639_n 0.0124085f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.175
cc_174 VPB N_A_779_380#_c_640_n 0.00923854f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_175 VPB N_A_779_380#_c_641_n 0.0341146f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_176 VPB N_A_779_380#_c_642_n 0.0036882f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_177 VPB N_A_779_380#_c_635_n 0.00636452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_596_81#_M1029_g 0.0449782f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_179 VPB N_A_596_81#_M1001_g 0.0233844f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.855
cc_180 VPB N_A_596_81#_c_721_n 0.0104002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_596_81#_c_739_n 0.00428261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_596_81#_c_730_n 0.00877385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_SET_B_M1016_g 0.0339288f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.02
cc_184 VPB N_SET_B_M1026_g 0.00278972f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.01
cc_185 VPB N_SET_B_M1014_g 0.0312145f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_186 VPB N_SET_B_c_880_n 0.0284959f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_187 VPB N_SET_B_c_891_n 0.0109698f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.02
cc_188 VPB N_SET_B_c_881_n 0.0176752f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_189 VPB N_SET_B_c_882_n 2.44984e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_SET_B_c_883_n 0.00209073f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_191 VPB SET_B 0.00142743f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_192 VPB N_SET_B_c_896_n 0.0400956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_SET_B_c_886_n 0.00347893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_225_74#_M1019_g 0.0197043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_225_74#_c_1035_n 0.0764525f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_196 VPB N_A_225_74#_c_1036_n 0.0600669f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.855
cc_197 VPB N_A_225_74#_c_1037_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_198 VPB N_A_225_74#_M1007_g 0.0350428f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_199 VPB N_A_225_74#_c_1039_n 0.236256f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_200 VPB N_A_225_74#_M1002_g 0.0193517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_225_74#_c_1025_n 0.0345476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_225_74#_c_1026_n 0.00758117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_225_74#_c_1028_n 7.74435e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_225_74#_c_1029_n 6.04301e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_225_74#_c_1030_n 0.00575231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_225_74#_c_1046_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_225_74#_c_1031_n 0.00240536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_225_74#_c_1048_n 0.0058961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_225_74#_c_1049_n 0.00519182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_225_74#_c_1050_n 0.00478803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_225_74#_c_1032_n 5.21083e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_225_74#_c_1052_n 7.70291e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1510_48#_M1010_g 0.0439167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1510_48#_c_1203_n 0.00685613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1510_48#_c_1204_n 3.23859e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1510_48#_c_1205_n 0.00468539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1510_48#_c_1199_n 0.00736865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1510_48#_c_1201_n 0.0304329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1358_377#_c_1311_n 0.0321219f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_220 VPB N_A_1358_377#_c_1324_n 0.0390121f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_221 VPB N_A_1358_377#_M1017_g 0.0308105f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.855
cc_222 VPB N_A_1358_377#_M1030_g 0.0269849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1358_377#_c_1319_n 0.00782321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1358_377#_c_1328_n 0.0325474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1358_377#_c_1329_n 0.003873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1358_377#_c_1330_n 0.00216924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1358_377#_c_1331_n 0.00538322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1358_377#_c_1332_n 0.00740771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1358_377#_c_1333_n 0.0192277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1358_377#_c_1334_n 0.00300004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1358_377#_c_1335_n 0.004488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1358_377#_c_1336_n 0.00109081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1358_377#_c_1337_n 0.00443161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1358_377#_c_1338_n 0.00401758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1358_377#_c_1339_n 0.0107693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2113_74#_M1027_g 0.0301333f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.61
cc_237 VPB N_A_2113_74#_c_1509_n 0.00968455f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.02
cc_238 VPB N_A_27_80#_c_1563_n 0.0249205f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.01
cc_239 VPB N_A_27_80#_c_1568_n 0.0275048f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.855
cc_240 VPB N_A_27_80#_c_1569_n 0.0259099f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.175
cc_241 VPB N_A_27_80#_c_1570_n 0.0151539f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_242 VPB N_A_27_80#_c_1564_n 0.00269752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_27_80#_c_1572_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1630_n 0.0138484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1631_n 0.00646119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1632_n 0.00583599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1633_n 0.00935928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1634_n 0.00802866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1635_n 0.00396654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1636_n 0.0118539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1637_n 0.0566956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1638_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1639_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1640_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1641_n 0.0500512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1642_n 0.029515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1643_n 0.0366076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1644_n 0.0325425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1645_n 0.0193106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1629_n 0.131094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1647_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1648_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1649_n 0.00523428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1650_n 0.00450185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1651_n 0.0063829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1652_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB Q_N 0.019404f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_268 VPB Q 0.0520162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_Q_c_1800_n 0.00750446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 N_D_c_270_n N_CLK_M1012_g 0.00427113f $X=0.61 $Y=1.825 $X2=0 $Y2=0
cc_271 N_D_c_270_n N_CLK_c_304_n 0.00572583f $X=0.61 $Y=1.825 $X2=0 $Y2=0
cc_272 N_D_c_272_n N_CLK_c_305_n 0.00207613f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_273 N_D_c_272_n N_A_225_74#_c_1031_n 0.00683059f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_274 N_D_c_273_n N_A_225_74#_c_1031_n 0.0532484f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_275 N_D_c_270_n N_A_225_74#_c_1049_n 0.00330843f $X=0.61 $Y=1.825 $X2=0 $Y2=0
cc_276 N_D_c_273_n N_A_225_74#_c_1049_n 0.0249554f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_277 N_D_M1003_g N_A_225_74#_c_1033_n 0.00630877f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_278 N_D_M1003_g N_A_27_80#_c_1562_n 0.00146243f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_279 N_D_M1003_g N_A_27_80#_c_1563_n 0.00600966f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_280 N_D_c_272_n N_A_27_80#_c_1563_n 0.0309478f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_281 N_D_c_273_n N_A_27_80#_c_1563_n 0.0697394f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_282 N_D_M1023_g N_A_27_80#_c_1568_n 0.0085308f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_283 N_D_M1023_g N_A_27_80#_c_1569_n 0.0217614f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_284 N_D_c_273_n N_A_27_80#_c_1569_n 0.0257673f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_285 N_D_c_277_n N_A_27_80#_c_1569_n 0.00145366f $X=0.64 $Y=1.855 $X2=0 $Y2=0
cc_286 N_D_M1023_g N_VPWR_c_1630_n 0.0135295f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_287 N_D_M1023_g N_VPWR_c_1639_n 0.00460063f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_288 N_D_M1023_g N_VPWR_c_1629_n 0.00912296f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_289 N_D_M1003_g N_VGND_c_1817_n 0.0138986f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_290 N_D_c_272_n N_VGND_c_1817_n 0.00175174f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_291 N_D_c_273_n N_VGND_c_1817_n 0.0220022f $X=0.64 $Y=1.175 $X2=0 $Y2=0
cc_292 N_D_M1003_g N_VGND_c_1828_n 0.00462012f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_293 N_D_M1003_g N_VGND_c_1833_n 0.00450456f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_294 CLK N_A_225_74#_M1013_g 0.00486292f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_295 N_CLK_c_304_n N_A_225_74#_M1013_g 0.014451f $X=1.465 $Y=1.385 $X2=0 $Y2=0
cc_296 N_CLK_c_305_n N_A_225_74#_M1013_g 0.0131347f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_297 N_CLK_M1012_g N_A_225_74#_c_1028_n 0.0524692f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_298 CLK N_A_225_74#_c_1028_n 9.33251e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_299 N_CLK_c_304_n N_A_225_74#_c_1028_n 0.00536051f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_300 N_CLK_M1012_g N_A_225_74#_c_1031_n 0.00354737f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_301 CLK N_A_225_74#_c_1031_n 0.0287772f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_302 N_CLK_c_304_n N_A_225_74#_c_1031_n 0.00297156f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_303 N_CLK_c_305_n N_A_225_74#_c_1031_n 0.00324692f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_304 N_CLK_c_304_n N_A_225_74#_c_1048_n 0.00313913f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_305 N_CLK_M1012_g N_A_225_74#_c_1050_n 0.009076f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_306 N_CLK_c_304_n N_A_225_74#_c_1050_n 5.60514e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_307 N_CLK_M1012_g N_A_225_74#_c_1032_n 8.01803e-19 $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_308 CLK N_A_225_74#_c_1032_n 0.0162663f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_309 CLK N_A_225_74#_c_1033_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_310 N_CLK_c_304_n N_A_225_74#_c_1033_n 0.00114511f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_311 N_CLK_c_305_n N_A_225_74#_c_1033_n 0.00765617f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_312 N_CLK_M1012_g N_A_225_74#_c_1052_n 0.00508679f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_313 CLK N_A_225_74#_c_1052_n 0.0368425f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_314 N_CLK_M1012_g N_A_27_80#_c_1569_n 0.0177479f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_315 N_CLK_M1012_g N_VPWR_c_1630_n 0.0116791f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_316 N_CLK_M1012_g N_VPWR_c_1631_n 0.0252424f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_317 N_CLK_M1012_g N_VPWR_c_1640_n 0.00540231f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_318 N_CLK_M1012_g N_VPWR_c_1629_n 0.00533457f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_319 N_CLK_c_305_n N_VGND_c_1817_n 0.00303096f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_320 N_CLK_c_305_n N_VGND_c_1818_n 0.00434272f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_321 CLK N_VGND_c_1819_n 0.0154902f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_322 N_CLK_c_305_n N_VGND_c_1819_n 0.00300619f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_323 N_CLK_c_305_n N_VGND_c_1833_n 0.00825157f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_324 N_A_398_74#_c_362_n N_A_779_380#_M1020_g 9.85524e-19 $X=3.03 $Y=2.105
+ $X2=0 $Y2=0
cc_325 N_A_398_74#_c_346_n N_A_779_380#_M1020_g 0.0068878f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_326 N_A_398_74#_c_369_n N_A_779_380#_M1020_g 0.00256901f $X=3.79 $Y=2.905
+ $X2=0 $Y2=0
cc_327 N_A_398_74#_c_370_n N_A_779_380#_M1020_g 0.0147373f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_328 N_A_398_74#_c_371_n N_A_779_380#_M1020_g 0.0034107f $X=4.695 $Y=2.905
+ $X2=0 $Y2=0
cc_329 N_A_398_74#_c_380_n N_A_779_380#_M1020_g 0.00467226f $X=3.825 $Y=2.25
+ $X2=0 $Y2=0
cc_330 N_A_398_74#_M1022_g N_A_779_380#_c_631_n 0.0419504f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_331 N_A_398_74#_c_370_n N_A_779_380#_c_638_n 0.0127912f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_332 N_A_398_74#_c_359_n N_A_779_380#_c_639_n 9.85524e-19 $X=3.03 $Y=1.94
+ $X2=0 $Y2=0
cc_333 N_A_398_74#_c_346_n N_A_779_380#_c_639_n 0.00757587f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_347_n N_A_779_380#_c_639_n 0.0066563f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_335 N_A_398_74#_c_347_n N_A_779_380#_c_633_n 5.49495e-19 $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_c_346_n N_A_779_380#_c_640_n 0.0117362f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_337 N_A_398_74#_c_370_n N_A_779_380#_c_640_n 0.0424712f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_338 N_A_398_74#_c_399_p N_A_779_380#_c_640_n 0.00122328f $X=5.95 $Y=2.125
+ $X2=0 $Y2=0
cc_339 N_A_398_74#_c_346_n N_A_779_380#_c_641_n 0.00274395f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_340 N_A_398_74#_c_370_n N_A_779_380#_c_642_n 0.0130883f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_341 N_A_398_74#_c_372_n N_A_779_380#_c_642_n 0.0168754f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_342 N_A_398_74#_c_374_n N_A_779_380#_c_642_n 0.0318347f $X=5.455 $Y=2.905
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_c_376_n N_A_779_380#_c_642_n 0.0139478f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_344 N_A_398_74#_c_399_p N_A_779_380#_c_642_n 0.00362126f $X=5.95 $Y=2.125
+ $X2=0 $Y2=0
cc_345 N_A_398_74#_c_346_n N_A_779_380#_c_635_n 0.00137731f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_346 N_A_398_74#_c_347_n N_A_779_380#_c_635_n 0.00875274f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_M1022_g N_A_779_380#_c_636_n 0.00279772f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_348 N_A_398_74#_c_343_n N_A_596_81#_M1004_d 2.28826e-19 $X=3.025 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_349 N_A_398_74#_c_352_n N_A_596_81#_M1004_d 0.00589878f $X=3.03 $Y=1.435
+ $X2=-0.19 $Y2=-0.245
cc_350 N_A_398_74#_c_370_n N_A_596_81#_M1029_g 0.00415215f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_351 N_A_398_74#_c_371_n N_A_596_81#_M1029_g 0.0121083f $X=4.695 $Y=2.905
+ $X2=0 $Y2=0
cc_352 N_A_398_74#_c_372_n N_A_596_81#_M1029_g 0.00396457f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_353 N_A_398_74#_c_374_n N_A_596_81#_M1029_g 6.25446e-19 $X=5.455 $Y=2.905
+ $X2=0 $Y2=0
cc_354 N_A_398_74#_c_374_n N_A_596_81#_M1001_g 8.97166e-19 $X=5.455 $Y=2.905
+ $X2=0 $Y2=0
cc_355 N_A_398_74#_c_375_n N_A_596_81#_M1001_g 0.00589206f $X=5.865 $Y=2.21
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_c_399_p N_A_596_81#_M1001_g 0.00879811f $X=5.95 $Y=2.125
+ $X2=0 $Y2=0
cc_357 N_A_398_74#_c_377_n N_A_596_81#_M1001_g 0.0168387f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_358 N_A_398_74#_c_349_n N_A_596_81#_M1001_g 0.00585685f $X=6.52 $Y=1.62 $X2=0
+ $Y2=0
cc_359 N_A_398_74#_M1022_g N_A_596_81#_c_722_n 0.0102403f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_360 N_A_398_74#_c_343_n N_A_596_81#_c_722_n 0.00340526f $X=3.025 $Y=0.34
+ $X2=0 $Y2=0
cc_361 N_A_398_74#_c_352_n N_A_596_81#_c_722_n 0.0344948f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_M1022_g N_A_596_81#_c_723_n 0.0134244f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_363 N_A_398_74#_c_346_n N_A_596_81#_c_723_n 0.012122f $X=3.825 $Y=1.525 $X2=0
+ $Y2=0
cc_364 N_A_398_74#_c_347_n N_A_596_81#_c_723_n 0.00250611f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_365 N_A_398_74#_M1022_g N_A_596_81#_c_724_n 0.00262599f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_366 N_A_398_74#_c_346_n N_A_596_81#_c_724_n 0.00546472f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_367 N_A_398_74#_c_347_n N_A_596_81#_c_724_n 6.63991e-19 $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_368 N_A_398_74#_c_346_n N_A_596_81#_c_726_n 0.0140304f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_369 N_A_398_74#_c_347_n N_A_596_81#_c_726_n 0.00182995f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_370 N_A_398_74#_c_370_n N_A_596_81#_c_726_n 0.00421951f $X=4.61 $Y=2.25 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_c_378_n N_A_596_81#_c_729_n 0.00241845f $X=6.035 $Y=1.705
+ $X2=0 $Y2=0
cc_372 N_A_398_74#_M1009_g N_A_596_81#_c_739_n 3.32291e-19 $X=3.065 $Y=2.525
+ $X2=0 $Y2=0
cc_373 N_A_398_74#_c_364_n N_A_596_81#_c_739_n 0.0232943f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_c_345_n N_A_596_81#_c_739_n 0.00142555f $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_375 N_A_398_74#_c_356_n N_A_596_81#_c_739_n 0.00439492f $X=3.59 $Y=1.525
+ $X2=0 $Y2=0
cc_376 N_A_398_74#_c_359_n N_A_596_81#_c_730_n 0.00688471f $X=3.03 $Y=1.94 $X2=0
+ $Y2=0
cc_377 N_A_398_74#_M1009_g N_A_596_81#_c_730_n 0.00298215f $X=3.065 $Y=2.525
+ $X2=0 $Y2=0
cc_378 N_A_398_74#_M1022_g N_A_596_81#_c_730_n 0.00867403f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_379 N_A_398_74#_c_346_n N_A_596_81#_c_730_n 0.0599451f $X=3.825 $Y=1.525
+ $X2=0 $Y2=0
cc_380 N_A_398_74#_c_352_n N_A_596_81#_c_730_n 0.0778256f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_381 N_A_398_74#_c_380_n N_A_596_81#_c_730_n 0.0129429f $X=3.825 $Y=2.25 $X2=0
+ $Y2=0
cc_382 N_A_398_74#_c_356_n N_A_596_81#_c_730_n 0.0188243f $X=3.59 $Y=1.525 $X2=0
+ $Y2=0
cc_383 N_A_398_74#_M1022_g N_A_596_81#_c_731_n 0.00408316f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_384 N_A_398_74#_c_352_n N_A_596_81#_c_731_n 0.0143574f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_356_n N_A_596_81#_c_731_n 0.0018726f $X=3.59 $Y=1.525 $X2=0
+ $Y2=0
cc_386 N_A_398_74#_c_377_n N_A_596_81#_c_732_n 0.014583f $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_387 N_A_398_74#_c_378_n N_A_596_81#_c_732_n 0.00671279f $X=6.035 $Y=1.705
+ $X2=0 $Y2=0
cc_388 N_A_398_74#_c_353_n N_A_596_81#_c_732_n 0.0267149f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_389 N_A_398_74#_c_354_n N_A_596_81#_c_732_n 3.11291e-19 $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_390 N_A_398_74#_c_377_n N_A_596_81#_c_733_n 0.00140448f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_391 N_A_398_74#_c_378_n N_A_596_81#_c_733_n 6.8465e-19 $X=6.035 $Y=1.705
+ $X2=0 $Y2=0
cc_392 N_A_398_74#_c_353_n N_A_596_81#_c_733_n 0.00226831f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_393 N_A_398_74#_c_354_n N_A_596_81#_c_733_n 0.0174522f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_394 N_A_398_74#_c_348_n N_A_596_81#_c_735_n 0.0078857f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_395 N_A_398_74#_c_351_n N_A_596_81#_c_735_n 0.00154379f $X=6.605 $Y=0.34
+ $X2=0 $Y2=0
cc_396 N_A_398_74#_c_357_n N_A_596_81#_c_735_n 0.0242288f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_c_372_n N_SET_B_M1016_g 0.00146714f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_398 N_A_398_74#_c_374_n N_SET_B_M1016_g 0.0181097f $X=5.455 $Y=2.905 $X2=0
+ $Y2=0
cc_399 N_A_398_74#_c_376_n N_SET_B_M1016_g 0.00825357f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_400 N_A_398_74#_c_399_p N_SET_B_M1016_g 0.00162872f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_401 N_A_398_74#_c_378_n N_SET_B_M1026_g 0.00119672f $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_402 N_A_398_74#_c_350_n N_SET_B_M1024_g 4.68011e-19 $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_403 N_A_398_74#_c_355_n N_SET_B_M1024_g 0.00193116f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_375_n N_SET_B_c_881_n 0.00636507f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_377_n N_SET_B_c_881_n 0.0372227f $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_378_n N_SET_B_c_881_n 0.0130627f $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_407 N_A_398_74#_c_349_n N_SET_B_c_881_n 0.0035869f $X=6.52 $Y=1.62 $X2=0
+ $Y2=0
cc_408 N_A_398_74#_c_353_n N_SET_B_c_881_n 0.0116123f $X=6.715 $Y=1.285 $X2=0
+ $Y2=0
cc_409 N_A_398_74#_c_354_n N_SET_B_c_881_n 0.00369024f $X=6.715 $Y=1.285 $X2=0
+ $Y2=0
cc_410 N_A_398_74#_c_381_n N_SET_B_c_881_n 0.00592462f $X=7.395 $Y=2.185 $X2=0
+ $Y2=0
cc_411 N_A_398_74#_c_382_n N_SET_B_c_881_n 2.64727e-19 $X=7.395 $Y=2.185 $X2=0
+ $Y2=0
cc_412 N_A_398_74#_c_355_n N_SET_B_c_881_n 0.0190815f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_413 N_A_398_74#_c_375_n N_SET_B_c_882_n 6.26369e-19 $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_414 N_A_398_74#_c_376_n N_SET_B_c_882_n 0.00191865f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_415 N_A_398_74#_c_378_n N_SET_B_c_882_n 3.52044e-19 $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_416 N_A_398_74#_c_375_n N_SET_B_c_883_n 0.0111106f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_417 N_A_398_74#_c_376_n N_SET_B_c_883_n 0.0104469f $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_418 N_A_398_74#_c_399_p N_SET_B_c_883_n 0.0120255f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_419 N_A_398_74#_c_378_n N_SET_B_c_883_n 0.0121378f $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_420 N_A_398_74#_c_375_n N_SET_B_c_896_n 0.00106941f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_421 N_A_398_74#_c_376_n N_SET_B_c_896_n 3.95737e-19 $X=5.54 $Y=2.21 $X2=0
+ $Y2=0
cc_422 N_A_398_74#_c_399_p N_SET_B_c_896_n 0.00131261f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_423 N_A_398_74#_c_342_n N_A_225_74#_M1013_g 0.00167653f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_424 N_A_398_74#_c_344_n N_A_225_74#_M1013_g 0.00266901f $X=2.295 $Y=0.34
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_365_n N_A_225_74#_M1019_g 0.00132039f $X=2.355 $Y=2.99
+ $X2=0 $Y2=0
cc_426 N_A_398_74#_c_359_n N_A_225_74#_c_1035_n 0.0130852f $X=3.03 $Y=1.94 $X2=0
+ $Y2=0
cc_427 N_A_398_74#_M1009_g N_A_225_74#_c_1035_n 0.0150675f $X=3.065 $Y=2.525
+ $X2=0 $Y2=0
cc_428 N_A_398_74#_c_363_n N_A_225_74#_c_1035_n 0.00725312f $X=2.19 $Y=2.565
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_c_364_n N_A_225_74#_c_1035_n 0.0116763f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_430 N_A_398_74#_c_345_n N_A_225_74#_c_1035_n 3.43168e-19 $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_431 N_A_398_74#_c_340_n N_A_225_74#_c_1023_n 0.00655065f $X=3.03 $Y=1.69
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_345_n N_A_225_74#_c_1023_n 8.57179e-19 $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_433 N_A_398_74#_M1009_g N_A_225_74#_c_1036_n 0.0105864f $X=3.065 $Y=2.525
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_c_364_n N_A_225_74#_c_1036_n 0.0142547f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_M1022_g N_A_225_74#_M1004_g 0.00834991f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_436 N_A_398_74#_c_342_n N_A_225_74#_M1004_g 0.00333039f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_437 N_A_398_74#_c_343_n N_A_225_74#_M1004_g 0.0158823f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_438 N_A_398_74#_c_352_n N_A_225_74#_M1004_g 0.00854965f $X=3.03 $Y=1.435
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_M1009_g N_A_225_74#_M1007_g 0.0109316f $X=3.065 $Y=2.525
+ $X2=0 $Y2=0
cc_440 N_A_398_74#_c_364_n N_A_225_74#_M1007_g 0.017774f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_441 N_A_398_74#_c_369_n N_A_225_74#_M1007_g 0.00617239f $X=3.79 $Y=2.905
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_380_n N_A_225_74#_M1007_g 0.00108428f $X=3.825 $Y=2.25
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_356_n N_A_225_74#_M1007_g 0.00563181f $X=3.59 $Y=1.525
+ $X2=0 $Y2=0
cc_444 N_A_398_74#_c_364_n N_A_225_74#_c_1039_n 0.00458792f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_372_n N_A_225_74#_c_1039_n 0.012039f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_446 N_A_398_74#_c_373_n N_A_225_74#_c_1039_n 0.00420304f $X=4.78 $Y=2.99
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_M1005_g N_A_225_74#_M1002_g 0.00608287f $X=7.51 $Y=2.75 $X2=0
+ $Y2=0
cc_448 N_A_398_74#_c_382_n N_A_225_74#_M1002_g 0.00408928f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_c_355_n N_A_225_74#_M1002_g 2.41977e-19 $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_381_n N_A_225_74#_c_1025_n 6.10091e-19 $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_382_n N_A_225_74#_c_1025_n 0.00534578f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_377_n N_A_225_74#_c_1026_n 0.00154931f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_353_n N_A_225_74#_c_1026_n 0.00134708f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_354_n N_A_225_74#_c_1026_n 0.0195395f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_349_n N_A_225_74#_M1031_g 7.76595e-19 $X=6.52 $Y=1.62 $X2=0
+ $Y2=0
cc_456 N_A_398_74#_c_350_n N_A_225_74#_M1031_g 0.0120073f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_457 N_A_398_74#_c_353_n N_A_225_74#_M1031_g 3.48236e-19 $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_458 N_A_398_74#_c_354_n N_A_225_74#_M1031_g 0.0149282f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_355_n N_A_225_74#_M1031_g 0.0115834f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_460 N_A_398_74#_c_357_n N_A_225_74#_M1031_g 0.0215718f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_461 N_A_398_74#_c_340_n N_A_225_74#_c_1029_n 0.0130852f $X=3.03 $Y=1.69 $X2=0
+ $Y2=0
cc_462 N_A_398_74#_c_342_n N_A_225_74#_c_1029_n 9.09054e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_343_n N_A_225_74#_c_1029_n 0.0034994f $X=3.025 $Y=0.34
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_345_n N_A_225_74#_c_1029_n 3.43168e-19 $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_465 N_A_398_74#_c_352_n N_A_225_74#_c_1029_n 7.05733e-19 $X=3.03 $Y=1.435
+ $X2=0 $Y2=0
cc_466 N_A_398_74#_c_342_n N_A_225_74#_c_1030_n 0.00168761f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_M1019_d N_A_225_74#_c_1050_n 0.00285614f $X=2.055 $Y=1.79
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_342_n N_A_225_74#_c_1032_n 0.0218452f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_c_350_n N_A_1510_48#_M1028_g 0.00449224f $X=7.39 $Y=0.34
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_355_n N_A_1510_48#_M1028_g 0.0218033f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_381_n N_A_1510_48#_M1010_g 4.62583e-19 $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_472 N_A_398_74#_c_382_n N_A_1510_48#_M1010_g 0.0549699f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_c_355_n N_A_1510_48#_M1010_g 0.00323148f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_474 N_A_398_74#_c_355_n N_A_1510_48#_c_1194_n 0.0541231f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_c_355_n N_A_1510_48#_c_1196_n 0.0117101f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_476 N_A_398_74#_c_382_n N_A_1510_48#_c_1201_n 0.00168634f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_477 N_A_398_74#_c_355_n N_A_1510_48#_c_1201_n 0.00609625f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_478 N_A_398_74#_c_350_n N_A_1358_377#_M1018_d 0.00260527f $X=7.39 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_479 N_A_398_74#_M1005_g N_A_1358_377#_c_1341_n 0.00247935f $X=7.51 $Y=2.75
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_381_n N_A_1358_377#_c_1341_n 0.0139926f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_481 N_A_398_74#_c_382_n N_A_1358_377#_c_1341_n 0.00278397f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_482 N_A_398_74#_c_381_n N_A_1358_377#_c_1329_n 0.0260174f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_382_n N_A_1358_377#_c_1329_n 0.00458462f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_484 N_A_398_74#_c_377_n N_A_1358_377#_c_1320_n 0.00151891f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_485 N_A_398_74#_c_348_n N_A_1358_377#_c_1320_n 0.0057326f $X=6.52 $Y=1.12
+ $X2=0 $Y2=0
cc_486 N_A_398_74#_c_349_n N_A_1358_377#_c_1320_n 0.00625163f $X=6.52 $Y=1.62
+ $X2=0 $Y2=0
cc_487 N_A_398_74#_c_353_n N_A_1358_377#_c_1320_n 0.025349f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_488 N_A_398_74#_c_354_n N_A_1358_377#_c_1320_n 0.00103124f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_489 N_A_398_74#_c_355_n N_A_1358_377#_c_1320_n 0.0536421f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_490 N_A_398_74#_c_357_n N_A_1358_377#_c_1320_n 0.00145074f $X=6.715 $Y=1.12
+ $X2=0 $Y2=0
cc_491 N_A_398_74#_c_377_n N_A_1358_377#_c_1335_n 0.00643961f $X=6.435 $Y=1.705
+ $X2=0 $Y2=0
cc_492 N_A_398_74#_c_353_n N_A_1358_377#_c_1335_n 0.0025166f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_493 N_A_398_74#_c_354_n N_A_1358_377#_c_1335_n 2.45275e-19 $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_494 N_A_398_74#_c_381_n N_A_1358_377#_c_1335_n 0.00406811f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_495 N_A_398_74#_c_382_n N_A_1358_377#_c_1335_n 5.29702e-19 $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_496 N_A_398_74#_c_355_n N_A_1358_377#_c_1335_n 0.0199168f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_497 N_A_398_74#_c_350_n N_A_1358_377#_c_1322_n 0.0232966f $X=7.39 $Y=0.34
+ $X2=0 $Y2=0
cc_498 N_A_398_74#_c_353_n N_A_1358_377#_c_1322_n 0.0051699f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_499 N_A_398_74#_c_354_n N_A_1358_377#_c_1322_n 0.00163857f $X=6.715 $Y=1.285
+ $X2=0 $Y2=0
cc_500 N_A_398_74#_c_355_n N_A_1358_377#_c_1322_n 0.0250923f $X=7.395 $Y=2.02
+ $X2=0 $Y2=0
cc_501 N_A_398_74#_c_357_n N_A_1358_377#_c_1322_n 0.0040576f $X=6.715 $Y=1.12
+ $X2=0 $Y2=0
cc_502 N_A_398_74#_M1005_g N_A_1358_377#_c_1336_n 0.0075732f $X=7.51 $Y=2.75
+ $X2=0 $Y2=0
cc_503 N_A_398_74#_M1005_g N_A_1358_377#_c_1337_n 0.0105624f $X=7.51 $Y=2.75
+ $X2=0 $Y2=0
cc_504 N_A_398_74#_c_381_n N_A_1358_377#_c_1338_n 0.0218418f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_505 N_A_398_74#_c_382_n N_A_1358_377#_c_1338_n 0.00671449f $X=7.395 $Y=2.185
+ $X2=0 $Y2=0
cc_506 N_A_398_74#_c_343_n N_A_27_80#_M1004_s 0.00233785f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_507 N_A_398_74#_M1019_d N_A_27_80#_c_1570_n 0.00449575f $X=2.055 $Y=1.79
+ $X2=0 $Y2=0
cc_508 N_A_398_74#_M1009_g N_A_27_80#_c_1570_n 0.00861167f $X=3.065 $Y=2.525
+ $X2=0 $Y2=0
cc_509 N_A_398_74#_c_362_n N_A_27_80#_c_1570_n 0.00113593f $X=3.03 $Y=2.105
+ $X2=0 $Y2=0
cc_510 N_A_398_74#_c_363_n N_A_27_80#_c_1570_n 0.046539f $X=2.19 $Y=2.565 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_364_n N_A_27_80#_c_1570_n 0.038146f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_512 N_A_398_74#_c_345_n N_A_27_80#_c_1570_n 0.0146617f $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_340_n N_A_27_80#_c_1564_n 0.00427076f $X=3.03 $Y=1.69 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_345_n N_A_27_80#_c_1564_n 0.0468227f $X=3.03 $Y=1.6 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_352_n N_A_27_80#_c_1564_n 0.0274015f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_342_n N_A_27_80#_c_1566_n 0.0340448f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_343_n N_A_27_80#_c_1566_n 0.0199805f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_352_n N_A_27_80#_c_1566_n 0.0100954f $X=3.03 $Y=1.435 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_370_n N_VPWR_M1020_d 0.0102694f $X=4.61 $Y=2.25 $X2=0 $Y2=0
cc_520 N_A_398_74#_c_371_n N_VPWR_M1020_d 0.0078004f $X=4.695 $Y=2.905 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_375_n N_VPWR_M1016_d 0.00600933f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_399_p N_VPWR_M1016_d 0.0096722f $X=5.95 $Y=2.125 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_377_n N_VPWR_M1016_d 2.54047e-19 $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_378_n N_VPWR_M1016_d 8.27891e-19 $X=6.035 $Y=1.705 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_365_n N_VPWR_c_1631_n 0.0125862f $X=2.355 $Y=2.99 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_364_n N_VPWR_c_1632_n 0.0152339f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_527 N_A_398_74#_c_369_n N_VPWR_c_1632_n 0.0219177f $X=3.79 $Y=2.905 $X2=0
+ $Y2=0
cc_528 N_A_398_74#_c_370_n N_VPWR_c_1632_n 0.027144f $X=4.61 $Y=2.25 $X2=0 $Y2=0
cc_529 N_A_398_74#_c_371_n N_VPWR_c_1632_n 0.0314631f $X=4.695 $Y=2.905 $X2=0
+ $Y2=0
cc_530 N_A_398_74#_c_373_n N_VPWR_c_1632_n 0.0152343f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_531 N_A_398_74#_c_372_n N_VPWR_c_1633_n 0.0150706f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_532 N_A_398_74#_c_374_n N_VPWR_c_1633_n 0.0242489f $X=5.455 $Y=2.905 $X2=0
+ $Y2=0
cc_533 N_A_398_74#_c_375_n N_VPWR_c_1633_n 0.0280035f $X=5.865 $Y=2.21 $X2=0
+ $Y2=0
cc_534 N_A_398_74#_c_377_n N_VPWR_c_1633_n 3.60079e-19 $X=6.435 $Y=1.705 $X2=0
+ $Y2=0
cc_535 N_A_398_74#_M1005_g N_VPWR_c_1637_n 0.00391275f $X=7.51 $Y=2.75 $X2=0
+ $Y2=0
cc_536 N_A_398_74#_c_364_n N_VPWR_c_1641_n 0.0975191f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_537 N_A_398_74#_c_365_n N_VPWR_c_1641_n 0.0179117f $X=2.355 $Y=2.99 $X2=0
+ $Y2=0
cc_538 N_A_398_74#_c_372_n N_VPWR_c_1642_n 0.0495251f $X=5.37 $Y=2.99 $X2=0
+ $Y2=0
cc_539 N_A_398_74#_c_373_n N_VPWR_c_1642_n 0.0115893f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_540 N_A_398_74#_M1005_g N_VPWR_c_1629_n 0.00499567f $X=7.51 $Y=2.75 $X2=0
+ $Y2=0
cc_541 N_A_398_74#_c_364_n N_VPWR_c_1629_n 0.0511446f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_542 N_A_398_74#_c_365_n N_VPWR_c_1629_n 0.00971754f $X=2.355 $Y=2.99 $X2=0
+ $Y2=0
cc_543 N_A_398_74#_c_372_n N_VPWR_c_1629_n 0.025655f $X=5.37 $Y=2.99 $X2=0 $Y2=0
cc_544 N_A_398_74#_c_373_n N_VPWR_c_1629_n 0.00583135f $X=4.78 $Y=2.99 $X2=0
+ $Y2=0
cc_545 N_A_398_74#_c_369_n A_731_463# 0.00145959f $X=3.79 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_546 N_A_398_74#_c_377_n A_1257_341# 0.00794982f $X=6.435 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_547 N_A_398_74#_c_344_n N_VGND_c_1819_n 0.0110038f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_548 N_A_398_74#_M1022_g N_VGND_c_1820_n 0.00147934f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_549 N_A_398_74#_c_348_n N_VGND_c_1821_n 0.0287935f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_550 N_A_398_74#_c_351_n N_VGND_c_1821_n 0.0106465f $X=6.605 $Y=0.34 $X2=0
+ $Y2=0
cc_551 N_A_398_74#_c_357_n N_VGND_c_1821_n 4.05806e-19 $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_552 N_A_398_74#_M1022_g N_VGND_c_1824_n 0.00527282f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_553 N_A_398_74#_c_343_n N_VGND_c_1824_n 0.0591538f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_554 N_A_398_74#_c_344_n N_VGND_c_1824_n 0.0179217f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_555 N_A_398_74#_c_350_n N_VGND_c_1830_n 0.0617884f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_556 N_A_398_74#_c_351_n N_VGND_c_1830_n 0.0121867f $X=6.605 $Y=0.34 $X2=0
+ $Y2=0
cc_557 N_A_398_74#_c_357_n N_VGND_c_1830_n 0.00278271f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_558 N_A_398_74#_M1022_g N_VGND_c_1833_n 0.00534666f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_559 N_A_398_74#_c_343_n N_VGND_c_1833_n 0.0340476f $X=3.025 $Y=0.34 $X2=0
+ $Y2=0
cc_560 N_A_398_74#_c_344_n N_VGND_c_1833_n 0.00971942f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_561 N_A_398_74#_c_350_n N_VGND_c_1833_n 0.0347045f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_562 N_A_398_74#_c_351_n N_VGND_c_1833_n 0.00660921f $X=6.605 $Y=0.34 $X2=0
+ $Y2=0
cc_563 N_A_398_74#_c_357_n N_VGND_c_1833_n 0.0035485f $X=6.715 $Y=1.12 $X2=0
+ $Y2=0
cc_564 N_A_398_74#_c_350_n N_VGND_c_1837_n 0.00587652f $X=7.39 $Y=0.34 $X2=0
+ $Y2=0
cc_565 N_A_398_74#_c_355_n N_VGND_c_1837_n 0.00763101f $X=7.395 $Y=2.02 $X2=0
+ $Y2=0
cc_566 N_A_398_74#_c_348_n A_1262_74# 0.00897986f $X=6.52 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_567 N_A_398_74#_c_351_n A_1262_74# 6.58104e-19 $X=6.605 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_568 N_A_398_74#_c_350_n A_1462_74# 8.39422e-19 $X=7.39 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_569 N_A_398_74#_c_355_n A_1462_74# 0.0034631f $X=7.395 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_570 N_A_779_380#_c_640_n N_A_596_81#_M1029_g 0.0174114f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_571 N_A_779_380#_c_641_n N_A_596_81#_M1029_g 0.0139263f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_572 N_A_779_380#_c_642_n N_A_596_81#_M1029_g 0.0163642f $X=5.115 $Y=2.515
+ $X2=0 $Y2=0
cc_573 N_A_779_380#_c_634_n N_A_596_81#_M1015_g 0.0153755f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_574 N_A_779_380#_c_636_n N_A_596_81#_M1015_g 0.00296272f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_575 N_A_779_380#_c_640_n N_A_596_81#_c_721_n 0.0036927f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_576 N_A_779_380#_c_634_n N_A_596_81#_c_721_n 7.42232e-19 $X=5.015 $Y=0.6
+ $X2=0 $Y2=0
cc_577 N_A_779_380#_c_635_n N_A_596_81#_c_721_n 0.0139263f $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_578 N_A_779_380#_c_631_n N_A_596_81#_c_722_n 0.00177919f $X=4.055 $Y=0.935
+ $X2=0 $Y2=0
cc_579 N_A_779_380#_c_631_n N_A_596_81#_c_723_n 0.0077045f $X=4.055 $Y=0.935
+ $X2=0 $Y2=0
cc_580 N_A_779_380#_c_632_n N_A_596_81#_c_723_n 0.00578861f $X=4.41 $Y=1.01
+ $X2=0 $Y2=0
cc_581 N_A_779_380#_c_633_n N_A_596_81#_c_723_n 0.00761441f $X=4.13 $Y=1.01
+ $X2=0 $Y2=0
cc_582 N_A_779_380#_c_634_n N_A_596_81#_c_723_n 0.0140413f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_583 N_A_779_380#_c_632_n N_A_596_81#_c_724_n 0.00406612f $X=4.41 $Y=1.01
+ $X2=0 $Y2=0
cc_584 N_A_779_380#_c_633_n N_A_596_81#_c_724_n 8.23249e-19 $X=4.13 $Y=1.01
+ $X2=0 $Y2=0
cc_585 N_A_779_380#_c_634_n N_A_596_81#_c_724_n 0.0156766f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_586 N_A_779_380#_c_636_n N_A_596_81#_c_724_n 0.00444456f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_587 N_A_779_380#_c_632_n N_A_596_81#_c_725_n 0.00237419f $X=4.41 $Y=1.01
+ $X2=0 $Y2=0
cc_588 N_A_779_380#_c_640_n N_A_596_81#_c_725_n 0.0704401f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_589 N_A_779_380#_c_641_n N_A_596_81#_c_725_n 0.00140465f $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_590 N_A_779_380#_c_634_n N_A_596_81#_c_725_n 0.0310993f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_591 N_A_779_380#_c_635_n N_A_596_81#_c_725_n 0.0123136f $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_592 N_A_779_380#_c_636_n N_A_596_81#_c_725_n 0.00126891f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_593 N_A_779_380#_c_638_n N_A_596_81#_c_726_n 0.00247902f $X=4.23 $Y=1.975
+ $X2=0 $Y2=0
cc_594 N_A_779_380#_c_640_n N_A_596_81#_c_726_n 0.00453512f $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_595 N_A_779_380#_c_641_n N_A_596_81#_c_726_n 6.72497e-19 $X=4.395 $Y=1.885
+ $X2=0 $Y2=0
cc_596 N_A_779_380#_c_634_n N_A_596_81#_c_727_n 0.0363901f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_597 N_A_779_380#_c_636_n N_A_596_81#_c_727_n 2.43226e-19 $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_598 N_A_779_380#_c_635_n N_A_596_81#_c_728_n 5.72749e-19 $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_599 N_A_779_380#_c_639_n N_A_596_81#_c_730_n 9.11465e-19 $X=4.075 $Y=1.975
+ $X2=0 $Y2=0
cc_600 N_A_779_380#_c_640_n N_A_596_81#_c_734_n 4.77624e-19 $X=4.95 $Y=1.885
+ $X2=0 $Y2=0
cc_601 N_A_779_380#_c_634_n N_A_596_81#_c_734_n 0.00223707f $X=5.015 $Y=0.6
+ $X2=0 $Y2=0
cc_602 N_A_779_380#_c_635_n N_A_596_81#_c_734_n 0.00869085f $X=4.395 $Y=1.72
+ $X2=0 $Y2=0
cc_603 N_A_779_380#_c_636_n N_A_596_81#_c_734_n 0.0136391f $X=4.575 $Y=1.01
+ $X2=0 $Y2=0
cc_604 N_A_779_380#_c_642_n N_SET_B_M1016_g 0.00434927f $X=5.115 $Y=2.515 $X2=0
+ $Y2=0
cc_605 N_A_779_380#_c_634_n N_SET_B_M1026_g 0.00137951f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_606 N_A_779_380#_c_640_n N_SET_B_c_883_n 0.0129984f $X=4.95 $Y=1.885 $X2=0
+ $Y2=0
cc_607 N_A_779_380#_c_640_n N_SET_B_c_896_n 0.00232552f $X=4.95 $Y=1.885 $X2=0
+ $Y2=0
cc_608 N_A_779_380#_M1020_g N_A_225_74#_M1007_g 0.0310413f $X=3.985 $Y=2.525
+ $X2=0 $Y2=0
cc_609 N_A_779_380#_M1020_g N_A_225_74#_c_1039_n 0.0123711f $X=3.985 $Y=2.525
+ $X2=0 $Y2=0
cc_610 N_A_779_380#_M1020_g N_VPWR_c_1632_n 0.00740427f $X=3.985 $Y=2.525 $X2=0
+ $Y2=0
cc_611 N_A_779_380#_M1020_g N_VPWR_c_1629_n 9.455e-19 $X=3.985 $Y=2.525 $X2=0
+ $Y2=0
cc_612 N_A_779_380#_c_631_n N_VGND_c_1820_n 0.0108567f $X=4.055 $Y=0.935 $X2=0
+ $Y2=0
cc_613 N_A_779_380#_c_632_n N_VGND_c_1820_n 0.00687895f $X=4.41 $Y=1.01 $X2=0
+ $Y2=0
cc_614 N_A_779_380#_c_634_n N_VGND_c_1820_n 0.0244437f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_615 N_A_779_380#_c_634_n N_VGND_c_1821_n 0.0122754f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_616 N_A_779_380#_c_631_n N_VGND_c_1824_n 0.0045897f $X=4.055 $Y=0.935 $X2=0
+ $Y2=0
cc_617 N_A_779_380#_c_634_n N_VGND_c_1829_n 0.0175574f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_618 N_A_779_380#_c_631_n N_VGND_c_1833_n 0.0044912f $X=4.055 $Y=0.935 $X2=0
+ $Y2=0
cc_619 N_A_779_380#_c_634_n N_VGND_c_1833_n 0.019759f $X=5.015 $Y=0.6 $X2=0
+ $Y2=0
cc_620 N_A_596_81#_M1001_g N_SET_B_M1016_g 0.010613f $X=6.195 $Y=2.205 $X2=0
+ $Y2=0
cc_621 N_A_596_81#_c_718_n N_SET_B_M1026_g 0.00527452f $X=5.025 $Y=1.57 $X2=0
+ $Y2=0
cc_622 N_A_596_81#_M1015_g N_SET_B_M1026_g 0.0611842f $X=5.23 $Y=0.58 $X2=0
+ $Y2=0
cc_623 N_A_596_81#_M1001_g N_SET_B_M1026_g 0.0142676f $X=6.195 $Y=2.205 $X2=0
+ $Y2=0
cc_624 N_A_596_81#_c_725_n N_SET_B_M1026_g 0.00301751f $X=4.95 $Y=1.52 $X2=0
+ $Y2=0
cc_625 N_A_596_81#_c_727_n N_SET_B_M1026_g 3.61773e-19 $X=5.092 $Y=1.29 $X2=0
+ $Y2=0
cc_626 N_A_596_81#_c_728_n N_SET_B_M1026_g 0.00154129f $X=5.092 $Y=1.435 $X2=0
+ $Y2=0
cc_627 N_A_596_81#_c_729_n N_SET_B_M1026_g 0.0148959f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_628 N_A_596_81#_c_732_n N_SET_B_M1026_g 0.00115306f $X=6.1 $Y=1.205 $X2=0
+ $Y2=0
cc_629 N_A_596_81#_c_733_n N_SET_B_M1026_g 0.0183335f $X=6.1 $Y=1.285 $X2=0
+ $Y2=0
cc_630 N_A_596_81#_c_735_n N_SET_B_M1026_g 0.0118733f $X=6.122 $Y=1.12 $X2=0
+ $Y2=0
cc_631 N_A_596_81#_M1001_g N_SET_B_c_881_n 0.0028286f $X=6.195 $Y=2.205 $X2=0
+ $Y2=0
cc_632 N_A_596_81#_c_729_n N_SET_B_c_881_n 0.00860328f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_633 N_A_596_81#_c_732_n N_SET_B_c_881_n 0.00789782f $X=6.1 $Y=1.205 $X2=0
+ $Y2=0
cc_634 N_A_596_81#_c_733_n N_SET_B_c_881_n 7.31285e-19 $X=6.1 $Y=1.285 $X2=0
+ $Y2=0
cc_635 N_A_596_81#_M1029_g N_SET_B_c_882_n 2.72666e-19 $X=4.89 $Y=2.525 $X2=0
+ $Y2=0
cc_636 N_A_596_81#_c_721_n N_SET_B_c_882_n 9.05772e-19 $X=5.025 $Y=1.645 $X2=0
+ $Y2=0
cc_637 N_A_596_81#_c_725_n N_SET_B_c_882_n 0.00172913f $X=4.95 $Y=1.52 $X2=0
+ $Y2=0
cc_638 N_A_596_81#_c_729_n N_SET_B_c_882_n 0.00314092f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_639 N_A_596_81#_M1029_g N_SET_B_c_883_n 6.13227e-19 $X=4.89 $Y=2.525 $X2=0
+ $Y2=0
cc_640 N_A_596_81#_M1001_g N_SET_B_c_883_n 7.12932e-19 $X=6.195 $Y=2.205 $X2=0
+ $Y2=0
cc_641 N_A_596_81#_c_721_n N_SET_B_c_883_n 0.00124776f $X=5.025 $Y=1.645 $X2=0
+ $Y2=0
cc_642 N_A_596_81#_c_725_n N_SET_B_c_883_n 0.00404118f $X=4.95 $Y=1.52 $X2=0
+ $Y2=0
cc_643 N_A_596_81#_c_729_n N_SET_B_c_883_n 0.0119231f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_644 N_A_596_81#_M1029_g N_SET_B_c_896_n 0.0256045f $X=4.89 $Y=2.525 $X2=0
+ $Y2=0
cc_645 N_A_596_81#_c_721_n N_SET_B_c_896_n 0.0065664f $X=5.025 $Y=1.645 $X2=0
+ $Y2=0
cc_646 N_A_596_81#_c_729_n N_SET_B_c_896_n 0.00385063f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_647 N_A_596_81#_c_722_n N_A_225_74#_M1004_g 8.37131e-19 $X=3.45 $Y=0.615
+ $X2=0 $Y2=0
cc_648 N_A_596_81#_c_739_n N_A_225_74#_M1007_g 0.0072187f $X=3.34 $Y=2.515 $X2=0
+ $Y2=0
cc_649 N_A_596_81#_c_730_n N_A_225_74#_M1007_g 0.00329404f $X=3.355 $Y=2.295
+ $X2=0 $Y2=0
cc_650 N_A_596_81#_M1029_g N_A_225_74#_c_1039_n 0.0105864f $X=4.89 $Y=2.525
+ $X2=0 $Y2=0
cc_651 N_A_596_81#_M1001_g N_A_225_74#_c_1039_n 0.0108881f $X=6.195 $Y=2.205
+ $X2=0 $Y2=0
cc_652 N_A_596_81#_M1001_g N_A_225_74#_c_1026_n 0.0437045f $X=6.195 $Y=2.205
+ $X2=0 $Y2=0
cc_653 N_A_596_81#_M1001_g N_A_1358_377#_c_1341_n 0.00184542f $X=6.195 $Y=2.205
+ $X2=0 $Y2=0
cc_654 N_A_596_81#_M1001_g N_A_1358_377#_c_1330_n 0.00164376f $X=6.195 $Y=2.205
+ $X2=0 $Y2=0
cc_655 N_A_596_81#_M1001_g N_A_1358_377#_c_1335_n 7.56949e-19 $X=6.195 $Y=2.205
+ $X2=0 $Y2=0
cc_656 N_A_596_81#_c_739_n N_A_27_80#_c_1570_n 0.0183821f $X=3.34 $Y=2.515 $X2=0
+ $Y2=0
cc_657 N_A_596_81#_c_730_n N_A_27_80#_c_1570_n 0.00583234f $X=3.355 $Y=2.295
+ $X2=0 $Y2=0
cc_658 N_A_596_81#_M1001_g N_VPWR_c_1633_n 0.00607807f $X=6.195 $Y=2.205 $X2=0
+ $Y2=0
cc_659 N_A_596_81#_M1001_g N_VPWR_c_1629_n 0.00113998f $X=6.195 $Y=2.205 $X2=0
+ $Y2=0
cc_660 N_A_596_81#_c_722_n N_VGND_c_1820_n 0.0102369f $X=3.45 $Y=0.615 $X2=0
+ $Y2=0
cc_661 N_A_596_81#_c_723_n N_VGND_c_1820_n 0.0136266f $X=4.115 $Y=0.97 $X2=0
+ $Y2=0
cc_662 N_A_596_81#_c_729_n N_VGND_c_1821_n 0.00656613f $X=5.935 $Y=1.205 $X2=0
+ $Y2=0
cc_663 N_A_596_81#_c_732_n N_VGND_c_1821_n 0.0179048f $X=6.1 $Y=1.205 $X2=0
+ $Y2=0
cc_664 N_A_596_81#_c_733_n N_VGND_c_1821_n 0.00159497f $X=6.1 $Y=1.285 $X2=0
+ $Y2=0
cc_665 N_A_596_81#_c_735_n N_VGND_c_1821_n 0.0113166f $X=6.122 $Y=1.12 $X2=0
+ $Y2=0
cc_666 N_A_596_81#_c_722_n N_VGND_c_1824_n 0.00962837f $X=3.45 $Y=0.615 $X2=0
+ $Y2=0
cc_667 N_A_596_81#_M1015_g N_VGND_c_1829_n 0.00434997f $X=5.23 $Y=0.58 $X2=0
+ $Y2=0
cc_668 N_A_596_81#_c_735_n N_VGND_c_1830_n 0.00383152f $X=6.122 $Y=1.12 $X2=0
+ $Y2=0
cc_669 N_A_596_81#_M1015_g N_VGND_c_1833_n 0.00824278f $X=5.23 $Y=0.58 $X2=0
+ $Y2=0
cc_670 N_A_596_81#_c_722_n N_VGND_c_1833_n 0.00894094f $X=3.45 $Y=0.615 $X2=0
+ $Y2=0
cc_671 N_A_596_81#_c_735_n N_VGND_c_1833_n 0.00758168f $X=6.122 $Y=1.12 $X2=0
+ $Y2=0
cc_672 N_SET_B_M1016_g N_A_225_74#_c_1039_n 0.0113188f $X=5.4 $Y=2.525 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_881_n N_A_225_74#_c_1025_n 0.00343552f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_881_n N_A_225_74#_c_1026_n 0.00710912f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_881_n N_A_225_74#_M1031_g 0.00409351f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_676 N_SET_B_M1024_g N_A_1510_48#_M1028_g 0.0563813f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_885_n N_A_1510_48#_M1028_g 0.00223551f $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_880_n N_A_1510_48#_M1010_g 0.0101099f $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_891_n N_A_1510_48#_M1010_g 0.026422f $X=8.39 $Y=2.305 $X2=0
+ $Y2=0
cc_680 N_SET_B_M1024_g N_A_1510_48#_c_1194_n 0.00739584f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_878_n N_A_1510_48#_c_1194_n 0.00256307f $X=8.34 $Y=1.3 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_879_n N_A_1510_48#_c_1194_n 0.00453006f $X=8.09 $Y=1.3 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_880_n N_A_1510_48#_c_1194_n 9.56134e-19 $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_881_n N_A_1510_48#_c_1194_n 0.025713f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_685 SET_B N_A_1510_48#_c_1194_n 0.00265164f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_686 N_SET_B_c_885_n N_A_1510_48#_c_1194_n 8.16272e-19 $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_886_n N_A_1510_48#_c_1194_n 0.0424843f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_878_n N_A_1510_48#_c_1195_n 0.0084215f $X=8.34 $Y=1.3 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_881_n N_A_1510_48#_c_1195_n 0.00472787f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_690 SET_B N_A_1510_48#_c_1195_n 0.00196951f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_691 N_SET_B_c_886_n N_A_1510_48#_c_1195_n 0.031422f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_692 N_SET_B_M1024_g N_A_1510_48#_c_1196_n 0.0108479f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_693 N_SET_B_M1014_g N_A_1510_48#_c_1203_n 8.10344e-19 $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_694 N_SET_B_M1014_g N_A_1510_48#_c_1205_n 7.2748e-19 $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_879_n N_A_1510_48#_c_1201_n 0.0104108f $X=8.09 $Y=1.3 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_880_n N_A_1510_48#_c_1201_n 0.0188382f $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_881_n N_A_1510_48#_c_1201_n 0.0105411f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_698 SET_B N_A_1510_48#_c_1201_n 8.64502e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_699 N_SET_B_c_886_n N_A_1510_48#_c_1201_n 9.42269e-19 $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_700 N_SET_B_M1024_g N_A_1358_377#_c_1309_n 0.00678433f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_886_n N_A_1358_377#_c_1310_n 0.00122225f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_891_n N_A_1358_377#_c_1311_n 0.00621639f $X=8.39 $Y=2.305 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_880_n N_A_1358_377#_c_1315_n 0.00621639f $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_885_n N_A_1358_377#_c_1315_n 0.0101337f $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_886_n N_A_1358_377#_c_1315_n 0.00368499f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_881_n N_A_1358_377#_c_1320_n 0.0130228f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_878_n N_A_1358_377#_c_1331_n 0.00442681f $X=8.34 $Y=1.3 $X2=0
+ $Y2=0
cc_708 N_SET_B_M1014_g N_A_1358_377#_c_1331_n 0.00824052f $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_880_n N_A_1358_377#_c_1331_n 0.00404324f $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_891_n N_A_1358_377#_c_1331_n 0.00462548f $X=8.39 $Y=2.305 $X2=0
+ $Y2=0
cc_711 N_SET_B_c_881_n N_A_1358_377#_c_1331_n 0.00672574f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_712 SET_B N_A_1358_377#_c_1331_n 0.00261165f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_713 N_SET_B_c_886_n N_A_1358_377#_c_1331_n 0.00628568f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_714 N_SET_B_M1014_g N_A_1358_377#_c_1332_n 0.00954469f $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_880_n N_A_1358_377#_c_1321_n 0.00158354f $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_716 SET_B N_A_1358_377#_c_1321_n 0.00118411f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_717 N_SET_B_c_885_n N_A_1358_377#_c_1321_n 0.00149353f $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_718 N_SET_B_c_886_n N_A_1358_377#_c_1321_n 0.0216237f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_719 N_SET_B_c_881_n N_A_1358_377#_c_1335_n 0.0266553f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_720 N_SET_B_M1014_g N_A_1358_377#_c_1338_n 4.5108e-19 $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_721 N_SET_B_c_881_n N_A_1358_377#_c_1338_n 0.00355761f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_722 N_SET_B_M1014_g N_A_1358_377#_c_1339_n 0.00399354f $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_880_n N_A_1358_377#_c_1339_n 0.00335406f $X=8.39 $Y=2.155 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_891_n N_A_1358_377#_c_1339_n 0.00409933f $X=8.39 $Y=2.305 $X2=0
+ $Y2=0
cc_725 SET_B N_A_1358_377#_c_1339_n 8.38169e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_726 N_SET_B_c_885_n N_A_1358_377#_c_1339_n 8.70886e-19 $X=8.505 $Y=1.3 $X2=0
+ $Y2=0
cc_727 N_SET_B_c_886_n N_A_1358_377#_c_1339_n 0.0129183f $X=8.505 $Y=1.39 $X2=0
+ $Y2=0
cc_728 N_SET_B_M1016_g N_VPWR_c_1633_n 0.00163772f $X=5.4 $Y=2.525 $X2=0 $Y2=0
cc_729 N_SET_B_M1014_g N_VPWR_c_1634_n 0.0027763f $X=8.38 $Y=2.75 $X2=0 $Y2=0
cc_730 N_SET_B_M1014_g N_VPWR_c_1643_n 0.005209f $X=8.38 $Y=2.75 $X2=0 $Y2=0
cc_731 N_SET_B_M1014_g N_VPWR_c_1629_n 0.00540654f $X=8.38 $Y=2.75 $X2=0 $Y2=0
cc_732 N_SET_B_M1026_g N_VGND_c_1821_n 0.0128389f $X=5.62 $Y=0.58 $X2=0 $Y2=0
cc_733 N_SET_B_M1026_g N_VGND_c_1829_n 0.00461464f $X=5.62 $Y=0.58 $X2=0 $Y2=0
cc_734 N_SET_B_M1024_g N_VGND_c_1830_n 0.00384553f $X=8.015 $Y=0.58 $X2=0 $Y2=0
cc_735 N_SET_B_M1026_g N_VGND_c_1833_n 0.00910593f $X=5.62 $Y=0.58 $X2=0 $Y2=0
cc_736 N_SET_B_M1024_g N_VGND_c_1833_n 0.00383468f $X=8.015 $Y=0.58 $X2=0 $Y2=0
cc_737 N_SET_B_M1024_g N_VGND_c_1837_n 0.0107673f $X=8.015 $Y=0.58 $X2=0 $Y2=0
cc_738 N_SET_B_c_878_n N_VGND_c_1837_n 2.20993e-19 $X=8.34 $Y=1.3 $X2=0 $Y2=0
cc_739 N_A_225_74#_M1031_g N_A_1510_48#_M1028_g 0.0378389f $X=7.235 $Y=0.58
+ $X2=0 $Y2=0
cc_740 N_A_225_74#_c_1025_n N_A_1510_48#_c_1201_n 0.039364f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_741 N_A_225_74#_M1002_g N_A_1358_377#_c_1341_n 0.00796309f $X=6.7 $Y=2.385
+ $X2=0 $Y2=0
cc_742 N_A_225_74#_c_1025_n N_A_1358_377#_c_1329_n 0.00139562f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_743 N_A_225_74#_M1002_g N_A_1358_377#_c_1330_n 0.0130962f $X=6.7 $Y=2.385
+ $X2=0 $Y2=0
cc_744 N_A_225_74#_c_1025_n N_A_1358_377#_c_1320_n 0.00327799f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_745 N_A_225_74#_M1031_g N_A_1358_377#_c_1320_n 0.0162403f $X=7.235 $Y=0.58
+ $X2=0 $Y2=0
cc_746 N_A_225_74#_M1002_g N_A_1358_377#_c_1335_n 0.00924922f $X=6.7 $Y=2.385
+ $X2=0 $Y2=0
cc_747 N_A_225_74#_c_1025_n N_A_1358_377#_c_1335_n 0.0170558f $X=7.16 $Y=1.735
+ $X2=0 $Y2=0
cc_748 N_A_225_74#_M1031_g N_A_1358_377#_c_1322_n 0.00979462f $X=7.235 $Y=0.58
+ $X2=0 $Y2=0
cc_749 N_A_225_74#_M1012_s N_A_27_80#_c_1569_n 0.0117593f $X=1.145 $Y=1.79 $X2=0
+ $Y2=0
cc_750 N_A_225_74#_c_1048_n N_A_27_80#_c_1569_n 0.0189258f $X=1.305 $Y=1.87
+ $X2=0 $Y2=0
cc_751 N_A_225_74#_c_1049_n N_A_27_80#_c_1569_n 0.0142272f $X=1.145 $Y=1.87
+ $X2=0 $Y2=0
cc_752 N_A_225_74#_c_1050_n N_A_27_80#_c_1569_n 0.00643406f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_753 N_A_225_74#_M1019_g N_A_27_80#_c_1570_n 0.0166103f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_754 N_A_225_74#_c_1035_n N_A_27_80#_c_1570_n 0.0298112f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_755 N_A_225_74#_c_1030_n N_A_27_80#_c_1570_n 6.87392e-19 $X=2.41 $Y=1.465
+ $X2=0 $Y2=0
cc_756 N_A_225_74#_c_1050_n N_A_27_80#_c_1570_n 0.0336256f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_757 N_A_225_74#_M1013_g N_A_27_80#_c_1564_n 8.15758e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_758 N_A_225_74#_M1019_g N_A_27_80#_c_1564_n 0.00102472f $X=1.965 $Y=2.35
+ $X2=0 $Y2=0
cc_759 N_A_225_74#_c_1035_n N_A_27_80#_c_1564_n 0.00927835f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_760 N_A_225_74#_c_1023_n N_A_27_80#_c_1564_n 0.0104106f $X=2.83 $Y=1.12 $X2=0
+ $Y2=0
cc_761 N_A_225_74#_M1004_g N_A_27_80#_c_1564_n 0.00434152f $X=2.905 $Y=0.615
+ $X2=0 $Y2=0
cc_762 N_A_225_74#_c_1029_n N_A_27_80#_c_1564_n 0.0147929f $X=2.485 $Y=1.12
+ $X2=0 $Y2=0
cc_763 N_A_225_74#_c_1050_n N_A_27_80#_c_1564_n 0.0137141f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_764 N_A_225_74#_c_1032_n N_A_27_80#_c_1564_n 0.0302853f $X=2.19 $Y=1.465
+ $X2=0 $Y2=0
cc_765 N_A_225_74#_M1019_g N_A_27_80#_c_1613_n 0.00329523f $X=1.965 $Y=2.35
+ $X2=0 $Y2=0
cc_766 N_A_225_74#_c_1050_n N_A_27_80#_c_1613_n 0.0100622f $X=2.025 $Y=1.805
+ $X2=0 $Y2=0
cc_767 N_A_225_74#_c_1023_n N_A_27_80#_c_1566_n 0.00467868f $X=2.83 $Y=1.12
+ $X2=0 $Y2=0
cc_768 N_A_225_74#_M1004_g N_A_27_80#_c_1566_n 0.00437989f $X=2.905 $Y=0.615
+ $X2=0 $Y2=0
cc_769 N_A_225_74#_c_1050_n N_VPWR_M1012_d 0.00164828f $X=2.025 $Y=1.805 $X2=0
+ $Y2=0
cc_770 N_A_225_74#_M1019_g N_VPWR_c_1631_n 0.00900773f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_771 N_A_225_74#_c_1035_n N_VPWR_c_1631_n 3.19321e-19 $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_772 N_A_225_74#_c_1037_n N_VPWR_c_1631_n 0.00272925f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_773 N_A_225_74#_M1007_g N_VPWR_c_1632_n 8.5651e-19 $X=3.565 $Y=2.525 $X2=0
+ $Y2=0
cc_774 N_A_225_74#_c_1039_n N_VPWR_c_1632_n 0.0290276f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_775 N_A_225_74#_c_1039_n N_VPWR_c_1633_n 0.0264687f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_776 N_A_225_74#_M1002_g N_VPWR_c_1633_n 0.00678774f $X=6.7 $Y=2.385 $X2=0
+ $Y2=0
cc_777 N_A_225_74#_c_1039_n N_VPWR_c_1637_n 0.0266989f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_778 N_A_225_74#_M1019_g N_VPWR_c_1641_n 0.00540231f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_779 N_A_225_74#_c_1037_n N_VPWR_c_1641_n 0.0376458f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_780 N_A_225_74#_c_1039_n N_VPWR_c_1642_n 0.0306837f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_781 N_A_225_74#_M1019_g N_VPWR_c_1629_n 0.00533457f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_782 N_A_225_74#_c_1036_n N_VPWR_c_1629_n 0.0215278f $X=3.475 $Y=3.15 $X2=0
+ $Y2=0
cc_783 N_A_225_74#_c_1037_n N_VPWR_c_1629_n 0.00604517f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_784 N_A_225_74#_c_1039_n N_VPWR_c_1629_n 0.0900942f $X=6.61 $Y=3.15 $X2=0
+ $Y2=0
cc_785 N_A_225_74#_c_1046_n N_VPWR_c_1629_n 0.00445015f $X=3.565 $Y=3.15 $X2=0
+ $Y2=0
cc_786 N_A_225_74#_c_1033_n N_VGND_c_1817_n 0.0387749f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_787 N_A_225_74#_c_1033_n N_VGND_c_1818_n 0.0203368f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_788 N_A_225_74#_M1013_g N_VGND_c_1819_n 0.0115714f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_789 N_A_225_74#_c_1033_n N_VGND_c_1819_n 0.0268179f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_790 N_A_225_74#_M1013_g N_VGND_c_1824_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_791 N_A_225_74#_M1004_g N_VGND_c_1824_n 9.15902e-19 $X=2.905 $Y=0.615 $X2=0
+ $Y2=0
cc_792 N_A_225_74#_M1031_g N_VGND_c_1830_n 0.00278271f $X=7.235 $Y=0.58 $X2=0
+ $Y2=0
cc_793 N_A_225_74#_M1013_g N_VGND_c_1833_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_794 N_A_225_74#_M1031_g N_VGND_c_1833_n 0.00353931f $X=7.235 $Y=0.58 $X2=0
+ $Y2=0
cc_795 N_A_225_74#_c_1033_n N_VGND_c_1833_n 0.0167889f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_796 N_A_1510_48#_c_1195_n N_A_1358_377#_c_1309_n 0.00361072f $X=8.925
+ $Y=0.925 $X2=0 $Y2=0
cc_797 N_A_1510_48#_c_1197_n N_A_1358_377#_c_1309_n 0.0116357f $X=9.09 $Y=0.58
+ $X2=0 $Y2=0
cc_798 N_A_1510_48#_c_1200_n N_A_1358_377#_c_1309_n 6.34661e-19 $X=9.09 $Y=0.925
+ $X2=0 $Y2=0
cc_799 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1311_n 0.0060783f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_800 N_A_1510_48#_c_1204_n N_A_1358_377#_c_1324_n 3.80361e-19 $X=9.565
+ $Y=2.475 $X2=0 $Y2=0
cc_801 N_A_1510_48#_c_1205_n N_A_1358_377#_c_1324_n 0.00203684f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_802 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1324_n 0.00447691f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_803 N_A_1510_48#_c_1203_n N_A_1358_377#_M1017_g 0.00846762f $X=9.165 $Y=2.75
+ $X2=0 $Y2=0
cc_804 N_A_1510_48#_c_1204_n N_A_1358_377#_M1017_g 0.0191381f $X=9.565 $Y=2.475
+ $X2=0 $Y2=0
cc_805 N_A_1510_48#_c_1197_n N_A_1358_377#_c_1312_n 0.0043971f $X=9.09 $Y=0.58
+ $X2=0 $Y2=0
cc_806 N_A_1510_48#_c_1198_n N_A_1358_377#_c_1312_n 0.00231095f $X=9.565
+ $Y=0.925 $X2=0 $Y2=0
cc_807 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1312_n 0.00225427f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_808 N_A_1510_48#_c_1204_n N_A_1358_377#_M1030_g 0.00180608f $X=9.565 $Y=2.475
+ $X2=0 $Y2=0
cc_809 N_A_1510_48#_c_1199_n N_A_1358_377#_M1030_g 0.00703389f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_810 N_A_1510_48#_c_1198_n N_A_1358_377#_c_1315_n 0.00745328f $X=9.565
+ $Y=0.925 $X2=0 $Y2=0
cc_811 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1315_n 0.0266131f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_812 N_A_1510_48#_c_1195_n N_A_1358_377#_c_1317_n 0.00925086f $X=8.925
+ $Y=0.925 $X2=0 $Y2=0
cc_813 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1317_n 0.00382379f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_814 N_A_1510_48#_c_1200_n N_A_1358_377#_c_1317_n 0.0207635f $X=9.09 $Y=0.925
+ $X2=0 $Y2=0
cc_815 N_A_1510_48#_M1028_g N_A_1358_377#_c_1320_n 6.67309e-19 $X=7.625 $Y=0.58
+ $X2=0 $Y2=0
cc_816 N_A_1510_48#_M1010_g N_A_1358_377#_c_1331_n 0.0145352f $X=7.93 $Y=2.75
+ $X2=0 $Y2=0
cc_817 N_A_1510_48#_c_1201_n N_A_1358_377#_c_1331_n 0.0019319f $X=7.93 $Y=1.75
+ $X2=0 $Y2=0
cc_818 N_A_1510_48#_M1010_g N_A_1358_377#_c_1332_n 5.32413e-19 $X=7.93 $Y=2.75
+ $X2=0 $Y2=0
cc_819 N_A_1510_48#_c_1203_n N_A_1358_377#_c_1332_n 0.0282823f $X=9.165 $Y=2.75
+ $X2=0 $Y2=0
cc_820 N_A_1510_48#_c_1205_n N_A_1358_377#_c_1332_n 0.00568936f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_821 N_A_1510_48#_c_1205_n N_A_1358_377#_c_1333_n 0.00538906f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_822 N_A_1510_48#_c_1204_n N_A_1358_377#_c_1334_n 0.00507721f $X=9.565
+ $Y=2.475 $X2=0 $Y2=0
cc_823 N_A_1510_48#_c_1205_n N_A_1358_377#_c_1334_n 0.0233648f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_824 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1334_n 0.0135838f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_825 N_A_1510_48#_c_1198_n N_A_1358_377#_c_1321_n 0.00978752f $X=9.565
+ $Y=0.925 $X2=0 $Y2=0
cc_826 N_A_1510_48#_c_1199_n N_A_1358_377#_c_1321_n 0.0615164f $X=9.65 $Y=2.39
+ $X2=0 $Y2=0
cc_827 N_A_1510_48#_c_1200_n N_A_1358_377#_c_1321_n 0.0140685f $X=9.09 $Y=0.925
+ $X2=0 $Y2=0
cc_828 N_A_1510_48#_M1028_g N_A_1358_377#_c_1322_n 2.73884e-19 $X=7.625 $Y=0.58
+ $X2=0 $Y2=0
cc_829 N_A_1510_48#_M1010_g N_A_1358_377#_c_1336_n 7.4227e-19 $X=7.93 $Y=2.75
+ $X2=0 $Y2=0
cc_830 N_A_1510_48#_M1010_g N_A_1358_377#_c_1338_n 0.0123678f $X=7.93 $Y=2.75
+ $X2=0 $Y2=0
cc_831 N_A_1510_48#_c_1194_n N_A_1358_377#_c_1338_n 0.0257755f $X=7.935 $Y=1.75
+ $X2=0 $Y2=0
cc_832 N_A_1510_48#_c_1201_n N_A_1358_377#_c_1338_n 0.00292111f $X=7.93 $Y=1.75
+ $X2=0 $Y2=0
cc_833 N_A_1510_48#_c_1205_n N_A_1358_377#_c_1339_n 0.00681171f $X=9.33 $Y=2.475
+ $X2=0 $Y2=0
cc_834 N_A_1510_48#_c_1204_n N_VPWR_M1017_d 0.00329098f $X=9.565 $Y=2.475 $X2=0
+ $Y2=0
cc_835 N_A_1510_48#_c_1199_n N_VPWR_M1017_d 0.0083441f $X=9.65 $Y=2.39 $X2=0
+ $Y2=0
cc_836 N_A_1510_48#_M1010_g N_VPWR_c_1634_n 0.00308998f $X=7.93 $Y=2.75 $X2=0
+ $Y2=0
cc_837 N_A_1510_48#_c_1203_n N_VPWR_c_1635_n 0.0080736f $X=9.165 $Y=2.75 $X2=0
+ $Y2=0
cc_838 N_A_1510_48#_c_1204_n N_VPWR_c_1635_n 0.00983167f $X=9.565 $Y=2.475 $X2=0
+ $Y2=0
cc_839 N_A_1510_48#_M1010_g N_VPWR_c_1637_n 0.0050156f $X=7.93 $Y=2.75 $X2=0
+ $Y2=0
cc_840 N_A_1510_48#_c_1203_n N_VPWR_c_1643_n 0.0144853f $X=9.165 $Y=2.75 $X2=0
+ $Y2=0
cc_841 N_A_1510_48#_M1010_g N_VPWR_c_1629_n 0.00540938f $X=7.93 $Y=2.75 $X2=0
+ $Y2=0
cc_842 N_A_1510_48#_c_1203_n N_VPWR_c_1629_n 0.0120561f $X=9.165 $Y=2.75 $X2=0
+ $Y2=0
cc_843 N_A_1510_48#_c_1204_n N_VPWR_c_1629_n 0.00788031f $X=9.565 $Y=2.475 $X2=0
+ $Y2=0
cc_844 N_A_1510_48#_c_1198_n N_Q_N_c_1769_n 0.00764487f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_845 N_A_1510_48#_c_1199_n Q_N 0.031214f $X=9.65 $Y=2.39 $X2=0 $Y2=0
cc_846 N_A_1510_48#_c_1198_n N_Q_N_c_1771_n 0.00277175f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_847 N_A_1510_48#_c_1199_n N_Q_N_c_1771_n 0.0148084f $X=9.65 $Y=2.39 $X2=0
+ $Y2=0
cc_848 N_A_1510_48#_c_1198_n N_VGND_M1008_s 0.00702554f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_849 N_A_1510_48#_c_1199_n N_VGND_M1008_s 0.00245883f $X=9.65 $Y=2.39 $X2=0
+ $Y2=0
cc_850 N_A_1510_48#_c_1197_n N_VGND_c_1822_n 0.0171919f $X=9.09 $Y=0.58 $X2=0
+ $Y2=0
cc_851 N_A_1510_48#_c_1198_n N_VGND_c_1822_n 0.0212677f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_852 N_A_1510_48#_c_1197_n N_VGND_c_1826_n 0.0102067f $X=9.09 $Y=0.58 $X2=0
+ $Y2=0
cc_853 N_A_1510_48#_M1028_g N_VGND_c_1830_n 0.00449242f $X=7.625 $Y=0.58 $X2=0
+ $Y2=0
cc_854 N_A_1510_48#_M1028_g N_VGND_c_1833_n 0.00871678f $X=7.625 $Y=0.58 $X2=0
+ $Y2=0
cc_855 N_A_1510_48#_c_1195_n N_VGND_c_1833_n 0.00709649f $X=8.925 $Y=0.925 $X2=0
+ $Y2=0
cc_856 N_A_1510_48#_c_1196_n N_VGND_c_1833_n 0.0108158f $X=8.1 $Y=0.925 $X2=0
+ $Y2=0
cc_857 N_A_1510_48#_c_1197_n N_VGND_c_1833_n 0.0114381f $X=9.09 $Y=0.58 $X2=0
+ $Y2=0
cc_858 N_A_1510_48#_c_1198_n N_VGND_c_1833_n 0.00883761f $X=9.565 $Y=0.925 $X2=0
+ $Y2=0
cc_859 N_A_1510_48#_M1028_g N_VGND_c_1837_n 0.00126877f $X=7.625 $Y=0.58 $X2=0
+ $Y2=0
cc_860 N_A_1510_48#_c_1195_n N_VGND_c_1837_n 0.0502316f $X=8.925 $Y=0.925 $X2=0
+ $Y2=0
cc_861 N_A_1510_48#_c_1196_n N_VGND_c_1837_n 0.00238625f $X=8.1 $Y=0.925 $X2=0
+ $Y2=0
cc_862 N_A_1358_377#_c_1318_n N_A_2113_74#_M1027_g 0.007876f $X=10.925 $Y=1.41
+ $X2=0 $Y2=0
cc_863 N_A_1358_377#_c_1328_n N_A_2113_74#_M1027_g 0.0162875f $X=10.965 $Y=1.94
+ $X2=0 $Y2=0
cc_864 N_A_1358_377#_c_1312_n N_A_2113_74#_c_1507_n 0.00119747f $X=9.935 $Y=1.21
+ $X2=0 $Y2=0
cc_865 N_A_1358_377#_M1025_g N_A_2113_74#_c_1507_n 0.00674464f $X=10.925
+ $Y=0.645 $X2=0 $Y2=0
cc_866 N_A_1358_377#_c_1312_n N_A_2113_74#_c_1508_n 3.90625e-19 $X=9.935 $Y=1.21
+ $X2=0 $Y2=0
cc_867 N_A_1358_377#_c_1314_n N_A_2113_74#_c_1508_n 0.00224708f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_868 N_A_1358_377#_M1025_g N_A_2113_74#_c_1508_n 0.0099886f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_869 N_A_1358_377#_c_1314_n N_A_2113_74#_c_1509_n 0.00487854f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_870 N_A_1358_377#_c_1319_n N_A_2113_74#_c_1509_n 0.0138825f $X=10.965 $Y=1.79
+ $X2=0 $Y2=0
cc_871 N_A_1358_377#_c_1328_n N_A_2113_74#_c_1509_n 0.0063108f $X=10.965 $Y=1.94
+ $X2=0 $Y2=0
cc_872 N_A_1358_377#_c_1318_n N_A_2113_74#_c_1510_n 0.0192f $X=10.925 $Y=1.41
+ $X2=0 $Y2=0
cc_873 N_A_1358_377#_c_1328_n N_A_2113_74#_c_1510_n 0.00290088f $X=10.965
+ $Y=1.94 $X2=0 $Y2=0
cc_874 N_A_1358_377#_c_1318_n N_A_2113_74#_c_1511_n 0.0169362f $X=10.925 $Y=1.41
+ $X2=0 $Y2=0
cc_875 N_A_1358_377#_c_1314_n N_A_2113_74#_c_1512_n 0.00533007f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_876 N_A_1358_377#_M1025_g N_A_2113_74#_c_1512_n 0.00377159f $X=10.925
+ $Y=0.645 $X2=0 $Y2=0
cc_877 N_A_1358_377#_c_1314_n N_A_2113_74#_c_1531_n 0.0110675f $X=10.85 $Y=1.41
+ $X2=0 $Y2=0
cc_878 N_A_1358_377#_c_1318_n N_A_2113_74#_c_1531_n 0.00192549f $X=10.925
+ $Y=1.41 $X2=0 $Y2=0
cc_879 N_A_1358_377#_M1025_g N_A_2113_74#_c_1513_n 0.0205551f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_880 N_A_1358_377#_c_1331_n N_VPWR_c_1634_n 0.0139684f $X=8.44 $Y=2.265 $X2=0
+ $Y2=0
cc_881 N_A_1358_377#_c_1332_n N_VPWR_c_1634_n 0.0115095f $X=8.605 $Y=2.75 $X2=0
+ $Y2=0
cc_882 N_A_1358_377#_M1017_g N_VPWR_c_1635_n 0.00918847f $X=9.475 $Y=2.75 $X2=0
+ $Y2=0
cc_883 N_A_1358_377#_M1030_g N_VPWR_c_1635_n 0.0107842f $X=9.98 $Y=2.4 $X2=0
+ $Y2=0
cc_884 N_A_1358_377#_c_1328_n N_VPWR_c_1636_n 0.0182547f $X=10.965 $Y=1.94 $X2=0
+ $Y2=0
cc_885 N_A_1358_377#_c_1329_n N_VPWR_c_1637_n 0.0133359f $X=7.238 $Y=2.692 $X2=0
+ $Y2=0
cc_886 N_A_1358_377#_c_1330_n N_VPWR_c_1637_n 0.00847891f $X=7.01 $Y=2.692 $X2=0
+ $Y2=0
cc_887 N_A_1358_377#_c_1337_n N_VPWR_c_1637_n 0.0062276f $X=7.73 $Y=2.35 $X2=0
+ $Y2=0
cc_888 N_A_1358_377#_M1017_g N_VPWR_c_1643_n 0.00536974f $X=9.475 $Y=2.75 $X2=0
+ $Y2=0
cc_889 N_A_1358_377#_c_1332_n N_VPWR_c_1643_n 0.014549f $X=8.605 $Y=2.75 $X2=0
+ $Y2=0
cc_890 N_A_1358_377#_M1030_g N_VPWR_c_1644_n 0.00490827f $X=9.98 $Y=2.4 $X2=0
+ $Y2=0
cc_891 N_A_1358_377#_c_1328_n N_VPWR_c_1644_n 0.00502645f $X=10.965 $Y=1.94
+ $X2=0 $Y2=0
cc_892 N_A_1358_377#_M1017_g N_VPWR_c_1629_n 0.00521875f $X=9.475 $Y=2.75 $X2=0
+ $Y2=0
cc_893 N_A_1358_377#_M1030_g N_VPWR_c_1629_n 0.009739f $X=9.98 $Y=2.4 $X2=0
+ $Y2=0
cc_894 N_A_1358_377#_c_1328_n N_VPWR_c_1629_n 0.00516335f $X=10.965 $Y=1.94
+ $X2=0 $Y2=0
cc_895 N_A_1358_377#_c_1329_n N_VPWR_c_1629_n 0.0150402f $X=7.238 $Y=2.692 $X2=0
+ $Y2=0
cc_896 N_A_1358_377#_c_1330_n N_VPWR_c_1629_n 0.0086556f $X=7.01 $Y=2.692 $X2=0
+ $Y2=0
cc_897 N_A_1358_377#_c_1331_n N_VPWR_c_1629_n 0.012403f $X=8.44 $Y=2.265 $X2=0
+ $Y2=0
cc_898 N_A_1358_377#_c_1332_n N_VPWR_c_1629_n 0.0119743f $X=8.605 $Y=2.75 $X2=0
+ $Y2=0
cc_899 N_A_1358_377#_c_1337_n N_VPWR_c_1629_n 0.0116125f $X=7.73 $Y=2.35 $X2=0
+ $Y2=0
cc_900 N_A_1358_377#_c_1337_n A_1520_508# 0.00131813f $X=7.73 $Y=2.35 $X2=-0.19
+ $Y2=-0.245
cc_901 N_A_1358_377#_c_1338_n A_1520_508# 0.00101432f $X=7.9 $Y=2.35 $X2=-0.19
+ $Y2=-0.245
cc_902 N_A_1358_377#_c_1312_n N_Q_N_c_1769_n 0.0141919f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_903 N_A_1358_377#_M1025_g N_Q_N_c_1769_n 0.00158934f $X=10.925 $Y=0.645 $X2=0
+ $Y2=0
cc_904 N_A_1358_377#_M1030_g Q_N 0.00759938f $X=9.98 $Y=2.4 $X2=0 $Y2=0
cc_905 N_A_1358_377#_c_1314_n Q_N 0.0254096f $X=10.85 $Y=1.41 $X2=0 $Y2=0
cc_906 N_A_1358_377#_c_1328_n Q_N 0.00375639f $X=10.965 $Y=1.94 $X2=0 $Y2=0
cc_907 N_A_1358_377#_c_1312_n N_Q_N_c_1771_n 0.00565895f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_908 N_A_1358_377#_c_1314_n N_Q_N_c_1771_n 0.0163549f $X=10.85 $Y=1.41 $X2=0
+ $Y2=0
cc_909 N_A_1358_377#_M1025_g N_Q_N_c_1771_n 0.00117107f $X=10.925 $Y=0.645 $X2=0
+ $Y2=0
cc_910 N_A_1358_377#_M1025_g N_Q_c_1798_n 6.13748e-19 $X=10.925 $Y=0.645 $X2=0
+ $Y2=0
cc_911 N_A_1358_377#_c_1328_n Q 0.00119838f $X=10.965 $Y=1.94 $X2=0 $Y2=0
cc_912 N_A_1358_377#_c_1309_n N_VGND_c_1822_n 0.00403474f $X=8.875 $Y=0.865
+ $X2=0 $Y2=0
cc_913 N_A_1358_377#_c_1312_n N_VGND_c_1822_n 0.0109009f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_914 N_A_1358_377#_c_1315_n N_VGND_c_1822_n 0.00184748f $X=10.07 $Y=1.41 $X2=0
+ $Y2=0
cc_915 N_A_1358_377#_M1025_g N_VGND_c_1823_n 0.00686847f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_916 N_A_1358_377#_c_1309_n N_VGND_c_1826_n 0.00435647f $X=8.875 $Y=0.865
+ $X2=0 $Y2=0
cc_917 N_A_1358_377#_c_1312_n N_VGND_c_1831_n 0.00434272f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_918 N_A_1358_377#_M1025_g N_VGND_c_1831_n 0.00434272f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_919 N_A_1358_377#_c_1309_n N_VGND_c_1833_n 0.00454088f $X=8.875 $Y=0.865
+ $X2=0 $Y2=0
cc_920 N_A_1358_377#_c_1312_n N_VGND_c_1833_n 0.00830058f $X=9.935 $Y=1.21 $X2=0
+ $Y2=0
cc_921 N_A_1358_377#_M1025_g N_VGND_c_1833_n 0.00826607f $X=10.925 $Y=0.645
+ $X2=0 $Y2=0
cc_922 N_A_1358_377#_c_1309_n N_VGND_c_1837_n 0.0074138f $X=8.875 $Y=0.865 $X2=0
+ $Y2=0
cc_923 N_A_2113_74#_M1027_g N_VPWR_c_1636_n 0.00607682f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_924 N_A_2113_74#_c_1509_n N_VPWR_c_1636_n 0.0302671f $X=10.765 $Y=2.16 $X2=0
+ $Y2=0
cc_925 N_A_2113_74#_c_1510_n N_VPWR_c_1636_n 0.0131129f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_926 N_A_2113_74#_c_1511_n N_VPWR_c_1636_n 0.00228579f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_927 N_A_2113_74#_c_1509_n N_VPWR_c_1644_n 0.00525601f $X=10.765 $Y=2.16 $X2=0
+ $Y2=0
cc_928 N_A_2113_74#_M1027_g N_VPWR_c_1645_n 0.005209f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_929 N_A_2113_74#_M1027_g N_VPWR_c_1629_n 0.00990581f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_930 N_A_2113_74#_c_1509_n N_VPWR_c_1629_n 0.00579841f $X=10.765 $Y=2.16 $X2=0
+ $Y2=0
cc_931 N_A_2113_74#_c_1507_n N_Q_N_c_1769_n 0.0397432f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_932 N_A_2113_74#_c_1508_n N_Q_N_c_1769_n 0.00113323f $X=10.777 $Y=1.22 $X2=0
+ $Y2=0
cc_933 N_A_2113_74#_c_1509_n Q_N 0.0793988f $X=10.765 $Y=2.16 $X2=0 $Y2=0
cc_934 N_A_2113_74#_c_1531_n Q_N 0.0126081f $X=10.777 $Y=1.385 $X2=0 $Y2=0
cc_935 N_A_2113_74#_c_1508_n N_Q_N_c_1771_n 0.0124563f $X=10.777 $Y=1.22 $X2=0
+ $Y2=0
cc_936 N_A_2113_74#_c_1531_n N_Q_N_c_1771_n 0.00696689f $X=10.777 $Y=1.385 $X2=0
+ $Y2=0
cc_937 N_A_2113_74#_c_1513_n N_Q_c_1798_n 0.00613596f $X=11.42 $Y=1.22 $X2=0
+ $Y2=0
cc_938 N_A_2113_74#_c_1513_n N_Q_c_1799_n 0.00402186f $X=11.42 $Y=1.22 $X2=0
+ $Y2=0
cc_939 N_A_2113_74#_M1027_g Q 0.0182443f $X=11.495 $Y=2.4 $X2=0 $Y2=0
cc_940 N_A_2113_74#_c_1510_n N_Q_c_1800_n 0.0256386f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_941 N_A_2113_74#_c_1511_n N_Q_c_1800_n 0.015816f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_942 N_A_2113_74#_c_1513_n N_Q_c_1800_n 0.00424967f $X=11.42 $Y=1.22 $X2=0
+ $Y2=0
cc_943 N_A_2113_74#_c_1507_n N_VGND_c_1823_n 0.022629f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_944 N_A_2113_74#_c_1510_n N_VGND_c_1823_n 0.0190052f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_945 N_A_2113_74#_c_1511_n N_VGND_c_1823_n 0.00278132f $X=11.42 $Y=1.385 $X2=0
+ $Y2=0
cc_946 N_A_2113_74#_c_1513_n N_VGND_c_1823_n 0.00691628f $X=11.42 $Y=1.22 $X2=0
+ $Y2=0
cc_947 N_A_2113_74#_c_1507_n N_VGND_c_1831_n 0.0145025f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_948 N_A_2113_74#_c_1513_n N_VGND_c_1832_n 0.00434272f $X=11.42 $Y=1.22 $X2=0
+ $Y2=0
cc_949 N_A_2113_74#_c_1507_n N_VGND_c_1833_n 0.0119747f $X=10.71 $Y=0.645 $X2=0
+ $Y2=0
cc_950 N_A_2113_74#_c_1513_n N_VGND_c_1833_n 0.00825042f $X=11.42 $Y=1.22 $X2=0
+ $Y2=0
cc_951 N_A_27_80#_c_1570_n N_VPWR_M1012_d 9.71305e-19 $X=2.525 $Y=2.145 $X2=0
+ $Y2=0
cc_952 N_A_27_80#_c_1613_n N_VPWR_M1012_d 0.00470031f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_953 N_A_27_80#_c_1568_n N_VPWR_c_1630_n 0.0135247f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_954 N_A_27_80#_c_1569_n N_VPWR_c_1630_n 0.0195559f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_955 N_A_27_80#_c_1569_n N_VPWR_c_1631_n 0.00216696f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_956 N_A_27_80#_c_1570_n N_VPWR_c_1631_n 0.00260316f $X=2.525 $Y=2.145 $X2=0
+ $Y2=0
cc_957 N_A_27_80#_c_1613_n N_VPWR_c_1631_n 0.0112212f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_958 N_A_27_80#_c_1568_n N_VPWR_c_1639_n 0.011066f $X=0.28 $Y=2.75 $X2=0 $Y2=0
cc_959 N_A_27_80#_c_1568_n N_VPWR_c_1629_n 0.00915947f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_960 N_A_27_80#_c_1562_n N_VGND_c_1817_n 0.0172562f $X=0.28 $Y=0.61 $X2=0
+ $Y2=0
cc_961 N_A_27_80#_c_1562_n N_VGND_c_1828_n 0.00978756f $X=0.28 $Y=0.61 $X2=0
+ $Y2=0
cc_962 N_A_27_80#_c_1562_n N_VGND_c_1833_n 0.00895297f $X=0.28 $Y=0.61 $X2=0
+ $Y2=0
cc_963 N_VPWR_c_1635_n Q_N 0.00867007f $X=9.735 $Y=2.815 $X2=0 $Y2=0
cc_964 N_VPWR_c_1636_n Q_N 0.00312645f $X=11.215 $Y=2.16 $X2=0 $Y2=0
cc_965 N_VPWR_c_1644_n Q_N 0.0139663f $X=11.05 $Y=3.33 $X2=0 $Y2=0
cc_966 N_VPWR_c_1629_n Q_N 0.0115601f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_967 N_VPWR_c_1636_n Q 0.0368843f $X=11.215 $Y=2.16 $X2=0 $Y2=0
cc_968 N_VPWR_c_1645_n Q 0.014549f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_969 N_VPWR_c_1629_n Q 0.0119743f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_970 N_Q_N_c_1769_n N_VGND_c_1822_n 0.0127977f $X=10.15 $Y=0.515 $X2=0 $Y2=0
cc_971 N_Q_N_c_1769_n N_VGND_c_1831_n 0.0145639f $X=10.15 $Y=0.515 $X2=0 $Y2=0
cc_972 N_Q_N_c_1769_n N_VGND_c_1833_n 0.0119984f $X=10.15 $Y=0.515 $X2=0 $Y2=0
cc_973 N_Q_c_1798_n N_VGND_c_1823_n 0.0228912f $X=11.72 $Y=0.515 $X2=0 $Y2=0
cc_974 N_Q_c_1798_n N_VGND_c_1832_n 0.0145787f $X=11.72 $Y=0.515 $X2=0 $Y2=0
cc_975 N_Q_c_1798_n N_VGND_c_1833_n 0.0120042f $X=11.72 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__or3_4.pxi.spice
* Created: Wed Sep  2 12:28:24 2020
* 
x_PM_SKY130_FD_SC_MS__OR3_4%A N_A_M1006_g N_A_M1013_g N_A_M1001_g N_A_c_96_n
+ N_A_c_97_n N_A_c_98_n N_A_c_99_n N_A_c_100_n A N_A_c_102_n N_A_c_103_n A
+ PM_SKY130_FD_SC_MS__OR3_4%A
x_PM_SKY130_FD_SC_MS__OR3_4%B N_B_M1009_g N_B_M1014_g N_B_M1015_g B B B B
+ N_B_c_184_n N_B_c_185_n N_B_c_186_n PM_SKY130_FD_SC_MS__OR3_4%B
x_PM_SKY130_FD_SC_MS__OR3_4%C N_C_M1003_g N_C_M1005_g N_C_c_243_n N_C_M1008_g
+ N_C_c_244_n C N_C_c_245_n N_C_c_246_n PM_SKY130_FD_SC_MS__OR3_4%C
x_PM_SKY130_FD_SC_MS__OR3_4%A_305_388# N_A_305_388#_M1008_s N_A_305_388#_M1015_d
+ N_A_305_388#_M1003_d N_A_305_388#_M1004_g N_A_305_388#_M1000_g
+ N_A_305_388#_M1007_g N_A_305_388#_M1002_g N_A_305_388#_M1011_g
+ N_A_305_388#_M1010_g N_A_305_388#_M1012_g N_A_305_388#_M1016_g
+ N_A_305_388#_c_302_n N_A_305_388#_c_318_n N_A_305_388#_c_322_n
+ N_A_305_388#_c_303_n N_A_305_388#_c_304_n N_A_305_388#_c_325_n
+ N_A_305_388#_c_305_n N_A_305_388#_c_306_n N_A_305_388#_c_395_p
+ N_A_305_388#_c_347_n N_A_305_388#_c_332_n N_A_305_388#_c_307_n
+ N_A_305_388#_c_308_n PM_SKY130_FD_SC_MS__OR3_4%A_305_388#
x_PM_SKY130_FD_SC_MS__OR3_4%VPWR N_VPWR_M1006_d N_VPWR_M1013_d N_VPWR_M1007_s
+ N_VPWR_M1012_s N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n
+ N_VPWR_c_462_n N_VPWR_c_463_n VPWR N_VPWR_c_464_n N_VPWR_c_465_n
+ N_VPWR_c_466_n N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_457_n
+ PM_SKY130_FD_SC_MS__OR3_4%VPWR
x_PM_SKY130_FD_SC_MS__OR3_4%A_119_388# N_A_119_388#_M1006_s N_A_119_388#_M1014_d
+ N_A_119_388#_c_526_n N_A_119_388#_c_524_n N_A_119_388#_c_533_n
+ N_A_119_388#_c_529_n N_A_119_388#_c_525_n N_A_119_388#_c_531_n
+ PM_SKY130_FD_SC_MS__OR3_4%A_119_388#
x_PM_SKY130_FD_SC_MS__OR3_4%A_209_388# N_A_209_388#_M1009_s N_A_209_388#_M1005_s
+ N_A_209_388#_c_556_n PM_SKY130_FD_SC_MS__OR3_4%A_209_388#
x_PM_SKY130_FD_SC_MS__OR3_4%X N_X_M1000_d N_X_M1010_d N_X_M1004_d N_X_M1011_d
+ N_X_c_570_n N_X_c_577_n N_X_c_571_n N_X_c_572_n N_X_c_578_n N_X_c_579_n
+ N_X_c_580_n N_X_c_573_n N_X_c_574_n N_X_c_581_n N_X_c_582_n N_X_c_575_n X X
+ PM_SKY130_FD_SC_MS__OR3_4%X
x_PM_SKY130_FD_SC_MS__OR3_4%VGND N_VGND_M1008_d N_VGND_M1001_d N_VGND_M1002_s
+ N_VGND_M1016_s N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n
+ N_VGND_c_653_n N_VGND_c_654_n VGND N_VGND_c_655_n N_VGND_c_656_n
+ N_VGND_c_657_n N_VGND_c_658_n N_VGND_c_659_n N_VGND_c_660_n N_VGND_c_661_n
+ PM_SKY130_FD_SC_MS__OR3_4%VGND
cc_1 VNB N_A_M1006_g 0.00241604f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.44
cc_2 VNB N_A_M1013_g 0.00642334f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=2.44
cc_3 VNB N_A_c_96_n 0.00249471f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_4 VNB N_A_c_97_n 0.156212f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_5 VNB N_A_c_98_n 0.0390478f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.195
cc_6 VNB N_A_c_99_n 0.00249596f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.195
cc_7 VNB N_A_c_100_n 0.0323079f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_8 VNB A 0.00692367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_c_102_n 0.0410223f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_A_c_103_n 0.0176807f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.22
cc_11 VNB A 0.00534102f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_12 VNB N_B_M1015_g 0.0292678f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=0.74
cc_13 VNB N_B_c_184_n 0.0192821f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_14 VNB N_B_c_185_n 0.0166162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_186_n 0.00863455f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.385
cc_16 VNB N_C_M1003_g 0.00649245f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.44
cc_17 VNB N_C_M1005_g 0.00671204f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=2.44
cc_18 VNB N_C_c_243_n 0.0167983f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=1.22
cc_19 VNB N_C_c_244_n 0.0571927f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_20 VNB N_C_c_245_n 0.0972169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_c_246_n 0.00245092f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.385
cc_22 VNB N_A_305_388#_M1004_g 0.00151688f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.11
cc_23 VNB N_A_305_388#_M1000_g 0.0204334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_305_388#_M1007_g 0.00154088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_305_388#_M1002_g 0.0211635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_305_388#_M1011_g 0.00154206f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.385
cc_27 VNB N_A_305_388#_M1010_g 0.02167f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_28 VNB N_A_305_388#_M1012_g 0.00167778f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_29 VNB N_A_305_388#_M1016_g 0.0232609f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.55
cc_30 VNB N_A_305_388#_c_302_n 0.00530233f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.33
cc_31 VNB N_A_305_388#_c_303_n 0.00124938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_305_388#_c_304_n 0.00279725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_305_388#_c_305_n 0.00113959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_305_388#_c_306_n 2.94743e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_305_388#_c_307_n 0.00237265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_305_388#_c_308_n 0.0824207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_457_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_570_n 0.0017961f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_39 VNB N_X_c_571_n 0.00311091f $X=-0.19 $Y=-0.245 $X2=2.92 $Y2=1.385
cc_40 VNB N_X_c_572_n 0.00138775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_573_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_42 VNB N_X_c_574_n 0.00874592f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.63
cc_43 VNB N_X_c_575_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_44 VNB X 0.0264101f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_45 VNB N_VGND_c_649_n 0.00595424f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.445
cc_46 VNB N_VGND_c_650_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.195
cc_47 VNB N_VGND_c_651_n 0.00499383f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.385
cc_48 VNB N_VGND_c_652_n 0.00425095f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_49 VNB N_VGND_c_653_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_654_n 0.0258474f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=0.445
cc_51 VNB N_VGND_c_655_n 0.0588809f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_52 VNB N_VGND_c_656_n 0.0153327f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.28
cc_53 VNB N_VGND_c_657_n 0.0191617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_658_n 0.00614151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_659_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_660_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_661_n 0.320708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VPB N_A_M1006_g 0.0355372f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.44
cc_59 VPB N_A_M1013_g 0.0294519f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=2.44
cc_60 VPB N_B_M1009_g 0.0213501f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.44
cc_61 VPB N_B_M1014_g 0.0221592f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=2.44
cc_62 VPB N_B_c_184_n 0.0113932f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.385
cc_63 VPB N_B_c_185_n 0.0107382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B_c_186_n 0.012713f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.385
cc_65 VPB N_C_M1003_g 0.0258167f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.44
cc_66 VPB N_C_M1005_g 0.0262533f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=2.44
cc_67 VPB N_A_305_388#_M1004_g 0.0223084f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.11
cc_68 VPB N_A_305_388#_M1007_g 0.0214493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_305_388#_M1011_g 0.0220562f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.385
cc_70 VPB N_A_305_388#_M1012_g 0.0240093f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_71 VPB N_A_305_388#_c_306_n 0.00182944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_458_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.445
cc_73 VPB N_VPWR_c_459_n 0.0535422f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.445
cc_74 VPB N_VPWR_c_460_n 0.00638034f $X=-0.19 $Y=1.66 $X2=2.905 $Y2=1.385
cc_75 VPB N_VPWR_c_461_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_76 VPB N_VPWR_c_462_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_463_n 0.0428715f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=0.445
cc_78 VPB N_VPWR_c_464_n 0.0707163f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_79 VPB N_VPWR_c_465_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.28
cc_80 VPB N_VPWR_c_466_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_467_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_468_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_457_n 0.0881585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_119_388#_c_524_n 0.00208201f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.445
cc_85 VPB N_A_119_388#_c_525_n 0.00283773f $X=-0.19 $Y=1.66 $X2=2.905 $Y2=1.195
cc_86 VPB N_A_209_388#_c_556_n 0.00780755f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=0.74
cc_87 VPB N_X_c_577_n 0.00179594f $X=-0.19 $Y=1.66 $X2=2.905 $Y2=1.195
cc_88 VPB N_X_c_578_n 0.00264443f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_89 VPB N_X_c_579_n 0.00156879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_X_c_580_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=0.445
cc_91 VPB N_X_c_581_n 0.00811587f $X=-0.19 $Y=1.66 $X2=2.92 $Y2=1.22
cc_92 VPB N_X_c_582_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.28
cc_93 VPB X 0.00682831f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_94 N_A_M1006_g N_B_M1009_g 0.0148372f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_95 N_A_M1013_g N_B_M1014_g 0.0260709f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_96 N_A_c_98_n N_B_M1015_g 0.010633f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_97 N_A_c_99_n N_B_M1015_g 0.00124415f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_98 N_A_c_100_n N_B_M1015_g 0.0127642f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_c_103_n N_B_M1015_g 0.0212043f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_100 N_A_c_98_n N_B_c_184_n 0.00665044f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_101 N_A_c_102_n N_B_c_184_n 0.0202782f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_102 N_A_M1013_g N_B_c_185_n 0.0108981f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_103 N_A_c_98_n N_B_c_185_n 0.00429179f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_104 N_A_c_100_n N_B_c_185_n 0.0063017f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_105 N_A_M1013_g N_B_c_186_n 0.00129203f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_106 N_A_c_98_n N_B_c_186_n 0.145451f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_107 N_A_c_99_n N_B_c_186_n 0.00662177f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_108 N_A_c_100_n N_B_c_186_n 3.44095e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_109 N_A_c_102_n N_B_c_186_n 0.00645036f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_110 A N_B_c_186_n 0.0150931f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_111 N_A_c_98_n N_C_c_243_n 0.00518557f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_112 N_A_c_98_n N_C_c_244_n 0.0255921f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_113 N_A_c_96_n N_C_c_245_n 0.00317605f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_c_97_n N_C_c_245_n 0.0259948f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_c_98_n N_C_c_245_n 0.0149653f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_116 N_A_c_96_n N_C_c_246_n 0.0170535f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_c_97_n N_C_c_246_n 0.00315685f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_118 N_A_c_98_n N_C_c_246_n 0.0249544f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_119 N_A_c_99_n N_A_305_388#_M1015_d 0.00108111f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_120 N_A_c_99_n N_A_305_388#_M1000_g 3.74191e-19 $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_121 N_A_c_100_n N_A_305_388#_M1000_g 0.0035568f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_122 N_A_c_103_n N_A_305_388#_M1000_g 0.0249349f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A_M1013_g N_A_305_388#_c_318_n 0.0183876f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_124 N_A_c_98_n N_A_305_388#_c_318_n 0.0055927f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_125 N_A_c_99_n N_A_305_388#_c_318_n 0.00927791f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_126 N_A_c_100_n N_A_305_388#_c_318_n 0.00116691f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_127 N_A_c_98_n N_A_305_388#_c_322_n 0.0424115f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_128 N_A_c_98_n N_A_305_388#_c_303_n 0.0243069f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_129 N_A_c_103_n N_A_305_388#_c_304_n 0.00627897f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_c_99_n N_A_305_388#_c_325_n 0.0112121f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_131 N_A_c_100_n N_A_305_388#_c_325_n 9.11899e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_132 N_A_c_103_n N_A_305_388#_c_325_n 0.00865712f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_c_99_n N_A_305_388#_c_305_n 0.014585f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_134 N_A_c_100_n N_A_305_388#_c_305_n 5.12525e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A_c_103_n N_A_305_388#_c_305_n 0.00373084f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_136 N_A_M1013_g N_A_305_388#_c_306_n 0.00627861f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_137 N_A_c_98_n N_A_305_388#_c_332_n 0.0157928f $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_138 N_A_c_99_n N_A_305_388#_c_332_n 0.0080232f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_139 N_A_c_100_n N_A_305_388#_c_332_n 4.47564e-19 $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_140 N_A_c_103_n N_A_305_388#_c_332_n 7.14557e-19 $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_141 N_A_M1013_g N_A_305_388#_c_307_n 9.95864e-19 $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_142 N_A_c_99_n N_A_305_388#_c_307_n 0.0209458f $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_143 N_A_c_100_n N_A_305_388#_c_307_n 0.00176886f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_144 N_A_M1013_g N_A_305_388#_c_308_n 0.035111f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_145 N_A_c_99_n N_A_305_388#_c_308_n 2.43886e-19 $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_146 N_A_c_100_n N_A_305_388#_c_308_n 0.0124829f $X=2.92 $Y=1.385 $X2=0 $Y2=0
cc_147 N_A_M1006_g N_VPWR_c_459_n 0.00586602f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_148 N_A_c_102_n N_VPWR_c_459_n 0.00182202f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_149 A N_VPWR_c_459_n 0.0148078f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_150 N_A_M1013_g N_VPWR_c_460_n 0.0067952f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_VPWR_c_464_n 0.00644749f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_152 N_A_M1013_g N_VPWR_c_464_n 0.00644749f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_153 N_A_M1006_g N_VPWR_c_457_n 0.00647345f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_154 N_A_M1013_g N_VPWR_c_457_n 0.00647345f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_155 N_A_M1006_g N_A_119_388#_c_526_n 0.0061092f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_156 N_A_c_98_n N_A_119_388#_c_526_n 8.3091e-19 $X=2.755 $Y=1.195 $X2=0 $Y2=0
cc_157 N_A_M1006_g N_A_119_388#_c_524_n 0.00570546f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_158 N_A_M1013_g N_A_119_388#_c_529_n 0.00345517f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_159 N_A_M1013_g N_A_119_388#_c_525_n 0.00559667f $X=2.89 $Y=2.44 $X2=0 $Y2=0
cc_160 N_A_M1006_g N_A_119_388#_c_531_n 0.00213632f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_161 N_A_c_99_n N_VGND_M1001_d 5.36408e-19 $X=2.905 $Y=1.195 $X2=0 $Y2=0
cc_162 N_A_c_103_n N_VGND_c_649_n 4.07914e-19 $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A_c_103_n N_VGND_c_650_n 0.00434272f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_c_103_n N_VGND_c_651_n 0.0030773f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_c_96_n N_VGND_c_655_n 0.0191905f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_c_97_n N_VGND_c_655_n 0.00793088f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A_c_96_n N_VGND_c_661_n 0.012382f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_c_97_n N_VGND_c_661_n 0.00575727f $X=0.27 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_c_103_n N_VGND_c_661_n 0.00431597f $X=2.92 $Y=1.22 $X2=0 $Y2=0
cc_170 N_B_M1009_g N_C_M1003_g 0.041734f $X=0.955 $Y=2.44 $X2=0 $Y2=0
cc_171 N_B_c_186_n N_C_M1003_g 0.0148463f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_172 N_B_M1014_g N_C_M1005_g 0.0392566f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_173 N_B_c_186_n N_C_M1005_g 0.0131094f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_174 N_B_M1015_g N_C_c_243_n 0.0303957f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B_M1015_g N_C_c_244_n 0.00483407f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B_c_184_n N_C_c_244_n 0.026692f $X=0.97 $Y=1.615 $X2=0 $Y2=0
cc_177 N_B_c_185_n N_C_c_244_n 0.0181091f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_178 N_B_c_186_n N_C_c_244_n 0.0172417f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_179 N_B_M1015_g N_A_305_388#_c_302_n 3.40036e-19 $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B_M1014_g N_A_305_388#_c_318_n 0.012748f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_181 N_B_c_185_n N_A_305_388#_c_318_n 0.00325088f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_182 N_B_M1015_g N_A_305_388#_c_322_n 0.0122153f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B_M1015_g N_A_305_388#_c_304_n 0.0022446f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B_M1009_g N_A_305_388#_c_347_n 0.00116219f $X=0.955 $Y=2.44 $X2=0 $Y2=0
cc_185 N_B_M1014_g N_A_305_388#_c_347_n 3.69339e-19 $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_186 N_B_c_186_n N_A_305_388#_c_347_n 0.068687f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_187 N_B_c_186_n N_A_305_388#_c_307_n 0.00244434f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_188 N_B_M1009_g N_VPWR_c_464_n 0.00643693f $X=0.955 $Y=2.44 $X2=0 $Y2=0
cc_189 N_B_M1014_g N_VPWR_c_464_n 0.00643693f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_190 N_B_M1009_g N_VPWR_c_457_n 0.00647345f $X=0.955 $Y=2.44 $X2=0 $Y2=0
cc_191 N_B_M1014_g N_VPWR_c_457_n 0.00647345f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_192 N_B_c_186_n N_A_119_388#_c_526_n 0.0157027f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_193 N_B_M1009_g N_A_119_388#_c_533_n 0.0134246f $X=0.955 $Y=2.44 $X2=0 $Y2=0
cc_194 N_B_M1014_g N_A_119_388#_c_533_n 0.0117288f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_195 N_B_c_184_n N_A_119_388#_c_533_n 0.00128059f $X=0.97 $Y=1.615 $X2=0 $Y2=0
cc_196 N_B_c_186_n N_A_119_388#_c_533_n 0.0166516f $X=2.38 $Y=1.615 $X2=0 $Y2=0
cc_197 N_B_M1009_g N_A_209_388#_c_556_n 0.00389644f $X=0.955 $Y=2.44 $X2=0 $Y2=0
cc_198 N_B_M1014_g N_A_209_388#_c_556_n 0.00376081f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_199 N_B_M1015_g N_VGND_c_649_n 0.0065526f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B_M1015_g N_VGND_c_650_n 0.00413917f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B_M1015_g N_VGND_c_661_n 0.00399073f $X=2.44 $Y=0.74 $X2=0 $Y2=0
cc_202 N_C_c_243_n N_A_305_388#_c_302_n 0.0064141f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_203 N_C_c_245_n N_A_305_388#_c_302_n 0.004172f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_204 N_C_c_246_n N_A_305_388#_c_302_n 0.0331922f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_205 N_C_M1005_g N_A_305_388#_c_318_n 0.00912051f $X=1.885 $Y=2.44 $X2=0 $Y2=0
cc_206 N_C_c_243_n N_A_305_388#_c_322_n 0.00871095f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_207 N_C_c_243_n N_A_305_388#_c_303_n 7.15561e-19 $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_208 N_C_c_244_n N_A_305_388#_c_303_n 0.00114784f $X=1.885 $Y=1.345 $X2=0
+ $Y2=0
cc_209 N_C_c_245_n N_A_305_388#_c_303_n 0.00179824f $X=1.215 $Y=0.435 $X2=0
+ $Y2=0
cc_210 N_C_c_246_n N_A_305_388#_c_303_n 0.0143345f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_211 N_C_M1003_g N_A_305_388#_c_347_n 0.00592243f $X=1.435 $Y=2.44 $X2=0 $Y2=0
cc_212 N_C_M1005_g N_A_305_388#_c_347_n 0.00284815f $X=1.885 $Y=2.44 $X2=0 $Y2=0
cc_213 N_C_c_244_n N_A_305_388#_c_347_n 3.55714e-19 $X=1.885 $Y=1.345 $X2=0
+ $Y2=0
cc_214 N_C_M1003_g N_VPWR_c_464_n 0.00481634f $X=1.435 $Y=2.44 $X2=0 $Y2=0
cc_215 N_C_M1005_g N_VPWR_c_464_n 0.00481634f $X=1.885 $Y=2.44 $X2=0 $Y2=0
cc_216 N_C_M1003_g N_VPWR_c_457_n 0.00647345f $X=1.435 $Y=2.44 $X2=0 $Y2=0
cc_217 N_C_M1005_g N_VPWR_c_457_n 0.00647345f $X=1.885 $Y=2.44 $X2=0 $Y2=0
cc_218 N_C_M1003_g N_A_119_388#_c_533_n 0.0137958f $X=1.435 $Y=2.44 $X2=0 $Y2=0
cc_219 N_C_M1005_g N_A_119_388#_c_533_n 0.0123969f $X=1.885 $Y=2.44 $X2=0 $Y2=0
cc_220 N_C_M1003_g N_A_209_388#_c_556_n 0.0116356f $X=1.435 $Y=2.44 $X2=0 $Y2=0
cc_221 N_C_M1005_g N_A_209_388#_c_556_n 0.0116502f $X=1.885 $Y=2.44 $X2=0 $Y2=0
cc_222 N_C_c_243_n N_VGND_c_649_n 0.00349022f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_223 N_C_c_246_n N_VGND_c_649_n 0.00220313f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_224 N_C_c_243_n N_VGND_c_655_n 0.00434272f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_225 N_C_c_245_n N_VGND_c_655_n 0.00637453f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_226 N_C_c_246_n N_VGND_c_655_n 0.0203268f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_227 N_C_c_243_n N_VGND_c_661_n 0.00436049f $X=1.93 $Y=1.185 $X2=0 $Y2=0
cc_228 N_C_c_245_n N_VGND_c_661_n 0.00418281f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_229 N_C_c_246_n N_VGND_c_661_n 0.0124484f $X=1.215 $Y=0.435 $X2=0 $Y2=0
cc_230 N_A_305_388#_c_318_n N_VPWR_M1013_d 0.00852767f $X=3.225 $Y=2.035 $X2=0
+ $Y2=0
cc_231 N_A_305_388#_c_306_n N_VPWR_M1013_d 0.0013373f $X=3.31 $Y=1.95 $X2=0
+ $Y2=0
cc_232 N_A_305_388#_M1004_g N_VPWR_c_460_n 0.0130024f $X=3.425 $Y=2.4 $X2=0
+ $Y2=0
cc_233 N_A_305_388#_M1007_g N_VPWR_c_460_n 5.41206e-19 $X=3.875 $Y=2.4 $X2=0
+ $Y2=0
cc_234 N_A_305_388#_c_318_n N_VPWR_c_460_n 0.022405f $X=3.225 $Y=2.035 $X2=0
+ $Y2=0
cc_235 N_A_305_388#_M1004_g N_VPWR_c_461_n 5.90862e-19 $X=3.425 $Y=2.4 $X2=0
+ $Y2=0
cc_236 N_A_305_388#_M1007_g N_VPWR_c_461_n 0.0152536f $X=3.875 $Y=2.4 $X2=0
+ $Y2=0
cc_237 N_A_305_388#_M1011_g N_VPWR_c_461_n 0.00349416f $X=4.325 $Y=2.4 $X2=0
+ $Y2=0
cc_238 N_A_305_388#_M1012_g N_VPWR_c_463_n 0.00742848f $X=4.775 $Y=2.4 $X2=0
+ $Y2=0
cc_239 N_A_305_388#_M1004_g N_VPWR_c_465_n 0.00460063f $X=3.425 $Y=2.4 $X2=0
+ $Y2=0
cc_240 N_A_305_388#_M1007_g N_VPWR_c_465_n 0.00460063f $X=3.875 $Y=2.4 $X2=0
+ $Y2=0
cc_241 N_A_305_388#_M1011_g N_VPWR_c_466_n 0.005209f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A_305_388#_M1012_g N_VPWR_c_466_n 0.005209f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_305_388#_M1004_g N_VPWR_c_457_n 0.00908554f $X=3.425 $Y=2.4 $X2=0
+ $Y2=0
cc_244 N_A_305_388#_M1007_g N_VPWR_c_457_n 0.00908554f $X=3.875 $Y=2.4 $X2=0
+ $Y2=0
cc_245 N_A_305_388#_M1011_g N_VPWR_c_457_n 0.00982266f $X=4.325 $Y=2.4 $X2=0
+ $Y2=0
cc_246 N_A_305_388#_M1012_g N_VPWR_c_457_n 0.00986008f $X=4.775 $Y=2.4 $X2=0
+ $Y2=0
cc_247 N_A_305_388#_c_318_n N_A_119_388#_M1014_d 0.00643546f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_248 N_A_305_388#_M1003_d N_A_119_388#_c_533_n 0.00329511f $X=1.525 $Y=1.94
+ $X2=0 $Y2=0
cc_249 N_A_305_388#_c_318_n N_A_119_388#_c_533_n 0.0279204f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_250 N_A_305_388#_c_347_n N_A_119_388#_c_533_n 0.0157867f $X=1.825 $Y=2.075
+ $X2=0 $Y2=0
cc_251 N_A_305_388#_c_318_n N_A_119_388#_c_529_n 0.01898f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_252 N_A_305_388#_c_318_n N_A_209_388#_M1005_s 0.0048549f $X=3.225 $Y=2.035
+ $X2=0 $Y2=0
cc_253 N_A_305_388#_M1003_d N_A_209_388#_c_556_n 0.00168223f $X=1.525 $Y=1.94
+ $X2=0 $Y2=0
cc_254 N_A_305_388#_M1000_g N_X_c_570_n 0.00492137f $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_305_388#_M1002_g N_X_c_570_n 3.97599e-19 $X=3.865 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_305_388#_c_325_n N_X_c_570_n 0.0133617f $X=3.225 $Y=0.855 $X2=0 $Y2=0
cc_257 N_A_305_388#_c_305_n N_X_c_570_n 0.00133388f $X=3.31 $Y=1.3 $X2=0 $Y2=0
cc_258 N_A_305_388#_M1004_g N_X_c_577_n 3.62369e-19 $X=3.425 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A_305_388#_M1007_g N_X_c_577_n 3.62369e-19 $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_305_388#_M1002_g N_X_c_571_n 0.0127819f $X=3.865 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_305_388#_M1010_g N_X_c_571_n 0.0114326f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_305_388#_c_395_p N_X_c_571_n 0.0492576f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_263 N_A_305_388#_c_308_n N_X_c_571_n 0.00386308f $X=4.785 $Y=1.465 $X2=0
+ $Y2=0
cc_264 N_A_305_388#_M1000_g N_X_c_572_n 7.34064e-19 $X=3.43 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_305_388#_c_305_n N_X_c_572_n 0.0134529f $X=3.31 $Y=1.3 $X2=0 $Y2=0
cc_266 N_A_305_388#_c_395_p N_X_c_572_n 0.014338f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_267 N_A_305_388#_c_308_n N_X_c_572_n 0.00250521f $X=4.785 $Y=1.465 $X2=0
+ $Y2=0
cc_268 N_A_305_388#_M1007_g N_X_c_578_n 0.0146056f $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A_305_388#_M1011_g N_X_c_578_n 0.0128923f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A_305_388#_c_395_p N_X_c_578_n 0.0475485f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_271 N_A_305_388#_c_308_n N_X_c_578_n 0.00201785f $X=4.785 $Y=1.465 $X2=0
+ $Y2=0
cc_272 N_A_305_388#_M1004_g N_X_c_579_n 3.24225e-19 $X=3.425 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_305_388#_c_306_n N_X_c_579_n 0.0068918f $X=3.31 $Y=1.95 $X2=0 $Y2=0
cc_274 N_A_305_388#_c_395_p N_X_c_579_n 0.0143383f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_275 N_A_305_388#_c_308_n N_X_c_579_n 0.00209661f $X=4.785 $Y=1.465 $X2=0
+ $Y2=0
cc_276 N_A_305_388#_M1007_g N_X_c_580_n 7.7208e-19 $X=3.875 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A_305_388#_M1011_g N_X_c_580_n 0.0145011f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A_305_388#_M1012_g N_X_c_580_n 0.019068f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A_305_388#_M1002_g N_X_c_573_n 7.04495e-19 $X=3.865 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_305_388#_M1010_g N_X_c_573_n 0.00953543f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_305_388#_M1016_g N_X_c_573_n 3.97481e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_305_388#_M1016_g N_X_c_574_n 0.0160626f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A_305_388#_c_395_p N_X_c_574_n 0.00221753f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_284 N_A_305_388#_M1012_g N_X_c_581_n 0.0165256f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_285 N_A_305_388#_M1011_g N_X_c_582_n 0.00135419f $X=4.325 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A_305_388#_M1012_g N_X_c_582_n 0.0017715f $X=4.775 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A_305_388#_c_395_p N_X_c_582_n 0.0251683f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_288 N_A_305_388#_c_308_n N_X_c_582_n 0.00215577f $X=4.785 $Y=1.465 $X2=0
+ $Y2=0
cc_289 N_A_305_388#_M1010_g N_X_c_575_n 9.7541e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_305_388#_c_395_p N_X_c_575_n 0.0209731f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_291 N_A_305_388#_c_308_n N_X_c_575_n 0.00242817f $X=4.785 $Y=1.465 $X2=0
+ $Y2=0
cc_292 N_A_305_388#_M1016_g X 0.0067245f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A_305_388#_c_395_p X 0.0206535f $X=4.52 $Y=1.465 $X2=0 $Y2=0
cc_294 N_A_305_388#_c_308_n X 0.0172466f $X=4.785 $Y=1.465 $X2=0 $Y2=0
cc_295 N_A_305_388#_c_322_n N_VGND_M1008_d 0.00507735f $X=2.55 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_296 N_A_305_388#_c_325_n N_VGND_M1001_d 0.00807426f $X=3.225 $Y=0.855 $X2=0
+ $Y2=0
cc_297 N_A_305_388#_c_305_n N_VGND_M1001_d 0.00203236f $X=3.31 $Y=1.3 $X2=0
+ $Y2=0
cc_298 N_A_305_388#_c_302_n N_VGND_c_649_n 0.0101711f $X=1.715 $Y=0.515 $X2=0
+ $Y2=0
cc_299 N_A_305_388#_c_322_n N_VGND_c_649_n 0.0204503f $X=2.55 $Y=0.855 $X2=0
+ $Y2=0
cc_300 N_A_305_388#_c_304_n N_VGND_c_649_n 0.0101711f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_301 N_A_305_388#_c_304_n N_VGND_c_650_n 0.014415f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_305_388#_M1000_g N_VGND_c_651_n 0.00690871f $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_305_388#_M1002_g N_VGND_c_651_n 4.02157e-19 $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_305_388#_c_304_n N_VGND_c_651_n 0.0101711f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_305 N_A_305_388#_c_325_n N_VGND_c_651_n 0.0211625f $X=3.225 $Y=0.855 $X2=0
+ $Y2=0
cc_306 N_A_305_388#_M1000_g N_VGND_c_652_n 4.57455e-19 $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_307 N_A_305_388#_M1002_g N_VGND_c_652_n 0.00897549f $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_308 N_A_305_388#_M1010_g N_VGND_c_652_n 0.00497505f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A_305_388#_M1010_g N_VGND_c_654_n 5.12327e-19 $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_310 N_A_305_388#_M1016_g N_VGND_c_654_n 0.0110492f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_311 N_A_305_388#_c_302_n N_VGND_c_655_n 0.014415f $X=1.715 $Y=0.515 $X2=0
+ $Y2=0
cc_312 N_A_305_388#_M1000_g N_VGND_c_656_n 0.00383152f $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_313 N_A_305_388#_M1002_g N_VGND_c_656_n 0.00383152f $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_314 N_A_305_388#_M1010_g N_VGND_c_657_n 0.00434272f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_315 N_A_305_388#_M1016_g N_VGND_c_657_n 0.00383152f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_A_305_388#_M1000_g N_VGND_c_661_n 0.00708259f $X=3.43 $Y=0.74 $X2=0
+ $Y2=0
cc_317 N_A_305_388#_M1002_g N_VGND_c_661_n 0.0075759f $X=3.865 $Y=0.74 $X2=0
+ $Y2=0
cc_318 N_A_305_388#_M1010_g N_VGND_c_661_n 0.00821839f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_305_388#_M1016_g N_VGND_c_661_n 0.0075754f $X=4.785 $Y=0.74 $X2=0
+ $Y2=0
cc_320 N_A_305_388#_c_302_n N_VGND_c_661_n 0.0119404f $X=1.715 $Y=0.515 $X2=0
+ $Y2=0
cc_321 N_A_305_388#_c_322_n N_VGND_c_661_n 0.0118074f $X=2.55 $Y=0.855 $X2=0
+ $Y2=0
cc_322 N_A_305_388#_c_304_n N_VGND_c_661_n 0.0119404f $X=2.715 $Y=0.515 $X2=0
+ $Y2=0
cc_323 N_A_305_388#_c_325_n N_VGND_c_661_n 0.00714277f $X=3.225 $Y=0.855 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_459_n N_A_119_388#_c_524_n 0.0139051f $X=0.28 $Y=2.085 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_464_n N_A_119_388#_c_524_n 0.0101587f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_457_n N_A_119_388#_c_524_n 0.00902356f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_457_n N_A_119_388#_c_533_n 0.0141151f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_460_n N_A_119_388#_c_525_n 0.0142276f $X=3.2 $Y=2.455 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_464_n N_A_119_388#_c_525_n 0.0134483f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_457_n N_A_119_388#_c_525_n 0.0119361f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_464_n N_A_209_388#_c_556_n 0.0493699f $X=3.035 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_457_n N_A_209_388#_c_556_n 0.046043f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_333 N_VPWR_c_460_n N_X_c_577_n 0.0233699f $X=3.2 $Y=2.455 $X2=0 $Y2=0
cc_334 N_VPWR_c_461_n N_X_c_577_n 0.0271589f $X=4.1 $Y=2.305 $X2=0 $Y2=0
cc_335 N_VPWR_c_465_n N_X_c_577_n 0.00749631f $X=3.935 $Y=3.33 $X2=0 $Y2=0
cc_336 N_VPWR_c_457_n N_X_c_577_n 0.0062048f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_337 N_VPWR_M1007_s N_X_c_578_n 0.00165831f $X=3.965 $Y=1.84 $X2=0 $Y2=0
cc_338 N_VPWR_c_461_n N_X_c_578_n 0.0148589f $X=4.1 $Y=2.305 $X2=0 $Y2=0
cc_339 N_VPWR_c_461_n N_X_c_580_n 0.0283501f $X=4.1 $Y=2.305 $X2=0 $Y2=0
cc_340 N_VPWR_c_463_n N_X_c_580_n 0.0283501f $X=5 $Y=2.305 $X2=0 $Y2=0
cc_341 N_VPWR_c_466_n N_X_c_580_n 0.0144623f $X=4.915 $Y=3.33 $X2=0 $Y2=0
cc_342 N_VPWR_c_457_n N_X_c_580_n 0.0118344f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_343 N_VPWR_M1012_s N_X_c_581_n 0.00315413f $X=4.865 $Y=1.84 $X2=0 $Y2=0
cc_344 N_VPWR_c_463_n N_X_c_581_n 0.0207257f $X=5 $Y=2.305 $X2=0 $Y2=0
cc_345 N_A_119_388#_c_533_n N_A_209_388#_M1009_s 0.00552585f $X=2.5 $Y=2.455
+ $X2=-0.19 $Y2=1.66
cc_346 N_A_119_388#_c_533_n N_A_209_388#_M1005_s 0.00484434f $X=2.5 $Y=2.455
+ $X2=0 $Y2=0
cc_347 N_A_119_388#_c_524_n N_A_209_388#_c_556_n 0.00980844f $X=0.73 $Y=2.795
+ $X2=0 $Y2=0
cc_348 N_A_119_388#_c_533_n N_A_209_388#_c_556_n 0.068494f $X=2.5 $Y=2.455 $X2=0
+ $Y2=0
cc_349 N_A_119_388#_c_525_n N_A_209_388#_c_556_n 0.0111988f $X=2.665 $Y=2.795
+ $X2=0 $Y2=0
cc_350 N_X_c_571_n N_VGND_M1002_s 0.00402642f $X=4.405 $Y=1.045 $X2=0 $Y2=0
cc_351 N_X_c_574_n N_VGND_M1016_s 0.00338075f $X=4.925 $Y=1.045 $X2=0 $Y2=0
cc_352 N_X_c_570_n N_VGND_c_651_n 0.0173183f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_353 N_X_c_570_n N_VGND_c_652_n 0.0157999f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_354 N_X_c_571_n N_VGND_c_652_n 0.0154151f $X=4.405 $Y=1.045 $X2=0 $Y2=0
cc_355 N_X_c_573_n N_VGND_c_652_n 0.0251662f $X=4.57 $Y=0.515 $X2=0 $Y2=0
cc_356 N_X_c_573_n N_VGND_c_654_n 0.0164981f $X=4.57 $Y=0.515 $X2=0 $Y2=0
cc_357 N_X_c_574_n N_VGND_c_654_n 0.023173f $X=4.925 $Y=1.045 $X2=0 $Y2=0
cc_358 N_X_c_570_n N_VGND_c_656_n 0.00749631f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_359 N_X_c_573_n N_VGND_c_657_n 0.0109942f $X=4.57 $Y=0.515 $X2=0 $Y2=0
cc_360 N_X_c_570_n N_VGND_c_661_n 0.0062048f $X=3.65 $Y=0.515 $X2=0 $Y2=0
cc_361 N_X_c_573_n N_VGND_c_661_n 0.00904371f $X=4.57 $Y=0.515 $X2=0 $Y2=0

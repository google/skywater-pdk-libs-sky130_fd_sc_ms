* File: sky130_fd_sc_ms__or2_4.pxi.spice
* Created: Fri Aug 28 18:06:31 2020
* 
x_PM_SKY130_FD_SC_MS__OR2_4%A_83_260# N_A_83_260#_M1004_d N_A_83_260#_M1007_d
+ N_A_83_260#_M1001_g N_A_83_260#_M1008_g N_A_83_260#_M1009_g
+ N_A_83_260#_M1002_g N_A_83_260#_M1012_g N_A_83_260#_M1003_g
+ N_A_83_260#_M1006_g N_A_83_260#_M1013_g N_A_83_260#_c_162_p N_A_83_260#_c_89_n
+ N_A_83_260#_c_90_n N_A_83_260#_c_91_n N_A_83_260#_c_108_p N_A_83_260#_c_100_n
+ N_A_83_260#_c_113_p N_A_83_260#_c_92_n N_A_83_260#_c_93_n N_A_83_260#_c_94_n
+ N_A_83_260#_c_95_n PM_SKY130_FD_SC_MS__OR2_4%A_83_260#
x_PM_SKY130_FD_SC_MS__OR2_4%A N_A_M1004_g N_A_M1005_g N_A_M1011_g N_A_c_235_n
+ N_A_c_216_n N_A_c_217_n A N_A_c_219_n PM_SKY130_FD_SC_MS__OR2_4%A
x_PM_SKY130_FD_SC_MS__OR2_4%B N_B_M1007_g N_B_M1000_g N_B_M1010_g B N_B_c_296_n
+ PM_SKY130_FD_SC_MS__OR2_4%B
x_PM_SKY130_FD_SC_MS__OR2_4%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1006_s
+ N_VPWR_M1011_s N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n VPWR
+ N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n N_VPWR_c_338_n
+ PM_SKY130_FD_SC_MS__OR2_4%VPWR
x_PM_SKY130_FD_SC_MS__OR2_4%X N_X_M1008_d N_X_M1012_d N_X_M1001_d N_X_M1003_d
+ N_X_c_397_n N_X_c_398_n N_X_c_404_n N_X_c_405_n N_X_c_399_n N_X_c_406_n
+ N_X_c_400_n N_X_c_407_n N_X_c_401_n N_X_c_408_n N_X_c_402_n N_X_c_409_n X X
+ PM_SKY130_FD_SC_MS__OR2_4%X
x_PM_SKY130_FD_SC_MS__OR2_4%A_496_388# N_A_496_388#_M1005_d N_A_496_388#_M1010_s
+ N_A_496_388#_c_483_n N_A_496_388#_c_473_n N_A_496_388#_c_474_n
+ N_A_496_388#_c_475_n PM_SKY130_FD_SC_MS__OR2_4%A_496_388#
x_PM_SKY130_FD_SC_MS__OR2_4%VGND N_VGND_M1008_s N_VGND_M1009_s N_VGND_M1013_s
+ N_VGND_M1000_d N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n N_VGND_c_505_n
+ N_VGND_c_506_n N_VGND_c_507_n VGND N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n PM_SKY130_FD_SC_MS__OR2_4%VGND
cc_1 VNB N_A_83_260#_M1001_g 0.00167778f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_260#_M1008_g 0.0224607f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_A_83_260#_M1009_g 0.0203442f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_A_83_260#_M1002_g 0.00154206f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_5 VNB N_A_83_260#_M1012_g 0.02196f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_6 VNB N_A_83_260#_M1003_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_7 VNB N_A_83_260#_M1006_g 0.00158577f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_8 VNB N_A_83_260#_M1013_g 0.0216596f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_9 VNB N_A_83_260#_c_89_n 0.00648005f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_10 VNB N_A_83_260#_c_90_n 0.0028029f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.515
cc_11 VNB N_A_83_260#_c_91_n 0.0303098f $X=-0.19 $Y=-0.245 $X2=4.065 $Y2=1.095
cc_12 VNB N_A_83_260#_c_92_n 0.0298057f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=2.29
cc_13 VNB N_A_83_260#_c_93_n 0.00625835f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.095
cc_14 VNB N_A_83_260#_c_94_n 0.00255036f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.095
cc_15 VNB N_A_83_260#_c_95_n 0.0827101f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.465
cc_16 VNB N_A_M1004_g 0.0256588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_c_216_n 0.00338952f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_18 VNB N_A_c_217_n 0.0260565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A 0.0080355f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_20 VNB N_A_c_219_n 0.0234792f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.3
cc_21 VNB N_B_M1000_g 0.0399583f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_22 VNB B 0.00357747f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_23 VNB N_B_c_296_n 0.0332168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_338_n 0.183584f $X=-0.19 $Y=-0.245 $X2=4.065 $Y2=2.375
cc_25 VNB N_X_c_397_n 9.41836e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_26 VNB N_X_c_398_n 0.00715794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_399_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.63
cc_28 VNB N_X_c_400_n 0.00485313f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.63
cc_29 VNB N_X_c_401_n 0.0025013f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_30 VNB N_X_c_402_n 0.0019324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB X 0.0264101f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.465
cc_32 VNB N_VGND_c_502_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_33 VNB N_VGND_c_503_n 0.0274133f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_34 VNB N_VGND_c_504_n 0.00497771f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.63
cc_35 VNB N_VGND_c_505_n 0.00571437f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.3
cc_36 VNB N_VGND_c_506_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_507_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.63
cc_38 VNB N_VGND_c_508_n 0.0196058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_509_n 0.0185359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_510_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_41 VNB N_VGND_c_511_n 0.070232f $X=-0.19 $Y=-0.245 $X2=3.105 $Y2=2.46
cc_42 VNB N_VGND_c_512_n 0.248241f $X=-0.19 $Y=-0.245 $X2=4.065 $Y2=2.375
cc_43 VPB N_A_83_260#_M1001_g 0.0240093f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_44 VPB N_A_83_260#_M1002_g 0.0220562f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_45 VPB N_A_83_260#_M1003_g 0.0220607f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_46 VPB N_A_83_260#_M1006_g 0.0237237f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_47 VPB N_A_83_260#_c_100_n 0.00863795f $X=-0.19 $Y=1.66 $X2=4.065 $Y2=2.375
cc_48 VPB N_A_83_260#_c_92_n 0.0255791f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=2.29
cc_49 VPB N_A_M1005_g 0.0241659f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_50 VPB N_A_M1011_g 0.0219077f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_51 VPB N_A_c_216_n 0.00317406f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_52 VPB N_A_c_217_n 0.0133814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB A 0.00202237f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_54 VPB N_A_c_219_n 0.00544607f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.3
cc_55 VPB N_B_M1007_g 0.0186912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_B_M1010_g 0.0201791f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_57 VPB B 8.34758e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_58 VPB N_B_c_296_n 0.0141172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_339_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_60 VPB N_VPWR_c_340_n 0.0428715f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_61 VPB N_VPWR_c_341_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.63
cc_62 VPB N_VPWR_c_342_n 0.0090227f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.3
cc_63 VPB N_VPWR_c_343_n 0.011133f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_64 VPB N_VPWR_c_344_n 0.0252905f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.63
cc_65 VPB N_VPWR_c_345_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_346_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.63
cc_67 VPB N_VPWR_c_347_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_348_n 0.0412895f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.465
cc_69 VPB N_VPWR_c_349_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=1.095
cc_70 VPB N_VPWR_c_338_n 0.0776071f $X=-0.19 $Y=1.66 $X2=4.065 $Y2=2.375
cc_71 VPB N_X_c_404_n 8.97027e-19 $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_72 VPB N_X_c_405_n 0.00721884f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_73 VPB N_X_c_406_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.3
cc_74 VPB N_X_c_407_n 0.00443716f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_75 VPB N_X_c_408_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_76 VPB N_X_c_409_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.465
cc_77 VPB X 0.00682831f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.465
cc_78 VPB N_A_496_388#_c_473_n 0.00467397f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_79 VPB N_A_496_388#_c_474_n 0.00244128f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_80 VPB N_A_496_388#_c_475_n 0.00265994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 N_A_83_260#_M1013_g N_A_M1004_g 0.0274315f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_82 N_A_83_260#_c_89_n N_A_M1004_g 0.0110153f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_83_260#_c_90_n N_A_M1004_g 0.00943664f $X=2.585 $Y=0.515 $X2=0 $Y2=0
cc_84 N_A_83_260#_c_93_n N_A_M1004_g 0.00344278f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_85 N_A_83_260#_c_94_n N_A_M1004_g 0.0016818f $X=2.585 $Y=1.095 $X2=0 $Y2=0
cc_86 N_A_83_260#_M1006_g N_A_M1005_g 0.0283699f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_83_260#_c_108_p N_A_M1011_g 7.27256e-19 $X=3.105 $Y=2.46 $X2=0 $Y2=0
cc_88 N_A_83_260#_c_100_n N_A_M1011_g 0.0178278f $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_89 N_A_83_260#_c_92_n N_A_M1011_g 0.00815828f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_90 N_A_83_260#_M1007_d N_A_c_235_n 0.00311147f $X=2.93 $Y=1.94 $X2=0 $Y2=0
cc_91 N_A_83_260#_c_100_n N_A_c_235_n 0.0391662f $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_92 N_A_83_260#_c_113_p N_A_c_235_n 0.0144741f $X=3.23 $Y=2.375 $X2=0 $Y2=0
cc_93 N_A_83_260#_c_91_n N_A_c_216_n 0.0170702f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_94 N_A_83_260#_c_92_n N_A_c_216_n 0.0375788f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_95 N_A_83_260#_c_91_n N_A_c_217_n 0.00280278f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_96 N_A_83_260#_c_100_n N_A_c_217_n 3.04749e-19 $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_97 N_A_83_260#_c_92_n N_A_c_217_n 0.00761916f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_98 N_A_83_260#_M1006_g A 0.00454408f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_83_260#_c_89_n A 0.0161138f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_100 N_A_83_260#_c_91_n A 3.8449e-19 $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_101 N_A_83_260#_c_93_n A 0.0219858f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_102 N_A_83_260#_c_94_n A 0.0301826f $X=2.585 $Y=1.095 $X2=0 $Y2=0
cc_103 N_A_83_260#_c_95_n A 2.95273e-19 $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_104 N_A_83_260#_c_89_n N_A_c_219_n 5.99205e-19 $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_105 N_A_83_260#_c_93_n N_A_c_219_n 8.67352e-19 $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_106 N_A_83_260#_c_94_n N_A_c_219_n 7.48593e-19 $X=2.585 $Y=1.095 $X2=0 $Y2=0
cc_107 N_A_83_260#_c_95_n N_A_c_219_n 0.0159136f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_108 N_A_83_260#_c_90_n N_B_M1000_g 4.78879e-19 $X=2.585 $Y=0.515 $X2=0 $Y2=0
cc_109 N_A_83_260#_c_91_n N_B_M1000_g 0.0200689f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_110 N_A_83_260#_c_108_p N_B_M1010_g 0.00511267f $X=3.105 $Y=2.46 $X2=0 $Y2=0
cc_111 N_A_83_260#_c_100_n N_B_M1010_g 0.0100353f $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_112 N_A_83_260#_c_113_p N_B_M1010_g 0.00109776f $X=3.23 $Y=2.375 $X2=0 $Y2=0
cc_113 N_A_83_260#_c_91_n B 0.0174918f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_114 N_A_83_260#_c_91_n N_B_c_296_n 0.00670847f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_115 N_A_83_260#_c_100_n N_VPWR_M1011_s 0.00867901f $X=4.065 $Y=2.375 $X2=0
+ $Y2=0
cc_116 N_A_83_260#_c_92_n N_VPWR_M1011_s 0.0057645f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_117 N_A_83_260#_M1001_g N_VPWR_c_340_n 0.00742848f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_118 N_A_83_260#_M1002_g N_VPWR_c_341_n 0.00329146f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_119 N_A_83_260#_M1003_g N_VPWR_c_341_n 0.00329146f $X=1.405 $Y=2.4 $X2=0
+ $Y2=0
cc_120 N_A_83_260#_M1006_g N_VPWR_c_342_n 0.00417147f $X=1.855 $Y=2.4 $X2=0
+ $Y2=0
cc_121 N_A_83_260#_c_93_n N_VPWR_c_342_n 0.00170784f $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_122 N_A_83_260#_c_100_n N_VPWR_c_344_n 0.022932f $X=4.065 $Y=2.375 $X2=0
+ $Y2=0
cc_123 N_A_83_260#_M1001_g N_VPWR_c_345_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_83_260#_M1002_g N_VPWR_c_345_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_83_260#_M1003_g N_VPWR_c_347_n 0.005209f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_83_260#_M1006_g N_VPWR_c_347_n 0.005209f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_83_260#_M1001_g N_VPWR_c_338_n 0.00986008f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_128 N_A_83_260#_M1002_g N_VPWR_c_338_n 0.00982266f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_129 N_A_83_260#_M1003_g N_VPWR_c_338_n 0.00982266f $X=1.405 $Y=2.4 $X2=0
+ $Y2=0
cc_130 N_A_83_260#_M1006_g N_VPWR_c_338_n 0.00987399f $X=1.855 $Y=2.4 $X2=0
+ $Y2=0
cc_131 N_A_83_260#_M1008_g N_X_c_397_n 0.0143395f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_83_260#_M1001_g N_X_c_404_n 0.0165252f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_83_260#_M1008_g N_X_c_399_n 0.0128625f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_83_260#_M1009_g N_X_c_399_n 3.97481e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_83_260#_M1001_g N_X_c_406_n 0.019068f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_83_260#_M1002_g N_X_c_406_n 0.0143027f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_83_260#_M1003_g N_X_c_406_n 6.97946e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_83_260#_M1009_g N_X_c_400_n 0.0124434f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_83_260#_M1012_g N_X_c_400_n 0.0121215f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_83_260#_M1013_g N_X_c_400_n 0.00257018f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_83_260#_c_162_p N_X_c_400_n 0.0695156f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_142 N_A_83_260#_c_93_n N_X_c_400_n 0.0095065f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_143 N_A_83_260#_c_95_n N_X_c_400_n 0.00696755f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_144 N_A_83_260#_M1002_g N_X_c_407_n 0.012931f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_83_260#_M1003_g N_X_c_407_n 0.0142852f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_83_260#_M1006_g N_X_c_407_n 0.00385266f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_83_260#_c_162_p N_X_c_407_n 0.0692143f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_148 N_A_83_260#_c_95_n N_X_c_407_n 0.00425236f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_149 N_A_83_260#_M1009_g N_X_c_401_n 6.70758e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_83_260#_M1012_g N_X_c_401_n 0.00887699f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_83_260#_M1013_g N_X_c_401_n 0.00731762f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_83_260#_M1002_g N_X_c_408_n 6.97946e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_83_260#_M1003_g N_X_c_408_n 0.0143027f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_83_260#_M1006_g N_X_c_408_n 0.0144734f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_83_260#_M1008_g N_X_c_402_n 0.00132305f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_83_260#_c_162_p N_X_c_402_n 0.0168687f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_157 N_A_83_260#_c_95_n N_X_c_402_n 0.00242817f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_158 N_A_83_260#_M1001_g N_X_c_409_n 0.00177079f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_83_260#_M1002_g N_X_c_409_n 0.00135419f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_83_260#_c_162_p N_X_c_409_n 0.0251683f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A_83_260#_c_95_n N_X_c_409_n 0.00215577f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A_83_260#_M1008_g X 0.0067245f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_83_260#_c_162_p X 0.0206535f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_164 N_A_83_260#_c_95_n X 0.0172466f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_165 N_A_83_260#_c_100_n N_A_496_388#_M1010_s 0.00431308f $X=4.065 $Y=2.375
+ $X2=0 $Y2=0
cc_166 N_A_83_260#_M1007_d N_A_496_388#_c_473_n 0.00165831f $X=2.93 $Y=1.94
+ $X2=0 $Y2=0
cc_167 N_A_83_260#_c_108_p N_A_496_388#_c_473_n 0.0134956f $X=3.105 $Y=2.46
+ $X2=0 $Y2=0
cc_168 N_A_83_260#_c_100_n N_A_496_388#_c_473_n 0.0046334f $X=4.065 $Y=2.375
+ $X2=0 $Y2=0
cc_169 N_A_83_260#_c_100_n N_A_496_388#_c_475_n 0.0182896f $X=4.065 $Y=2.375
+ $X2=0 $Y2=0
cc_170 N_A_83_260#_c_89_n N_VGND_M1013_s 0.0023395f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_171 N_A_83_260#_c_93_n N_VGND_M1013_s 6.54518e-19 $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_172 N_A_83_260#_c_91_n N_VGND_M1000_d 0.0186685f $X=4.065 $Y=1.095 $X2=0
+ $Y2=0
cc_173 N_A_83_260#_M1008_g N_VGND_c_503_n 0.00409307f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_83_260#_M1008_g N_VGND_c_504_n 5.05592e-19 $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_83_260#_M1009_g N_VGND_c_504_n 0.008885f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_83_260#_M1012_g N_VGND_c_504_n 0.00307459f $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_83_260#_M1012_g N_VGND_c_505_n 7.0576e-19 $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_83_260#_M1013_g N_VGND_c_505_n 0.0114822f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_83_260#_c_89_n N_VGND_c_505_n 0.016109f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_180 N_A_83_260#_c_90_n N_VGND_c_505_n 0.0191765f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_181 N_A_83_260#_c_93_n N_VGND_c_505_n 0.00528841f $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_182 N_A_83_260#_M1008_g N_VGND_c_506_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_83_260#_M1009_g N_VGND_c_506_n 0.00383152f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_83_260#_M1012_g N_VGND_c_508_n 0.00434272f $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A_83_260#_M1013_g N_VGND_c_508_n 0.00383152f $X=1.87 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_83_260#_c_90_n N_VGND_c_509_n 0.0145639f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_187 N_A_83_260#_c_90_n N_VGND_c_511_n 0.0214346f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_83_260#_c_91_n N_VGND_c_511_n 0.101081f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_189 N_A_83_260#_M1008_g N_VGND_c_512_n 0.00823942f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_83_260#_M1009_g N_VGND_c_512_n 0.0075754f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_83_260#_M1012_g N_VGND_c_512_n 0.00821072f $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_83_260#_M1013_g N_VGND_c_512_n 0.00758328f $X=1.87 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_83_260#_c_90_n N_VGND_c_512_n 0.0119984f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_194 N_A_c_235_n N_B_M1007_g 0.0191126f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_195 A N_B_M1007_g 0.00670077f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A_M1004_g N_B_M1000_g 0.0160308f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_197 A N_B_M1000_g 0.00466058f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A_c_219_n N_B_M1000_g 0.0144774f $X=2.375 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A_M1011_g N_B_M1010_g 0.0367438f $X=3.79 $Y=2.44 $X2=0 $Y2=0
cc_200 N_A_c_235_n N_B_M1010_g 0.0151741f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_201 N_A_c_216_n N_B_M1010_g 0.0038244f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_202 A N_B_M1010_g 7.6463e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_c_235_n B 0.0200424f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_204 N_A_c_216_n B 0.0142939f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_205 N_A_c_217_n B 0.00116857f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_206 A B 0.0266673f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A_M1005_g N_B_c_296_n 0.033055f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_208 N_A_c_235_n N_B_c_296_n 6.34453e-19 $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_209 N_A_c_216_n N_B_c_296_n 0.00142915f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_210 N_A_c_217_n N_B_c_296_n 0.0161869f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_211 A N_B_c_296_n 0.00393808f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A_c_219_n N_B_c_296_n 0.00325514f $X=2.375 $Y=1.515 $X2=0 $Y2=0
cc_213 A N_VPWR_M1006_s 0.0018048f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A_M1005_g N_VPWR_c_342_n 0.00558205f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_215 A N_VPWR_c_342_n 0.00294797f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_216 N_A_M1011_g N_VPWR_c_344_n 0.00307938f $X=3.79 $Y=2.44 $X2=0 $Y2=0
cc_217 N_A_M1005_g N_VPWR_c_348_n 0.00582583f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_218 N_A_M1011_g N_VPWR_c_348_n 0.005857f $X=3.79 $Y=2.44 $X2=0 $Y2=0
cc_219 N_A_M1005_g N_VPWR_c_338_n 0.00539454f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_220 N_A_M1011_g N_VPWR_c_338_n 0.0054305f $X=3.79 $Y=2.44 $X2=0 $Y2=0
cc_221 N_A_M1005_g N_X_c_407_n 2.29539e-19 $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_222 A N_X_c_407_n 0.00651558f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A_M1005_g N_X_c_408_n 9.08651e-19 $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_224 A N_A_496_388#_M1005_d 0.00172633f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_225 N_A_c_235_n N_A_496_388#_M1010_s 0.00799597f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_226 N_A_M1005_g N_A_496_388#_c_483_n 0.00805456f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_227 N_A_c_235_n N_A_496_388#_c_483_n 0.00179416f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_228 A N_A_496_388#_c_483_n 0.0158107f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_229 N_A_M1005_g N_A_496_388#_c_474_n 0.00390371f $X=2.39 $Y=2.44 $X2=0 $Y2=0
cc_230 N_A_M1011_g N_A_496_388#_c_475_n 0.0077794f $X=3.79 $Y=2.44 $X2=0 $Y2=0
cc_231 N_A_M1004_g N_VGND_c_505_n 0.00432719f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_M1004_g N_VGND_c_509_n 0.00434272f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_M1004_g N_VGND_c_511_n 4.84975e-19 $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_M1004_g N_VGND_c_512_n 0.00821358f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B_M1007_g N_VPWR_c_348_n 0.00117044f $X=2.84 $Y=2.44 $X2=0 $Y2=0
cc_236 N_B_M1010_g N_VPWR_c_348_n 0.00115138f $X=3.29 $Y=2.44 $X2=0 $Y2=0
cc_237 N_B_M1007_g N_A_496_388#_c_483_n 0.00898288f $X=2.84 $Y=2.44 $X2=0 $Y2=0
cc_238 N_B_M1010_g N_A_496_388#_c_483_n 6.69226e-19 $X=3.29 $Y=2.44 $X2=0 $Y2=0
cc_239 N_B_M1007_g N_A_496_388#_c_473_n 0.0128118f $X=2.84 $Y=2.44 $X2=0 $Y2=0
cc_240 N_B_M1010_g N_A_496_388#_c_473_n 0.0115928f $X=3.29 $Y=2.44 $X2=0 $Y2=0
cc_241 N_B_M1007_g N_A_496_388#_c_474_n 0.00234159f $X=2.84 $Y=2.44 $X2=0 $Y2=0
cc_242 N_B_M1010_g N_A_496_388#_c_475_n 4.70101e-19 $X=3.29 $Y=2.44 $X2=0 $Y2=0
cc_243 N_B_M1000_g N_VGND_c_509_n 0.00429299f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B_M1000_g N_VGND_c_511_n 0.0126649f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B_M1000_g N_VGND_c_512_n 0.00843495f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_246 N_VPWR_M1001_s N_X_c_405_n 0.00315413f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_247 N_VPWR_c_340_n N_X_c_405_n 0.0207257f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_248 N_VPWR_c_340_n N_X_c_406_n 0.0283501f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_249 N_VPWR_c_341_n N_X_c_406_n 0.0283117f $X=1.18 $Y=2.305 $X2=0 $Y2=0
cc_250 N_VPWR_c_345_n N_X_c_406_n 0.0144623f $X=1.095 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_c_338_n N_X_c_406_n 0.0118344f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_M1002_s N_X_c_407_n 0.00165831f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_253 N_VPWR_c_341_n N_X_c_407_n 0.0126919f $X=1.18 $Y=2.305 $X2=0 $Y2=0
cc_254 N_VPWR_c_341_n N_X_c_408_n 0.0283117f $X=1.18 $Y=2.305 $X2=0 $Y2=0
cc_255 N_VPWR_c_342_n N_X_c_408_n 0.029009f $X=2.08 $Y=2.285 $X2=0 $Y2=0
cc_256 N_VPWR_c_347_n N_X_c_408_n 0.0144623f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_338_n N_X_c_408_n 0.0118344f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_258 N_VPWR_c_348_n N_A_496_388#_c_473_n 0.0399102f $X=3.93 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_338_n N_A_496_388#_c_473_n 0.0233066f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_342_n N_A_496_388#_c_474_n 0.0108854f $X=2.08 $Y=2.285 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_348_n N_A_496_388#_c_474_n 0.0236566f $X=3.93 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_338_n N_A_496_388#_c_474_n 0.0128296f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_344_n N_A_496_388#_c_475_n 0.019519f $X=4.025 $Y=2.795 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_348_n N_A_496_388#_c_475_n 0.0227798f $X=3.93 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_338_n N_A_496_388#_c_475_n 0.0126147f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_266 N_X_c_398_n N_VGND_M1008_s 0.00330634f $X=0.355 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_267 N_X_c_400_n N_VGND_M1009_s 0.00176461f $X=1.405 $Y=1.045 $X2=0 $Y2=0
cc_268 N_X_c_397_n N_VGND_c_503_n 6.14392e-19 $X=0.545 $Y=1.045 $X2=0 $Y2=0
cc_269 N_X_c_398_n N_VGND_c_503_n 0.0207726f $X=0.355 $Y=1.045 $X2=0 $Y2=0
cc_270 N_X_c_399_n N_VGND_c_503_n 0.0158413f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_271 N_X_c_399_n N_VGND_c_504_n 0.0158413f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_272 N_X_c_400_n N_VGND_c_504_n 0.0153337f $X=1.405 $Y=1.045 $X2=0 $Y2=0
cc_273 N_X_c_401_n N_VGND_c_504_n 0.0162297f $X=1.59 $Y=0.515 $X2=0 $Y2=0
cc_274 N_X_c_401_n N_VGND_c_505_n 0.0309614f $X=1.59 $Y=0.515 $X2=0 $Y2=0
cc_275 N_X_c_399_n N_VGND_c_506_n 0.0109942f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_276 N_X_c_401_n N_VGND_c_508_n 0.0130022f $X=1.59 $Y=0.515 $X2=0 $Y2=0
cc_277 N_X_c_399_n N_VGND_c_512_n 0.00904371f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_278 N_X_c_401_n N_VGND_c_512_n 0.0107057f $X=1.59 $Y=0.515 $X2=0 $Y2=0

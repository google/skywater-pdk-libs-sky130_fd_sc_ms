* File: sky130_fd_sc_ms__nand4b_1.spice
* Created: Wed Sep  2 12:14:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4b_1.pex.spice"
.subckt sky130_fd_sc_ms__nand4b_1  VNB VPB A_N D C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_N_M1006_g N_A_27_112#_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.114946 AS=0.2695 PD=0.963566 PS=2.08 NRD=23.988 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1008 A_263_74# N_D_M1008_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.154654 PD=0.98 PS=1.29643 NRD=10.536 NRS=0.804 M=1 R=4.93333 SA=75000.8
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1009 A_341_74# N_C_M1009_g A_263_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1332
+ AS=0.0888 PD=1.1 PS=0.98 NRD=20.268 NRS=10.536 M=1 R=4.93333 SA=75001.2
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1002 A_443_74# N_B_M1002_g A_341_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.1332 PD=1.13 PS=1.1 NRD=22.692 NRS=20.268 M=1 R=4.93333 SA=75001.7
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_A_27_112#_M1003_g A_443_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.3404 AS=0.1443 PD=2.4 PS=1.13 NRD=15.396 NRS=22.692 M=1 R=4.93333
+ SA=75002.2 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_27_112#_M1004_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1854 AS=0.2352 PD=1.30714 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1005 N_Y_M1005_d N_D_M1005_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2472 PD=1.39 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_C_M1007_g N_Y_M1005_d VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1512 PD=1.51 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90001.3
+ A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2184 PD=1.39 PS=1.51 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90001.7 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_27_112#_M1001_g N_Y_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__nand4b_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sedfxtp_2.pex.spice
* Created: Wed Sep  2 12:32:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%D 3 7 11 12 17 18 20 22
c39 22 0 2.2081e-19 $X=0.525 $Y=1.99
c40 17 0 1.59585e-19 $X=0.525 $Y=1.145
r41 20 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.825
+ $X2=0.525 $Y2=1.99
r42 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.825 $X2=0.525 $Y2=1.825
r43 17 20 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.525 $Y=1.145
+ $X2=0.525 $Y2=1.825
r44 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.145 $X2=0.525 $Y2=1.145
r45 12 21 4.85239 $w=3.78e-07 $l=1.6e-07 $layer=LI1_cond $X=0.615 $Y=1.665
+ $X2=0.615 $Y2=1.825
r46 11 12 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.665
r47 11 18 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.145
r48 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=0.98
+ $X2=0.525 $Y2=1.145
r49 7 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.615 $Y=0.58 $X2=0.615
+ $Y2=0.98
r50 3 22 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=0.57 $Y=2.64 $X2=0.57
+ $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_180_290# 1 2 9 13 16 20 21 22 23 24 25
+ 28 32 34 36 46
c106 46 0 1.26127e-19 $X=2.425 $Y=1.685
c107 36 0 7.02076e-20 $X=2.22 $Y=1.685
c108 34 0 7.48038e-20 $X=2.22 $Y=1.95
c109 25 0 3.52195e-20 $X=1.305 $Y=2.035
c110 23 0 1.59585e-19 $X=1.305 $Y=1.065
c111 21 0 1.74672e-19 $X=1.14 $Y=1.615
r112 37 46 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.22 $Y=1.685
+ $X2=2.425 $Y2=1.685
r113 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.685 $X2=2.22 $Y2=1.685
r114 34 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.22 $Y=2.035
+ $X2=1.895 $Y2=2.035
r115 34 36 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=1.95
+ $X2=2.22 $Y2=1.685
r116 30 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=2.12
+ $X2=1.895 $Y2=2.035
r117 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.895 $Y=2.12
+ $X2=1.895 $Y2=2.515
r118 26 28 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.74 $Y=0.98
+ $X2=1.74 $Y2=0.775
r119 24 39 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=2.035
+ $X2=1.895 $Y2=2.035
r120 24 25 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.81 $Y=2.035
+ $X2=1.305 $Y2=2.035
r121 22 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=1.74 $Y2=0.98
r122 22 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=1.305 $Y2=1.065
r123 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.615 $X2=1.14 $Y2=1.615
r124 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.305 $Y2=2.035
r125 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.14 $Y2=1.615
r126 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.305 $Y2=1.065
r127 17 20 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.14 $Y2=1.615
r128 15 21 41.6085 $w=4.05e-07 $l=3.03e-07 $layer=POLY_cond $X=1.102 $Y=1.918
+ $X2=1.102 $Y2=1.615
r129 15 16 45.1538 $w=4.05e-07 $l=2.02e-07 $layer=POLY_cond $X=1.102 $Y=1.918
+ $X2=1.102 $Y2=2.12
r130 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=1.52
+ $X2=2.425 $Y2=1.685
r131 11 13 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=2.425 $Y=1.52
+ $X2=2.425 $Y2=0.775
r132 9 16 202.129 $w=1.8e-07 $l=5.2e-07 $layer=POLY_cond $X=0.99 $Y=2.64
+ $X2=0.99 $Y2=2.12
r133 2 32 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.315 $X2=1.895 $Y2=2.515
r134 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.635
+ $Y=0.565 $X2=1.78 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%DE 3 5 6 10 11 12 13 15 16 18 19 21 23 25
+ 27 28 31 32 33
c92 33 0 7.48038e-20 $X=1.68 $Y=1.65
c93 32 0 1.3237e-19 $X=1.68 $Y=1.485
c94 25 0 7.02076e-20 $X=1.995 $Y=1.135
r95 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.485
+ $X2=1.68 $Y2=1.65
r96 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.485 $X2=1.68 $Y2=1.485
r97 28 32 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.485
r98 21 23 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.8 $Y=2.24 $X2=2.8
+ $Y2=2.635
r99 20 27 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.21 $Y=2.165 $X2=2.12
+ $Y2=2.165
r100 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.71 $Y=2.165
+ $X2=2.8 $Y2=2.24
r101 19 20 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.71 $Y=2.165
+ $X2=2.21 $Y2=2.165
r102 16 27 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=2.24
+ $X2=2.12 $Y2=2.165
r103 16 18 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.12 $Y=2.24
+ $X2=2.12 $Y2=2.635
r104 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.995 $Y=1.06
+ $X2=1.995 $Y2=1.135
r105 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.995 $Y=1.06
+ $X2=1.995 $Y2=0.775
r106 11 27 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.03 $Y=2.165
+ $X2=2.12 $Y2=2.165
r107 11 12 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.03 $Y=2.165
+ $X2=1.815 $Y2=2.165
r108 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.815 $Y2=2.165
r109 10 33 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.74 $Y2=1.65
r110 7 25 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.68 $Y=1.135
+ $X2=1.995 $Y2=1.135
r111 7 31 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.68 $Y=1.21
+ $X2=1.68 $Y2=1.485
r112 5 7 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.135
+ $X2=1.68 $Y2=1.135
r113 5 6 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.515 $Y=1.135
+ $X2=1.08 $Y2=1.135
r114 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.005 $Y=1.06
+ $X2=1.08 $Y2=1.135
r115 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.005 $Y=1.06
+ $X2=1.005 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_548_87# 1 2 9 13 15 17 18 19 22 26 30 35
+ 37 39 40 45 47 49 50 51 57 58 64 65 68
c246 68 0 3.76658e-20 $X=13.675 $Y=2.05
c247 50 0 1.56582e-19 $X=14.975 $Y=1.665
c248 49 0 1.70806e-19 $X=14.665 $Y=1.665
c249 39 0 1.30289e-19 $X=13.675 $Y=2.215
c250 13 0 3.18376e-19 $X=3.19 $Y=2.635
r251 63 65 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.905 $Y=1.68
+ $X2=3.19 $Y2=1.68
r252 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.68 $X2=2.905 $Y2=1.68
r253 60 63 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.815 $Y=1.68
+ $X2=2.905 $Y2=1.68
r254 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=1.665
+ $X2=15.12 $Y2=1.665
r255 54 64 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.64 $Y=1.68
+ $X2=2.905 $Y2=1.68
r256 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r257 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r258 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=15.12 $Y2=1.665
r259 50 51 15.0866 $w=1.4e-07 $l=1.219e-05 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=2.785 $Y2=1.665
r260 48 58 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=14.75 $Y=1.665
+ $X2=15.12 $Y2=1.665
r261 48 49 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.75 $Y=1.665
+ $X2=14.665 $Y2=1.665
r262 44 45 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.532 $Y=1.12
+ $X2=14.532 $Y2=1.29
r263 40 69 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.675 $Y=2.215
+ $X2=13.675 $Y2=2.38
r264 40 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.675 $Y=2.215
+ $X2=13.675 $Y2=2.05
r265 39 42 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=13.675 $Y=2.215
+ $X2=13.675 $Y2=2.385
r266 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.675
+ $Y=2.215 $X2=13.675 $Y2=2.215
r267 37 47 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=14.665 $Y=2.3
+ $X2=14.575 $Y2=2.385
r268 36 49 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=14.665 $Y=1.78
+ $X2=14.665 $Y2=1.665
r269 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=14.665 $Y=1.78
+ $X2=14.665 $Y2=2.3
r270 35 49 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=14.665 $Y=1.55
+ $X2=14.665 $Y2=1.665
r271 35 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=14.665 $Y=1.55
+ $X2=14.665 $Y2=1.29
r272 30 44 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=14.48 $Y=0.58
+ $X2=14.48 $Y2=1.12
r273 27 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.84 $Y=2.385
+ $X2=13.675 $Y2=2.385
r274 26 47 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=14.4 $Y=2.385
+ $X2=14.575 $Y2=2.385
r275 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=14.4 $Y=2.385
+ $X2=13.84 $Y2=2.385
r276 24 68 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.765 $Y=1.015
+ $X2=13.765 $Y2=2.05
r277 22 69 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=13.63 $Y=2.75
+ $X2=13.63 $Y2=2.38
r278 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.69 $Y=0.94
+ $X2=13.765 $Y2=1.015
r279 18 19 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=13.69 $Y=0.94
+ $X2=13.235 $Y2=0.94
r280 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.16 $Y=0.865
+ $X2=13.235 $Y2=0.94
r281 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.16 $Y=0.865
+ $X2=13.16 $Y2=0.58
r282 11 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.845
+ $X2=3.19 $Y2=1.68
r283 11 13 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=3.19 $Y=1.845
+ $X2=3.19 $Y2=2.635
r284 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.515
+ $X2=2.815 $Y2=1.68
r285 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.815 $Y=1.515
+ $X2=2.815 $Y2=0.775
r286 2 47 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=14.43
+ $Y=2.32 $X2=14.565 $Y2=2.465
r287 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.34
+ $Y=0.37 $X2=14.48 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_663_87# 1 2 7 9 10 11 14 18 20 23 24 29
+ 30 32 33 37 38 43 45 49
c109 43 0 1.05969e-19 $X=4.55 $Y=0.805
r110 46 49 5.10825 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=4.21 $Y=2.495
+ $X2=4.415 $Y2=2.495
r111 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.785
+ $Y=1.58 $X2=5.785 $Y2=1.58
r112 35 37 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=5.752 $Y=1.915
+ $X2=5.752 $Y2=1.58
r113 34 45 2.40986 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.295 $Y=2
+ $X2=4.152 $Y2=2
r114 33 35 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.62 $Y=2
+ $X2=5.752 $Y2=1.915
r115 33 34 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=5.62 $Y=2
+ $X2=4.295 $Y2=2
r116 32 46 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.21 $Y=2.255
+ $X2=4.21 $Y2=2.495
r117 31 45 4.02809 $w=2.27e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.21 $Y=2.085
+ $X2=4.152 $Y2=2
r118 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.21 $Y=2.085
+ $X2=4.21 $Y2=2.255
r119 29 30 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.13
+ $Y=1.78 $X2=4.13 $Y2=1.78
r120 27 45 4.02809 $w=2.27e-07 $l=8.5e-08 $layer=LI1_cond $X=4.152 $Y=1.915
+ $X2=4.152 $Y2=2
r121 27 29 5.45894 $w=2.83e-07 $l=1.35e-07 $layer=LI1_cond $X=4.152 $Y=1.915
+ $X2=4.152 $Y2=1.78
r122 26 29 31.1362 $w=2.83e-07 $l=7.7e-07 $layer=LI1_cond $X=4.152 $Y=1.01
+ $X2=4.152 $Y2=1.78
r123 23 24 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.13
+ $Y=0.42 $X2=4.13 $Y2=0.42
r124 21 43 11.3252 $w=4.03e-07 $l=3.98e-07 $layer=LI1_cond $X=4.152 $Y=0.807
+ $X2=4.55 $Y2=0.807
r125 21 26 2.81058 $w=2.85e-07 $l=2.03e-07 $layer=LI1_cond $X=4.152 $Y=0.807
+ $X2=4.152 $Y2=1.01
r126 21 23 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=4.152 $Y=0.605
+ $X2=4.152 $Y2=0.42
r127 19 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.785 $Y=1.92
+ $X2=5.785 $Y2=1.58
r128 19 20 37.308 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.785 $Y=1.92
+ $X2=5.785 $Y2=2.085
r129 17 30 99.6709 $w=3.3e-07 $l=5.7e-07 $layer=POLY_cond $X=4.13 $Y=1.21
+ $X2=4.13 $Y2=1.78
r130 17 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.13 $Y=1.21
+ $X2=4.13 $Y2=1.135
r131 16 24 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=4.13 $Y=1.06
+ $X2=4.13 $Y2=0.42
r132 16 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.13 $Y=1.06
+ $X2=4.13 $Y2=1.135
r133 14 20 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=5.74 $Y=2.595
+ $X2=5.74 $Y2=2.085
r134 10 18 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.135
+ $X2=4.13 $Y2=1.135
r135 10 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.965 $Y=1.135
+ $X2=3.465 $Y2=1.135
r136 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=1.06
+ $X2=3.465 $Y2=1.135
r137 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.39 $Y=1.06 $X2=3.39
+ $Y2=0.775
r138 2 49 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=2.275 $X2=4.415 $Y2=2.495
r139 1 43 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=4.405
+ $Y=0.625 $X2=4.55 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%SCD 3 7 9 12
c39 12 0 8.67074e-20 $X=5.245 $Y=1.58
c40 3 0 3.01793e-19 $X=5.265 $Y=0.835
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.58
+ $X2=5.245 $Y2=1.745
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.58
+ $X2=5.245 $Y2=1.415
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.245
+ $Y=1.58 $X2=5.245 $Y2=1.58
r44 9 13 7.49192 $w=4.53e-07 $l=2.85e-07 $layer=LI1_cond $X=5.182 $Y=1.295
+ $X2=5.182 $Y2=1.58
r45 7 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.32 $Y=2.595
+ $X2=5.32 $Y2=1.745
r46 3 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.265 $Y=0.835
+ $X2=5.265 $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%SCE 1 3 4 5 9 13 14 15 18 20 23 24
c76 24 0 2.82531e-19 $X=4.67 $Y=1.345
c77 18 0 1.9935e-19 $X=5.625 $Y=0.835
c78 1 0 1.43862e-19 $X=3.64 $Y=3.03
r79 23 26 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.672 $Y=1.345
+ $X2=4.672 $Y2=1.51
r80 23 25 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.672 $Y=1.345
+ $X2=4.672 $Y2=1.18
r81 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.67
+ $Y=1.345 $X2=4.67 $Y2=1.345
r82 20 24 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.56 $Y=1.345
+ $X2=4.67 $Y2=1.345
r83 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.625 $Y=0.255
+ $X2=5.625 $Y2=0.835
r84 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.55 $Y=0.18
+ $X2=5.625 $Y2=0.255
r85 14 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.55 $Y=0.18
+ $X2=4.84 $Y2=0.18
r86 13 25 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.765 $Y=0.835
+ $X2=4.765 $Y2=1.18
r87 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.765 $Y=0.255
+ $X2=4.84 $Y2=0.18
r88 10 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.765 $Y=0.255
+ $X2=4.765 $Y2=0.835
r89 9 26 421.75 $w=1.8e-07 $l=1.085e-06 $layer=POLY_cond $X=4.64 $Y=2.595
+ $X2=4.64 $Y2=1.51
r90 7 9 169.089 $w=1.8e-07 $l=4.35e-07 $layer=POLY_cond $X=4.64 $Y=3.03 $X2=4.64
+ $Y2=2.595
r91 4 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.55 $Y=3.105
+ $X2=4.64 $Y2=3.03
r92 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4.55 $Y=3.105 $X2=3.73
+ $Y2=3.105
r93 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.64 $Y=3.03
+ $X2=3.73 $Y2=3.105
r94 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.64 $Y=3.03 $X2=3.64
+ $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%CLK 1 3 6 8 15
c38 15 0 2.59911e-20 $X=6.755 $Y=1.385
c39 8 0 1.22168e-20 $X=6.48 $Y=1.295
r40 14 15 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=6.625 $Y=1.385
+ $X2=6.755 $Y2=1.385
r41 11 14 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=6.56 $Y=1.385
+ $X2=6.625 $Y2=1.385
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.56
+ $Y=1.385 $X2=6.56 $Y2=1.385
r43 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.56 $Y=1.295 $X2=6.56
+ $Y2=1.385
r44 4 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.755 $Y=1.55
+ $X2=6.755 $Y2=1.385
r45 4 6 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=6.755 $Y=1.55
+ $X2=6.755 $Y2=2.38
r46 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.625 $Y=1.22
+ $X2=6.625 $Y2=1.385
r47 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.625 $Y=1.22 $X2=6.625
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_1538_74# 1 2 9 11 13 16 20 24 26 27 28
+ 33 34 38 41 42 43 45 46 47 49 52 53 55 57 58 61 62 63 66 68 69 73
c231 73 0 2.65373e-20 $X=13.285 $Y=1.42
c232 61 0 1.50148e-19 $X=8.84 $Y=2.185
c233 53 0 1.80054e-19 $X=12.205 $Y=1.635
c234 33 0 1.39112e-19 $X=8.73 $Y=1.82
c235 20 0 1.46653e-19 $X=13.21 $Y=2.75
r236 73 86 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.285 $Y=1.42
+ $X2=13.285 $Y2=1.585
r237 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.285
+ $Y=1.42 $X2=13.285 $Y2=1.42
r238 69 72 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=13.285 $Y=1.275
+ $X2=13.285 $Y2=1.42
r239 66 77 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.49 $Y=1.18
+ $X2=9.285 $Y2=1.18
r240 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.49
+ $Y=1.18 $X2=9.49 $Y2=1.18
r241 62 65 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.49 $Y=0.935
+ $X2=9.49 $Y2=1.18
r242 62 63 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.49 $Y=0.935
+ $X2=9.49 $Y2=0.85
r243 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.84
+ $Y=2.185 $X2=8.84 $Y2=2.185
r244 58 60 3.16509 $w=4.24e-07 $l=1.1e-07 $layer=LI1_cond $X=8.73 $Y=2.085
+ $X2=8.84 $Y2=2.085
r245 56 68 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.37 $Y=1.275
+ $X2=12.205 $Y2=1.275
r246 55 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.12 $Y=1.275
+ $X2=13.285 $Y2=1.275
r247 55 56 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=13.12 $Y=1.275
+ $X2=12.37 $Y2=1.275
r248 53 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.205 $Y=1.635
+ $X2=12.205 $Y2=1.47
r249 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.205
+ $Y=1.635 $X2=12.205 $Y2=1.635
r250 50 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.205 $Y=1.36
+ $X2=12.205 $Y2=1.275
r251 50 52 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.205 $Y=1.36
+ $X2=12.205 $Y2=1.635
r252 49 68 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=12.125 $Y=1.19
+ $X2=12.205 $Y2=1.275
r253 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=12.125 $Y=1.02
+ $X2=12.125 $Y2=1.19
r254 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.04 $Y=0.935
+ $X2=12.125 $Y2=1.02
r255 46 47 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=12.04 $Y=0.935
+ $X2=11.465 $Y2=0.935
r256 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.38 $Y=0.85
+ $X2=11.465 $Y2=0.935
r257 44 45 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=11.38 $Y=0.425
+ $X2=11.38 $Y2=0.85
r258 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.295 $Y=0.34
+ $X2=11.38 $Y2=0.425
r259 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.295 $Y=0.34
+ $X2=10.705 $Y2=0.34
r260 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.62 $Y=0.425
+ $X2=10.705 $Y2=0.34
r261 40 41 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.62 $Y=0.425
+ $X2=10.62 $Y2=0.85
r262 39 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.655 $Y=0.935
+ $X2=9.49 $Y2=0.935
r263 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.535 $Y=0.935
+ $X2=10.62 $Y2=0.85
r264 38 39 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=10.535 $Y=0.935
+ $X2=9.655 $Y2=0.935
r265 36 63 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.41 $Y=0.425
+ $X2=9.41 $Y2=0.85
r266 35 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=0.34
+ $X2=8.73 $Y2=0.34
r267 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.325 $Y=0.34
+ $X2=9.41 $Y2=0.425
r268 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.325 $Y=0.34
+ $X2=8.815 $Y2=0.34
r269 33 58 6.13403 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=8.73 $Y=1.82
+ $X2=8.73 $Y2=2.085
r270 32 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.73 $Y=0.425
+ $X2=8.73 $Y2=0.34
r271 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.73 $Y=0.425
+ $X2=8.73 $Y2=1.82
r272 28 58 2.60462 $w=4.24e-07 $l=1.16619e-07 $layer=LI1_cond $X=8.645 $Y=2.01
+ $X2=8.73 $Y2=2.085
r273 28 30 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=8.645 $Y=2.01
+ $X2=8.37 $Y2=2.01
r274 26 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.645 $Y=0.34
+ $X2=8.73 $Y2=0.34
r275 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.645 $Y=0.34
+ $X2=7.995 $Y2=0.34
r276 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.83 $Y=0.425
+ $X2=7.995 $Y2=0.34
r277 22 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.83 $Y=0.425
+ $X2=7.83 $Y2=0.515
r278 20 86 452.847 $w=1.8e-07 $l=1.165e-06 $layer=POLY_cond $X=13.21 $Y=2.75
+ $X2=13.21 $Y2=1.585
r279 16 82 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.295 $Y=0.69
+ $X2=12.295 $Y2=1.47
r280 11 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.285 $Y=1.015
+ $X2=9.285 $Y2=1.18
r281 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.285 $Y=1.015
+ $X2=9.285 $Y2=0.695
r282 7 61 59.7756 $w=2.54e-07 $l=3.88844e-07 $layer=POLY_cond $X=9.155 $Y=2.35
+ $X2=8.84 $Y2=2.185
r283 7 9 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=9.155 $Y=2.35 $X2=9.155
+ $Y2=2.75
r284 2 30 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=8.235
+ $Y=1.84 $X2=8.37 $Y2=2.01
r285 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.69
+ $Y=0.37 $X2=7.83 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_1340_74# 1 2 11 13 15 17 18 22 24 30 34
+ 38 40 41 44 47 48 51 52 57 58 61 62 67 68 72
c193 72 0 1.39112e-19 $X=9.68 $Y=2.02
c194 61 0 1.50148e-19 $X=9.69 $Y=2.185
c195 58 0 1.22168e-20 $X=7.45 $Y=1.695
c196 48 0 1.46653e-19 $X=12.56 $Y=2.475
r197 68 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.745 $Y=1.635
+ $X2=12.745 $Y2=1.8
r198 68 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.745 $Y=1.635
+ $X2=12.745 $Y2=1.47
r199 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.745
+ $Y=1.635 $X2=12.745 $Y2=1.635
r200 64 67 5.12197 $w=2.23e-07 $l=1e-07 $layer=LI1_cond $X=12.645 $Y=1.642
+ $X2=12.745 $Y2=1.642
r201 62 73 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.68 $Y=2.185
+ $X2=9.68 $Y2=2.35
r202 62 72 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.68 $Y=2.185
+ $X2=9.68 $Y2=2.02
r203 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=2.185 $X2=9.69 $Y2=2.185
r204 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.45
+ $Y=1.695 $X2=7.45 $Y2=1.695
r205 55 57 8.3904 $w=6.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.98 $Y=1.865
+ $X2=7.45 $Y2=1.865
r206 50 64 2.38091 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=12.645 $Y=1.755
+ $X2=12.645 $Y2=1.642
r207 50 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.645 $Y=1.755
+ $X2=12.645 $Y2=2.39
r208 49 61 12.3706 $w=2.86e-07 $l=3.69188e-07 $layer=LI1_cond $X=9.885 $Y=2.475
+ $X2=9.705 $Y2=2.185
r209 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.56 $Y=2.475
+ $X2=12.645 $Y2=2.39
r210 48 49 174.519 $w=1.68e-07 $l=2.675e-06 $layer=LI1_cond $X=12.56 $Y=2.475
+ $X2=9.885 $Y2=2.475
r211 47 55 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=6.98 $Y=1.53
+ $X2=6.98 $Y2=1.865
r212 47 52 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.98 $Y=1.53
+ $X2=6.98 $Y2=1.01
r213 42 52 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=6.87 $Y=0.815
+ $X2=6.87 $Y2=1.01
r214 42 44 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=6.87 $Y=0.815
+ $X2=6.87 $Y2=0.515
r215 38 75 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=12.77 $Y=0.58
+ $X2=12.77 $Y2=1.47
r216 34 76 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=12.67 $Y=2.46
+ $X2=12.67 $Y2=1.8
r217 30 73 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=9.605 $Y=2.75
+ $X2=9.605 $Y2=2.35
r218 26 72 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=9.58 $Y=1.765
+ $X2=9.58 $Y2=2.02
r219 25 41 17.0838 $w=1.85e-07 $l=9.08295e-08 $layer=POLY_cond $X=8.68 $Y=1.69
+ $X2=8.605 $Y2=1.655
r220 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.505 $Y=1.69
+ $X2=9.58 $Y2=1.765
r221 24 25 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=9.505 $Y=1.69
+ $X2=8.68 $Y2=1.69
r222 20 41 8.32657 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=8.605 $Y=1.545
+ $X2=8.605 $Y2=1.655
r223 20 22 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=8.605 $Y=1.545
+ $X2=8.605 $Y2=0.695
r224 19 40 17.2177 $w=2.2e-07 $l=9e-08 $layer=POLY_cond $X=8.235 $Y=1.655
+ $X2=8.145 $Y2=1.655
r225 18 41 17.0838 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=8.53 $Y=1.655
+ $X2=8.605 $Y2=1.655
r226 18 19 86.0483 $w=2.2e-07 $l=2.95e-07 $layer=POLY_cond $X=8.53 $Y=1.655
+ $X2=8.235 $Y2=1.655
r227 15 40 8.19472 $w=1.8e-07 $l=1.1e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=1.655
r228 15 17 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=2.4
r229 14 58 8.65449 $w=2.2e-07 $l=2.06961e-07 $layer=POLY_cond $X=7.69 $Y=1.655
+ $X2=7.487 $Y2=1.647
r230 13 40 17.2177 $w=2.2e-07 $l=9e-08 $layer=POLY_cond $X=8.055 $Y=1.655
+ $X2=8.145 $Y2=1.655
r231 13 14 106.467 $w=2.2e-07 $l=3.65e-07 $layer=POLY_cond $X=8.055 $Y=1.655
+ $X2=7.69 $Y2=1.655
r232 9 58 16.755 $w=2.77e-07 $l=1.77088e-07 $layer=POLY_cond $X=7.615 $Y=1.53
+ $X2=7.487 $Y2=1.647
r233 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.615 $Y=1.53
+ $X2=7.615 $Y2=0.74
r234 2 55 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.82 $X2=6.98 $Y2=2
r235 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.7
+ $Y=0.37 $X2=6.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_1979_71# 1 2 9 13 17 19 21 23 24 28 31
+ 34 35 41 45 47 51
c104 34 0 1.80054e-19 $X=11.635 $Y=1.355
r105 43 45 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.915 $Y=2.135
+ $X2=11.04 $Y2=2.135
r106 39 51 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.08 $Y=1.34
+ $X2=10.155 $Y2=1.34
r107 39 48 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=10.08 $Y=1.34
+ $X2=9.97 $Y2=1.34
r108 38 41 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=10.08 $Y=1.34
+ $X2=10.245 $Y2=1.34
r109 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.08
+ $Y=1.34 $X2=10.08 $Y2=1.34
r110 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.635
+ $Y=1.355 $X2=11.635 $Y2=1.355
r111 32 47 2.53577 $w=3.3e-07 $l=3.22102e-07 $layer=LI1_cond $X=11.125 $Y=1.355
+ $X2=10.875 $Y2=1.19
r112 32 34 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=11.125 $Y=1.355
+ $X2=11.635 $Y2=1.355
r113 31 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.04 $Y=2.05
+ $X2=11.04 $Y2=2.135
r114 30 47 3.59786 $w=1.7e-07 $l=4.04166e-07 $layer=LI1_cond $X=11.04 $Y=1.52
+ $X2=10.875 $Y2=1.19
r115 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.04 $Y=1.52
+ $X2=11.04 $Y2=2.05
r116 26 47 3.59786 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=11 $Y=1.19
+ $X2=10.875 $Y2=1.19
r117 26 28 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=11 $Y=1.19 $X2=11
+ $Y2=0.81
r118 24 47 2.53577 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.875 $Y=1.275
+ $X2=10.875 $Y2=1.19
r119 24 41 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.875 $Y=1.275
+ $X2=10.245 $Y2=1.275
r120 21 23 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=11.935 $Y=1.11
+ $X2=11.935 $Y2=0.69
r121 17 21 40.1667 $w=2.7e-07 $l=3.76032e-07 $layer=POLY_cond $X=11.71 $Y=1.39
+ $X2=11.935 $Y2=1.11
r122 17 35 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=11.71 $Y=1.39
+ $X2=11.635 $Y2=1.39
r123 17 19 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=11.71 $Y=1.52
+ $X2=11.71 $Y2=2.46
r124 11 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.155 $Y=1.505
+ $X2=10.155 $Y2=1.34
r125 11 13 483.944 $w=1.8e-07 $l=1.245e-06 $layer=POLY_cond $X=10.155 $Y=1.505
+ $X2=10.155 $Y2=2.75
r126 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.97 $Y=1.175
+ $X2=9.97 $Y2=1.34
r127 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.97 $Y=1.175
+ $X2=9.97 $Y2=0.695
r128 2 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.78
+ $Y=1.99 $X2=10.915 $Y2=2.135
r129 1 28 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=10.82
+ $Y=0.37 $X2=10.96 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_1736_97# 1 2 9 13 17 21 22 27 28 31 32
r88 32 38 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.637 $Y=1.665
+ $X2=10.637 $Y2=1.83
r89 32 37 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.637 $Y=1.665
+ $X2=10.637 $Y2=1.5
r90 31 34 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.62 $Y=1.665
+ $X2=10.62 $Y2=1.745
r91 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.62
+ $Y=1.665 $X2=10.62 $Y2=1.665
r92 27 28 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=9.365 $Y=2.75
+ $X2=9.365 $Y2=2.52
r93 23 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.07 $Y=1.745 $X2=9.27
+ $Y2=1.745
r94 22 25 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=1.745
+ $X2=9.27 $Y2=1.745
r95 21 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.455 $Y=1.745
+ $X2=10.62 $Y2=1.745
r96 21 22 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=10.455 $Y=1.745
+ $X2=9.355 $Y2=1.745
r97 19 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=1.83
+ $X2=9.27 $Y2=1.745
r98 19 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.27 $Y=1.83 $X2=9.27
+ $Y2=2.52
r99 15 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.07 $Y=1.66
+ $X2=9.07 $Y2=1.745
r100 15 17 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=9.07 $Y=1.66 $X2=9.07
+ $Y2=0.76
r101 13 37 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.745 $Y=0.69
+ $X2=10.745 $Y2=1.5
r102 9 38 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=10.69 $Y=2.41
+ $X2=10.69 $Y2=1.83
r103 2 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=9.245
+ $Y=2.54 $X2=9.38 $Y2=2.75
r104 1 17 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=8.68
+ $Y=0.485 $X2=9.07 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_2474_74# 1 2 9 13 15 19 23 27 31 34 36
+ 39 43 45 46 49 51 52 54 55 58 60 61
c166 45 0 3.76658e-20 $X=13.62 $Y=0.935
c167 36 0 1.30289e-19 $X=14.255 $Y=2.13
r168 60 63 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=14.245 $Y=1.625
+ $X2=14.245 $Y2=1.84
r169 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.245
+ $Y=1.625 $X2=14.245 $Y2=1.625
r170 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.79 $Y=1.84
+ $X2=13.705 $Y2=1.84
r171 55 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.08 $Y=1.84
+ $X2=14.245 $Y2=1.84
r172 55 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=14.08 $Y=1.84
+ $X2=13.79 $Y2=1.84
r173 54 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=1.755
+ $X2=13.705 $Y2=1.84
r174 53 54 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=13.705 $Y=1.02
+ $X2=13.705 $Y2=1.755
r175 51 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.62 $Y=1.84
+ $X2=13.705 $Y2=1.84
r176 51 52 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.62 $Y=1.84
+ $X2=13.25 $Y2=1.84
r177 47 52 9.70699 $w=2.57e-07 $l=2.14126e-07 $layer=LI1_cond $X=13.075 $Y=1.927
+ $X2=13.25 $Y2=1.84
r178 47 49 21.4025 $w=3.48e-07 $l=6.5e-07 $layer=LI1_cond $X=13.075 $Y=2.1
+ $X2=13.075 $Y2=2.75
r179 45 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.62 $Y=0.935
+ $X2=13.705 $Y2=1.02
r180 45 46 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=13.62 $Y=0.935
+ $X2=12.72 $Y2=0.935
r181 41 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.555 $Y=0.85
+ $X2=12.72 $Y2=0.935
r182 41 43 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=12.555 $Y=0.85
+ $X2=12.555 $Y2=0.58
r183 39 40 12.1513 $w=2.38e-07 $l=6e-08 $layer=POLY_cond $X=15.755 $Y=1.485
+ $X2=15.815 $Y2=1.485
r184 38 39 82.021 $w=2.38e-07 $l=4.05e-07 $layer=POLY_cond $X=15.35 $Y=1.485
+ $X2=15.755 $Y2=1.485
r185 37 38 5.06302 $w=2.38e-07 $l=2.5e-08 $layer=POLY_cond $X=15.325 $Y=1.485
+ $X2=15.35 $Y2=1.485
r186 35 61 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=14.255 $Y=1.955
+ $X2=14.255 $Y2=1.625
r187 35 36 42.4214 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=14.255 $Y=1.955
+ $X2=14.255 $Y2=2.13
r188 33 61 2.47304 $w=3.5e-07 $l=1.5e-08 $layer=POLY_cond $X=14.255 $Y=1.61
+ $X2=14.255 $Y2=1.625
r189 33 34 20.4101 $w=2.5e-07 $l=2.38485e-07 $layer=POLY_cond $X=14.255 $Y=1.61
+ $X2=14.08 $Y2=1.46
r190 29 40 9.38375 $w=1.8e-07 $l=1.25e-07 $layer=POLY_cond $X=15.815 $Y=1.61
+ $X2=15.815 $Y2=1.485
r191 29 31 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=15.815 $Y=1.61
+ $X2=15.815 $Y2=2.4
r192 25 39 13.5836 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=15.755 $Y=1.36
+ $X2=15.755 $Y2=1.485
r193 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.755 $Y=1.36
+ $X2=15.755 $Y2=0.74
r194 21 38 9.38375 $w=1.8e-07 $l=1.25e-07 $layer=POLY_cond $X=15.35 $Y=1.61
+ $X2=15.35 $Y2=1.485
r195 21 23 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=15.35 $Y=1.61
+ $X2=15.35 $Y2=2.4
r196 17 37 13.5836 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=15.325 $Y=1.36
+ $X2=15.325 $Y2=1.485
r197 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.325 $Y=1.36
+ $X2=15.325 $Y2=0.74
r198 16 34 5.30422 $w=2.5e-07 $l=3.62284e-07 $layer=POLY_cond $X=14.43 $Y=1.485
+ $X2=14.08 $Y2=1.46
r199 15 37 14.6161 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.25 $Y=1.485
+ $X2=15.325 $Y2=1.485
r200 15 16 203.732 $w=2.5e-07 $l=8.2e-07 $layer=POLY_cond $X=15.25 $Y=1.485
+ $X2=14.43 $Y2=1.485
r201 13 36 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=14.34 $Y=2.64
+ $X2=14.34 $Y2=2.13
r202 7 34 20.4101 $w=2.5e-07 $l=2.29619e-07 $layer=POLY_cond $X=14.265 $Y=1.36
+ $X2=14.08 $Y2=1.46
r203 7 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=14.265 $Y=1.36
+ $X2=14.265 $Y2=0.58
r204 2 49 600 $w=1.7e-07 $l=8.95461e-07 $layer=licon1_PDIFF $count=1 $X=12.76
+ $Y=1.96 $X2=12.985 $Y2=2.75
r205 1 43 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=12.37
+ $Y=0.37 $X2=12.555 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_40_464# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 30 33 36 40 42 46 50 52
c121 33 0 1.43862e-19 $X=3.415 $Y=2.46
c122 19 0 1.8559e-19 $X=1.47 $Y=2.375
r123 48 50 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.255 $Y=1.26
+ $X2=3.415 $Y2=1.26
r124 44 46 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.1 $Y=0.84
+ $X2=3.255 $Y2=0.84
r125 37 40 5.98039 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.17 $Y=0.58
+ $X2=0.4 $Y2=0.58
r126 36 52 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.415 $Y=2.29
+ $X2=3.375 $Y2=2.375
r127 35 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.345
+ $X2=3.415 $Y2=1.26
r128 35 36 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.415 $Y=1.345
+ $X2=3.415 $Y2=2.29
r129 33 52 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=2.46
+ $X2=3.375 $Y2=2.375
r130 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.255 $Y=1.175
+ $X2=3.255 $Y2=1.26
r131 29 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=1.005
+ $X2=3.255 $Y2=0.84
r132 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.255 $Y=1.005
+ $X2=3.255 $Y2=1.175
r133 27 52 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.25 $Y=2.375
+ $X2=3.375 $Y2=2.375
r134 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.25 $Y=2.375
+ $X2=2.32 $Y2=2.375
r135 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.235 $Y=2.46
+ $X2=2.32 $Y2=2.375
r136 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.235 $Y=2.46
+ $X2=2.235 $Y2=2.905
r137 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.15 $Y=2.99
+ $X2=2.235 $Y2=2.905
r138 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.15 $Y=2.99
+ $X2=1.64 $Y2=2.99
r139 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=2.905
+ $X2=1.64 $Y2=2.99
r140 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.555 $Y=2.46
+ $X2=1.555 $Y2=2.905
r141 20 42 3.41642 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.51 $Y=2.375
+ $X2=0.297 $Y2=2.375
r142 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.47 $Y=2.375
+ $X2=1.555 $Y2=2.46
r143 19 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.47 $Y=2.375
+ $X2=0.51 $Y2=2.375
r144 15 42 3.17288 $w=2.97e-07 $l=8.5e-08 $layer=LI1_cond $X=0.297 $Y=2.46
+ $X2=0.297 $Y2=2.375
r145 15 17 0.135582 $w=4.23e-07 $l=5e-09 $layer=LI1_cond $X=0.297 $Y=2.46
+ $X2=0.297 $Y2=2.465
r146 14 42 3.17288 $w=2.97e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.297 $Y2=2.375
r147 13 37 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.17 $Y=0.81 $X2=0.17
+ $Y2=0.58
r148 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.29
r149 4 33 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=2.315 $X2=3.415 $Y2=2.46
r150 3 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=2.32 $X2=0.345 $Y2=2.465
r151 2 44 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.565 $X2=3.1 $Y2=0.84
r152 1 40 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.37 $X2=0.4 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 53 57 61 65 69 71 74 75 77 78 79 81 86 91 96 101 106 124 128 134 137 140 143
+ 146 149 152 156
c183 65 0 1.04054e-19 $X=15.125 $Y=2.035
c184 3 0 9.48608e-20 $X=4.73 $Y=2.275
r185 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r186 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r187 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r188 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r189 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 140 141 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r191 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 132 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.08 $Y2=3.33
r194 132 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=15.12 $Y2=3.33
r195 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r196 129 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.29 $Y=3.33
+ $X2=15.125 $Y2=3.33
r197 129 131 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=15.29 $Y=3.33
+ $X2=15.6 $Y2=3.33
r198 128 155 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.875 $Y=3.33
+ $X2=16.097 $Y2=3.33
r199 128 131 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.875 $Y=3.33
+ $X2=15.6 $Y2=3.33
r200 127 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r201 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r202 124 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.96 $Y=3.33
+ $X2=15.125 $Y2=3.33
r203 124 126 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=14.96 $Y=3.33
+ $X2=14.64 $Y2=3.33
r204 123 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r205 122 123 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r206 120 123 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r207 119 122 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r208 119 120 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r209 117 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 117 150 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r211 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r212 114 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.545 $Y=3.33
+ $X2=10.38 $Y2=3.33
r213 114 116 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=10.545 $Y=3.33
+ $X2=11.28 $Y2=3.33
r214 113 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r215 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r216 110 113 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r217 109 112 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r218 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r219 107 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=7.92 $Y2=3.33
r220 107 109 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=8.4 $Y2=3.33
r221 106 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.215 $Y=3.33
+ $X2=10.38 $Y2=3.33
r222 106 112 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.215 $Y=3.33
+ $X2=9.84 $Y2=3.33
r223 105 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 105 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r225 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r226 102 143 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.527 $Y2=3.33
r227 102 104 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r228 101 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.92 $Y2=3.33
r229 101 104 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.44 $Y2=3.33
r230 100 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r231 100 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r232 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r233 97 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.135 $Y2=3.33
r234 97 99 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.26 $Y=3.33 $X2=6
+ $Y2=3.33
r235 96 143 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=6.36 $Y=3.33
+ $X2=6.527 $Y2=3.33
r236 96 99 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6
+ $Y2=3.33
r237 95 141 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r238 95 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r239 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r240 92 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.615 $Y2=3.33
r241 92 94 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=3.12 $Y2=3.33
r242 91 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=5.135 $Y2=3.33
r243 91 94 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=3.12 $Y2=3.33
r244 90 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r245 90 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r246 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r247 87 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.175 $Y2=3.33
r248 87 89 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=2.16
+ $Y2=3.33
r249 86 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.615 $Y2=3.33
r250 86 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.16 $Y2=3.33
r251 84 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r252 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r253 81 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=1.175 $Y2=3.33
r254 81 83 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 79 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=8.4 $Y2=3.33
r256 79 147 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 77 122 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=13.69 $Y=3.33
+ $X2=13.68 $Y2=3.33
r258 77 78 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=13.69 $Y=3.33
+ $X2=13.96 $Y2=3.33
r259 76 126 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=14.23 $Y=3.33
+ $X2=14.64 $Y2=3.33
r260 76 78 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=14.23 $Y=3.33
+ $X2=13.96 $Y2=3.33
r261 74 116 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=11.31 $Y=3.33
+ $X2=11.28 $Y2=3.33
r262 74 75 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.31 $Y=3.33
+ $X2=11.48 $Y2=3.33
r263 73 119 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.76 $Y2=3.33
r264 73 75 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.48 $Y2=3.33
r265 69 155 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=16.04 $Y=3.245
+ $X2=16.097 $Y2=3.33
r266 69 71 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=16.04 $Y=3.245
+ $X2=16.04 $Y2=2.405
r267 65 68 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=15.125 $Y=2.035
+ $X2=15.125 $Y2=2.815
r268 63 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.125 $Y=3.245
+ $X2=15.125 $Y2=3.33
r269 63 68 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.125 $Y=3.245
+ $X2=15.125 $Y2=2.815
r270 59 78 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=13.96 $Y=3.245
+ $X2=13.96 $Y2=3.33
r271 59 61 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=13.96 $Y=3.245
+ $X2=13.96 $Y2=2.815
r272 55 75 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=11.48 $Y=3.245
+ $X2=11.48 $Y2=3.33
r273 55 57 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=11.48 $Y=3.245
+ $X2=11.48 $Y2=2.815
r274 51 149 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.38 $Y=3.245
+ $X2=10.38 $Y2=3.33
r275 51 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.38 $Y=3.245
+ $X2=10.38 $Y2=2.815
r276 47 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r277 47 49 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.805
r278 43 143 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.527 $Y=3.245
+ $X2=6.527 $Y2=3.33
r279 43 45 15.4806 $w=3.33e-07 $l=4.5e-07 $layer=LI1_cond $X=6.527 $Y=3.245
+ $X2=6.527 $Y2=2.795
r280 39 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.135 $Y=3.245
+ $X2=5.135 $Y2=3.33
r281 39 41 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=5.135 $Y=3.245
+ $X2=5.135 $Y2=2.765
r282 35 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=3.33
r283 35 37 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=2.8
r284 31 134 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=3.245
+ $X2=1.175 $Y2=3.33
r285 31 33 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.175 $Y=3.245
+ $X2=1.175 $Y2=2.805
r286 10 71 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=15.905
+ $Y=1.84 $X2=16.04 $Y2=2.405
r287 9 68 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=14.98
+ $Y=1.84 $X2=15.125 $Y2=2.815
r288 9 65 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=14.98
+ $Y=1.84 $X2=15.125 $Y2=2.035
r289 8 61 600 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_PDIFF $count=1 $X=13.72
+ $Y=2.54 $X2=13.96 $Y2=2.815
r290 7 57 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=11.33
+ $Y=1.96 $X2=11.48 $Y2=2.815
r291 6 53 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=10.245
+ $Y=2.54 $X2=10.38 $Y2=2.815
r292 5 49 600 $w=1.7e-07 $l=1.03496e-06 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.92 $Y2=2.805
r293 4 45 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.82 $X2=6.525 $Y2=2.795
r294 3 41 600 $w=1.7e-07 $l=6.47263e-07 $layer=licon1_PDIFF $count=1 $X=4.73
+ $Y=2.275 $X2=5.095 $Y2=2.765
r295 2 37 600 $w=1.7e-07 $l=6.42067e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=2.315 $X2=2.575 $Y2=2.8
r296 1 33 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=2.32 $X2=1.215 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%A_693_113# 1 2 3 4 5 6 21 24 25 26 28 29
+ 30 35 38 39 40 41 45 47 51 54 57 59 62 65 67 68
c169 57 0 1.92249e-19 $X=3.81 $Y=2.295
c170 25 0 9.48608e-20 $X=4.67 $Y=2.99
r171 68 70 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.34 $Y=2.455
+ $X2=8.34 $Y2=2.605
r172 64 65 0.949071 $w=4.23e-07 $l=3.5e-08 $layer=LI1_cond $X=6.012 $Y=2.42
+ $X2=6.012 $Y2=2.455
r173 56 57 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=3.755 $Y=1.005
+ $X2=3.755 $Y2=2.295
r174 54 56 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.675 $Y=0.775
+ $X2=3.675 $Y2=1.005
r175 49 51 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=8.89 $Y=2.69 $X2=8.89
+ $Y2=2.75
r176 48 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=2.605
+ $X2=8.34 $Y2=2.605
r177 47 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.765 $Y=2.605
+ $X2=8.89 $Y2=2.69
r178 47 48 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.765 $Y=2.605
+ $X2=8.425 $Y2=2.605
r179 43 45 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.35 $Y=1.48
+ $X2=8.35 $Y2=0.76
r180 42 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.035 $Y=2.455
+ $X2=7.95 $Y2=2.455
r181 41 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.255 $Y=2.455
+ $X2=8.34 $Y2=2.455
r182 41 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.255 $Y=2.455
+ $X2=8.035 $Y2=2.455
r183 39 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.225 $Y=1.565
+ $X2=8.35 $Y2=1.48
r184 39 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=8.225 $Y=1.565
+ $X2=8.035 $Y2=1.565
r185 38 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.95 $Y=2.37
+ $X2=7.95 $Y2=2.455
r186 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.95 $Y=1.65
+ $X2=8.035 $Y2=1.565
r187 37 38 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.95 $Y=1.65
+ $X2=7.95 $Y2=2.37
r188 36 65 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=6.225 $Y=2.455
+ $X2=6.012 $Y2=2.455
r189 35 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=2.455
+ $X2=7.95 $Y2=2.455
r190 35 36 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=7.865 $Y=2.455
+ $X2=6.225 $Y2=2.455
r191 33 59 10.6395 $w=3.44e-07 $l=3.98748e-07 $layer=LI1_cond $X=6.14 $Y=1.065
+ $X2=5.84 $Y2=0.835
r192 33 62 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=6.14 $Y=1.065
+ $X2=6.14 $Y2=2.255
r193 29 64 2.1693 $w=4.23e-07 $l=8e-08 $layer=LI1_cond $X=6.012 $Y=2.34
+ $X2=6.012 $Y2=2.42
r194 29 62 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=6.012 $Y=2.34
+ $X2=6.012 $Y2=2.255
r195 29 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.8 $Y=2.34 $X2=4.84
+ $Y2=2.34
r196 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.755 $Y=2.425
+ $X2=4.84 $Y2=2.34
r197 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.755 $Y=2.425
+ $X2=4.755 $Y2=2.905
r198 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.67 $Y=2.99
+ $X2=4.755 $Y2=2.905
r199 25 26 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.67 $Y=2.99
+ $X2=3.95 $Y2=2.99
r200 22 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.95 $Y2=2.99
r201 22 24 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.46
r202 21 57 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.81 $Y=2.435
+ $X2=3.81 $Y2=2.295
r203 21 24 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.81 $Y=2.435
+ $X2=3.81 $Y2=2.46
r204 6 51 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=2.54 $X2=8.93 $Y2=2.75
r205 5 64 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.83
+ $Y=2.275 $X2=5.965 $Y2=2.42
r206 4 24 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.73
+ $Y=2.315 $X2=3.865 $Y2=2.46
r207 3 45 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.245
+ $Y=0.485 $X2=8.39 $Y2=0.76
r208 2 59 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.625 $X2=5.84 $Y2=0.835
r209 1 54 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.565 $X2=3.675 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%Q 1 2 9 12 15 17 18 19
r33 23 25 0.0398693 $w=5.98e-07 $l=2e-09 $layer=LI1_cond $X=15.58 $Y=1.85
+ $X2=15.582 $Y2=1.85
r34 18 19 9.56863 $w=5.98e-07 $l=4.8e-07 $layer=LI1_cond $X=15.6 $Y=1.85
+ $X2=16.08 $Y2=1.85
r35 18 25 0.358824 $w=5.98e-07 $l=1.8e-08 $layer=LI1_cond $X=15.6 $Y=1.85
+ $X2=15.582 $Y2=1.85
r36 13 25 6.03242 $w=2.45e-07 $l=3e-07 $layer=LI1_cond $X=15.582 $Y=2.15
+ $X2=15.582 $Y2=1.85
r37 13 15 12.23 $w=2.43e-07 $l=2.6e-07 $layer=LI1_cond $X=15.582 $Y=2.15
+ $X2=15.582 $Y2=2.41
r38 12 25 6.03242 $w=2.45e-07 $l=3e-07 $layer=LI1_cond $X=15.582 $Y=1.55
+ $X2=15.582 $Y2=1.85
r39 12 17 19.7562 $w=2.43e-07 $l=4.2e-07 $layer=LI1_cond $X=15.582 $Y=1.55
+ $X2=15.582 $Y2=1.13
r40 7 17 6.55101 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.54 $Y=0.965
+ $X2=15.54 $Y2=1.13
r41 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=15.54 $Y=0.965
+ $X2=15.54 $Y2=0.515
r42 2 23 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.44
+ $Y=1.84 $X2=15.58 $Y2=1.985
r43 2 15 300 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_PDIFF $count=2 $X=15.44
+ $Y=1.84 $X2=15.58 $Y2=2.41
r44 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.4
+ $Y=0.37 $X2=15.54 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_2%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49
+ 53 57 61 63 65 68 69 70 72 77 82 94 98 103 116 121 127 130 133 136 139 142 147
+ 150 152 156
c186 45 0 1.9935e-19 $X=6.405 $Y=0.515
c187 33 0 1.74672e-19 $X=1.22 $Y=0.58
r188 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r189 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r190 149 150 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=13.98 $Y=0.297
+ $X2=14.145 $Y2=0.297
r191 145 149 4.6905 $w=7.63e-07 $l=3e-07 $layer=LI1_cond $X=13.68 $Y=0.297
+ $X2=13.98 $Y2=0.297
r192 145 147 15.9858 $w=7.63e-07 $l=4.7e-07 $layer=LI1_cond $X=13.68 $Y=0.297
+ $X2=13.21 $Y2=0.297
r193 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r194 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r195 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r196 136 137 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r197 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r198 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r199 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r200 125 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.08 $Y2=0
r201 125 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=15.12 $Y2=0
r202 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r203 122 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.205 $Y=0
+ $X2=15.04 $Y2=0
r204 122 124 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=15.205 $Y=0
+ $X2=15.6 $Y2=0
r205 121 155 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.875 $Y=0
+ $X2=16.097 $Y2=0
r206 121 124 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.875 $Y=0
+ $X2=15.6 $Y2=0
r207 120 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r208 120 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=13.68 $Y2=0
r209 119 150 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=14.64 $Y=0
+ $X2=14.145 $Y2=0
r210 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r211 116 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.875 $Y=0
+ $X2=15.04 $Y2=0
r212 116 119 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=14.875 $Y=0
+ $X2=14.64 $Y2=0
r213 115 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r214 114 147 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=13.2 $Y=0
+ $X2=13.21 $Y2=0
r215 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r216 112 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r217 112 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r218 111 114 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r219 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r220 109 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.885 $Y=0
+ $X2=11.76 $Y2=0
r221 109 111 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.885 $Y=0
+ $X2=12.24 $Y2=0
r222 107 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r223 107 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r224 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r225 104 139 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=10.232 $Y2=0
r226 104 106 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=10.365 $Y=0
+ $X2=11.28 $Y2=0
r227 103 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.76 $Y2=0
r228 103 106 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.28 $Y2=0
r229 102 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r230 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r231 99 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=0
+ $X2=7.36 $Y2=0
r232 99 101 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=7.485 $Y=0
+ $X2=9.84 $Y2=0
r233 98 139 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=10.1 $Y=0
+ $X2=10.232 $Y2=0
r234 98 101 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.1 $Y=0 $X2=9.84
+ $Y2=0
r235 97 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r236 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r237 94 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=0
+ $X2=7.36 $Y2=0
r238 94 96 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=0
+ $X2=6.96 $Y2=0
r239 93 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r240 93 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r241 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r242 90 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=5.05 $Y2=0
r243 90 92 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=6
+ $Y2=0
r244 89 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r245 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r246 86 89 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r247 86 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r248 85 88 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r249 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r250 83 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.21 $Y2=0
r251 83 85 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.64 $Y2=0
r252 82 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=0
+ $X2=5.05 $Y2=0
r253 82 88 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.885 $Y=0
+ $X2=4.56 $Y2=0
r254 81 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r255 81 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r256 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r257 78 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.22 $Y2=0
r258 78 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r259 77 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.21 $Y2=0
r260 77 80 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r261 75 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r262 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r263 72 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=1.22 $Y2=0
r264 72 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r265 70 102 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=9.84 $Y2=0
r266 70 137 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=7.44 $Y2=0
r267 68 92 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6
+ $Y2=0
r268 68 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.235 $Y=0 $X2=6.365
+ $Y2=0
r269 67 96 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.495 $Y=0
+ $X2=6.96 $Y2=0
r270 67 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.495 $Y=0 $X2=6.365
+ $Y2=0
r271 63 155 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=16.04 $Y=0.085
+ $X2=16.097 $Y2=0
r272 63 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=16.04 $Y=0.085
+ $X2=16.04 $Y2=0.515
r273 59 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.04 $Y=0.085
+ $X2=15.04 $Y2=0
r274 59 61 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.04 $Y=0.085
+ $X2=15.04 $Y2=0.515
r275 55 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.76 $Y2=0
r276 55 57 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.76 $Y2=0.515
r277 51 139 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.232 $Y=0.085
+ $X2=10.232 $Y2=0
r278 51 53 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=10.232 $Y=0.085
+ $X2=10.232 $Y2=0.515
r279 47 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r280 47 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.515
r281 43 69 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0
r282 43 45 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0.515
r283 39 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0
r284 39 41 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0.805
r285 35 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r286 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.775
r287 31 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r288 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.58
r289 10 65 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=15.83
+ $Y=0.37 $X2=16.04 $Y2=0.515
r290 9 61 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=14.895
+ $Y=0.37 $X2=15.04 $Y2=0.515
r291 8 149 91 $w=1.7e-07 $l=8.14279e-07 $layer=licon1_NDIFF $count=2 $X=13.235
+ $Y=0.37 $X2=13.98 $Y2=0.515
r292 7 57 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.72 $Y2=0.515
r293 6 53 182 $w=1.7e-07 $l=2.39531e-07 $layer=licon1_NDIFF $count=1 $X=10.045
+ $Y=0.485 $X2=10.27 $Y2=0.515
r294 5 49 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.255
+ $Y=0.37 $X2=7.4 $Y2=0.515
r295 4 45 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.37 $X2=6.405 $Y2=0.515
r296 3 41 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.625 $X2=5.05 $Y2=0.805
r297 2 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.565 $X2=2.21 $Y2=0.775
r298 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.37 $X2=1.22 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__dlclkp_1.pxi.spice
* Created: Fri Aug 28 17:25:54 2020
* 
x_PM_SKY130_FD_SC_MS__DLCLKP_1%A_83_260# N_A_83_260#_M1019_d N_A_83_260#_M1003_d
+ N_A_83_260#_M1006_g N_A_83_260#_M1017_g N_A_83_260#_c_126_n
+ N_A_83_260#_c_127_n N_A_83_260#_c_128_n N_A_83_260#_c_135_p
+ N_A_83_260#_c_198_p N_A_83_260#_c_129_n N_A_83_260#_c_136_p
+ N_A_83_260#_c_194_p N_A_83_260#_c_155_p N_A_83_260#_c_137_p
+ N_A_83_260#_c_156_p N_A_83_260#_c_130_n PM_SKY130_FD_SC_MS__DLCLKP_1%A_83_260#
x_PM_SKY130_FD_SC_MS__DLCLKP_1%GATE N_GATE_M1000_g N_GATE_M1018_g GATE
+ N_GATE_c_222_n PM_SKY130_FD_SC_MS__DLCLKP_1%GATE
x_PM_SKY130_FD_SC_MS__DLCLKP_1%A_315_54# N_A_315_54#_M1002_s N_A_315_54#_M1008_s
+ N_A_315_54#_c_264_n N_A_315_54#_M1019_g N_A_315_54#_M1007_g
+ N_A_315_54#_M1014_g N_A_315_54#_M1004_g N_A_315_54#_c_266_n
+ N_A_315_54#_c_267_n N_A_315_54#_c_274_n N_A_315_54#_c_292_n
+ N_A_315_54#_c_275_n N_A_315_54#_c_276_n N_A_315_54#_c_277_n
+ N_A_315_54#_c_268_n N_A_315_54#_c_279_n N_A_315_54#_c_280_n
+ N_A_315_54#_c_269_n N_A_315_54#_c_270_n N_A_315_54#_c_351_p
+ PM_SKY130_FD_SC_MS__DLCLKP_1%A_315_54#
x_PM_SKY130_FD_SC_MS__DLCLKP_1%A_309_338# N_A_309_338#_M1004_d
+ N_A_309_338#_M1014_d N_A_309_338#_c_392_n N_A_309_338#_M1003_g
+ N_A_309_338#_c_393_n N_A_309_338#_c_394_n N_A_309_338#_M1001_g
+ N_A_309_338#_c_385_n N_A_309_338#_c_386_n N_A_309_338#_c_387_n
+ N_A_309_338#_c_388_n N_A_309_338#_c_389_n N_A_309_338#_c_390_n
+ N_A_309_338#_c_398_n N_A_309_338#_c_391_n
+ PM_SKY130_FD_SC_MS__DLCLKP_1%A_309_338#
x_PM_SKY130_FD_SC_MS__DLCLKP_1%CLK N_CLK_c_470_n N_CLK_M1008_g N_CLK_c_466_n
+ N_CLK_M1002_g N_CLK_M1012_g N_CLK_c_471_n N_CLK_M1015_g CLK CLK N_CLK_c_469_n
+ PM_SKY130_FD_SC_MS__DLCLKP_1%CLK
x_PM_SKY130_FD_SC_MS__DLCLKP_1%A_27_74# N_A_27_74#_M1017_s N_A_27_74#_M1006_s
+ N_A_27_74#_M1016_g N_A_27_74#_M1010_g N_A_27_74#_c_511_n N_A_27_74#_M1009_g
+ N_A_27_74#_M1011_g N_A_27_74#_c_514_n N_A_27_74#_c_515_n N_A_27_74#_c_527_n
+ N_A_27_74#_c_516_n N_A_27_74#_c_517_n N_A_27_74#_c_528_n N_A_27_74#_c_535_n
+ N_A_27_74#_c_539_n N_A_27_74#_c_518_n N_A_27_74#_c_519_n N_A_27_74#_c_529_n
+ N_A_27_74#_c_520_n N_A_27_74#_c_521_n N_A_27_74#_c_522_n N_A_27_74#_c_523_n
+ PM_SKY130_FD_SC_MS__DLCLKP_1%A_27_74#
x_PM_SKY130_FD_SC_MS__DLCLKP_1%A_990_393# N_A_990_393#_M1009_d
+ N_A_990_393#_M1015_d N_A_990_393#_M1005_g N_A_990_393#_M1013_g
+ N_A_990_393#_c_646_n N_A_990_393#_c_647_n N_A_990_393#_c_648_n
+ N_A_990_393#_c_649_n N_A_990_393#_c_650_n N_A_990_393#_c_654_n
+ N_A_990_393#_c_659_n N_A_990_393#_c_651_n
+ PM_SKY130_FD_SC_MS__DLCLKP_1%A_990_393#
x_PM_SKY130_FD_SC_MS__DLCLKP_1%VPWR N_VPWR_M1006_d N_VPWR_M1010_d N_VPWR_M1008_d
+ N_VPWR_M1011_d N_VPWR_c_708_n N_VPWR_c_709_n N_VPWR_c_710_n N_VPWR_c_711_n
+ N_VPWR_c_712_n N_VPWR_c_713_n VPWR N_VPWR_c_714_n N_VPWR_c_715_n
+ N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_707_n N_VPWR_c_719_n N_VPWR_c_720_n
+ N_VPWR_c_721_n PM_SKY130_FD_SC_MS__DLCLKP_1%VPWR
x_PM_SKY130_FD_SC_MS__DLCLKP_1%GCLK N_GCLK_M1013_d N_GCLK_M1005_d N_GCLK_c_794_n
+ GCLK GCLK GCLK GCLK N_GCLK_c_797_n PM_SKY130_FD_SC_MS__DLCLKP_1%GCLK
x_PM_SKY130_FD_SC_MS__DLCLKP_1%VGND N_VGND_M1017_d N_VGND_M1016_d N_VGND_M1002_d
+ N_VGND_M1013_s N_VGND_c_813_n N_VGND_c_828_n N_VGND_c_814_n N_VGND_c_815_n
+ N_VGND_c_816_n N_VGND_c_817_n N_VGND_c_818_n VGND N_VGND_c_819_n
+ N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n N_VGND_c_824_n
+ N_VGND_c_825_n N_VGND_c_826_n PM_SKY130_FD_SC_MS__DLCLKP_1%VGND
cc_1 VNB N_A_83_260#_M1006_g 0.00187581f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_260#_M1017_g 0.030146f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_A_83_260#_c_126_n 0.00759181f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.63
cc_4 VNB N_A_83_260#_c_127_n 4.07393e-19 $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.97
cc_5 VNB N_A_83_260#_c_128_n 0.0146521f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.215
cc_6 VNB N_A_83_260#_c_129_n 0.00159251f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.13
cc_7 VNB N_A_83_260#_c_130_n 0.0356685f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_8 VNB N_GATE_M1018_g 0.0345308f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_9 VNB GATE 0.00166024f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_10 VNB N_GATE_c_222_n 0.0205978f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_A_315_54#_c_264_n 0.0180708f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_12 VNB N_A_315_54#_M1004_g 0.0207868f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.055
cc_13 VNB N_A_315_54#_c_266_n 0.00535921f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.55
cc_14 VNB N_A_315_54#_c_267_n 0.0395251f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.815
cc_15 VNB N_A_315_54#_c_268_n 0.0132392f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.3
cc_16 VNB N_A_315_54#_c_269_n 0.00584675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_315_54#_c_270_n 0.0254205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_309_338#_M1001_g 0.0339887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_309_338#_c_385_n 0.00319078f $X=-0.19 $Y=-0.245 $X2=0.785
+ $Y2=1.215
cc_20 VNB N_A_309_338#_c_386_n 0.0165635f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=2.055
cc_21 VNB N_A_309_338#_c_387_n 0.0152503f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=0.98
cc_22 VNB N_A_309_338#_c_388_n 0.00748342f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.13
cc_23 VNB N_A_309_338#_c_389_n 0.0105451f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.815
cc_24 VNB N_A_309_338#_c_390_n 0.00878008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_309_338#_c_391_n 0.00173862f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_26 VNB N_CLK_c_466_n 0.0187791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_CLK_M1012_g 0.0209903f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB CLK 0.0101706f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.63
cc_29 VNB N_CLK_c_469_n 0.0418771f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.14
cc_30 VNB N_A_27_74#_M1016_g 0.0108504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_511_n 0.184715f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.215
cc_32 VNB N_A_27_74#_M1009_g 0.0294989f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.13
cc_33 VNB N_A_27_74#_M1011_g 0.0092132f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.815
cc_34 VNB N_A_27_74#_c_514_n 0.015735f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.715
cc_35 VNB N_A_27_74#_c_515_n 0.0271016f $X=-0.19 $Y=-0.245 $X2=1.99 $Y2=2.715
cc_36 VNB N_A_27_74#_c_516_n 0.0136991f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_37 VNB N_A_27_74#_c_517_n 0.0199695f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_38 VNB N_A_27_74#_c_518_n 0.0022869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_519_n 0.019497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_520_n 0.0245895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_521_n 0.00496022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_522_n 0.025466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_523_n 0.0493903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_990_393#_M1005_g 0.00225585f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_45 VNB N_A_990_393#_M1013_g 0.0293558f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_46 VNB N_A_990_393#_c_646_n 0.038908f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.63
cc_47 VNB N_A_990_393#_c_647_n 0.0221319f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.97
cc_48 VNB N_A_990_393#_c_648_n 0.00849579f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=0.98
cc_49 VNB N_A_990_393#_c_649_n 3.54303e-19 $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.55
cc_50 VNB N_A_990_393#_c_650_n 0.00663381f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.815
cc_51 VNB N_A_990_393#_c_651_n 0.00656085f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_52 VNB N_VPWR_c_707_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_GCLK_c_794_n 0.0505628f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_54 VNB GCLK 0.00521116f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_55 VNB N_VGND_c_813_n 0.00805223f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.63
cc_56 VNB N_VGND_c_814_n 0.0115327f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.13
cc_57 VNB N_VGND_c_815_n 0.0153007f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=0.815
cc_58 VNB N_VGND_c_816_n 0.0196172f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.715
cc_59 VNB N_VGND_c_817_n 0.0517199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_818_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.215
cc_61 VNB N_VGND_c_819_n 0.0193135f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.465
cc_62 VNB N_VGND_c_820_n 0.0310734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_821_n 0.0332986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_822_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_823_n 0.364249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_824_n 0.00478372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_825_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_826_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VPB N_A_83_260#_M1006_g 0.0308699f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_70 VPB N_A_83_260#_c_127_n 0.00292534f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.97
cc_71 VPB N_GATE_M1000_g 0.0244225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB GATE 0.00137271f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_73 VPB N_GATE_c_222_n 0.0151473f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_74 VPB N_A_315_54#_M1007_g 0.0246333f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_75 VPB N_A_315_54#_M1014_g 0.0266196f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.97
cc_76 VPB N_A_315_54#_c_266_n 0.0092089f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.55
cc_77 VPB N_A_315_54#_c_274_n 0.0231456f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=0.815
cc_78 VPB N_A_315_54#_c_275_n 0.0308098f $X=-0.19 $Y=1.66 $X2=1.99 $Y2=2.715
cc_79 VPB N_A_315_54#_c_276_n 0.00294598f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.215
cc_80 VPB N_A_315_54#_c_277_n 0.0196829f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_81 VPB N_A_315_54#_c_268_n 0.00322662f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.3
cc_82 VPB N_A_315_54#_c_279_n 0.00226897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_315_54#_c_280_n 0.00334762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_315_54#_c_269_n 0.00100914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_315_54#_c_270_n 0.00749977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_309_338#_c_392_n 0.0213414f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_87 VPB N_A_309_338#_c_393_n 0.0321781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_309_338#_c_394_n 0.00944475f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_89 VPB N_A_309_338#_c_385_n 0.00243131f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.215
cc_90 VPB N_A_309_338#_c_386_n 0.0146979f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=2.055
cc_91 VPB N_A_309_338#_c_390_n 0.00512842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_309_338#_c_398_n 0.0029141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_CLK_c_470_n 0.0213481f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=0.4
cc_94 VPB N_CLK_c_471_n 0.0175878f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_95 VPB CLK 0.00294547f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.63
cc_96 VPB N_CLK_c_469_n 0.0156772f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.14
cc_97 VPB N_A_27_74#_M1010_g 0.0306188f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_98 VPB N_A_27_74#_M1011_g 0.0325626f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=0.815
cc_99 VPB N_A_27_74#_c_515_n 0.0214684f $X=-0.19 $Y=1.66 $X2=1.99 $Y2=2.715
cc_100 VPB N_A_27_74#_c_527_n 0.0104331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_74#_c_528_n 0.0411673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_74#_c_529_n 0.0130047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_74#_c_520_n 0.00743101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_990_393#_M1005_g 0.0311589f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_105 VPB N_A_990_393#_c_649_n 0.00362665f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.55
cc_106 VPB N_A_990_393#_c_654_n 0.00309112f $X=-0.19 $Y=1.66 $X2=1.99 $Y2=2.715
cc_107 VPB N_VPWR_c_708_n 0.00992799f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.63
cc_108 VPB N_VPWR_c_709_n 0.0114049f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=2.055
cc_109 VPB N_VPWR_c_710_n 0.0228463f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.14
cc_110 VPB N_VPWR_c_711_n 0.0160668f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=0.815
cc_111 VPB N_VPWR_c_712_n 0.0281191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_713_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.215
cc_113 VPB N_VPWR_c_714_n 0.0189953f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.465
cc_114 VPB N_VPWR_c_715_n 0.0541479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_716_n 0.03837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_717_n 0.0208322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_707_n 0.116293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_719_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_720_n 0.00613689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_721_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB GCLK 0.00406323f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_122 VPB N_GCLK_c_797_n 0.0545086f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.13
cc_123 N_A_83_260#_M1006_g N_GATE_M1000_g 0.0152222f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_83_260#_c_127_n N_GATE_M1000_g 0.00319185f $X=0.7 $Y=1.97 $X2=0 $Y2=0
cc_125 N_A_83_260#_c_135_p N_GATE_M1000_g 0.0179185f $X=1.385 $Y=2.055 $X2=0
+ $Y2=0
cc_126 N_A_83_260#_c_136_p N_GATE_M1000_g 0.00616963f $X=1.47 $Y=2.55 $X2=0
+ $Y2=0
cc_127 N_A_83_260#_c_137_p N_GATE_M1000_g 0.0039889f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_128 N_A_83_260#_M1017_g N_GATE_M1018_g 0.0146085f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_83_260#_c_126_n N_GATE_M1018_g 0.00326474f $X=0.7 $Y=1.63 $X2=0 $Y2=0
cc_130 N_A_83_260#_c_128_n N_GATE_M1018_g 0.0146591f $X=1.385 $Y=1.215 $X2=0
+ $Y2=0
cc_131 N_A_83_260#_c_129_n N_GATE_M1018_g 0.00229553f $X=1.47 $Y=1.13 $X2=0
+ $Y2=0
cc_132 N_A_83_260#_c_130_n N_GATE_M1018_g 0.00413511f $X=0.6 $Y=1.465 $X2=0
+ $Y2=0
cc_133 N_A_83_260#_c_126_n GATE 0.0105342f $X=0.7 $Y=1.63 $X2=0 $Y2=0
cc_134 N_A_83_260#_c_127_n GATE 0.0105003f $X=0.7 $Y=1.97 $X2=0 $Y2=0
cc_135 N_A_83_260#_c_128_n GATE 0.0242156f $X=1.385 $Y=1.215 $X2=0 $Y2=0
cc_136 N_A_83_260#_c_135_p GATE 0.0207679f $X=1.385 $Y=2.055 $X2=0 $Y2=0
cc_137 N_A_83_260#_M1006_g N_GATE_c_222_n 0.0037308f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_83_260#_c_126_n N_GATE_c_222_n 9.81638e-19 $X=0.7 $Y=1.63 $X2=0 $Y2=0
cc_139 N_A_83_260#_c_127_n N_GATE_c_222_n 0.00128824f $X=0.7 $Y=1.97 $X2=0 $Y2=0
cc_140 N_A_83_260#_c_128_n N_GATE_c_222_n 0.00125621f $X=1.385 $Y=1.215 $X2=0
+ $Y2=0
cc_141 N_A_83_260#_c_135_p N_GATE_c_222_n 7.14516e-19 $X=1.385 $Y=2.055 $X2=0
+ $Y2=0
cc_142 N_A_83_260#_c_130_n N_GATE_c_222_n 0.00850882f $X=0.6 $Y=1.465 $X2=0
+ $Y2=0
cc_143 N_A_83_260#_c_128_n N_A_315_54#_c_264_n 0.00202048f $X=1.385 $Y=1.215
+ $X2=0 $Y2=0
cc_144 N_A_83_260#_c_129_n N_A_315_54#_c_264_n 0.00239048f $X=1.47 $Y=1.13 $X2=0
+ $Y2=0
cc_145 N_A_83_260#_c_155_p N_A_315_54#_c_264_n 0.0220414f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_146 N_A_83_260#_c_156_p N_A_315_54#_M1007_g 0.0132521f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_147 N_A_83_260#_M1003_d N_A_315_54#_c_266_n 2.77692e-19 $X=1.725 $Y=1.96
+ $X2=0 $Y2=0
cc_148 N_A_83_260#_c_128_n N_A_315_54#_c_266_n 0.0124767f $X=1.385 $Y=1.215
+ $X2=0 $Y2=0
cc_149 N_A_83_260#_c_155_p N_A_315_54#_c_266_n 0.0198287f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_150 N_A_83_260#_c_155_p N_A_315_54#_c_267_n 0.00184334f $X=1.98 $Y=0.815
+ $X2=0 $Y2=0
cc_151 N_A_83_260#_c_156_p N_A_315_54#_c_274_n 0.0206825f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_152 N_A_83_260#_M1003_d N_A_315_54#_c_292_n 0.00523972f $X=1.725 $Y=1.96
+ $X2=0 $Y2=0
cc_153 N_A_83_260#_c_135_p N_A_315_54#_c_292_n 0.00761858f $X=1.385 $Y=2.055
+ $X2=0 $Y2=0
cc_154 N_A_83_260#_c_136_p N_A_315_54#_c_292_n 0.018248f $X=1.47 $Y=2.55 $X2=0
+ $Y2=0
cc_155 N_A_83_260#_c_156_p N_A_315_54#_c_292_n 0.0181287f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_156 N_A_83_260#_c_156_p N_A_315_54#_c_275_n 0.0025882f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_157 N_A_83_260#_c_135_p N_A_309_338#_c_392_n 0.00413034f $X=1.385 $Y=2.055
+ $X2=0 $Y2=0
cc_158 N_A_83_260#_c_136_p N_A_309_338#_c_392_n 0.0127294f $X=1.47 $Y=2.55 $X2=0
+ $Y2=0
cc_159 N_A_83_260#_c_137_p N_A_309_338#_c_392_n 0.00266167f $X=1.555 $Y=2.715
+ $X2=0 $Y2=0
cc_160 N_A_83_260#_c_156_p N_A_309_338#_c_392_n 0.0217063f $X=1.99 $Y=2.715
+ $X2=0 $Y2=0
cc_161 N_A_83_260#_c_128_n N_A_309_338#_c_394_n 2.57525e-19 $X=1.385 $Y=1.215
+ $X2=0 $Y2=0
cc_162 N_A_83_260#_c_155_p N_A_309_338#_M1001_g 0.0121375f $X=1.98 $Y=0.815
+ $X2=0 $Y2=0
cc_163 N_A_83_260#_c_155_p N_A_309_338#_c_388_n 0.00324967f $X=1.98 $Y=0.815
+ $X2=0 $Y2=0
cc_164 N_A_83_260#_c_155_p N_A_27_74#_M1016_g 0.00109152f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_165 N_A_83_260#_c_156_p N_A_27_74#_M1010_g 0.00127449f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_166 N_A_83_260#_M1017_g N_A_27_74#_c_517_n 0.00835019f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_83_260#_M1006_g N_A_27_74#_c_528_n 0.0150068f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_168 N_A_83_260#_M1017_g N_A_27_74#_c_535_n 0.0110265f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_83_260#_c_126_n N_A_27_74#_c_535_n 0.0198027f $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_170 N_A_83_260#_c_128_n N_A_27_74#_c_535_n 0.030488f $X=1.385 $Y=1.215 $X2=0
+ $Y2=0
cc_171 N_A_83_260#_c_130_n N_A_27_74#_c_535_n 6.82831e-19 $X=0.6 $Y=1.465 $X2=0
+ $Y2=0
cc_172 N_A_83_260#_M1017_g N_A_27_74#_c_539_n 0.00154004f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_173 N_A_83_260#_M1017_g N_A_27_74#_c_519_n 0.0096554f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_83_260#_c_126_n N_A_27_74#_c_519_n 7.22171e-19 $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_175 N_A_83_260#_c_130_n N_A_27_74#_c_519_n 2.41927e-19 $X=0.6 $Y=1.465 $X2=0
+ $Y2=0
cc_176 N_A_83_260#_M1006_g N_A_27_74#_c_529_n 0.00355858f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_177 N_A_83_260#_c_126_n N_A_27_74#_c_529_n 6.59918e-19 $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_178 N_A_83_260#_c_127_n N_A_27_74#_c_529_n 0.00639411f $X=0.7 $Y=1.97 $X2=0
+ $Y2=0
cc_179 N_A_83_260#_M1017_g N_A_27_74#_c_520_n 0.00256037f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_A_83_260#_c_126_n N_A_27_74#_c_520_n 0.0311509f $X=0.7 $Y=1.63 $X2=0
+ $Y2=0
cc_181 N_A_83_260#_c_127_n N_A_27_74#_c_520_n 0.00635205f $X=0.7 $Y=1.97 $X2=0
+ $Y2=0
cc_182 N_A_83_260#_c_130_n N_A_27_74#_c_520_n 0.0107748f $X=0.6 $Y=1.465 $X2=0
+ $Y2=0
cc_183 N_A_83_260#_M1019_d N_A_27_74#_c_522_n 0.00241797f $X=1.725 $Y=0.4 $X2=0
+ $Y2=0
cc_184 N_A_83_260#_c_194_p N_A_27_74#_c_522_n 0.00750924f $X=1.555 $Y=0.815
+ $X2=0 $Y2=0
cc_185 N_A_83_260#_c_155_p N_A_27_74#_c_522_n 0.0336011f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_186 N_A_83_260#_c_127_n N_VPWR_M1006_d 0.002662f $X=0.7 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_83_260#_c_135_p N_VPWR_M1006_d 0.0127562f $X=1.385 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_83_260#_c_198_p N_VPWR_M1006_d 0.00271221f $X=0.785 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_189 N_A_83_260#_M1006_g N_VPWR_c_708_n 0.00369882f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_190 N_A_83_260#_c_135_p N_VPWR_c_708_n 0.0128995f $X=1.385 $Y=2.055 $X2=0
+ $Y2=0
cc_191 N_A_83_260#_c_198_p N_VPWR_c_708_n 0.0119464f $X=0.785 $Y=2.055 $X2=0
+ $Y2=0
cc_192 N_A_83_260#_c_136_p N_VPWR_c_708_n 0.00905618f $X=1.47 $Y=2.55 $X2=0
+ $Y2=0
cc_193 N_A_83_260#_c_137_p N_VPWR_c_708_n 0.0138666f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_194 N_A_83_260#_c_130_n N_VPWR_c_708_n 3.92061e-19 $X=0.6 $Y=1.465 $X2=0
+ $Y2=0
cc_195 N_A_83_260#_c_156_p N_VPWR_c_709_n 0.00451947f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_196 N_A_83_260#_M1006_g N_VPWR_c_714_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_83_260#_c_137_p N_VPWR_c_715_n 0.00438733f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_198 N_A_83_260#_c_156_p N_VPWR_c_715_n 0.019514f $X=1.99 $Y=2.715 $X2=0 $Y2=0
cc_199 N_A_83_260#_M1006_g N_VPWR_c_707_n 0.00987422f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_200 N_A_83_260#_c_137_p N_VPWR_c_707_n 0.00583745f $X=1.555 $Y=2.715 $X2=0
+ $Y2=0
cc_201 N_A_83_260#_c_156_p N_VPWR_c_707_n 0.0235795f $X=1.99 $Y=2.715 $X2=0
+ $Y2=0
cc_202 N_A_83_260#_c_135_p A_261_392# 0.00334039f $X=1.385 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_83_260#_c_136_p A_261_392# 0.00476493f $X=1.47 $Y=2.55 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_83_260#_c_137_p A_261_392# 0.00563595f $X=1.555 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_83_260#_M1017_g N_VGND_c_813_n 0.00578197f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_83_260#_c_155_p N_VGND_c_828_n 0.00866412f $X=1.98 $Y=0.815 $X2=0
+ $Y2=0
cc_207 N_A_83_260#_M1017_g N_VGND_c_819_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A_83_260#_M1017_g N_VGND_c_823_n 0.00443309f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_83_260#_c_194_p A_267_80# 0.00151363f $X=1.555 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_210 N_GATE_M1018_g N_A_315_54#_c_264_n 0.0312233f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_211 N_GATE_M1018_g N_A_315_54#_c_266_n 9.40021e-19 $X=1.26 $Y=0.72 $X2=0
+ $Y2=0
cc_212 GATE N_A_315_54#_c_266_n 0.0133585f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_213 N_GATE_c_222_n N_A_315_54#_c_266_n 0.00437665f $X=1.17 $Y=1.635 $X2=0
+ $Y2=0
cc_214 N_GATE_c_222_n N_A_315_54#_c_267_n 0.0312233f $X=1.17 $Y=1.635 $X2=0
+ $Y2=0
cc_215 N_GATE_M1000_g N_A_309_338#_c_394_n 0.0677517f $X=1.215 $Y=2.46 $X2=0
+ $Y2=0
cc_216 GATE N_A_309_338#_c_394_n 4.953e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_217 N_GATE_c_222_n N_A_309_338#_c_394_n 0.00734855f $X=1.17 $Y=1.635 $X2=0
+ $Y2=0
cc_218 N_GATE_M1000_g N_A_27_74#_c_528_n 8.20057e-19 $X=1.215 $Y=2.46 $X2=0
+ $Y2=0
cc_219 N_GATE_M1018_g N_A_27_74#_c_535_n 0.00554112f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_220 N_GATE_M1018_g N_A_27_74#_c_539_n 0.00991337f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_221 N_GATE_M1018_g N_A_27_74#_c_518_n 0.00285373f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_222 N_GATE_M1018_g N_A_27_74#_c_522_n 0.010234f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_223 N_GATE_M1000_g N_VPWR_c_708_n 0.0120729f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_224 N_GATE_M1000_g N_VPWR_c_715_n 0.00553757f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_225 N_GATE_M1000_g N_VPWR_c_707_n 0.0109166f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_226 N_GATE_M1018_g N_VGND_c_813_n 0.0010533f $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_227 N_GATE_M1018_g N_VGND_c_817_n 9.48944e-19 $X=1.26 $Y=0.72 $X2=0 $Y2=0
cc_228 N_A_315_54#_c_277_n N_A_309_338#_M1014_d 0.00751807f $X=3.945 $Y=2.475
+ $X2=0 $Y2=0
cc_229 N_A_315_54#_M1007_g N_A_309_338#_c_392_n 0.0167739f $X=2.345 $Y=2.75
+ $X2=0 $Y2=0
cc_230 N_A_315_54#_c_266_n N_A_309_338#_c_392_n 0.00720012f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_231 N_A_315_54#_c_292_n N_A_309_338#_c_392_n 0.0036824f $X=1.995 $Y=2.215
+ $X2=0 $Y2=0
cc_232 N_A_315_54#_c_275_n N_A_309_338#_c_392_n 0.00884923f $X=2.3 $Y=2.215
+ $X2=0 $Y2=0
cc_233 N_A_315_54#_c_266_n N_A_309_338#_c_393_n 0.0168228f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_234 N_A_315_54#_c_274_n N_A_309_338#_c_393_n 0.00542654f $X=3.03 $Y=2.215
+ $X2=0 $Y2=0
cc_235 N_A_315_54#_c_275_n N_A_309_338#_c_393_n 0.0215521f $X=2.3 $Y=2.215 $X2=0
+ $Y2=0
cc_236 N_A_315_54#_c_267_n N_A_309_338#_c_394_n 0.0299681f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_237 N_A_315_54#_c_264_n N_A_309_338#_M1001_g 0.0150689f $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_238 N_A_315_54#_c_266_n N_A_309_338#_M1001_g 6.52036e-19 $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_239 N_A_315_54#_c_267_n N_A_309_338#_M1001_g 0.0177805f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_240 N_A_315_54#_c_266_n N_A_309_338#_c_385_n 0.0334095f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_241 N_A_315_54#_c_267_n N_A_309_338#_c_385_n 9.37391e-19 $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_242 N_A_315_54#_c_274_n N_A_309_338#_c_385_n 0.0223796f $X=3.03 $Y=2.215
+ $X2=0 $Y2=0
cc_243 N_A_315_54#_c_275_n N_A_309_338#_c_385_n 0.00100046f $X=2.3 $Y=2.215
+ $X2=0 $Y2=0
cc_244 N_A_315_54#_c_276_n N_A_309_338#_c_385_n 3.35121e-19 $X=3.115 $Y=2.05
+ $X2=0 $Y2=0
cc_245 N_A_315_54#_c_269_n N_A_309_338#_c_385_n 0.0118744f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_246 N_A_315_54#_c_266_n N_A_309_338#_c_386_n 0.00398033f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_247 N_A_315_54#_c_274_n N_A_309_338#_c_386_n 8.18206e-19 $X=3.03 $Y=2.215
+ $X2=0 $Y2=0
cc_248 N_A_315_54#_M1004_g N_A_309_338#_c_387_n 0.0122329f $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_249 N_A_315_54#_c_269_n N_A_309_338#_c_387_n 0.0268373f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_250 N_A_315_54#_c_270_n N_A_309_338#_c_387_n 0.00350773f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_251 N_A_315_54#_c_266_n N_A_309_338#_c_388_n 0.0120735f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_252 N_A_315_54#_c_267_n N_A_309_338#_c_388_n 0.00116112f $X=1.83 $Y=1.315
+ $X2=0 $Y2=0
cc_253 N_A_315_54#_M1004_g N_A_309_338#_c_389_n 5.39498e-19 $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_254 N_A_315_54#_c_268_n N_A_309_338#_c_389_n 0.00850585f $X=4.115 $Y=1.22
+ $X2=0 $Y2=0
cc_255 N_A_315_54#_M1014_g N_A_309_338#_c_390_n 0.00367497f $X=3.31 $Y=2.41
+ $X2=0 $Y2=0
cc_256 N_A_315_54#_M1004_g N_A_309_338#_c_390_n 0.00513868f $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_257 N_A_315_54#_c_276_n N_A_309_338#_c_390_n 0.00771021f $X=3.115 $Y=2.05
+ $X2=0 $Y2=0
cc_258 N_A_315_54#_c_268_n N_A_309_338#_c_390_n 0.0560683f $X=4.115 $Y=1.22
+ $X2=0 $Y2=0
cc_259 N_A_315_54#_c_269_n N_A_309_338#_c_390_n 0.0251647f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_260 N_A_315_54#_c_270_n N_A_309_338#_c_390_n 0.00231223f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_261 N_A_315_54#_M1014_g N_A_309_338#_c_398_n 0.0027501f $X=3.31 $Y=2.41 $X2=0
+ $Y2=0
cc_262 N_A_315_54#_c_277_n N_A_309_338#_c_398_n 0.0253127f $X=3.945 $Y=2.475
+ $X2=0 $Y2=0
cc_263 N_A_315_54#_c_279_n N_A_309_338#_c_398_n 0.014183f $X=4.102 $Y=2.102
+ $X2=0 $Y2=0
cc_264 N_A_315_54#_c_269_n N_A_309_338#_c_398_n 0.00278437f $X=3.27 $Y=1.665
+ $X2=0 $Y2=0
cc_265 N_A_315_54#_c_268_n N_A_309_338#_c_391_n 0.0147863f $X=4.115 $Y=1.22
+ $X2=0 $Y2=0
cc_266 N_A_315_54#_c_277_n N_CLK_c_470_n 0.00755872f $X=3.945 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A_315_54#_c_279_n N_CLK_c_470_n 0.00382838f $X=4.102 $Y=2.102 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_315_54#_c_280_n N_CLK_c_470_n 0.00490916f $X=4.095 $Y=2.11 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_315_54#_c_268_n N_CLK_c_466_n 0.00445076f $X=4.115 $Y=1.22 $X2=0
+ $Y2=0
cc_270 N_A_315_54#_c_279_n N_CLK_c_471_n 2.03939e-19 $X=4.102 $Y=2.102 $X2=0
+ $Y2=0
cc_271 N_A_315_54#_c_268_n CLK 0.0209126f $X=4.115 $Y=1.22 $X2=0 $Y2=0
cc_272 N_A_315_54#_c_268_n N_CLK_c_469_n 0.0173356f $X=4.115 $Y=1.22 $X2=0 $Y2=0
cc_273 N_A_315_54#_M1004_g N_A_27_74#_M1016_g 0.0131462f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_315_54#_M1007_g N_A_27_74#_M1010_g 0.0387775f $X=2.345 $Y=2.75 $X2=0
+ $Y2=0
cc_275 N_A_315_54#_M1014_g N_A_27_74#_M1010_g 0.0167945f $X=3.31 $Y=2.41 $X2=0
+ $Y2=0
cc_276 N_A_315_54#_c_274_n N_A_27_74#_M1010_g 0.0138346f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_277 N_A_315_54#_c_351_p N_A_27_74#_M1010_g 0.00504885f $X=3.115 $Y=2.305
+ $X2=0 $Y2=0
cc_278 N_A_315_54#_M1004_g N_A_27_74#_c_511_n 0.00889043f $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_279 N_A_315_54#_M1004_g N_A_27_74#_c_514_n 0.0138204f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_315_54#_M1014_g N_A_27_74#_c_515_n 0.0122425f $X=3.31 $Y=2.41 $X2=0
+ $Y2=0
cc_281 N_A_315_54#_c_274_n N_A_27_74#_c_515_n 0.00820717f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_282 N_A_315_54#_c_275_n N_A_27_74#_c_515_n 0.00134234f $X=2.3 $Y=2.215 $X2=0
+ $Y2=0
cc_283 N_A_315_54#_c_276_n N_A_27_74#_c_515_n 0.00472182f $X=3.115 $Y=2.05 $X2=0
+ $Y2=0
cc_284 N_A_315_54#_c_269_n N_A_27_74#_c_515_n 0.00331054f $X=3.27 $Y=1.665 $X2=0
+ $Y2=0
cc_285 N_A_315_54#_c_270_n N_A_27_74#_c_515_n 0.0194451f $X=3.27 $Y=1.665 $X2=0
+ $Y2=0
cc_286 N_A_315_54#_c_274_n N_A_27_74#_c_527_n 0.00789146f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_287 N_A_315_54#_c_275_n N_A_27_74#_c_527_n 0.0193895f $X=2.3 $Y=2.215 $X2=0
+ $Y2=0
cc_288 N_A_315_54#_c_264_n N_A_27_74#_c_539_n 0.00124375f $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_289 N_A_315_54#_c_264_n N_A_27_74#_c_522_n 0.0119481f $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_290 N_A_315_54#_M1004_g N_A_27_74#_c_523_n 6.13725e-19 $X=3.335 $Y=0.995
+ $X2=0 $Y2=0
cc_291 N_A_315_54#_c_274_n N_VPWR_M1010_d 0.0033399f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_292 N_A_315_54#_c_276_n N_VPWR_M1010_d 8.64634e-19 $X=3.115 $Y=2.05 $X2=0
+ $Y2=0
cc_293 N_A_315_54#_c_351_p N_VPWR_M1010_d 0.00471146f $X=3.115 $Y=2.305 $X2=0
+ $Y2=0
cc_294 N_A_315_54#_M1007_g N_VPWR_c_709_n 0.00142492f $X=2.345 $Y=2.75 $X2=0
+ $Y2=0
cc_295 N_A_315_54#_M1014_g N_VPWR_c_709_n 0.0042229f $X=3.31 $Y=2.41 $X2=0 $Y2=0
cc_296 N_A_315_54#_c_274_n N_VPWR_c_709_n 0.00824218f $X=3.03 $Y=2.215 $X2=0
+ $Y2=0
cc_297 N_A_315_54#_c_351_p N_VPWR_c_709_n 0.0115793f $X=3.115 $Y=2.305 $X2=0
+ $Y2=0
cc_298 N_A_315_54#_c_277_n N_VPWR_c_710_n 0.0178842f $X=3.945 $Y=2.475 $X2=0
+ $Y2=0
cc_299 N_A_315_54#_M1007_g N_VPWR_c_715_n 0.00522399f $X=2.345 $Y=2.75 $X2=0
+ $Y2=0
cc_300 N_A_315_54#_M1014_g N_VPWR_c_716_n 0.00585197f $X=3.31 $Y=2.41 $X2=0
+ $Y2=0
cc_301 N_A_315_54#_c_277_n N_VPWR_c_716_n 0.00851122f $X=3.945 $Y=2.475 $X2=0
+ $Y2=0
cc_302 N_A_315_54#_M1007_g N_VPWR_c_707_n 0.00984518f $X=2.345 $Y=2.75 $X2=0
+ $Y2=0
cc_303 N_A_315_54#_M1014_g N_VPWR_c_707_n 0.00606454f $X=3.31 $Y=2.41 $X2=0
+ $Y2=0
cc_304 N_A_315_54#_c_277_n N_VPWR_c_707_n 0.0372005f $X=3.945 $Y=2.475 $X2=0
+ $Y2=0
cc_305 N_A_315_54#_c_351_p N_VPWR_c_707_n 0.00202923f $X=3.115 $Y=2.305 $X2=0
+ $Y2=0
cc_306 N_A_315_54#_M1004_g N_VGND_c_828_n 0.00774033f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_315_54#_M1004_g N_VGND_c_814_n 0.00779576f $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_315_54#_c_264_n N_VGND_c_817_n 9.29978e-19 $X=1.65 $Y=1.15 $X2=0
+ $Y2=0
cc_309 N_A_315_54#_M1004_g N_VGND_c_823_n 7.34656e-19 $X=3.335 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_A_309_338#_c_389_n N_CLK_c_466_n 0.00722606f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_311 N_A_309_338#_c_389_n N_A_27_74#_c_511_n 0.0061136f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_312 N_A_309_338#_c_387_n N_A_27_74#_c_514_n 0.0119084f $X=3.465 $Y=1.245
+ $X2=0 $Y2=0
cc_313 N_A_309_338#_M1001_g N_A_27_74#_c_515_n 0.0072772f $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_314 N_A_309_338#_c_385_n N_A_27_74#_c_515_n 0.00526915f $X=2.37 $Y=1.675
+ $X2=0 $Y2=0
cc_315 N_A_309_338#_c_386_n N_A_27_74#_c_515_n 0.02065f $X=2.37 $Y=1.675 $X2=0
+ $Y2=0
cc_316 N_A_309_338#_c_387_n N_A_27_74#_c_515_n 0.00932416f $X=3.465 $Y=1.245
+ $X2=0 $Y2=0
cc_317 N_A_309_338#_c_387_n N_A_27_74#_c_521_n 0.00285995f $X=3.465 $Y=1.245
+ $X2=0 $Y2=0
cc_318 N_A_309_338#_M1001_g N_A_27_74#_c_522_n 0.00658236f $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_319 N_A_309_338#_M1001_g N_A_27_74#_c_523_n 0.0418981f $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_320 N_A_309_338#_c_392_n N_VPWR_c_715_n 0.00365603f $X=1.635 $Y=1.84 $X2=0
+ $Y2=0
cc_321 N_A_309_338#_c_392_n N_VPWR_c_707_n 0.00448802f $X=1.635 $Y=1.84 $X2=0
+ $Y2=0
cc_322 N_A_309_338#_c_387_n N_VGND_M1016_d 0.00469367f $X=3.465 $Y=1.245 $X2=0
+ $Y2=0
cc_323 N_A_309_338#_M1001_g N_VGND_c_828_n 7.00177e-19 $X=2.31 $Y=0.83 $X2=0
+ $Y2=0
cc_324 N_A_309_338#_c_387_n N_VGND_c_828_n 0.0279461f $X=3.465 $Y=1.245 $X2=0
+ $Y2=0
cc_325 N_A_309_338#_c_389_n N_VGND_c_814_n 0.00346039f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_326 N_A_309_338#_c_389_n N_VGND_c_815_n 0.0134733f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_327 N_A_309_338#_c_389_n N_VGND_c_820_n 0.00663535f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_328 N_A_309_338#_c_389_n N_VGND_c_823_n 0.00833855f $X=3.55 $Y=0.77 $X2=0
+ $Y2=0
cc_329 N_CLK_c_466_n N_A_27_74#_c_511_n 0.00894529f $X=4.335 $Y=1.475 $X2=0
+ $Y2=0
cc_330 N_CLK_M1012_g N_A_27_74#_c_511_n 0.00907339f $X=4.845 $Y=0.945 $X2=0
+ $Y2=0
cc_331 N_CLK_M1012_g N_A_27_74#_M1009_g 0.0253528f $X=4.845 $Y=0.945 $X2=0 $Y2=0
cc_332 CLK N_A_27_74#_M1011_g 0.00281729f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_333 N_CLK_c_469_n N_A_27_74#_M1011_g 0.0314654f $X=4.845 $Y=1.677 $X2=0 $Y2=0
cc_334 N_CLK_c_469_n N_A_27_74#_c_516_n 0.0253528f $X=4.845 $Y=1.677 $X2=0 $Y2=0
cc_335 N_CLK_M1012_g N_A_990_393#_c_648_n 0.00151317f $X=4.845 $Y=0.945 $X2=0
+ $Y2=0
cc_336 CLK N_A_990_393#_c_649_n 0.0120025f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_337 N_CLK_c_469_n N_A_990_393#_c_649_n 0.00101064f $X=4.845 $Y=1.677 $X2=0
+ $Y2=0
cc_338 N_CLK_c_471_n N_A_990_393#_c_654_n 0.00930083f $X=4.86 $Y=1.88 $X2=0
+ $Y2=0
cc_339 N_CLK_c_471_n N_A_990_393#_c_659_n 0.00211055f $X=4.86 $Y=1.88 $X2=0
+ $Y2=0
cc_340 CLK N_A_990_393#_c_659_n 0.0153044f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_341 N_CLK_M1012_g N_A_990_393#_c_651_n 0.0010598f $X=4.845 $Y=0.945 $X2=0
+ $Y2=0
cc_342 CLK N_A_990_393#_c_651_n 0.0116912f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_343 N_CLK_c_470_n N_VPWR_c_710_n 0.00420746f $X=4.32 $Y=1.88 $X2=0 $Y2=0
cc_344 N_CLK_c_471_n N_VPWR_c_710_n 0.0042704f $X=4.86 $Y=1.88 $X2=0 $Y2=0
cc_345 CLK N_VPWR_c_710_n 0.0228784f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_346 N_CLK_c_469_n N_VPWR_c_710_n 0.00478242f $X=4.845 $Y=1.677 $X2=0 $Y2=0
cc_347 N_CLK_c_471_n N_VPWR_c_712_n 0.00551389f $X=4.86 $Y=1.88 $X2=0 $Y2=0
cc_348 N_CLK_c_470_n N_VPWR_c_716_n 0.00542625f $X=4.32 $Y=1.88 $X2=0 $Y2=0
cc_349 N_CLK_c_470_n N_VPWR_c_707_n 0.00597552f $X=4.32 $Y=1.88 $X2=0 $Y2=0
cc_350 N_CLK_c_471_n N_VPWR_c_707_n 0.00597552f $X=4.86 $Y=1.88 $X2=0 $Y2=0
cc_351 N_CLK_c_466_n N_VGND_c_815_n 0.0200484f $X=4.335 $Y=1.475 $X2=0 $Y2=0
cc_352 N_CLK_M1012_g N_VGND_c_815_n 0.00730266f $X=4.845 $Y=0.945 $X2=0 $Y2=0
cc_353 CLK N_VGND_c_815_n 0.0212606f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_354 N_CLK_c_469_n N_VGND_c_815_n 0.00436753f $X=4.845 $Y=1.677 $X2=0 $Y2=0
cc_355 N_CLK_c_466_n N_VGND_c_823_n 7.97988e-19 $X=4.335 $Y=1.475 $X2=0 $Y2=0
cc_356 N_CLK_M1012_g N_VGND_c_823_n 9.49986e-19 $X=4.845 $Y=0.945 $X2=0 $Y2=0
cc_357 N_A_27_74#_M1011_g N_A_990_393#_M1005_g 0.00923223f $X=5.32 $Y=2.385
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_M1009_g N_A_990_393#_c_646_n 9.88035e-19 $X=5.235 $Y=0.945
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_516_n N_A_990_393#_c_646_n 0.012306f $X=5.285 $Y=1.49 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_M1009_g N_A_990_393#_c_648_n 0.0100958f $X=5.235 $Y=0.945
+ $X2=0 $Y2=0
cc_361 N_A_27_74#_M1011_g N_A_990_393#_c_649_n 0.0101259f $X=5.32 $Y=2.385 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_M1011_g N_A_990_393#_c_654_n 0.0149168f $X=5.32 $Y=2.385 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_M1011_g N_A_990_393#_c_659_n 0.0177339f $X=5.32 $Y=2.385 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_516_n N_A_990_393#_c_659_n 0.00137716f $X=5.285 $Y=1.49
+ $X2=0 $Y2=0
cc_365 N_A_27_74#_M1009_g N_A_990_393#_c_651_n 0.00624269f $X=5.235 $Y=0.945
+ $X2=0 $Y2=0
cc_366 N_A_27_74#_M1011_g N_A_990_393#_c_651_n 0.003544f $X=5.32 $Y=2.385 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_516_n N_A_990_393#_c_651_n 0.00927666f $X=5.285 $Y=1.49
+ $X2=0 $Y2=0
cc_368 N_A_27_74#_c_528_n N_VPWR_c_708_n 0.0261579f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_369 N_A_27_74#_M1010_g N_VPWR_c_709_n 0.0098771f $X=2.765 $Y=2.75 $X2=0 $Y2=0
cc_370 N_A_27_74#_M1011_g N_VPWR_c_711_n 0.0102738f $X=5.32 $Y=2.385 $X2=0 $Y2=0
cc_371 N_A_27_74#_M1011_g N_VPWR_c_712_n 0.00543421f $X=5.32 $Y=2.385 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_528_n N_VPWR_c_714_n 0.0154414f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_373 N_A_27_74#_M1010_g N_VPWR_c_715_n 0.00490827f $X=2.765 $Y=2.75 $X2=0
+ $Y2=0
cc_374 N_A_27_74#_M1010_g N_VPWR_c_707_n 0.00968584f $X=2.765 $Y=2.75 $X2=0
+ $Y2=0
cc_375 N_A_27_74#_M1011_g N_VPWR_c_707_n 0.00597552f $X=5.32 $Y=2.385 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_528_n N_VPWR_c_707_n 0.0127129f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_377 N_A_27_74#_c_535_n N_VGND_M1017_d 0.0132019f $X=1.045 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_378 N_A_27_74#_c_539_n N_VGND_M1017_d 0.00441864f $X=1.13 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_379 N_A_27_74#_c_518_n N_VGND_M1017_d 2.44449e-19 $X=1.215 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_74#_c_517_n N_VGND_c_813_n 0.0104927f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_535_n N_VGND_c_813_n 0.0196232f $X=1.045 $Y=0.875 $X2=0
+ $Y2=0
cc_382 N_A_27_74#_c_539_n N_VGND_c_813_n 0.0145482f $X=1.13 $Y=0.79 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_518_n N_VGND_c_813_n 0.0145354f $X=1.215 $Y=0.34 $X2=0 $Y2=0
cc_384 N_A_27_74#_M1016_g N_VGND_c_828_n 0.00917897f $X=2.7 $Y=0.83 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_511_n N_VGND_c_828_n 0.00138507f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_514_n N_VGND_c_828_n 0.00126939f $X=2.82 $Y=1.19 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_521_n N_VGND_c_828_n 0.0122171f $X=2.79 $Y=0.345 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_523_n N_VGND_c_828_n 0.00251883f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_389 N_A_27_74#_M1016_g N_VGND_c_814_n 0.00316397f $X=2.7 $Y=0.83 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_511_n N_VGND_c_814_n 0.0163869f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_521_n N_VGND_c_814_n 0.0198501f $X=2.79 $Y=0.345 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_523_n N_VGND_c_814_n 0.00172991f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_511_n N_VGND_c_815_n 0.0257165f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_394 N_A_27_74#_M1009_g N_VGND_c_815_n 0.00806567f $X=5.235 $Y=0.945 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_511_n N_VGND_c_816_n 0.0111053f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_396 N_A_27_74#_M1009_g N_VGND_c_816_n 8.98699e-19 $X=5.235 $Y=0.945 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_c_518_n N_VGND_c_817_n 0.0122203f $X=1.215 $Y=0.34 $X2=0 $Y2=0
cc_398 N_A_27_74#_c_522_n N_VGND_c_817_n 0.111626f $X=2.625 $Y=0.382 $X2=0 $Y2=0
cc_399 N_A_27_74#_c_523_n N_VGND_c_817_n 0.0121847f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_400 N_A_27_74#_c_517_n N_VGND_c_819_n 0.0154563f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_401 N_A_27_74#_c_511_n N_VGND_c_820_n 0.0350534f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_402 N_A_27_74#_c_511_n N_VGND_c_821_n 0.0215943f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_403 N_A_27_74#_c_511_n N_VGND_c_823_n 0.0817763f $X=5.16 $Y=0.18 $X2=0 $Y2=0
cc_404 N_A_27_74#_c_517_n N_VGND_c_823_n 0.012737f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_405 N_A_27_74#_c_535_n N_VGND_c_823_n 0.0126469f $X=1.045 $Y=0.875 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_518_n N_VGND_c_823_n 0.00661553f $X=1.215 $Y=0.34 $X2=0
+ $Y2=0
cc_407 N_A_27_74#_c_522_n N_VGND_c_823_n 0.0640172f $X=2.625 $Y=0.382 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_523_n N_VGND_c_823_n 0.0102842f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_522_n A_267_80# 0.00151475f $X=2.625 $Y=0.382 $X2=-0.19
+ $Y2=-0.245
cc_410 N_A_990_393#_c_649_n N_VPWR_M1011_d 2.93405e-19 $X=5.45 $Y=1.975 $X2=0
+ $Y2=0
cc_411 N_A_990_393#_c_659_n N_VPWR_M1011_d 0.00441497f $X=5.45 $Y=2.06 $X2=0
+ $Y2=0
cc_412 N_A_990_393#_c_654_n N_VPWR_c_710_n 0.0263057f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_413 N_A_990_393#_M1005_g N_VPWR_c_711_n 0.00534567f $X=6.145 $Y=2.4 $X2=0
+ $Y2=0
cc_414 N_A_990_393#_c_646_n N_VPWR_c_711_n 0.00687408f $X=6.055 $Y=1.465 $X2=0
+ $Y2=0
cc_415 N_A_990_393#_c_649_n N_VPWR_c_711_n 0.00234978f $X=5.45 $Y=1.975 $X2=0
+ $Y2=0
cc_416 N_A_990_393#_c_650_n N_VPWR_c_711_n 0.0158782f $X=5.87 $Y=1.465 $X2=0
+ $Y2=0
cc_417 N_A_990_393#_c_654_n N_VPWR_c_711_n 0.0251355f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_418 N_A_990_393#_c_659_n N_VPWR_c_711_n 0.0141779f $X=5.45 $Y=2.06 $X2=0
+ $Y2=0
cc_419 N_A_990_393#_c_654_n N_VPWR_c_712_n 0.00883445f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_420 N_A_990_393#_M1005_g N_VPWR_c_717_n 0.005209f $X=6.145 $Y=2.4 $X2=0 $Y2=0
cc_421 N_A_990_393#_M1005_g N_VPWR_c_707_n 0.00990688f $X=6.145 $Y=2.4 $X2=0
+ $Y2=0
cc_422 N_A_990_393#_c_654_n N_VPWR_c_707_n 0.0108836f $X=5.095 $Y=2.14 $X2=0
+ $Y2=0
cc_423 N_A_990_393#_M1013_g N_GCLK_c_794_n 0.0179032f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_424 N_A_990_393#_c_647_n N_GCLK_c_794_n 0.00953446f $X=6.055 $Y=1.3 $X2=0
+ $Y2=0
cc_425 N_A_990_393#_c_650_n N_GCLK_c_794_n 0.0154371f $X=5.87 $Y=1.465 $X2=0
+ $Y2=0
cc_426 N_A_990_393#_c_651_n N_GCLK_c_794_n 0.00478285f $X=5.285 $Y=1.12 $X2=0
+ $Y2=0
cc_427 N_A_990_393#_M1005_g GCLK 0.00530566f $X=6.145 $Y=2.4 $X2=0 $Y2=0
cc_428 N_A_990_393#_c_647_n GCLK 0.00661996f $X=6.055 $Y=1.3 $X2=0 $Y2=0
cc_429 N_A_990_393#_c_649_n GCLK 0.0083676f $X=5.45 $Y=1.975 $X2=0 $Y2=0
cc_430 N_A_990_393#_c_650_n GCLK 0.00638763f $X=5.87 $Y=1.465 $X2=0 $Y2=0
cc_431 N_A_990_393#_M1005_g N_GCLK_c_797_n 0.020296f $X=6.145 $Y=2.4 $X2=0 $Y2=0
cc_432 N_A_990_393#_c_648_n N_VGND_c_815_n 0.0074529f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_433 N_A_990_393#_c_651_n N_VGND_c_815_n 0.00326799f $X=5.285 $Y=1.12 $X2=0
+ $Y2=0
cc_434 N_A_990_393#_M1013_g N_VGND_c_816_n 0.00647412f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_435 N_A_990_393#_c_646_n N_VGND_c_816_n 0.00715849f $X=6.055 $Y=1.465 $X2=0
+ $Y2=0
cc_436 N_A_990_393#_c_648_n N_VGND_c_816_n 0.0339721f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_437 N_A_990_393#_c_650_n N_VGND_c_816_n 0.015939f $X=5.87 $Y=1.465 $X2=0
+ $Y2=0
cc_438 N_A_990_393#_c_651_n N_VGND_c_816_n 6.6261e-19 $X=5.285 $Y=1.12 $X2=0
+ $Y2=0
cc_439 N_A_990_393#_c_648_n N_VGND_c_821_n 0.00702137f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_440 N_A_990_393#_M1013_g N_VGND_c_822_n 0.00434272f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A_990_393#_M1013_g N_VGND_c_823_n 0.00828941f $X=6.225 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_990_393#_c_648_n N_VGND_c_823_n 0.0100521f $X=5.45 $Y=0.77 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_711_n N_GCLK_c_797_n 0.0407863f $X=5.87 $Y=2.11 $X2=0 $Y2=0
cc_444 N_VPWR_c_717_n N_GCLK_c_797_n 0.0176724f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_445 N_VPWR_c_707_n N_GCLK_c_797_n 0.0145596f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_446 N_GCLK_c_794_n N_VGND_c_816_n 0.0294122f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_447 N_GCLK_c_794_n N_VGND_c_822_n 0.0145639f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_448 N_GCLK_c_794_n N_VGND_c_823_n 0.0119984f $X=6.44 $Y=0.515 $X2=0 $Y2=0

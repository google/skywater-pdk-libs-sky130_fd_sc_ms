* File: sky130_fd_sc_ms__o21ba_4.pex.spice
* Created: Wed Sep  2 12:22:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21BA_4%B1_N 3 7 8 11 13
r33 11 14 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.385
+ $X2=0.585 $Y2=1.55
r34 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.385
+ $X2=0.585 $Y2=1.22
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.385 $X2=0.59 $Y2=1.385
r36 8 12 4.04912 $w=3.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.59 $Y2=1.365
r37 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.525 $Y=0.74
+ $X2=0.525 $Y2=1.22
r38 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%A_193_48# 1 2 3 12 16 20 24 28 32 36 40 42
+ 51 52 53 54 60 63 64 66 68 70 72 83
c158 66 0 8.37567e-20 $X=5.06 $Y=2.3
c159 54 0 9.42363e-21 $X=3.66 $Y=1.375
c160 36 0 7.8786e-20 $X=2.34 $Y=0.74
c161 12 0 1.76934e-19 $X=1.04 $Y=0.74
r162 83 84 10.1392 $w=3.09e-07 $l=6.5e-08 $layer=POLY_cond $X=2.34 $Y=1.455
+ $X2=2.405 $Y2=1.455
r163 80 81 7.01942 $w=3.09e-07 $l=4.5e-08 $layer=POLY_cond $X=1.91 $Y=1.455
+ $X2=1.955 $Y2=1.455
r164 77 78 3.89968 $w=3.09e-07 $l=2.5e-08 $layer=POLY_cond $X=1.48 $Y=1.455
+ $X2=1.505 $Y2=1.455
r165 66 74 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.06 $Y=2.3
+ $X2=5.06 $Y2=2.125
r166 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.06 $Y=2.3 $X2=5.06
+ $Y2=2.57
r167 65 72 0.414005 $w=3.5e-07 $l=3.42491e-07 $layer=LI1_cond $X=3.83 $Y=2.125
+ $X2=3.49 $Y2=2.13
r168 64 74 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=2.125
+ $X2=5.06 $Y2=2.125
r169 64 65 37.7014 $w=3.48e-07 $l=1.145e-06 $layer=LI1_cond $X=4.975 $Y=2.125
+ $X2=3.83 $Y2=2.125
r170 63 72 7.71803 $w=2.1e-07 $l=3.33054e-07 $layer=LI1_cond $X=3.745 $Y=1.95
+ $X2=3.49 $Y2=2.13
r171 62 63 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.745 $Y=1.46
+ $X2=3.745 $Y2=1.95
r172 58 60 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.665 $Y=0.425
+ $X2=3.665 $Y2=0.615
r173 55 70 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.98 $Y=1.375
+ $X2=2.895 $Y2=1.455
r174 54 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.66 $Y=1.375
+ $X2=3.745 $Y2=1.46
r175 54 55 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.66 $Y=1.375
+ $X2=2.98 $Y2=1.375
r176 52 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.5 $Y=0.34
+ $X2=3.665 $Y2=0.425
r177 52 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.5 $Y=0.34
+ $X2=2.98 $Y2=0.34
r178 51 70 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=1.29
+ $X2=2.895 $Y2=1.455
r179 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.895 $Y=0.425
+ $X2=2.98 $Y2=0.34
r180 50 51 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.895 $Y=0.425
+ $X2=2.895 $Y2=1.29
r181 49 83 1.55987 $w=3.09e-07 $l=1e-08 $layer=POLY_cond $X=2.33 $Y=1.455
+ $X2=2.34 $Y2=1.455
r182 49 81 58.4951 $w=3.09e-07 $l=3.75e-07 $layer=POLY_cond $X=2.33 $Y=1.455
+ $X2=1.955 $Y2=1.455
r183 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.455 $X2=2.33 $Y2=1.455
r184 45 80 40.5566 $w=3.09e-07 $l=2.6e-07 $layer=POLY_cond $X=1.65 $Y=1.455
+ $X2=1.91 $Y2=1.455
r185 45 78 22.6181 $w=3.09e-07 $l=1.45e-07 $layer=POLY_cond $X=1.65 $Y=1.455
+ $X2=1.505 $Y2=1.455
r186 44 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.65 $Y=1.455
+ $X2=2.33 $Y2=1.455
r187 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.455 $X2=1.65 $Y2=1.455
r188 42 70 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=1.455
+ $X2=2.895 $Y2=1.455
r189 42 48 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.81 $Y=1.455
+ $X2=2.33 $Y2=1.455
r190 38 84 15.404 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.62
+ $X2=2.405 $Y2=1.455
r191 38 40 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=2.405 $Y=1.62
+ $X2=2.405 $Y2=2.4
r192 34 83 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.29
+ $X2=2.34 $Y2=1.455
r193 34 36 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.34 $Y=1.29
+ $X2=2.34 $Y2=0.74
r194 30 81 15.404 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.62
+ $X2=1.955 $Y2=1.455
r195 30 32 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=1.955 $Y=1.62
+ $X2=1.955 $Y2=2.4
r196 26 80 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.29
+ $X2=1.91 $Y2=1.455
r197 26 28 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.91 $Y=1.29
+ $X2=1.91 $Y2=0.74
r198 22 78 15.404 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.62
+ $X2=1.505 $Y2=1.455
r199 22 24 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=1.505 $Y=1.62
+ $X2=1.505 $Y2=2.4
r200 18 77 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=1.29
+ $X2=1.48 $Y2=1.455
r201 18 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.48 $Y=1.29
+ $X2=1.48 $Y2=0.74
r202 14 77 66.2945 $w=3.09e-07 $l=4.25e-07 $layer=POLY_cond $X=1.055 $Y=1.455
+ $X2=1.48 $Y2=1.455
r203 14 75 2.33981 $w=3.09e-07 $l=1.5e-08 $layer=POLY_cond $X=1.055 $Y=1.455
+ $X2=1.04 $Y2=1.455
r204 14 16 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.055 $Y=1.55
+ $X2=1.055 $Y2=2.4
r205 10 75 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.29
+ $X2=1.04 $Y2=1.455
r206 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.04 $Y=1.29
+ $X2=1.04 $Y2=0.74
r207 3 74 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.96 $X2=5.06 $Y2=2.115
r208 3 68 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.96 $X2=5.06 $Y2=2.57
r209 2 72 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.44
+ $Y=2.12 $X2=3.575 $Y2=2.295
r210 1 60 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.47 $X2=3.665 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%A_27_368# 1 2 9 13 17 21 25 30 33 35 38 39
+ 41 42 43 47 53
c95 25 0 1.76934e-19 $X=0.31 $Y=0.515
r96 53 54 12.2413 $w=3.15e-07 $l=8e-08 $layer=POLY_cond $X=3.8 $Y=1.795 $X2=3.88
+ $Y2=1.795
r97 52 53 53.5556 $w=3.15e-07 $l=3.5e-07 $layer=POLY_cond $X=3.45 $Y=1.795
+ $X2=3.8 $Y2=1.795
r98 51 52 15.3016 $w=3.15e-07 $l=1e-07 $layer=POLY_cond $X=3.35 $Y=1.795
+ $X2=3.45 $Y2=1.795
r99 48 51 3.8254 $w=3.15e-07 $l=2.5e-08 $layer=POLY_cond $X=3.325 $Y=1.795
+ $X2=3.35 $Y2=1.795
r100 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.325
+ $Y=1.795 $X2=3.325 $Y2=1.795
r101 44 47 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.235 $Y=1.795
+ $X2=3.325 $Y2=1.795
r102 41 42 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=1.82
r103 39 42 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.17 $Y=1.01
+ $X2=0.17 $Y2=1.82
r104 37 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=1.96
+ $X2=3.235 $Y2=1.795
r105 37 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.235 $Y=1.96
+ $X2=3.235 $Y2=2.39
r106 36 43 4.14084 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.475
+ $X2=0.265 $Y2=2.475
r107 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.15 $Y=2.475
+ $X2=3.235 $Y2=2.39
r108 35 36 176.476 $w=1.68e-07 $l=2.705e-06 $layer=LI1_cond $X=3.15 $Y=2.475
+ $X2=0.445 $Y2=2.475
r109 31 43 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.56
+ $X2=0.265 $Y2=2.475
r110 31 33 8.16314 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.265 $Y=2.56
+ $X2=0.265 $Y2=2.815
r111 30 43 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.265 $Y2=2.475
r112 29 41 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=1.985
r113 29 30 12.4848 $w=3.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=2.39
r114 23 39 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=0.28 $Y=0.815
+ $X2=0.28 $Y2=1.01
r115 23 25 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=0.28 $Y=0.815
+ $X2=0.28 $Y2=0.515
r116 19 54 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.88 $Y=1.63
+ $X2=3.88 $Y2=1.795
r117 19 21 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.88 $Y=1.63
+ $X2=3.88 $Y2=0.79
r118 15 53 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.96 $X2=3.8
+ $Y2=1.795
r119 15 17 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.8 $Y=1.96 $X2=3.8
+ $Y2=2.54
r120 11 52 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.45 $Y=1.63
+ $X2=3.45 $Y2=1.795
r121 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.45 $Y=1.63
+ $X2=3.45 $Y2=0.79
r122 7 51 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.96 $X2=3.35
+ $Y2=1.795
r123 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.35 $Y=1.96 $X2=3.35
+ $Y2=2.54
r124 2 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r125 2 33 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r126 1 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%A2 3 7 11 15 17 18 19 28
c53 28 0 5.14477e-20 $X=5.285 $Y=1.615
c54 15 0 1.44963e-19 $X=5.31 $Y=0.945
c55 11 0 8.37567e-20 $X=5.285 $Y=2.46
c56 7 0 7.82385e-20 $X=4.88 $Y=0.945
r57 28 29 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.285 $Y=1.615
+ $X2=5.31 $Y2=1.615
r58 26 28 40.5352 $w=3.27e-07 $l=2.75e-07 $layer=POLY_cond $X=5.01 $Y=1.615
+ $X2=5.285 $Y2=1.615
r59 24 26 19.1621 $w=3.27e-07 $l=1.3e-07 $layer=POLY_cond $X=4.88 $Y=1.615
+ $X2=5.01 $Y2=1.615
r60 23 24 6.63303 $w=3.27e-07 $l=4.5e-08 $layer=POLY_cond $X=4.835 $Y=1.615
+ $X2=4.88 $Y2=1.615
r61 18 19 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.615 $X2=6
+ $Y2=1.615
r62 17 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.01 $Y=1.615
+ $X2=5.52 $Y2=1.615
r63 17 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.615 $X2=5.01 $Y2=1.615
r64 13 29 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.45
+ $X2=5.31 $Y2=1.615
r65 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.31 $Y=1.45
+ $X2=5.31 $Y2=0.945
r66 9 28 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.78
+ $X2=5.285 $Y2=1.615
r67 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.285 $Y=1.78
+ $X2=5.285 $Y2=2.46
r68 5 24 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.45
+ $X2=4.88 $Y2=1.615
r69 5 7 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.88 $Y=1.45 $X2=4.88
+ $Y2=0.945
r70 1 23 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.78
+ $X2=4.835 $Y2=1.615
r71 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=4.835 $Y=1.78
+ $X2=4.835 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%A1 3 8 9 10 11 13 18 20 23
c70 23 0 9.42363e-21 $X=4.34 $Y=1.615
c71 8 0 4.38187e-20 $X=4.38 $Y=0.945
r72 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.34 $Y=1.615
+ $X2=4.34 $Y2=1.78
r73 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.34 $Y=1.615
+ $X2=4.34 $Y2=1.45
r74 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.34
+ $Y=1.615 $X2=4.34 $Y2=1.615
r75 20 24 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.34 $Y2=1.615
r76 18 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.74 $Y=0.945
+ $X2=5.74 $Y2=1.34
r77 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.74 $Y=0.255
+ $X2=5.74 $Y2=0.945
r78 11 19 36.2738 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.735 $Y=1.43
+ $X2=5.735 $Y2=1.34
r79 11 13 400.371 $w=1.8e-07 $l=1.03e-06 $layer=POLY_cond $X=5.735 $Y=1.43
+ $X2=5.735 $Y2=2.46
r80 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.665 $Y=0.18
+ $X2=5.74 $Y2=0.255
r81 9 10 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.665 $Y=0.18
+ $X2=4.455 $Y2=0.18
r82 8 25 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.38 $Y=0.945
+ $X2=4.38 $Y2=1.45
r83 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.38 $Y=0.255
+ $X2=4.455 $Y2=0.18
r84 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.38 $Y=0.255 $X2=4.38
+ $Y2=0.945
r85 3 26 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=4.385 $Y=2.46
+ $X2=4.385 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%VPWR 1 2 3 4 5 18 22 26 28 30 34 36 41 51 56
+ 65 68 72 76 78 82
r78 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r79 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 74 76 9.31175 $w=6.83e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=3.072
+ $X2=3.205 $Y2=3.072
r81 71 74 1.39688 $w=6.83e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=3.072 $X2=3.12
+ $Y2=3.072
r82 71 72 17.8676 $w=6.83e-07 $l=5.75e-07 $layer=LI1_cond $X=3.04 $Y=3.072
+ $X2=2.465 $Y2=3.072
r83 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r86 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r87 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r90 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.11 $Y2=3.33
r92 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 56 81 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=5.875 $Y=3.33
+ $X2=6.057 $Y2=3.33
r94 56 62 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.875 $Y=3.33
+ $X2=5.52 $Y2=3.33
r95 55 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 54 76 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=3.205 $Y2=3.33
r97 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r98 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.11 $Y2=3.33
r99 51 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r100 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 49 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.465 $Y2=3.33
r102 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=1.73 $Y2=3.33
r104 47 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 45 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 45 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r108 42 65 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.805 $Y2=3.33
r109 42 44 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 41 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.73 $Y2=3.33
r111 41 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 39 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r114 36 65 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.805 $Y2=3.33
r115 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r116 34 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 34 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 34 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 30 33 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=6 $Y=2.115 $X2=6
+ $Y2=2.815
r120 28 81 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=6 $Y=3.245
+ $X2=6.057 $Y2=3.33
r121 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6 $Y=3.245 $X2=6
+ $Y2=2.815
r122 24 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r123 24 26 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.635
r124 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=3.33
r125 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=2.815
r126 16 65 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r127 16 18 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.815
r128 5 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.96 $X2=5.96 $Y2=2.815
r129 5 30 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.96 $X2=5.96 $Y2=2.115
r130 4 26 600 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=2.12 $X2=4.11 $Y2=2.635
r131 3 71 300 $w=1.7e-07 $l=1.21737e-06 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=3.04 $Y2=2.815
r132 2 22 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.73 $Y2=2.815
r133 1 18 600 $w=1.7e-07 $l=1.07488e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.805 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%X 1 2 3 4 15 21 23 27 29 30 31 36 38 41
c52 30 0 4.78765e-20 $X=1.115 $Y=1.58
c53 23 0 7.8786e-20 $X=1.96 $Y=1.035
r54 31 36 4.75094 $w=2.3e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.2
+ $Y2=1.82
r55 30 38 2.15457 $w=2.28e-07 $l=4.3e-08 $layer=LI1_cond $X=1.2 $Y=1.622 $X2=1.2
+ $Y2=1.665
r56 30 41 4.41536 $w=2.28e-07 $l=7.2e-08 $layer=LI1_cond $X=1.2 $Y=1.622 $X2=1.2
+ $Y2=1.55
r57 30 36 5.662 $w=2.28e-07 $l=1.13e-07 $layer=LI1_cond $X=1.2 $Y=1.707 $X2=1.2
+ $Y2=1.82
r58 30 38 2.10446 $w=2.28e-07 $l=4.2e-08 $layer=LI1_cond $X=1.2 $Y=1.707 $X2=1.2
+ $Y2=1.665
r59 25 27 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.085 $Y=0.95
+ $X2=2.085 $Y2=0.515
r60 24 29 1.59926 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.34 $Y=1.035
+ $X2=1.242 $Y2=1.035
r61 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.96 $Y=1.035
+ $X2=2.085 $Y2=0.95
r62 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.96 $Y=1.035
+ $X2=1.34 $Y2=1.035
r63 19 31 2.73179 $w=4e-07 $l=1.15e-07 $layer=LI1_cond $X=1.315 $Y=2.02 $X2=1.2
+ $Y2=2.02
r64 19 21 24.9216 $w=3.98e-07 $l=8.65e-07 $layer=LI1_cond $X=1.315 $Y=2.02
+ $X2=2.18 $Y2=2.02
r65 17 29 4.86787 $w=1.82e-07 $l=9.0802e-08 $layer=LI1_cond $X=1.23 $Y=1.12
+ $X2=1.242 $Y2=1.035
r66 17 41 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.23 $Y=1.12
+ $X2=1.23 $Y2=1.55
r67 13 29 4.86787 $w=1.82e-07 $l=8.5e-08 $layer=LI1_cond $X=1.242 $Y=0.95
+ $X2=1.242 $Y2=1.035
r68 13 15 24.7413 $w=1.93e-07 $l=4.35e-07 $layer=LI1_cond $X=1.242 $Y=0.95
+ $X2=1.242 $Y2=0.515
r69 4 21 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.84 $X2=2.18 $Y2=2.02
r70 3 31 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.28 $Y2=2.02
r71 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.985
+ $Y=0.37 $X2=2.125 $Y2=0.515
r72 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.115
+ $Y=0.37 $X2=1.255 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%A_895_392# 1 2 9 11 12 15
c28 15 0 5.14477e-20 $X=5.51 $Y=2.115
r29 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.51 $Y=2.115 $X2=5.51
+ $Y2=2.815
r30 13 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.51 $Y=2.905 $X2=5.51
+ $Y2=2.815
r31 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.345 $Y=2.99
+ $X2=5.51 $Y2=2.905
r32 11 12 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.345 $Y=2.99
+ $X2=4.775 $Y2=2.99
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.61 $Y=2.905
+ $X2=4.775 $Y2=2.99
r34 7 9 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.61 $Y=2.905 $X2=4.61
+ $Y2=2.635
r35 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=1.96 $X2=5.51 $Y2=2.815
r36 2 15 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=1.96 $X2=5.51 $Y2=2.115
r37 1 9 600 $w=1.7e-07 $l=7.39425e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.96 $X2=4.61 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%VGND 1 2 3 4 5 20 24 28 32 36 39 40 41 43 52
+ 56 63 64 67 70 73 76
r91 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r94 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 64 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r97 61 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.485
+ $Y2=0
r98 61 63 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=6
+ $Y2=0
r99 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r100 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r101 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 57 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.625
+ $Y2=0
r103 57 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=5.04
+ $Y2=0
r104 56 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.485
+ $Y2=0
r105 56 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.04
+ $Y2=0
r106 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r107 52 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.625
+ $Y2=0
r108 52 54 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=4.5 $Y=0 $X2=2.64
+ $Y2=0
r109 51 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r110 51 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r111 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 48 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.655
+ $Y2=0
r113 48 50 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r115 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.81
+ $Y2=0
r118 44 46 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.2
+ $Y2=0
r119 43 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.655
+ $Y2=0
r120 43 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.2
+ $Y2=0
r121 41 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.56 $Y2=0
r122 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r123 40 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=0 $X2=2.64
+ $Y2=0
r124 39 50 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.16
+ $Y2=0
r125 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.515
+ $Y2=0
r126 34 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=0.085
+ $X2=5.485 $Y2=0
r127 34 36 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.485 $Y=0.085
+ $X2=5.485 $Y2=0.77
r128 30 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0
r129 30 32 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=4.625 $Y=0.085
+ $X2=4.625 $Y2=0.77
r130 26 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0
r131 26 28 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0.515
r132 22 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0
r133 22 24 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0.565
r134 18 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0
r135 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0.495
r136 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.625 $X2=5.525 $Y2=0.77
r137 4 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.625 $X2=4.665 $Y2=0.77
r138 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.415
+ $Y=0.37 $X2=2.555 $Y2=0.515
r139 2 24 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.37 $X2=1.695 $Y2=0.565
r140 1 20 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.37 $X2=0.81 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_4%A_618_94# 1 2 3 4 15 17 18 19 22 26 28 32 34
+ 37
c61 34 0 7.82385e-20 $X=4.165 $Y=1.035
c62 26 0 1.44963e-19 $X=5.095 $Y=0.77
c63 17 0 4.38187e-20 $X=4 $Y=1.035
r64 34 35 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.165 $Y=1.035
+ $X2=4.165 $Y2=1.195
r65 30 32 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=5.957 $Y=1.11
+ $X2=5.957 $Y2=0.77
r66 29 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.18 $Y=1.195
+ $X2=5.055 $Y2=1.195
r67 28 30 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=5.79 $Y=1.195
+ $X2=5.957 $Y2=1.11
r68 28 29 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.79 $Y=1.195
+ $X2=5.18 $Y2=1.195
r69 24 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=1.11
+ $X2=5.055 $Y2=1.195
r70 24 26 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.055 $Y=1.11
+ $X2=5.055 $Y2=0.77
r71 23 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=1.195
+ $X2=4.165 $Y2=1.195
r72 22 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.93 $Y=1.195
+ $X2=5.055 $Y2=1.195
r73 22 23 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.93 $Y=1.195 $X2=4.33
+ $Y2=1.195
r74 19 34 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.95
+ $X2=4.165 $Y2=1.035
r75 19 21 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.95
+ $X2=4.165 $Y2=0.865
r76 17 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=1.035 $X2=4.165
+ $Y2=1.035
r77 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4 $Y=1.035 $X2=3.32
+ $Y2=1.035
r78 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.235 $Y=0.95
+ $X2=3.32 $Y2=1.035
r79 13 15 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.235 $Y=0.95
+ $X2=3.235 $Y2=0.855
r80 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.815
+ $Y=0.625 $X2=5.955 $Y2=0.77
r81 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.955
+ $Y=0.625 $X2=5.095 $Y2=0.77
r82 2 21 182 $w=1.7e-07 $l=4.88851e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.47 $X2=4.165 $Y2=0.865
r83 1 15 182 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.47 $X2=3.235 $Y2=0.855
.ends


* File: sky130_fd_sc_ms__inv_16.pxi.spice
* Created: Wed Sep  2 12:10:43 2020
* 
x_PM_SKY130_FD_SC_MS__INV_16%A N_A_M1004_g N_A_M1000_g N_A_M1006_g N_A_M1001_g
+ N_A_M1007_g N_A_M1002_g N_A_M1008_g N_A_M1003_g N_A_M1009_g N_A_M1005_g
+ N_A_M1011_g N_A_M1010_g N_A_M1012_g N_A_M1013_g N_A_M1014_g N_A_M1015_g
+ N_A_M1016_g N_A_M1019_g N_A_M1017_g N_A_M1020_g N_A_M1018_g N_A_M1023_g
+ N_A_M1021_g N_A_M1025_g N_A_M1022_g N_A_M1026_g N_A_M1024_g N_A_M1027_g
+ N_A_M1030_g N_A_M1028_g N_A_M1031_g N_A_M1029_g N_A_c_150_n N_A_c_151_n A
+ N_A_c_152_n N_A_c_153_n N_A_c_154_n N_A_c_155_n N_A_c_156_n N_A_c_157_n
+ N_A_c_158_n N_A_c_159_n N_A_c_186_n A PM_SKY130_FD_SC_MS__INV_16%A
x_PM_SKY130_FD_SC_MS__INV_16%VPWR N_VPWR_M1004_s N_VPWR_M1006_s N_VPWR_M1008_s
+ N_VPWR_M1011_s N_VPWR_M1015_s N_VPWR_M1020_s N_VPWR_M1025_s N_VPWR_M1027_s
+ N_VPWR_M1029_s N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n
+ N_VPWR_c_476_n N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n
+ N_VPWR_c_481_n N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n
+ N_VPWR_c_486_n VPWR N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_471_n
+ PM_SKY130_FD_SC_MS__INV_16%VPWR
x_PM_SKY130_FD_SC_MS__INV_16%Y N_Y_M1000_d N_Y_M1002_d N_Y_M1005_d N_Y_M1013_d
+ N_Y_M1016_d N_Y_M1018_d N_Y_M1022_d N_Y_M1030_d N_Y_M1004_d N_Y_M1007_d
+ N_Y_M1009_d N_Y_M1012_d N_Y_M1019_d N_Y_M1023_d N_Y_M1026_d N_Y_M1028_d
+ N_Y_c_618_n N_Y_c_632_n N_Y_c_619_n N_Y_c_634_n N_Y_c_620_n N_Y_c_621_n
+ N_Y_c_636_n N_Y_c_622_n N_Y_c_623_n N_Y_c_624_n N_Y_c_625_n N_Y_c_626_n
+ N_Y_c_702_n N_Y_c_627_n N_Y_c_628_n N_Y_c_629_n Y N_Y_c_637_n N_Y_c_630_n
+ N_Y_c_639_n N_Y_c_640_n N_Y_c_631_n N_Y_c_749_n N_Y_c_772_n N_Y_c_775_n
+ N_Y_c_778_n PM_SKY130_FD_SC_MS__INV_16%Y
x_PM_SKY130_FD_SC_MS__INV_16%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1003_s
+ N_VGND_M1010_s N_VGND_M1014_s N_VGND_M1017_s N_VGND_M1021_s N_VGND_M1024_s
+ N_VGND_M1031_s N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n
+ N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n
+ N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n
+ N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n VGND N_VGND_c_883_n
+ N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n
+ PM_SKY130_FD_SC_MS__INV_16%VGND
cc_1 VNB N_A_M1000_g 0.0298158f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_2 VNB N_A_M1001_g 0.0244831f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_M1002_g 0.0236443f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_4 VNB N_A_M1003_g 0.0246673f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_5 VNB N_A_M1005_g 0.0236422f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_6 VNB N_A_M1010_g 0.0236401f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.74
cc_7 VNB N_A_M1013_g 0.023639f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=0.74
cc_8 VNB N_A_M1014_g 0.0236474f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.74
cc_9 VNB N_A_M1016_g 0.0230083f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.74
cc_10 VNB N_A_M1017_g 0.0236404f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.74
cc_11 VNB N_A_M1018_g 0.024294f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=0.74
cc_12 VNB N_A_M1021_g 0.0245364f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=0.74
cc_13 VNB N_A_M1022_g 0.0251803f $X=-0.19 $Y=-0.245 $X2=6.145 $Y2=0.74
cc_14 VNB N_A_M1024_g 0.0247749f $X=-0.19 $Y=-0.245 $X2=6.575 $Y2=0.74
cc_15 VNB N_A_M1030_g 0.0256095f $X=-0.19 $Y=-0.245 $X2=7.165 $Y2=0.74
cc_16 VNB N_A_M1031_g 0.0298291f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=0.74
cc_17 VNB N_A_c_150_n 0.0185028f $X=-0.19 $Y=-0.245 $X2=7.09 $Y2=1.515
cc_18 VNB N_A_c_151_n 0.0448647f $X=-0.19 $Y=-0.245 $X2=7.655 $Y2=1.515
cc_19 VNB N_A_c_152_n 0.277968f $X=-0.19 $Y=-0.245 $X2=6.745 $Y2=1.515
cc_20 VNB N_A_c_153_n 0.0023355f $X=-0.19 $Y=-0.245 $X2=6.925 $Y2=1.515
cc_21 VNB N_A_c_154_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.515
cc_22 VNB N_A_c_155_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.515
cc_23 VNB N_A_c_156_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=1.515
cc_24 VNB N_A_c_157_n 0.00101987f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=1.515
cc_25 VNB N_A_c_158_n 0.00173377f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=1.515
cc_26 VNB N_A_c_159_n 0.0022845f $X=-0.19 $Y=-0.245 $X2=5.93 $Y2=1.515
cc_27 VNB N_VPWR_c_471_n 0.342803f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.515
cc_28 VNB N_Y_c_618_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=2.4
cc_29 VNB N_Y_c_619_n 0.00468918f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.68
cc_30 VNB N_Y_c_620_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=4.255 $Y2=1.68
cc_31 VNB N_Y_c_621_n 0.00417093f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=1.35
cc_32 VNB N_Y_c_622_n 0.00219079f $X=-0.19 $Y=-0.245 $X2=4.705 $Y2=2.4
cc_33 VNB N_Y_c_623_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=1.35
cc_34 VNB N_Y_c_624_n 0.00237467f $X=-0.19 $Y=-0.245 $X2=5.145 $Y2=0.74
cc_35 VNB N_Y_c_625_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=5.175 $Y2=1.68
cc_36 VNB N_Y_c_626_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=1.35
cc_37 VNB N_Y_c_627_n 0.00169784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_628_n 0.00142546f $X=-0.19 $Y=-0.245 $X2=5.655 $Y2=1.68
cc_39 VNB N_Y_c_629_n 0.00101819f $X=-0.19 $Y=-0.245 $X2=6.145 $Y2=1.35
cc_40 VNB N_Y_c_630_n 0.00473182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_631_n 0.00203504f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=1.515
cc_42 VNB N_VGND_c_866_n 0.0131032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_867_n 0.0502481f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_44 VNB N_VGND_c_868_n 0.00986225f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=2.4
cc_45 VNB N_VGND_c_869_n 0.0103371f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=0.74
cc_46 VNB N_VGND_c_870_n 0.0100559f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=2.4
cc_47 VNB N_VGND_c_871_n 0.00669123f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=0.74
cc_48 VNB N_VGND_c_872_n 0.0105034f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=2.4
cc_49 VNB N_VGND_c_873_n 0.012516f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=0.74
cc_50 VNB N_VGND_c_874_n 0.0121504f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.74
cc_51 VNB N_VGND_c_875_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_876_n 0.0567567f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=2.4
cc_53 VNB N_VGND_c_877_n 0.0181599f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=1.35
cc_54 VNB N_VGND_c_878_n 0.00482535f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.74
cc_55 VNB N_VGND_c_879_n 0.0173725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_880_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.255 $Y2=1.68
cc_57 VNB N_VGND_c_881_n 0.0191493f $X=-0.19 $Y=-0.245 $X2=4.255 $Y2=2.4
cc_58 VNB N_VGND_c_882_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_883_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=4.645 $Y2=0.74
cc_60 VNB N_VGND_c_884_n 0.0183708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_885_n 0.018851f $X=-0.19 $Y=-0.245 $X2=5.175 $Y2=1.68
cc_62 VNB N_VGND_c_886_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_887_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_888_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=7.165 $Y2=1.35
cc_65 VNB N_VGND_c_889_n 0.00538573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_890_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=7.205 $Y2=2.4
cc_67 VNB N_VGND_c_891_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=7.595 $Y2=0.74
cc_68 VNB N_VGND_c_892_n 0.436313f $X=-0.19 $Y=-0.245 $X2=7.655 $Y2=2.4
cc_69 VPB N_A_M1004_g 0.0256794f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_70 VPB N_A_M1006_g 0.0211046f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_71 VPB N_A_M1007_g 0.0210512f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_72 VPB N_A_M1008_g 0.0208015f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=2.4
cc_73 VPB N_A_M1009_g 0.0208028f $X=-0.19 $Y=1.66 $X2=2.405 $Y2=2.4
cc_74 VPB N_A_M1011_g 0.020801f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=2.4
cc_75 VPB N_A_M1012_g 0.0207998f $X=-0.19 $Y=1.66 $X2=3.355 $Y2=2.4
cc_76 VPB N_A_M1015_g 0.0205756f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=2.4
cc_77 VPB N_A_M1019_g 0.0202363f $X=-0.19 $Y=1.66 $X2=4.255 $Y2=2.4
cc_78 VPB N_A_M1020_g 0.0207175f $X=-0.19 $Y=1.66 $X2=4.705 $Y2=2.4
cc_79 VPB N_A_M1023_g 0.0205593f $X=-0.19 $Y=1.66 $X2=5.175 $Y2=2.4
cc_80 VPB N_A_M1025_g 0.0216787f $X=-0.19 $Y=1.66 $X2=5.655 $Y2=2.4
cc_81 VPB N_A_M1026_g 0.021322f $X=-0.19 $Y=1.66 $X2=6.205 $Y2=2.4
cc_82 VPB N_A_M1027_g 0.0213216f $X=-0.19 $Y=1.66 $X2=6.655 $Y2=2.4
cc_83 VPB N_A_M1028_g 0.0216776f $X=-0.19 $Y=1.66 $X2=7.205 $Y2=2.4
cc_84 VPB N_A_M1029_g 0.0273126f $X=-0.19 $Y=1.66 $X2=7.655 $Y2=2.4
cc_85 VPB N_A_c_150_n 0.00615867f $X=-0.19 $Y=1.66 $X2=7.09 $Y2=1.515
cc_86 VPB N_A_c_151_n 0.00506647f $X=-0.19 $Y=1.66 $X2=7.655 $Y2=1.515
cc_87 VPB N_A_c_152_n 0.0565484f $X=-0.19 $Y=1.66 $X2=6.745 $Y2=1.515
cc_88 VPB N_A_c_153_n 0.00200161f $X=-0.19 $Y=1.66 $X2=6.925 $Y2=1.515
cc_89 VPB N_A_c_154_n 0.00179173f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.515
cc_90 VPB N_A_c_155_n 0.00198947f $X=-0.19 $Y=1.66 $X2=2.17 $Y2=1.515
cc_91 VPB N_A_c_156_n 0.00178763f $X=-0.19 $Y=1.66 $X2=3.11 $Y2=1.515
cc_92 VPB N_A_c_157_n 0.00157069f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.515
cc_93 VPB N_A_c_158_n 0.00145671f $X=-0.19 $Y=1.66 $X2=4.935 $Y2=1.515
cc_94 VPB N_A_c_159_n 0.00185727f $X=-0.19 $Y=1.66 $X2=5.93 $Y2=1.515
cc_95 VPB N_A_c_186_n 0.00893936f $X=-0.19 $Y=1.66 $X2=6.925 $Y2=1.665
cc_96 VPB N_VPWR_c_472_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_473_n 0.0645074f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_98 VPB N_VPWR_c_474_n 0.00917612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_475_n 0.00884785f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=2.4
cc_100 VPB N_VPWR_c_476_n 0.0081889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_477_n 0.00741052f $X=-0.19 $Y=1.66 $X2=3.355 $Y2=0.74
cc_102 VPB N_VPWR_c_478_n 0.00488809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_479_n 0.00836214f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=0.74
cc_104 VPB N_VPWR_c_480_n 0.00824466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_481_n 0.0116305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_482_n 0.0645306f $X=-0.19 $Y=1.66 $X2=4.705 $Y2=2.4
cc_107 VPB N_VPWR_c_483_n 0.0189682f $X=-0.19 $Y=1.66 $X2=5.145 $Y2=0.74
cc_108 VPB N_VPWR_c_484_n 0.00449427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_485_n 0.0186691f $X=-0.19 $Y=1.66 $X2=5.175 $Y2=2.4
cc_110 VPB N_VPWR_c_486_n 0.00528033f $X=-0.19 $Y=1.66 $X2=5.175 $Y2=2.4
cc_111 VPB N_VPWR_c_487_n 0.0193352f $X=-0.19 $Y=1.66 $X2=5.575 $Y2=0.74
cc_112 VPB N_VPWR_c_488_n 0.0196495f $X=-0.19 $Y=1.66 $X2=5.655 $Y2=2.4
cc_113 VPB N_VPWR_c_489_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_490_n 0.0186412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_491_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_492_n 0.0179727f $X=-0.19 $Y=1.66 $X2=7.595 $Y2=1.35
cc_117 VPB N_VPWR_c_493_n 0.00555219f $X=-0.19 $Y=1.66 $X2=7.165 $Y2=1.515
cc_118 VPB N_VPWR_c_494_n 0.0047828f $X=-0.19 $Y=1.66 $X2=7.655 $Y2=1.515
cc_119 VPB N_VPWR_c_495_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_496_n 0.00632158f $X=-0.19 $Y=1.66 $X2=6.925 $Y2=1.515
cc_121 VPB N_VPWR_c_497_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_471_n 0.0771804f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.515
cc_123 VPB N_Y_c_632_n 0.00231613f $X=-0.19 $Y=1.66 $X2=3.785 $Y2=1.35
cc_124 VPB N_Y_c_619_n 9.14116e-19 $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.68
cc_125 VPB N_Y_c_634_n 0.00231613f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=1.35
cc_126 VPB N_Y_c_621_n 9.14222e-19 $X=-0.19 $Y=1.66 $X2=4.645 $Y2=1.35
cc_127 VPB N_Y_c_636_n 0.00231613f $X=-0.19 $Y=1.66 $X2=4.705 $Y2=1.68
cc_128 VPB N_Y_c_637_n 0.00225767f $X=-0.19 $Y=1.66 $X2=6.205 $Y2=1.68
cc_129 VPB N_Y_c_630_n 0.00333766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_Y_c_639_n 0.00367812f $X=-0.19 $Y=1.66 $X2=7.205 $Y2=2.4
cc_131 VPB N_Y_c_640_n 0.00231613f $X=-0.19 $Y=1.66 $X2=7.655 $Y2=1.68
cc_132 VPB N_Y_c_631_n 0.00375772f $X=-0.19 $Y=1.66 $X2=7.595 $Y2=1.515
cc_133 N_A_M1004_g N_VPWR_c_473_n 0.00622149f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A_M1006_g N_VPWR_c_474_n 0.00331759f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_M1007_g N_VPWR_c_474_n 0.00356293f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_c_152_n N_VPWR_c_474_n 7.49127e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A_c_154_n N_VPWR_c_474_n 0.0186213f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_186_n N_VPWR_c_474_n 8.28135e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_139 N_A_M1008_g N_VPWR_c_475_n 0.00337371f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_M1009_g N_VPWR_c_475_n 0.00347237f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_c_152_n N_VPWR_c_475_n 7.50577e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_c_155_n N_VPWR_c_475_n 0.017259f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_c_186_n N_VPWR_c_475_n 7.92963e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_144 N_A_M1011_g N_VPWR_c_476_n 0.00337371f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_M1012_g N_VPWR_c_476_n 0.00216006f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_c_152_n N_VPWR_c_476_n 7.5094e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A_c_156_n N_VPWR_c_476_n 0.017259f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_c_186_n N_VPWR_c_476_n 7.92963e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_149 N_A_M1015_g N_VPWR_c_477_n 0.00211108f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1019_g N_VPWR_c_477_n 0.00209433f $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_c_152_n N_VPWR_c_477_n 4.80934e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A_c_157_n N_VPWR_c_477_n 0.0155724f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A_c_186_n N_VPWR_c_477_n 7.45001e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_154 N_A_M1020_g N_VPWR_c_478_n 0.00217407f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_M1023_g N_VPWR_c_478_n 0.0134216f $X=5.175 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_M1025_g N_VPWR_c_478_n 6.67972e-19 $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_c_152_n N_VPWR_c_478_n 5.88936e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A_c_158_n N_VPWR_c_478_n 0.0181297f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A_c_186_n N_VPWR_c_478_n 0.00102938f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_160 N_A_M1025_g N_VPWR_c_479_n 0.00236601f $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_M1026_g N_VPWR_c_479_n 0.00233698f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_c_152_n N_VPWR_c_479_n 0.00101587f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A_c_159_n N_VPWR_c_479_n 0.0222679f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A_c_186_n N_VPWR_c_479_n 0.00106883f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_165 N_A_M1027_g N_VPWR_c_480_n 0.00233698f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_M1028_g N_VPWR_c_480_n 0.00229781f $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A_c_150_n N_VPWR_c_480_n 0.00101732f $X=7.09 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A_c_153_n N_VPWR_c_480_n 0.0219612f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A_c_186_n N_VPWR_c_480_n 9.92096e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_170 N_A_M1028_g N_VPWR_c_482_n 6.87624e-19 $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_M1029_g N_VPWR_c_482_n 0.0184536f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_M1012_g N_VPWR_c_483_n 0.005209f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A_M1015_g N_VPWR_c_483_n 0.00553757f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_M1019_g N_VPWR_c_485_n 0.00549225f $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_M1020_g N_VPWR_c_485_n 0.00537895f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A_M1004_g N_VPWR_c_487_n 0.00520504f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_M1006_g N_VPWR_c_487_n 0.00531971f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A_M1007_g N_VPWR_c_488_n 0.005209f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_M1008_g N_VPWR_c_488_n 0.005209f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_M1009_g N_VPWR_c_489_n 0.005209f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_M1011_g N_VPWR_c_489_n 0.005209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_M1023_g N_VPWR_c_490_n 0.00521592f $X=5.175 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_M1025_g N_VPWR_c_490_n 0.00537895f $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_M1026_g N_VPWR_c_491_n 0.005209f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A_M1027_g N_VPWR_c_491_n 0.005209f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A_M1028_g N_VPWR_c_492_n 0.005209f $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_M1029_g N_VPWR_c_492_n 0.00521592f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_M1004_g N_VPWR_c_471_n 0.00985724f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_M1006_g N_VPWR_c_471_n 0.0101836f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_M1007_g N_VPWR_c_471_n 0.00982082f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_M1008_g N_VPWR_c_471_n 0.00982754f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_M1009_g N_VPWR_c_471_n 0.00982082f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_M1011_g N_VPWR_c_471_n 0.00982754f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_M1012_g N_VPWR_c_471_n 0.00982082f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_M1015_g N_VPWR_c_471_n 0.0108799f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_M1019_g N_VPWR_c_471_n 0.0106941f $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_M1020_g N_VPWR_c_471_n 0.0103671f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_M1023_g N_VPWR_c_471_n 0.0102928f $X=5.175 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_M1025_g N_VPWR_c_471_n 0.0103785f $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_M1026_g N_VPWR_c_471_n 0.00982526f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_M1027_g N_VPWR_c_471_n 0.00982526f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_M1028_g N_VPWR_c_471_n 0.00982526f $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_M1029_g N_VPWR_c_471_n 0.0102898f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_M1000_g N_Y_c_618_n 0.00772833f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_M1001_g N_Y_c_618_n 0.00746162f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_M1007_g N_Y_c_632_n 0.0103361f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_M1008_g N_Y_c_632_n 0.0109404f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_M1001_g N_Y_c_619_n 8.65347e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_M1007_g N_Y_c_619_n 0.00176373f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_M1002_g N_Y_c_619_n 0.0151729f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_M1008_g N_Y_c_619_n 0.00556477f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_M1003_g N_Y_c_619_n 0.00396849f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_M1009_g N_Y_c_619_n 8.86537e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_c_152_n N_Y_c_619_n 0.0213664f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A_c_154_n N_Y_c_619_n 0.0286379f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A_c_155_n N_Y_c_619_n 0.0285602f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_c_186_n N_Y_c_619_n 0.0319887f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_218 N_A_M1009_g N_Y_c_634_n 0.0108027f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_M1011_g N_Y_c_634_n 0.0114071f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_M1008_g N_Y_c_620_n 5.01231e-19 $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A_M1003_g N_Y_c_620_n 8.58503e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_M1009_g N_Y_c_620_n 0.00554828f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_M1005_g N_Y_c_620_n 0.015703f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_M1011_g N_Y_c_620_n 0.00584779f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_M1010_g N_Y_c_620_n 0.0156374f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_M1012_g N_Y_c_620_n 8.82859e-19 $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_M1013_g N_Y_c_620_n 8.54281e-19 $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_c_152_n N_Y_c_620_n 0.0219828f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A_c_155_n N_Y_c_620_n 0.0286379f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_230 N_A_c_156_n N_Y_c_620_n 0.0285726f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_231 N_A_c_186_n N_Y_c_620_n 0.033789f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_232 N_A_M1015_g N_Y_c_621_n 9.04147e-19 $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_M1016_g N_Y_c_621_n 0.00354167f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_M1019_g N_Y_c_621_n 0.00503491f $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_M1017_g N_Y_c_621_n 0.0154727f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_M1020_g N_Y_c_621_n 0.0016976f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_M1018_g N_Y_c_621_n 8.71251e-19 $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_c_152_n N_Y_c_621_n 0.0202692f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A_c_157_n N_Y_c_621_n 0.0283691f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A_c_158_n N_Y_c_621_n 0.0284993f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A_c_186_n N_Y_c_621_n 0.0286815f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_242 N_A_M1019_g N_Y_c_636_n 0.00945159f $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_M1020_g N_Y_c_636_n 0.0100453f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_M1018_g N_Y_c_622_n 0.00526964f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_M1021_g N_Y_c_622_n 0.0110561f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_M1022_g N_Y_c_622_n 9.81084e-19 $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_c_152_n N_Y_c_622_n 0.007852f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A_c_158_n N_Y_c_622_n 0.00658047f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A_c_159_n N_Y_c_622_n 0.00676348f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_250 N_A_c_186_n N_Y_c_622_n 0.00205475f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_251 N_A_M1018_g N_Y_c_623_n 0.00722691f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_M1021_g N_Y_c_623_n 0.00830039f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_M1022_g N_Y_c_624_n 0.00815379f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_M1024_g N_Y_c_624_n 0.0120406f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_M1030_g N_Y_c_624_n 9.51769e-19 $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_c_152_n N_Y_c_624_n 0.00846048f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_257 N_A_c_153_n N_Y_c_624_n 0.00735182f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_258 N_A_c_159_n N_Y_c_624_n 0.00737762f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_259 N_A_c_186_n N_Y_c_624_n 0.00280382f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_260 N_A_M1022_g N_Y_c_625_n 0.0080359f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_M1024_g N_Y_c_625_n 0.00821155f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_M1030_g N_Y_c_626_n 0.00753493f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_M1031_g N_Y_c_626_n 0.00772833f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_M1000_g N_Y_c_702_n 0.00362234f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_c_152_n N_Y_c_702_n 0.0145286f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_266 N_A_c_154_n N_Y_c_702_n 0.0279825f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_267 N_A_M1000_g N_Y_c_627_n 0.0102796f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_M1001_g N_Y_c_627_n 0.00319122f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_M1000_g N_Y_c_628_n 0.00198651f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_M1001_g N_Y_c_628_n 0.0031608f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_M1030_g N_Y_c_629_n 0.0031805f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A_M1031_g N_Y_c_629_n 0.00198651f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_M1004_g N_Y_c_637_n 0.0239154f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_274 N_A_M1006_g N_Y_c_637_n 0.0177678f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A_M1007_g N_Y_c_637_n 8.28785e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A_c_152_n N_Y_c_637_n 0.0184221f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_277 N_A_c_186_n N_Y_c_637_n 0.00187673f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_278 N_A_M1011_g N_Y_c_630_n 8.3139e-19 $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A_M1010_g N_Y_c_630_n 8.44821e-19 $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_M1012_g N_Y_c_630_n 0.0175554f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A_M1013_g N_Y_c_630_n 0.0148554f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_M1014_g N_Y_c_630_n 0.00398243f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A_M1015_g N_Y_c_630_n 0.00252788f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A_c_152_n N_Y_c_630_n 0.0214323f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_285 N_A_c_156_n N_Y_c_630_n 0.0293067f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_286 N_A_c_157_n N_Y_c_630_n 0.0285407f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_287 N_A_c_186_n N_Y_c_630_n 0.0324168f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_288 N_A_M1023_g N_Y_c_639_n 0.00223303f $X=5.175 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A_M1025_g N_Y_c_639_n 0.0170218f $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A_M1026_g N_Y_c_639_n 0.0010986f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A_c_152_n N_Y_c_639_n 0.0150997f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_292 N_A_c_158_n N_Y_c_639_n 0.021723f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_293 N_A_c_159_n N_Y_c_639_n 0.0220708f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_294 N_A_c_186_n N_Y_c_639_n 0.0340778f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_295 N_A_M1025_g N_Y_c_640_n 0.00110853f $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A_M1026_g N_Y_c_640_n 0.0183475f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A_M1027_g N_Y_c_640_n 0.0182438f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A_M1028_g N_Y_c_640_n 8.06796e-19 $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A_c_152_n N_Y_c_640_n 0.0141736f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_300 N_A_c_153_n N_Y_c_640_n 0.0214823f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_301 N_A_c_159_n N_Y_c_640_n 0.0215141f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_302 N_A_c_186_n N_Y_c_640_n 0.0352047f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_303 N_A_M1027_g N_Y_c_631_n 7.61077e-19 $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A_M1030_g N_Y_c_631_n 0.0051716f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_M1028_g N_Y_c_631_n 0.0180168f $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A_M1031_g N_Y_c_631_n 0.0113953f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_M1029_g N_Y_c_631_n 0.00474937f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_308 N_A_c_151_n N_Y_c_631_n 0.0316196f $X=7.655 $Y=1.515 $X2=0 $Y2=0
cc_309 N_A_c_153_n N_Y_c_631_n 0.0291941f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_310 N_A_c_186_n N_Y_c_631_n 0.00184883f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_311 N_A_M1006_g N_Y_c_749_n 0.0137675f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A_M1007_g N_Y_c_749_n 0.00797362f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A_M1008_g N_Y_c_749_n 0.00779332f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_314 N_A_M1009_g N_Y_c_749_n 0.0079486f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_315 N_A_M1011_g N_Y_c_749_n 0.00779332f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A_M1012_g N_Y_c_749_n 0.00777271f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_317 N_A_M1015_g N_Y_c_749_n 0.00926785f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_318 N_A_M1019_g N_Y_c_749_n 0.00906816f $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_319 N_A_M1020_g N_Y_c_749_n 0.00858409f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_320 N_A_M1023_g N_Y_c_749_n 0.00887943f $X=5.175 $Y=2.4 $X2=0 $Y2=0
cc_321 N_A_M1025_g N_Y_c_749_n 0.00854998f $X=5.655 $Y=2.4 $X2=0 $Y2=0
cc_322 N_A_M1026_g N_Y_c_749_n 0.00777271f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_323 N_A_M1027_g N_Y_c_749_n 0.00777271f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_324 N_A_M1028_g N_Y_c_749_n 0.0129071f $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A_M1029_g N_Y_c_749_n 0.00276416f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_326 N_A_c_153_n N_Y_c_749_n 0.00153204f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_327 N_A_c_154_n N_Y_c_749_n 0.00164778f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_328 N_A_c_155_n N_Y_c_749_n 0.00112367f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_329 N_A_c_156_n N_Y_c_749_n 0.00100926f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_330 N_A_c_157_n N_Y_c_749_n 0.00119042f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_331 N_A_c_158_n N_Y_c_749_n 0.00142273f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_332 N_A_c_159_n N_Y_c_749_n 0.0011424f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_333 N_A_c_186_n N_Y_c_749_n 0.592639f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_334 N_A_M1007_g N_Y_c_772_n 0.00201241f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A_M1008_g N_Y_c_772_n 0.00142298f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A_c_186_n N_Y_c_772_n 5.77561e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_337 N_A_M1009_g N_Y_c_775_n 0.00179794f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_338 N_A_M1011_g N_Y_c_775_n 0.00142298f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_339 N_A_c_186_n N_Y_c_775_n 3.38351e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_340 N_A_M1019_g N_Y_c_778_n 9.98284e-19 $X=4.255 $Y=2.4 $X2=0 $Y2=0
cc_341 N_A_M1020_g N_Y_c_778_n 0.00137743f $X=4.705 $Y=2.4 $X2=0 $Y2=0
cc_342 N_A_M1023_g N_Y_c_778_n 3.51193e-19 $X=5.175 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A_c_186_n N_Y_c_778_n 3.82569e-19 $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_344 N_A_M1000_g N_VGND_c_867_n 0.00525456f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A_c_152_n N_VGND_c_867_n 0.00132967f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_346 N_A_M1001_g N_VGND_c_868_n 0.00583652f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A_M1002_g N_VGND_c_868_n 0.00227436f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A_c_152_n N_VGND_c_868_n 0.00129886f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_349 N_A_c_154_n N_VGND_c_868_n 0.0167206f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_350 N_A_c_186_n N_VGND_c_868_n 0.00144887f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_351 N_A_M1003_g N_VGND_c_869_n 0.00238904f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_352 N_A_M1005_g N_VGND_c_869_n 0.00586329f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_c_152_n N_VGND_c_869_n 0.00130048f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_354 N_A_c_155_n N_VGND_c_869_n 0.018017f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_355 N_A_c_186_n N_VGND_c_869_n 0.00156118f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_356 N_A_M1010_g N_VGND_c_870_n 0.00230839f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A_M1013_g N_VGND_c_870_n 0.00231837f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A_c_152_n N_VGND_c_870_n 0.00130088f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_359 N_A_c_156_n N_VGND_c_870_n 0.0173688f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_360 N_A_c_186_n N_VGND_c_870_n 0.00150502f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_361 N_A_M1014_g N_VGND_c_871_n 0.00214082f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A_M1016_g N_VGND_c_871_n 0.0116992f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_M1017_g N_VGND_c_871_n 6.07804e-19 $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A_c_152_n N_VGND_c_871_n 7.63823e-19 $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_365 N_A_c_157_n N_VGND_c_871_n 0.0166865f $X=4.025 $Y=1.515 $X2=0 $Y2=0
cc_366 N_A_c_186_n N_VGND_c_871_n 0.00144416f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_367 N_A_M1017_g N_VGND_c_872_n 0.00214733f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A_M1018_g N_VGND_c_872_n 0.00353535f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A_c_152_n N_VGND_c_872_n 0.00129725f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_370 N_A_c_158_n N_VGND_c_872_n 0.0163965f $X=4.935 $Y=1.515 $X2=0 $Y2=0
cc_371 N_A_c_186_n N_VGND_c_872_n 0.00161813f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_372 N_A_M1021_g N_VGND_c_873_n 0.00789946f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A_M1022_g N_VGND_c_873_n 0.00803145f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A_c_152_n N_VGND_c_873_n 0.00244453f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_375 N_A_c_159_n N_VGND_c_873_n 0.0173678f $X=5.93 $Y=1.515 $X2=0 $Y2=0
cc_376 N_A_c_186_n N_VGND_c_873_n 0.00347842f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_377 N_A_M1024_g N_VGND_c_874_n 0.00814162f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A_M1030_g N_VGND_c_874_n 0.00688674f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A_c_150_n N_VGND_c_874_n 0.00175046f $X=7.09 $Y=1.515 $X2=0 $Y2=0
cc_380 N_A_c_152_n N_VGND_c_874_n 0.00139845f $X=6.745 $Y=1.515 $X2=0 $Y2=0
cc_381 N_A_c_153_n N_VGND_c_874_n 0.0176918f $X=6.925 $Y=1.515 $X2=0 $Y2=0
cc_382 N_A_c_186_n N_VGND_c_874_n 0.00408288f $X=6.925 $Y=1.665 $X2=0 $Y2=0
cc_383 N_A_M1031_g N_VGND_c_876_n 0.00532106f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A_c_151_n N_VGND_c_876_n 0.00132967f $X=7.655 $Y=1.515 $X2=0 $Y2=0
cc_385 N_A_M1013_g N_VGND_c_877_n 0.00445602f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A_M1014_g N_VGND_c_877_n 0.00461464f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A_M1016_g N_VGND_c_879_n 0.00429299f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A_M1017_g N_VGND_c_879_n 0.00434272f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_389 N_A_M1018_g N_VGND_c_881_n 0.00456932f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_390 N_A_M1021_g N_VGND_c_881_n 0.00434272f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A_M1000_g N_VGND_c_883_n 0.00434272f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A_M1001_g N_VGND_c_883_n 0.00434272f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A_M1002_g N_VGND_c_884_n 0.00445602f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A_M1003_g N_VGND_c_884_n 0.00461464f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A_M1005_g N_VGND_c_885_n 0.00445602f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A_M1010_g N_VGND_c_885_n 0.00445602f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A_M1022_g N_VGND_c_886_n 0.00434272f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_398 N_A_M1024_g N_VGND_c_886_n 0.00434272f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A_M1030_g N_VGND_c_887_n 0.00434272f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A_M1031_g N_VGND_c_887_n 0.00434272f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A_M1000_g N_VGND_c_892_n 0.00823934f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A_M1001_g N_VGND_c_892_n 0.00820718f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A_M1002_g N_VGND_c_892_n 0.00857405f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A_M1003_g N_VGND_c_892_n 0.00908319f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A_M1005_g N_VGND_c_892_n 0.00857405f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_M1010_g N_VGND_c_892_n 0.00857405f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A_M1013_g N_VGND_c_892_n 0.00857181f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_408 N_A_M1014_g N_VGND_c_892_n 0.00907773f $X=3.785 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A_M1016_g N_VGND_c_892_n 0.00847524f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_410 N_A_M1017_g N_VGND_c_892_n 0.00820718f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_411 N_A_M1018_g N_VGND_c_892_n 0.00890307f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_412 N_A_M1021_g N_VGND_c_892_n 0.00821518f $X=5.575 $Y=0.74 $X2=0 $Y2=0
cc_413 N_A_M1022_g N_VGND_c_892_n 0.00821294f $X=6.145 $Y=0.74 $X2=0 $Y2=0
cc_414 N_A_M1024_g N_VGND_c_892_n 0.00821668f $X=6.575 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A_M1030_g N_VGND_c_892_n 0.00821444f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A_M1031_g N_VGND_c_892_n 0.00823934f $X=7.595 $Y=0.74 $X2=0 $Y2=0
cc_417 N_VPWR_c_488_n N_Y_c_632_n 0.0144623f $X=2.045 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_471_n N_Y_c_632_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_419 N_VPWR_c_489_n N_Y_c_634_n 0.0144623f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_471_n N_Y_c_634_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_c_485_n N_Y_c_636_n 0.012797f $X=4.81 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_471_n N_Y_c_636_n 0.01055f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_423 N_VPWR_c_473_n N_Y_c_637_n 0.0404146f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_424 N_VPWR_c_474_n N_Y_c_637_n 0.0435605f $X=1.18 $Y=2.105 $X2=0 $Y2=0
cc_425 N_VPWR_c_487_n N_Y_c_637_n 0.0149495f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_426 N_VPWR_c_471_n N_Y_c_637_n 0.0116197f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_c_476_n N_Y_c_630_n 0.0419652f $X=3.08 $Y=2.105 $X2=0 $Y2=0
cc_428 N_VPWR_c_477_n N_Y_c_630_n 0.00758344f $X=4.03 $Y=2.105 $X2=0 $Y2=0
cc_429 N_VPWR_c_483_n N_Y_c_630_n 0.0129872f $X=3.915 $Y=3.33 $X2=0 $Y2=0
cc_430 N_VPWR_c_471_n N_Y_c_630_n 0.0106816f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_431 N_VPWR_c_478_n N_Y_c_639_n 0.0770296f $X=4.93 $Y=2.105 $X2=0 $Y2=0
cc_432 N_VPWR_c_479_n N_Y_c_639_n 0.0393523f $X=5.93 $Y=2.105 $X2=0 $Y2=0
cc_433 N_VPWR_c_490_n N_Y_c_639_n 0.0139245f $X=5.765 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_471_n N_Y_c_639_n 0.0114926f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_435 N_VPWR_c_479_n N_Y_c_640_n 0.0425672f $X=5.93 $Y=2.105 $X2=0 $Y2=0
cc_436 N_VPWR_c_480_n N_Y_c_640_n 0.0425672f $X=6.93 $Y=2.105 $X2=0 $Y2=0
cc_437 N_VPWR_c_491_n N_Y_c_640_n 0.0144623f $X=6.765 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_471_n N_Y_c_640_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_c_480_n N_Y_c_631_n 0.0417838f $X=6.93 $Y=2.105 $X2=0 $Y2=0
cc_440 N_VPWR_c_482_n N_Y_c_631_n 0.0427611f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_441 N_VPWR_c_492_n N_Y_c_631_n 0.0123179f $X=7.735 $Y=3.33 $X2=0 $Y2=0
cc_442 N_VPWR_c_471_n N_Y_c_631_n 0.0101276f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_443 N_VPWR_M1006_s N_Y_c_749_n 0.00334902f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_444 N_VPWR_M1008_s N_Y_c_749_n 0.00411448f $X=1.995 $Y=1.84 $X2=0 $Y2=0
cc_445 N_VPWR_M1011_s N_Y_c_749_n 0.00417089f $X=2.945 $Y=1.84 $X2=0 $Y2=0
cc_446 N_VPWR_M1015_s N_Y_c_749_n 0.00239084f $X=3.895 $Y=1.84 $X2=0 $Y2=0
cc_447 N_VPWR_M1020_s N_Y_c_749_n 0.00175943f $X=4.795 $Y=1.84 $X2=0 $Y2=0
cc_448 N_VPWR_M1025_s N_Y_c_749_n 0.00315275f $X=5.745 $Y=1.84 $X2=0 $Y2=0
cc_449 N_VPWR_M1027_s N_Y_c_749_n 0.00407615f $X=6.745 $Y=1.84 $X2=0 $Y2=0
cc_450 N_VPWR_c_473_n N_Y_c_749_n 0.00161913f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_451 N_VPWR_c_474_n N_Y_c_749_n 0.0278681f $X=1.18 $Y=2.105 $X2=0 $Y2=0
cc_452 N_VPWR_c_475_n N_Y_c_749_n 0.0246664f $X=2.13 $Y=2.105 $X2=0 $Y2=0
cc_453 N_VPWR_c_476_n N_Y_c_749_n 0.0246664f $X=3.08 $Y=2.105 $X2=0 $Y2=0
cc_454 N_VPWR_c_477_n N_Y_c_749_n 0.0236853f $X=4.03 $Y=2.105 $X2=0 $Y2=0
cc_455 N_VPWR_c_478_n N_Y_c_749_n 0.027209f $X=4.93 $Y=2.105 $X2=0 $Y2=0
cc_456 N_VPWR_c_479_n N_Y_c_749_n 0.0311183f $X=5.93 $Y=2.105 $X2=0 $Y2=0
cc_457 N_VPWR_c_480_n N_Y_c_749_n 0.0310485f $X=6.93 $Y=2.105 $X2=0 $Y2=0
cc_458 N_VPWR_c_482_n N_Y_c_749_n 0.00683675f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_459 N_VPWR_c_474_n N_Y_c_772_n 0.0425039f $X=1.18 $Y=2.105 $X2=0 $Y2=0
cc_460 N_VPWR_c_475_n N_Y_c_772_n 0.0369073f $X=2.13 $Y=2.105 $X2=0 $Y2=0
cc_461 N_VPWR_c_475_n N_Y_c_775_n 0.0424691f $X=2.13 $Y=2.105 $X2=0 $Y2=0
cc_462 N_VPWR_c_476_n N_Y_c_775_n 0.0369073f $X=3.08 $Y=2.105 $X2=0 $Y2=0
cc_463 N_VPWR_c_477_n N_Y_c_778_n 0.0379955f $X=4.03 $Y=2.105 $X2=0 $Y2=0
cc_464 N_VPWR_c_478_n N_Y_c_778_n 0.0398555f $X=4.93 $Y=2.105 $X2=0 $Y2=0
cc_465 N_Y_c_618_n N_VGND_c_867_n 0.0307549f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_466 N_Y_c_618_n N_VGND_c_868_n 0.0307549f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_467 N_Y_c_619_n N_VGND_c_868_n 0.028873f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_468 N_Y_c_619_n N_VGND_c_869_n 0.00297007f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_469 N_Y_c_620_n N_VGND_c_869_n 0.029171f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_470 N_Y_c_620_n N_VGND_c_870_n 0.0291629f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_471 N_Y_c_630_n N_VGND_c_870_n 0.0303029f $X=3.57 $Y=0.515 $X2=0 $Y2=0
cc_472 N_Y_c_621_n N_VGND_c_871_n 0.0272179f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_473 N_Y_c_630_n N_VGND_c_871_n 0.0296712f $X=3.57 $Y=0.515 $X2=0 $Y2=0
cc_474 N_Y_c_621_n N_VGND_c_872_n 0.0296586f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_475 N_Y_c_622_n N_VGND_c_872_n 0.00429585f $X=5.37 $Y=1.025 $X2=0 $Y2=0
cc_476 N_Y_c_623_n N_VGND_c_872_n 0.0236187f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_477 N_Y_c_622_n N_VGND_c_873_n 0.00450652f $X=5.37 $Y=1.025 $X2=0 $Y2=0
cc_478 N_Y_c_623_n N_VGND_c_873_n 0.0246826f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_479 N_Y_c_624_n N_VGND_c_873_n 0.0051297f $X=6.36 $Y=1.015 $X2=0 $Y2=0
cc_480 N_Y_c_625_n N_VGND_c_873_n 0.0257017f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_481 N_Y_c_624_n N_VGND_c_874_n 0.00490968f $X=6.36 $Y=1.015 $X2=0 $Y2=0
cc_482 N_Y_c_625_n N_VGND_c_874_n 0.0245613f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_483 N_Y_c_626_n N_VGND_c_874_n 0.0308181f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_484 N_Y_c_626_n N_VGND_c_876_n 0.0308109f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_485 N_Y_c_630_n N_VGND_c_877_n 0.0130321f $X=3.57 $Y=0.515 $X2=0 $Y2=0
cc_486 N_Y_c_621_n N_VGND_c_879_n 0.0112174f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_487 N_Y_c_623_n N_VGND_c_881_n 0.0136595f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_488 N_Y_c_618_n N_VGND_c_883_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_489 N_Y_c_619_n N_VGND_c_884_n 0.012809f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_490 N_Y_c_620_n N_VGND_c_885_n 0.0136595f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_491 N_Y_c_625_n N_VGND_c_886_n 0.0144922f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_492 N_Y_c_626_n N_VGND_c_887_n 0.0144922f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_493 N_Y_c_618_n N_VGND_c_892_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_494 N_Y_c_619_n N_VGND_c_892_n 0.0105693f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_495 N_Y_c_620_n N_VGND_c_892_n 0.0112404f $X=2.64 $Y=0.515 $X2=0 $Y2=0
cc_496 N_Y_c_621_n N_VGND_c_892_n 0.00922837f $X=4.43 $Y=0.515 $X2=0 $Y2=0
cc_497 N_Y_c_623_n N_VGND_c_892_n 0.0112404f $X=5.36 $Y=0.515 $X2=0 $Y2=0
cc_498 N_Y_c_625_n N_VGND_c_892_n 0.0118826f $X=6.36 $Y=0.515 $X2=0 $Y2=0
cc_499 N_Y_c_626_n N_VGND_c_892_n 0.0118826f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_500 N_Y_c_630_n N_VGND_c_892_n 0.0107539f $X=3.57 $Y=0.515 $X2=0 $Y2=0

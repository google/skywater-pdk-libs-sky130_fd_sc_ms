# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.825000 2.025000 2.155000 2.355000 ;
        RECT 1.985000 1.125000 2.375000 1.780000 ;
        RECT 1.985000 1.780000 2.155000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.145000 0.370000 8.450000 1.550000 ;
        RECT 8.145000 1.550000 8.515000 2.070000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.140000 1.820000 10.505000 2.980000 ;
        RECT 10.165000 0.350000 10.505000 1.130000 ;
        RECT 10.335000 1.130000 10.505000 1.820000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.585000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 0.730000 ;
      RECT  0.115000  0.730000  2.530000 0.900000 ;
      RECT  0.115000  0.900000  1.100000 1.010000 ;
      RECT  0.115000  1.720000  0.925000 1.890000 ;
      RECT  0.115000  1.890000  0.445000 2.980000 ;
      RECT  0.625000  0.085000  1.010000 0.560000 ;
      RECT  0.645000  2.060000  0.895000 3.245000 ;
      RECT  0.755000  1.010000  1.100000 1.550000 ;
      RECT  0.755000  1.550000  0.925000 1.720000 ;
      RECT  1.095000  1.815000  1.440000 2.625000 ;
      RECT  1.095000  2.625000  5.205000 2.795000 ;
      RECT  1.095000  2.795000  1.345000 2.980000 ;
      RECT  1.270000  1.070000  1.600000 1.485000 ;
      RECT  1.270000  1.485000  1.815000 1.815000 ;
      RECT  1.575000  2.965000  2.035000 3.245000 ;
      RECT  1.860000  0.085000  2.190000 0.560000 ;
      RECT  2.325000  2.205000  2.715000 2.455000 ;
      RECT  2.360000  0.255000  3.640000 0.425000 ;
      RECT  2.360000  0.425000  2.530000 0.730000 ;
      RECT  2.545000  1.070000  2.870000 1.240000 ;
      RECT  2.545000  1.240000  2.715000 2.205000 ;
      RECT  2.700000  0.595000  2.870000 1.070000 ;
      RECT  2.885000  1.410000  3.300000 1.580000 ;
      RECT  2.885000  1.580000  3.055000 2.285000 ;
      RECT  2.885000  2.285000  4.325000 2.455000 ;
      RECT  3.050000  0.595000  3.300000 1.410000 ;
      RECT  3.225000  1.750000  3.640000 2.065000 ;
      RECT  3.470000  0.425000  3.640000 0.780000 ;
      RECT  3.470000  0.780000  4.815000 0.950000 ;
      RECT  3.470000  0.950000  3.640000 1.750000 ;
      RECT  3.810000  1.120000  4.815000 1.450000 ;
      RECT  4.000000  2.965000  4.330000 3.245000 ;
      RECT  4.030000  0.085000  4.370000 0.610000 ;
      RECT  4.155000  1.630000  4.475000 1.960000 ;
      RECT  4.155000  1.960000  4.325000 2.285000 ;
      RECT  4.535000  2.180000  4.865000 2.455000 ;
      RECT  4.645000  0.255000  6.240000 0.530000 ;
      RECT  4.645000  0.530000  4.815000 0.780000 ;
      RECT  4.645000  1.450000  4.815000 2.180000 ;
      RECT  4.985000  1.120000  5.275000 1.450000 ;
      RECT  5.035000  1.450000  5.205000 2.625000 ;
      RECT  5.035000  2.795000  6.205000 2.965000 ;
      RECT  5.375000  1.620000  6.545000 1.670000 ;
      RECT  5.375000  1.670000  7.585000 1.790000 ;
      RECT  5.375000  1.790000  5.705000 2.625000 ;
      RECT  5.445000  0.530000  5.615000 1.170000 ;
      RECT  5.445000  1.170000  5.845000 1.450000 ;
      RECT  5.785000  0.700000  6.185000 0.950000 ;
      RECT  5.875000  1.960000  6.205000 2.795000 ;
      RECT  6.015000  0.950000  6.185000 1.620000 ;
      RECT  6.375000  1.790000  7.585000 1.960000 ;
      RECT  6.600000  2.375000  6.930000 3.245000 ;
      RECT  6.655000  0.085000  6.985000 1.000000 ;
      RECT  6.715000  1.170000  7.465000 1.330000 ;
      RECT  6.715000  1.330000  7.925000 1.500000 ;
      RECT  7.160000  2.130000  7.925000 2.240000 ;
      RECT  7.160000  2.240000  9.015000 2.410000 ;
      RECT  7.160000  2.410000  7.490000 2.980000 ;
      RECT  7.215000  0.370000  7.465000 1.170000 ;
      RECT  7.645000  0.085000  7.975000 1.150000 ;
      RECT  7.695000  2.580000  8.025000 3.245000 ;
      RECT  7.755000  1.500000  7.925000 2.130000 ;
      RECT  8.595000  2.580000  8.925000 3.245000 ;
      RECT  8.620000  0.085000  8.950000 1.150000 ;
      RECT  8.685000  1.320000  9.015000 2.240000 ;
      RECT  9.235000  0.540000  9.510000 1.300000 ;
      RECT  9.235000  1.300000 10.165000 1.630000 ;
      RECT  9.235000  1.630000  9.485000 2.860000 ;
      RECT  9.690000  1.820000  9.940000 3.245000 ;
      RECT  9.735000  0.085000  9.985000 1.130000 ;
      RECT 10.675000  0.085000 10.925000 1.130000 ;
      RECT 10.675000  1.820000 10.925000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_ms__dfxbp_2

* File: sky130_fd_sc_ms__xor3_4.pex.spice
* Created: Fri Aug 28 18:19:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_74_294# 1 2 3 4 15 19 23 24 26 27 31 34 35
+ 38 41 45 48 49 54
c116 38 0 3.89081e-20 $X=1.54 $Y=1.085
r117 52 54 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.08 $Y=1.1 $X2=4.24
+ $Y2=1.1
r118 48 50 19.8947 $w=6.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.99 $Y=2.07
+ $X2=3.99 $Y2=2.755
r119 48 49 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=2.07
+ $X2=3.99 $Y2=1.905
r120 42 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=1.265
+ $X2=4.24 $Y2=1.1
r121 42 49 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.24 $Y=1.265
+ $X2=4.24 $Y2=1.905
r122 41 50 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.74 $Y=2.905
+ $X2=3.74 $Y2=2.755
r123 36 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.84
+ $X2=1.54 $Y2=1.925
r124 36 38 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.54 $Y=1.84
+ $X2=1.54 $Y2=1.085
r125 34 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=2.99
+ $X2=3.74 $Y2=2.905
r126 34 35 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=3.655 $Y=2.99
+ $X2=1.395 $Y2=2.99
r127 31 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.23 $Y=2.105
+ $X2=1.23 $Y2=2.815
r128 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.395 $Y2=2.99
r129 29 33 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.815
r130 28 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.23 $Y=1.925
+ $X2=1.54 $Y2=1.925
r131 28 31 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.23 $Y=2.01
+ $X2=1.23 $Y2=2.105
r132 26 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=1.925
+ $X2=1.23 $Y2=1.925
r133 26 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.065 $Y=1.925
+ $X2=0.7 $Y2=1.925
r134 24 58 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.635
+ $X2=0.535 $Y2=1.8
r135 24 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.635
+ $X2=0.535 $Y2=1.47
r136 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.535
+ $Y=1.635 $X2=0.535 $Y2=1.635
r137 21 27 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=0.562 $Y=1.84
+ $X2=0.7 $Y2=1.925
r138 21 23 8.59094 $w=2.73e-07 $l=2.05e-07 $layer=LI1_cond $X=0.562 $Y=1.84
+ $X2=0.562 $Y2=1.635
r139 19 57 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=0.91
+ $X2=0.495 $Y2=1.47
r140 15 58 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=2.46
+ $X2=0.505 $Y2=1.8
r141 4 48 300 $w=1.7e-07 $l=5.25262e-07 $layer=licon1_PDIFF $count=2 $X=3.295
+ $Y=1.895 $X2=3.74 $Y2=2.07
r142 3 33 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.96 $X2=1.23 $Y2=2.815
r143 3 31 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.96 $X2=1.23 $Y2=2.105
r144 2 52 182 $w=1.7e-07 $l=6.10635e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.625 $X2=4.08 $Y2=1.1
r145 1 38 182 $w=1.7e-07 $l=6.27316e-07 $layer=licon1_NDIFF $count=1 $X=1.24
+ $Y=0.59 $X2=1.54 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A 3 7 8 11 13
c40 13 0 1.02266e-19 $X=1.075 $Y=1.34
r41 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.505
+ $X2=1.075 $Y2=1.67
r42 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.505
+ $X2=1.075 $Y2=1.34
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.505 $X2=1.075 $Y2=1.505
r44 8 12 6.45368 $w=3.73e-07 $l=2.1e-07 $layer=LI1_cond $X=1.097 $Y=1.295
+ $X2=1.097 $Y2=1.505
r45 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.165 $Y=0.91
+ $X2=1.165 $Y2=1.34
r46 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.005 $Y=2.46
+ $X2=1.005 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_397_320# 1 2 9 11 12 15 17 21 23 27 29 30
+ 32 33 34 38 41 48 49 51
c111 32 0 4.26801e-20 $X=3.74 $Y=1.435
c112 27 0 9.37054e-20 $X=3.695 $Y=0.945
c113 9 0 3.89081e-20 $X=2.075 $Y=2.28
r114 49 53 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.802 $Y=1.57
+ $X2=3.802 $Y2=1.405
r115 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.82
+ $Y=1.57 $X2=3.82 $Y2=1.57
r116 45 48 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=3.74 $Y=1.585
+ $X2=3.82 $Y2=1.585
r117 41 43 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.62 $Y=1.985
+ $X2=4.62 $Y2=2.815
r118 41 51 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.62 $Y=1.985
+ $X2=4.62 $Y2=1.13
r119 36 51 5.87448 $w=2.03e-07 $l=1.02e-07 $layer=LI1_cond $X=4.637 $Y=1.028
+ $X2=4.637 $Y2=1.13
r120 36 38 9.08914 $w=2.03e-07 $l=1.68e-07 $layer=LI1_cond $X=4.637 $Y=1.028
+ $X2=4.637 $Y2=0.86
r121 35 38 5.13969 $w=2.03e-07 $l=9.5e-08 $layer=LI1_cond $X=4.637 $Y=0.765
+ $X2=4.637 $Y2=0.86
r122 33 35 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=4.535 $Y=0.68
+ $X2=4.637 $Y2=0.765
r123 33 34 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.535 $Y=0.68
+ $X2=3.825 $Y2=0.68
r124 32 45 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.74 $Y=1.435 $X2=3.74
+ $Y2=1.585
r125 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.74 $Y=0.765
+ $X2=3.825 $Y2=0.68
r126 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.74 $Y=0.765
+ $X2=3.74 $Y2=1.435
r127 27 53 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.695 $Y=0.945
+ $X2=3.695 $Y2=1.405
r128 24 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.295 $Y=1.675
+ $X2=3.205 $Y2=1.675
r129 23 49 16.5998 $w=3.65e-07 $l=1.05e-07 $layer=POLY_cond $X=3.802 $Y=1.675
+ $X2=3.802 $Y2=1.57
r130 23 24 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.62 $Y=1.675
+ $X2=3.295 $Y2=1.675
r131 19 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.205 $Y=1.75
+ $X2=3.205 $Y2=1.675
r132 19 21 219.621 $w=1.8e-07 $l=5.65e-07 $layer=POLY_cond $X=3.205 $Y=1.75
+ $X2=3.205 $Y2=2.315
r133 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.675
+ $X2=2.505 $Y2=1.675
r134 17 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.115 $Y=1.675
+ $X2=3.205 $Y2=1.675
r135 17 18 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.115 $Y=1.675
+ $X2=2.58 $Y2=1.675
r136 13 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=1.6
+ $X2=2.505 $Y2=1.675
r137 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.505 $Y=1.6
+ $X2=2.505 $Y2=1.02
r138 11 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.43 $Y=1.675
+ $X2=2.505 $Y2=1.675
r139 11 12 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.43 $Y=1.675
+ $X2=2.165 $Y2=1.675
r140 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.075 $Y=1.75
+ $X2=2.165 $Y2=1.675
r141 7 9 206.016 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=2.075 $Y=1.75
+ $X2=2.075 $Y2=2.28
r142 2 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.84 $X2=4.62 $Y2=2.815
r143 2 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.84 $X2=4.62 $Y2=1.985
r144 1 38 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.37 $X2=4.655 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%B 3 5 6 9 11 12 15 17 21 23 26 28 33 35 37 38
+ 39 40 41 44 47
c133 47 0 2.09006e-20 $X=5.075 $Y=1.385
c134 40 0 1.36386e-19 $X=4.345 $Y=1.475
c135 21 0 1.77022e-19 $X=3.105 $Y=0.91
c136 9 0 1.59849e-19 $X=2.005 $Y=0.91
r137 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.075
+ $Y=1.385 $X2=5.075 $Y2=1.385
r138 45 47 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.87 $Y=1.385
+ $X2=5.075 $Y2=1.385
r139 43 45 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=4.845 $Y=1.385
+ $X2=4.87 $Y2=1.385
r140 43 44 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.845 $Y=1.385
+ $X2=4.755 $Y2=1.385
r141 41 48 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.075 $Y=1.295
+ $X2=5.075 $Y2=1.385
r142 35 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=1.22
+ $X2=4.87 $Y2=1.385
r143 35 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.87 $Y=1.22
+ $X2=4.87 $Y2=0.74
r144 31 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.55
+ $X2=4.845 $Y2=1.385
r145 31 33 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.845 $Y=1.55
+ $X2=4.845 $Y2=2.4
r146 30 40 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=4.44 $Y=1.475
+ $X2=4.345 $Y2=1.475
r147 30 44 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.44 $Y=1.475
+ $X2=4.755 $Y2=1.475
r148 28 40 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.365 $Y=1.4
+ $X2=4.345 $Y2=1.475
r149 27 28 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=4.365 $Y=0.255
+ $X2=4.365 $Y2=1.4
r150 25 40 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.325 $Y=1.55
+ $X2=4.345 $Y2=1.475
r151 25 26 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=4.325 $Y=1.55
+ $X2=4.325 $Y2=3.075
r152 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=0.18
+ $X2=3.105 $Y2=0.18
r153 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.29 $Y=0.18
+ $X2=4.365 $Y2=0.255
r154 23 24 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=4.29 $Y=0.18
+ $X2=3.18 $Y2=0.18
r155 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=0.255
+ $X2=3.105 $Y2=0.18
r156 19 21 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.105 $Y=0.255
+ $X2=3.105 $Y2=0.91
r157 18 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.76 $Y=3.15 $X2=2.67
+ $Y2=3.15
r158 17 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.25 $Y=3.15
+ $X2=4.325 $Y2=3.075
r159 17 18 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=4.25 $Y=3.15
+ $X2=2.76 $Y2=3.15
r160 13 38 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=3.075
+ $X2=2.67 $Y2=3.15
r161 13 15 258.492 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=2.67 $Y=3.075
+ $X2=2.67 $Y2=2.41
r162 11 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.03 $Y=0.18
+ $X2=3.105 $Y2=0.18
r163 11 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.03 $Y=0.18
+ $X2=2.08 $Y2=0.18
r164 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.08 $Y2=0.18
r165 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.005 $Y2=0.91
r166 5 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.58 $Y=3.15 $X2=2.67
+ $Y2=3.15
r167 5 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.58 $Y=3.15 $X2=1.63
+ $Y2=3.15
r168 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.54 $Y=3.075
+ $X2=1.63 $Y2=3.15
r169 1 3 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=1.54 $Y=3.075
+ $X2=1.54 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_1155_284# 1 2 9 13 16 17 18 20 25 27 30 31
+ 36
c91 36 0 6.08064e-20 $X=7.985 $Y=0.58
r92 33 36 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=7.665 $Y=0.58
+ $X2=7.985 $Y2=0.58
r93 30 32 11.2061 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=7.54 $Y=2.455
+ $X2=7.54 $Y2=2.71
r94 30 31 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=2.455
+ $X2=7.54 $Y2=2.29
r95 25 40 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.585
+ $X2=5.97 $Y2=1.75
r96 25 39 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.585
+ $X2=5.97 $Y2=1.42
r97 24 27 4.37134 $w=2.88e-07 $l=1.1e-07 $layer=LI1_cond $X=5.94 $Y=1.605
+ $X2=6.05 $Y2=1.605
r98 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.94
+ $Y=1.585 $X2=5.94 $Y2=1.585
r99 21 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0.745
+ $X2=7.665 $Y2=0.58
r100 21 31 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=7.665 $Y=0.745
+ $X2=7.665 $Y2=2.29
r101 20 32 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.415 $Y=2.905
+ $X2=7.415 $Y2=2.71
r102 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.33 $Y=2.99
+ $X2=7.415 $Y2=2.905
r103 17 18 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=7.33 $Y=2.99
+ $X2=6.135 $Y2=2.99
r104 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.05 $Y=2.905
+ $X2=6.135 $Y2=2.99
r105 15 27 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.05 $Y=1.75
+ $X2=6.05 $Y2=1.605
r106 15 16 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=6.05 $Y=1.75
+ $X2=6.05 $Y2=2.905
r107 13 39 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.09 $Y=0.935
+ $X2=6.09 $Y2=1.42
r108 9 40 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.015 $Y=2.36
+ $X2=6.015 $Y2=1.75
r109 2 30 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=7.35
+ $Y=2.05 $X2=7.495 $Y2=2.455
r110 1 36 182 $w=1.7e-07 $l=4.58121e-07 $layer=licon1_NDIFF $count=1 $X=7.62
+ $Y=0.37 $X2=7.985 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%C 3 7 10 11 12 13 15 17 18 20 22 23 24 25
c80 24 0 1.82049e-20 $X=7.28 $Y=1.712
c81 22 0 8.51369e-20 $X=6.725 $Y=1.615
r82 25 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.94
+ $Y=1.615 $X2=6.94 $Y2=1.615
r83 23 28 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=7.205 $Y=1.615
+ $X2=6.94 $Y2=1.615
r84 23 24 13.5877 $w=2.4e-07 $l=1.29167e-07 $layer=POLY_cond $X=7.205 $Y=1.615
+ $X2=7.28 $Y2=1.712
r85 21 28 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.845 $Y=1.615
+ $X2=6.94 $Y2=1.615
r86 21 22 3.90195 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=6.845 $Y=1.615
+ $X2=6.725 $Y2=1.615
r87 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.2 $Y=0.865 $X2=8.2
+ $Y2=0.58
r88 15 17 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.72 $Y=1.975
+ $X2=7.72 $Y2=2.37
r89 14 24 13.5877 $w=2.4e-07 $l=2.2236e-07 $layer=POLY_cond $X=7.355 $Y=1.9
+ $X2=7.28 $Y2=1.712
r90 13 15 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.63 $Y=1.9
+ $X2=7.72 $Y2=1.975
r91 13 14 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.63 $Y=1.9
+ $X2=7.355 $Y2=1.9
r92 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.125 $Y=0.94
+ $X2=8.2 $Y2=0.865
r93 11 12 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=8.125 $Y=0.94
+ $X2=7.355 $Y2=0.94
r94 10 24 12.1617 $w=1.5e-07 $l=2.62e-07 $layer=POLY_cond $X=7.28 $Y=1.45
+ $X2=7.28 $Y2=1.712
r95 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.28 $Y=1.015
+ $X2=7.355 $Y2=0.94
r96 9 10 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.28 $Y=1.015
+ $X2=7.28 $Y2=1.45
r97 5 22 34.7346 $w=1.65e-07 $l=1.86145e-07 $layer=POLY_cond $X=6.77 $Y=1.45
+ $X2=6.725 $Y2=1.615
r98 5 7 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.77 $Y=1.45 $X2=6.77
+ $Y2=0.935
r99 1 22 34.7346 $w=1.65e-07 $l=1.79374e-07 $layer=POLY_cond $X=6.695 $Y=1.78
+ $X2=6.725 $Y2=1.615
r100 1 3 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.695 $Y=1.78
+ $X2=6.695 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_1221_388# 1 2 9 13 17 21 25 29 33 37 43 45
+ 53 56 57 60 63 64 66 77
c144 66 0 6.08064e-20 $X=8.535 $Y=1.42
c145 60 0 1.82049e-20 $X=6.48 $Y=2.035
c146 57 0 1.54548e-19 $X=6.625 $Y=2.035
r147 76 77 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=10.055 $Y=1.42
+ $X2=10.07 $Y2=1.42
r148 75 76 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=9.64 $Y=1.42
+ $X2=10.055 $Y2=1.42
r149 74 75 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.605 $Y=1.42
+ $X2=9.64 $Y2=1.42
r150 73 74 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=9.21 $Y=1.42
+ $X2=9.605 $Y2=1.42
r151 72 73 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=9.075 $Y=1.42
+ $X2=9.21 $Y2=1.42
r152 71 72 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=8.78 $Y=1.42
+ $X2=9.075 $Y2=1.42
r153 66 69 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.535 $Y=1.42
+ $X2=8.625 $Y2=1.42
r154 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r155 60 82 6.74607 $w=3.33e-07 $l=1.15e-07 $layer=LI1_cond $X=6.472 $Y=2.035
+ $X2=6.472 $Y2=1.92
r156 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=2.035
+ $X2=6.48 $Y2=2.035
r157 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=2.035
+ $X2=6.48 $Y2=2.035
r158 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r159 56 57 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=6.625 $Y2=2.035
r160 54 71 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=8.695 $Y=1.42
+ $X2=8.78 $Y2=1.42
r161 54 69 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.695 $Y=1.42
+ $X2=8.625 $Y2=1.42
r162 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.695
+ $Y=1.42 $X2=8.695 $Y2=1.42
r163 51 64 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.4 $Y=1.585
+ $X2=8.4 $Y2=2.035
r164 50 53 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.4 $Y=1.42
+ $X2=8.695 $Y2=1.42
r165 50 51 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.4 $Y=1.42 $X2=8.4
+ $Y2=1.585
r166 48 66 90.9279 $w=3.3e-07 $l=5.2e-07 $layer=POLY_cond $X=8.015 $Y=1.42
+ $X2=8.535 $Y2=1.42
r167 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.015
+ $Y=1.42 $X2=8.015 $Y2=1.42
r168 45 50 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.285 $Y=1.42
+ $X2=8.4 $Y2=1.42
r169 45 47 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.285 $Y=1.42
+ $X2=8.015 $Y2=1.42
r170 43 82 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.555 $Y=1.105
+ $X2=6.555 $Y2=1.92
r171 35 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.07 $Y=1.255
+ $X2=10.07 $Y2=1.42
r172 35 37 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=10.07 $Y=1.255
+ $X2=10.07 $Y2=0.74
r173 31 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.055 $Y=1.585
+ $X2=10.055 $Y2=1.42
r174 31 33 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=10.055 $Y=1.585
+ $X2=10.055 $Y2=2.4
r175 27 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.64 $Y=1.255
+ $X2=9.64 $Y2=1.42
r176 27 29 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=9.64 $Y=1.255
+ $X2=9.64 $Y2=0.74
r177 23 74 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.585
+ $X2=9.605 $Y2=1.42
r178 23 25 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=9.605 $Y=1.585
+ $X2=9.605 $Y2=2.4
r179 19 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=1.255
+ $X2=9.21 $Y2=1.42
r180 19 21 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=9.21 $Y=1.255
+ $X2=9.21 $Y2=0.74
r181 15 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.075 $Y=1.585
+ $X2=9.075 $Y2=1.42
r182 15 17 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=9.075 $Y=1.585
+ $X2=9.075 $Y2=2.4
r183 11 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.78 $Y=1.255
+ $X2=8.78 $Y2=1.42
r184 11 13 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=8.78 $Y=1.255
+ $X2=8.78 $Y2=0.74
r185 7 69 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.585
+ $X2=8.625 $Y2=1.42
r186 7 9 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=8.625 $Y=1.585
+ $X2=8.625 $Y2=2.4
r187 2 60 300 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.94 $X2=6.47 $Y2=2.085
r188 1 43 182 $w=1.7e-07 $l=6.56658e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.615 $X2=6.555 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_27_118# 1 2 3 4 13 14 17 19 21 24 27 29 31
+ 35 36
c84 35 0 5.90733e-20 $X=0.265 $Y=1.25
c85 29 0 1.18804e-19 $X=2.68 $Y=1.42
c86 13 0 4.31925e-20 $X=0.265 $Y=0.75
r87 35 36 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.17 $Y=1.25
+ $X2=0.17 $Y2=2.18
r88 29 31 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=2.68 $Y=1.42 $X2=2.68
+ $Y2=1.02
r89 25 29 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.26 $Y=1.505
+ $X2=2.68 $Y2=1.505
r90 25 37 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=1.505
+ $X2=1.88 $Y2=1.505
r91 25 27 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=2.26 $Y=1.59
+ $X2=2.26 $Y2=2.21
r92 24 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=1.42
+ $X2=1.88 $Y2=1.505
r93 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.88 $Y=0.75
+ $X2=1.88 $Y2=1.42
r94 22 34 5.39736 $w=1.7e-07 $l=1.82483e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=0.265 $Y2=0.66
r95 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=0.665
+ $X2=1.88 $Y2=0.75
r96 21 22 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=1.795 $Y=0.665
+ $X2=0.445 $Y2=0.665
r97 17 36 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=2.32
+ $X2=0.225 $Y2=2.18
r98 17 19 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.225 $Y=2.32
+ $X2=0.225 $Y2=2.345
r99 14 35 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1.07
+ $X2=0.265 $Y2=1.25
r100 13 34 2.62574 $w=3.6e-07 $l=9e-08 $layer=LI1_cond $X=0.265 $Y=0.75
+ $X2=0.265 $Y2=0.66
r101 13 14 10.2439 $w=3.58e-07 $l=3.2e-07 $layer=LI1_cond $X=0.265 $Y=0.75
+ $X2=0.265 $Y2=1.07
r102 4 27 600 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.96 $X2=2.3 $Y2=2.21
r103 3 19 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.345
r104 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.81 $X2=2.72 $Y2=1.02
r105 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.59 $X2=0.28 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%VPWR 1 2 3 4 5 18 22 28 31 32 36 40 42 47 49
+ 51 56 64 72 78 81 84 87 91
r114 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r115 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r117 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r118 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 76 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r121 76 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r122 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r123 73 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.38 $Y2=3.33
r124 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.84 $Y2=3.33
r125 72 90 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.377 $Y2=3.33
r126 72 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=9.84 $Y2=3.33
r127 71 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r129 68 71 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r130 67 70 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r132 65 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=3.33
+ $X2=5.07 $Y2=3.33
r133 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.235 $Y=3.33
+ $X2=5.52 $Y2=3.33
r134 64 84 12.0118 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=7.945 $Y=3.33
+ $X2=8.222 $Y2=3.33
r135 64 70 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.945 $Y=3.33
+ $X2=7.92 $Y2=3.33
r136 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r137 62 63 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 60 63 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 59 62 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 59 60 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r143 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 56 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.07 $Y2=3.33
r145 56 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r149 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r150 49 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r151 49 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r152 47 48 9.86413 $w=5.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.222 $Y=2.495
+ $X2=8.222 $Y2=2.33
r153 42 45 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.32 $Y=1.985
+ $X2=10.32 $Y2=2.815
r154 40 90 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.377 $Y2=3.33
r155 40 45 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.32 $Y2=2.815
r156 36 39 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.38 $Y=1.985
+ $X2=9.38 $Y2=2.815
r157 34 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=3.33
r158 34 39 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=2.815
r159 33 84 12.0118 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=8.5 $Y=3.33
+ $X2=8.222 $Y2=3.33
r160 32 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=9.38 $Y2=3.33
r161 32 33 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=8.5 $Y2=3.33
r162 31 84 2.33542 $w=5.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.222 $Y=3.245
+ $X2=8.222 $Y2=3.33
r163 30 47 2.41371 $w=5.53e-07 $l=1.12e-07 $layer=LI1_cond $X=8.222 $Y=2.607
+ $X2=8.222 $Y2=2.495
r164 30 31 13.7495 $w=5.53e-07 $l=6.38e-07 $layer=LI1_cond $X=8.222 $Y=2.607
+ $X2=8.222 $Y2=3.245
r165 28 48 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.03 $Y=1.985
+ $X2=8.03 $Y2=2.33
r166 22 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.07 $Y=1.985
+ $X2=5.07 $Y2=2.815
r167 20 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=3.33
r168 20 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=2.815
r169 16 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r170 16 18 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.345
r171 5 45 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.145
+ $Y=1.84 $X2=10.28 $Y2=2.815
r172 5 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.145
+ $Y=1.84 $X2=10.28 $Y2=1.985
r173 4 39 400 $w=1.7e-07 $l=1.07715e-06 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.84 $X2=9.38 $Y2=2.815
r174 4 36 400 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.84 $X2=9.38 $Y2=1.985
r175 3 47 200 $w=1.7e-07 $l=7.81441e-07 $layer=licon1_PDIFF $count=3 $X=7.81
+ $Y=2.05 $X2=8.4 $Y2=2.495
r176 3 28 300 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=2 $X=7.81
+ $Y=2.05 $X2=8.03 $Y2=1.985
r177 2 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.84 $X2=5.07 $Y2=2.815
r178 2 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.84 $X2=5.07 $Y2=1.985
r179 1 18 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_326_392# 1 2 3 4 13 15 17 22 23 24 26 27 28
+ 32 33 34 38 42 44
c121 38 0 1.54548e-19 $X=7.325 $Y=1.95
c122 13 0 1.12299e-19 $X=1.765 $Y=2.565
r123 42 44 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.92 $Y=2.035
+ $X2=7.325 $Y2=2.035
r124 38 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=1.95
+ $X2=7.325 $Y2=2.035
r125 37 38 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=7.325 $Y=0.425
+ $X2=7.325 $Y2=1.95
r126 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.24 $Y=0.34
+ $X2=7.325 $Y2=0.425
r127 33 34 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=7.24 $Y=0.34
+ $X2=5.96 $Y2=0.34
r128 30 32 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=5.835 $Y=0.78
+ $X2=5.835 $Y2=0.77
r129 29 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.835 $Y=0.425
+ $X2=5.96 $Y2=0.34
r130 29 32 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.835 $Y=0.425
+ $X2=5.835 $Y2=0.77
r131 27 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.71 $Y=0.865
+ $X2=5.835 $Y2=0.78
r132 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.71 $Y=0.865
+ $X2=5.08 $Y2=0.865
r133 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.995 $Y=0.78
+ $X2=5.08 $Y2=0.865
r134 25 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.995 $Y=0.425
+ $X2=4.995 $Y2=0.78
r135 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.91 $Y=0.34
+ $X2=4.995 $Y2=0.425
r136 23 24 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=4.91 $Y=0.34
+ $X2=3.485 $Y2=0.34
r137 20 22 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=3.4 $Y=2.565
+ $X2=3.4 $Y2=0.735
r138 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.4 $Y=0.425
+ $X2=3.485 $Y2=0.34
r139 19 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.4 $Y=0.425
+ $X2=3.4 $Y2=0.735
r140 18 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=2.65
+ $X2=1.765 $Y2=2.65
r141 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.315 $Y=2.65
+ $X2=3.4 $Y2=2.565
r142 17 18 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=3.315 $Y=2.65
+ $X2=1.93 $Y2=2.65
r143 13 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=2.565
+ $X2=1.765 $Y2=2.65
r144 13 15 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.765 $Y=2.565
+ $X2=1.765 $Y2=2.265
r145 4 42 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.785
+ $Y=1.94 $X2=6.92 $Y2=2.115
r146 3 40 600 $w=1.7e-07 $l=7.54487e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.96 $X2=1.765 $Y2=2.65
r147 3 15 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.96 $X2=1.765 $Y2=2.265
r148 2 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.74
+ $Y=0.615 $X2=5.875 $Y2=0.77
r149 1 22 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=3.18
+ $Y=0.59 $X2=3.4 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%A_416_118# 1 2 3 4 15 19 20 22 27 28 30 31 32
+ 36 37 38 44 45 51 54
c123 51 0 3.34966e-20 $X=3.06 $Y=2.135
c124 37 0 2.8323e-19 $X=5.375 $Y=2.035
c125 31 0 8.51369e-20 $X=6.82 $Y=0.68
c126 15 0 1.59849e-19 $X=2.22 $Y=0.735
r127 50 51 1.84012 $w=5.18e-07 $l=8e-08 $layer=LI1_cond $X=2.98 $Y=2.135
+ $X2=3.06 $Y2=2.135
r128 45 54 7.13013 $w=3.88e-07 $l=1.15e-07 $layer=LI1_cond $X=5.6 $Y=2.035
+ $X2=5.6 $Y2=1.92
r129 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r130 41 50 7.82051 $w=5.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.64 $Y=2.135
+ $X2=2.98 $Y2=2.135
r131 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=2.035
+ $X2=2.64 $Y2=2.035
r132 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=2.035
+ $X2=2.64 $Y2=2.035
r133 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r134 37 38 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=2.785 $Y2=2.035
r135 31 36 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.82 $Y=0.68
+ $X2=6.945 $Y2=0.68
r136 31 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.82 $Y=0.68
+ $X2=6.3 $Y2=0.68
r137 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.215 $Y=0.765
+ $X2=6.3 $Y2=0.68
r138 29 30 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.215 $Y=0.765
+ $X2=6.215 $Y2=1.12
r139 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.13 $Y=1.205
+ $X2=6.215 $Y2=1.12
r140 27 28 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.13 $Y=1.205
+ $X2=5.605 $Y2=1.205
r141 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.52 $Y=1.29
+ $X2=5.605 $Y2=1.205
r142 25 54 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.52 $Y=1.29
+ $X2=5.52 $Y2=1.92
r143 22 51 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.06 $Y=1.875
+ $X2=3.06 $Y2=2.135
r144 21 22 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=3.06 $Y=0.62
+ $X2=3.06 $Y2=1.875
r145 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.975 $Y=0.535
+ $X2=3.06 $Y2=0.62
r146 19 20 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.975 $Y=0.535
+ $X2=2.385 $Y2=0.535
r147 15 17 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=2.26 $Y=0.735
+ $X2=2.26 $Y2=1.085
r148 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.26 $Y=0.62
+ $X2=2.385 $Y2=0.535
r149 13 15 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.26 $Y=0.62
+ $X2=2.26 $Y2=0.735
r150 4 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.485
+ $Y=1.94 $X2=5.63 $Y2=2.085
r151 3 50 600 $w=1.7e-07 $l=2.73496e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.09 $X2=2.98 $Y2=2.21
r152 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.615 $X2=6.985 $Y2=0.76
r153 1 17 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.59 $X2=2.22 $Y2=1.085
r154 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.59 $X2=2.22 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%X 1 2 3 4 15 19 22 25 29 32 33 34 35 36 37 38
+ 39 45 59
r65 45 59 2.00531 $w=3.3e-07 $l=5e-08 $layer=LI1_cond $X=9.83 $Y=1.715 $X2=9.83
+ $Y2=1.665
r66 38 39 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.83 $Y=2.405
+ $X2=9.83 $Y2=2.775
r67 37 38 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.83 $Y=1.985
+ $X2=9.83 $Y2=2.405
r68 36 59 0.741892 $w=2.96e-07 $l=1.8e-08 $layer=LI1_cond $X=9.83 $Y=1.647
+ $X2=9.83 $Y2=1.665
r69 36 56 10.7986 $w=2.96e-07 $l=2.62e-07 $layer=LI1_cond $X=9.83 $Y=1.647
+ $X2=9.83 $Y2=1.385
r70 36 37 8.8354 $w=3.28e-07 $l=2.53e-07 $layer=LI1_cond $X=9.83 $Y=1.732
+ $X2=9.83 $Y2=1.985
r71 36 45 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=9.83 $Y=1.732
+ $X2=9.83 $Y2=1.715
r72 32 33 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.905 $Y=1.985
+ $X2=8.905 $Y2=1.82
r73 27 56 3.83342 $w=2.96e-07 $l=9.21954e-08 $layer=LI1_cond $X=9.815 $Y=1.3
+ $X2=9.83 $Y2=1.385
r74 27 29 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=9.815 $Y=1.3
+ $X2=9.815 $Y2=0.515
r75 26 35 1.69765 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=9.16 $Y=1.385
+ $X2=9.057 $Y2=1.385
r76 25 56 3.98214 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=1.385
+ $X2=9.83 $Y2=1.385
r77 25 26 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=9.665 $Y=1.385
+ $X2=9.16 $Y2=1.385
r78 23 35 4.7579 $w=1.87e-07 $l=9.31128e-08 $layer=LI1_cond $X=9.04 $Y=1.47
+ $X2=9.057 $Y2=1.385
r79 23 33 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.04 $Y=1.47
+ $X2=9.04 $Y2=1.82
r80 22 35 4.7579 $w=1.87e-07 $l=8.5e-08 $layer=LI1_cond $X=9.057 $Y=1.3
+ $X2=9.057 $Y2=1.385
r81 22 34 11.6319 $w=2.03e-07 $l=2.15e-07 $layer=LI1_cond $X=9.057 $Y=1.3
+ $X2=9.057 $Y2=1.085
r82 17 34 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.995 $Y=0.92
+ $X2=8.995 $Y2=1.085
r83 17 19 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=8.995 $Y=0.92
+ $X2=8.995 $Y2=0.515
r84 13 32 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=8.905 $Y=2.04
+ $X2=8.905 $Y2=1.985
r85 13 15 20.2987 $w=4.38e-07 $l=7.75e-07 $layer=LI1_cond $X=8.905 $Y=2.04
+ $X2=8.905 $Y2=2.815
r86 4 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.695
+ $Y=1.84 $X2=9.83 $Y2=2.815
r87 4 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.695
+ $Y=1.84 $X2=9.83 $Y2=1.985
r88 3 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.85 $Y2=1.985
r89 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.85 $Y2=2.815
r90 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.715
+ $Y=0.37 $X2=9.855 $Y2=0.515
r91 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.855
+ $Y=0.37 $X2=8.995 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_4%VGND 1 2 3 4 5 18 22 24 28 30 32 35 36 37 39
+ 51 55 62 68 71 75
r89 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0 $X2=10.32
+ $Y2=0
r90 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r91 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r92 68 69 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r93 62 65 9.13522 $w=4.08e-07 $l=3.25e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.83
+ $Y2=0.325
r94 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 59 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.32
+ $Y2=0
r96 59 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r97 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r98 56 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.51 $Y=0 $X2=9.425
+ $Y2=0
r99 56 58 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.51 $Y=0 $X2=9.84
+ $Y2=0
r100 55 74 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=10.12 $Y=0 $X2=10.34
+ $Y2=0
r101 55 58 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.12 $Y=0 $X2=9.84
+ $Y2=0
r102 54 69 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=8.4
+ $Y2=0
r103 53 54 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r104 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.33 $Y=0 $X2=8.495
+ $Y2=0
r105 51 53 183.326 $w=1.68e-07 $l=2.81e-06 $layer=LI1_cond $X=8.33 $Y=0 $X2=5.52
+ $Y2=0
r106 49 50 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r107 47 50 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r108 47 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 46 49 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r110 46 47 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r111 44 62 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.83
+ $Y2=0
r112 44 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r113 42 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r114 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 39 62 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.83
+ $Y2=0
r116 39 41 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r117 37 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r118 37 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r119 35 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.04
+ $Y2=0
r120 35 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.375
+ $Y2=0
r121 34 53 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=5.5 $Y=0 $X2=5.52
+ $Y2=0
r122 34 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.5 $Y=0 $X2=5.375
+ $Y2=0
r123 30 74 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.34 $Y2=0
r124 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.515
r125 26 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.425 $Y=0.085
+ $X2=9.425 $Y2=0
r126 26 28 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.425 $Y=0.085
+ $X2=9.425 $Y2=0.515
r127 25 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.66 $Y=0 $X2=8.495
+ $Y2=0
r128 24 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=0 $X2=9.425
+ $Y2=0
r129 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.34 $Y=0 $X2=8.66
+ $Y2=0
r130 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.495 $Y=0.085
+ $X2=8.495 $Y2=0
r131 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.495 $Y=0.085
+ $X2=8.495 $Y2=0.515
r132 16 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0
r133 16 18 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0.445
r134 5 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.145
+ $Y=0.37 $X2=10.285 $Y2=0.515
r135 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.285
+ $Y=0.37 $X2=9.425 $Y2=0.515
r136 3 22 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=8.275
+ $Y=0.37 $X2=8.495 $Y2=0.515
r137 2 18 182 $w=1.7e-07 $l=4.25852e-07 $layer=licon1_NDIFF $count=1 $X=4.945
+ $Y=0.37 $X2=5.335 $Y2=0.445
r138 1 65 182 $w=1.7e-07 $l=3.72995e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.59 $X2=0.83 $Y2=0.325
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
M1000 a_856_294# a_714_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=7.5e+11p pd=3.5e+06u as=1.65038e+12p ps=1.553e+07u
M1001 a_1266_119# a_510_74# a_856_294# VPB pshort w=1e+06u l=180000u
+  ad=4.264e+11p pd=3.34e+06u as=0p ps=0u
M1002 VGND a_1598_93# a_1550_119# VNB nlowvt w=420000u l=150000u
+  ad=1.2824e+12p pd=1.089e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_510_74# a_300_347# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1004 a_1598_93# a_1266_119# a_1736_119# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1005 VPWR a_856_294# a_820_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_714_119# a_510_74# a_33_74# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=2.31e+11p ps=2.78e+06u
M1007 a_1266_119# a_300_347# a_856_294# VNB nlowvt w=740000u l=150000u
+  ad=6.134e+11p pd=4.02e+06u as=2.146e+11p ps=2.06e+06u
M1008 VPWR a_1598_93# a_1550_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1009 VGND RESET_B a_922_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 a_1736_119# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_74# a_300_347# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.257e+11p pd=2.09e+06u as=0p ps=0u
M1012 a_714_119# a_300_347# a_33_74# VPB pshort w=420000u l=180000u
+  ad=2.226e+11p pd=2.74e+06u as=2.31e+11p ps=2.78e+06u
M1013 VGND CLK_N a_300_347# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.442e+11p ps=2.14e+06u
M1014 a_820_457# a_510_74# a_714_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1598_93# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1016 a_922_119# a_856_294# a_850_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 VPWR CLK_N a_300_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9575e+11p ps=2.65e+06u
M1018 a_714_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_850_119# a_300_347# a_714_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_856_294# a_714_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1266_119# a_1934_94# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1022 a_1550_119# a_510_74# a_1266_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1266_119# a_1598_93# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND RESET_B a_120_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VPWR a_1266_119# a_1934_94# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1026 Q a_1934_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 Q a_1934_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=0p ps=0u
M1028 a_120_74# D a_33_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1550_508# a_300_347# a_1266_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_33_74# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR RESET_B a_33_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__sdfxtp_4.spice
* Created: Fri Aug 28 18:14:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfxtp_4.pex.spice"
.subckt sky130_fd_sc_ms__sdfxtp_4  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1036 N_VGND_M1036_d N_SCE_M1036_g N_A_36_74#_M1036_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1022 A_223_74# N_A_36_74#_M1022_g N_VGND_M1036_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_301_74#_M1023_d N_D_M1023_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.12705 AS=0.0504 PD=1.025 PS=0.66 NRD=45.708 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 A_452_74# N_SCE_M1011_g N_A_301_74#_M1023_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.12705 PD=0.66 PS=1.025 NRD=18.564 NRS=47.136 M=1 R=2.8
+ SA=75001.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_SCD_M1010_g A_452_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_630_74#_M1003_d N_CLK_M1003_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_A_828_74#_M1021_d N_A_630_74#_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_1026_100#_M1027_d N_A_630_74#_M1027_g N_A_301_74#_M1027_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1012 A_1162_100# N_A_828_74#_M1012_g N_A_1026_100#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.09975 AS=0.1113 PD=0.895 PS=0.95 NRD=52.14 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_1257_74#_M1034_g A_1162_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.179149 AS=0.09975 PD=1.14309 PS=0.895 NRD=24.276 NRS=52.14 M=1 R=2.8
+ SA=75001.5 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1035 N_A_1257_74#_M1035_d N_A_1026_100#_M1035_g N_VGND_M1034_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.11825 AS=0.234601 PD=0.98 PS=1.49691 NRD=13.08 NRS=89.448
+ M=1 R=3.66667 SA=75002 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1032 N_A_1587_74#_M1032_d N_A_828_74#_M1032_g N_A_1257_74#_M1035_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.226804 AS=0.11825 PD=1.46856 PS=0.98 NRD=84 NRS=19.632 M=1
+ R=3.66667 SA=75002.6 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1020 A_1766_74# N_A_630_74#_M1020_g N_A_1587_74#_M1032_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.173196 PD=0.66 PS=1.12144 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75003.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1814_48#_M1018_g A_1766_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_A_1587_74#_M1030_g N_A_1814_48#_M1030_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.12025 AS=0.2109 PD=1.065 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1030_d N_A_1814_48#_M1004_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.13505 PD=1.065 PS=1.105 NRD=7.296 NRS=13.776 M=1 R=4.93333
+ SA=75000.7 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_1814_48#_M1016_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.13505 PD=1.02 PS=1.105 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1016_d N_A_1814_48#_M1019_g N_Q_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1031_d N_A_1814_48#_M1031_g N_Q_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_SCE_M1015_g N_A_36_74#_M1015_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.1792 PD=0.96 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.8 A=0.1152 P=1.64 MULT=1
MM1013 A_241_464# N_SCE_M1013_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90002.3 A=0.1152 P=1.64 MULT=1
MM1026 N_A_301_74#_M1026_d N_D_M1026_g A_241_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.1
+ SB=90001.9 A=0.1152 P=1.64 MULT=1
MM1029 A_415_464# N_A_36_74#_M1029_g N_A_301_74#_M1026_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1152 AS=0.0864 PD=1 PS=0.91 NRD=38.4741 NRS=0 M=1 R=3.55556
+ SA=90001.6 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1000 N_VPWR_M1000_d N_SCD_M1000_g A_415_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.173964 AS=0.1152 PD=1.22182 PS=1 NRD=43.0839 NRS=38.4741 M=1 R=3.55556
+ SA=90002.1 SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1001 N_A_630_74#_M1001_d N_CLK_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.304436 PD=2.8 PS=2.13818 NRD=0 NRS=24.625 M=1 R=6.22222
+ SA=90001.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1025 N_A_828_74#_M1025_d N_A_630_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.6048 PD=2.8 PS=3.32 NRD=0 NRS=21.9852 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1002 N_A_1026_100#_M1002_d N_A_828_74#_M1002_g N_A_301_74#_M1002_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90005.3 A=0.0756 P=1.2 MULT=1
MM1006 A_1217_506# N_A_630_74#_M1006_g N_A_1026_100#_M1002_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0756 AS=0.0567 PD=0.78 PS=0.69 NRD=58.6272 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90004.8 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_A_1257_74#_M1009_g A_1217_506# VPB PSHORT L=0.18 W=0.42
+ AD=0.117092 AS=0.0756 PD=0.993333 PS=0.78 NRD=39.8531 NRS=58.6272 M=1
+ R=2.33333 SA=90001.2 SB=90004.3 A=0.0756 P=1.2 MULT=1
MM1037 N_A_1257_74#_M1037_d N_A_1026_100#_M1037_g N_VPWR_M1009_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.3654 AS=0.234183 PD=1.71 PS=1.98667 NRD=5.2599 NRS=52.4808
+ M=1 R=4.66667 SA=90001 SB=90003.1 A=0.1512 P=2.04 MULT=1
MM1033 N_A_1587_74#_M1033_d N_A_630_74#_M1033_g N_A_1257_74#_M1037_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1806 AS=0.3654 PD=1.6 PS=1.71 NRD=0 NRS=114.91 M=1
+ R=4.66667 SA=90002 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1038 A_1767_476# N_A_828_74#_M1038_g N_A_1587_74#_M1033_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0903 PD=0.66 PS=0.8 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90002.8 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_1814_48#_M1007_g A_1767_476# VPB PSHORT L=0.18 W=0.42
+ AD=0.0805 AS=0.0504 PD=0.776667 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333
+ SA=90003.2 SB=90003 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1007_d N_A_1587_74#_M1008_g N_A_1814_48#_M1008_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.161 AS=0.1134 PD=1.55333 PS=1.11 NRD=11.7215 NRS=0 M=1
+ R=4.66667 SA=90001.9 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1028 N_VPWR_M1028_d N_A_1587_74#_M1028_g N_A_1814_48#_M1008_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.1134 PD=1.23857 PS=1.11 NRD=9.3772 NRS=0 M=1
+ R=4.66667 SA=90002.4 SB=90002 A=0.1512 P=2.04 MULT=1
MM1005 N_Q_M1005_d N_A_1814_48#_M1005_g N_VPWR_M1028_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196 PD=1.39 PS=1.65143 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90002.2 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1014 N_Q_M1005_d N_A_1814_48#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.7
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1017 N_Q_M1017_d N_A_1814_48#_M1017_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1024 N_Q_M1017_d N_A_1814_48#_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX39_noxref VNB VPB NWDIODE A=23.9196 P=29.44
c_145 VNB 0 1.73925e-19 $X=0 $Y=0
c_248 VPB 0 2.97017e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__sdfxtp_4.pxi.spice"
*
.ends
*
*

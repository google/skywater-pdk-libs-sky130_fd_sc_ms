* File: sky130_fd_sc_ms__o22a_1.pex.spice
* Created: Fri Aug 28 17:57:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O22A_1%A_83_260# 1 2 9 13 16 17 22 25 27 31 35 36 41
c77 36 0 1.80886e-19 $X=2.26 $Y=1.202
c78 31 0 4.2886e-20 $X=0.93 $Y=1.465
c79 22 0 1.51466e-19 $X=2.26 $Y=1.97
r80 38 41 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.26 $Y=2.055 $X2=2.56
+ $Y2=2.055
r81 34 36 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.09 $Y=1.202 $X2=2.26
+ $Y2=1.202
r82 34 35 10.7338 $w=1.93e-07 $l=1.85e-07 $layer=LI1_cond $X=2.09 $Y=1.202
+ $X2=1.905 $Y2=1.202
r83 25 41 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.56 $Y=2.815
+ $X2=2.56 $Y2=2.14
r84 22 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=1.97
+ $X2=2.26 $Y2=2.055
r85 21 36 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=2.26 $Y=1.3 $X2=2.26
+ $Y2=1.202
r86 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.26 $Y=1.3 $X2=2.26
+ $Y2=1.97
r87 20 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=1.215
+ $X2=1.01 $Y2=1.215
r88 20 35 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.095 $Y=1.215
+ $X2=1.905 $Y2=1.215
r89 17 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.465 $X2=0.93 $Y2=1.465
r90 17 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.01 $Y=1.465
+ $X2=1.01 $Y2=1.215
r91 15 31 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=0.595 $Y=1.465
+ $X2=0.93 $Y2=1.465
r92 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.465
+ $X2=0.505 $Y2=1.465
r93 11 16 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.505 $Y2=1.465
r94 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
r95 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r96 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
r97 2 41 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.96 $X2=2.56 $Y2=2.135
r98 2 25 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.96 $X2=2.56 $Y2=2.815
r99 1 34 182 $w=1.7e-07 $l=5.69408e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.695 $X2=2.09 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%B1 5 9 11 14 15
r37 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.84
+ $Y=1.635 $X2=1.84 $Y2=1.635
r38 11 15 0.535558 $w=6.68e-07 $l=3e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.635
r39 7 14 34.7346 $w=1.65e-07 $l=1.76125e-07 $layer=POLY_cond $X=1.915 $Y=1.8
+ $X2=1.892 $Y2=1.635
r40 7 9 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.915 $Y=1.8 $X2=1.915
+ $Y2=2.46
r41 3 14 34.7346 $w=1.65e-07 $l=1.82565e-07 $layer=POLY_cond $X=1.855 $Y=1.47
+ $X2=1.892 $Y2=1.635
r42 3 5 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.855 $Y=1.47
+ $X2=1.855 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%B2 1 3 8 12 13 15 23
c46 23 0 4.2886e-20 $X=1.305 $Y=0.462
c47 12 0 6.69395e-20 $X=2.305 $Y=0.42
r48 15 23 3.43205 $w=4.13e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=0.462
+ $X2=1.305 $Y2=0.462
r49 13 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.42
+ $X2=2.305 $Y2=0.585
r50 12 23 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=2.305 $Y=0.42
+ $X2=1.305 $Y2=0.42
r51 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=0.42 $X2=2.305 $Y2=0.42
r52 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.325 $Y=1.015
+ $X2=2.325 $Y2=1.41
r53 8 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.325 $Y=1.015
+ $X2=2.325 $Y2=0.585
r54 1 9 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.5 $X2=2.335
+ $Y2=1.41
r55 1 3 373.161 $w=1.8e-07 $l=9.6e-07 $layer=POLY_cond $X=2.335 $Y=1.5 $X2=2.335
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%A2 3 7 9 12 13
c40 3 0 2.47825e-19 $X=2.755 $Y=1.015
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.635
+ $X2=2.83 $Y2=1.8
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.635
+ $X2=2.83 $Y2=1.47
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.635 $X2=2.83 $Y2=1.635
r44 9 13 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.635
+ $X2=2.83 $Y2=1.635
r45 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.785 $Y=2.46
+ $X2=2.785 $Y2=1.8
r46 3 14 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.755 $Y=1.015
+ $X2=2.755 $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%A1 3 7 9 12
r27 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.635
+ $X2=3.4 $Y2=1.8
r28 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.635
+ $X2=3.4 $Y2=1.47
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.635 $X2=3.4 $Y2=1.635
r30 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.635 $X2=3.4
+ $Y2=1.635
r31 7 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.345 $Y=0.97 $X2=3.345
+ $Y2=1.47
r32 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.325 $Y=2.46
+ $X2=3.325 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%X 1 2 9 13 14 15 16 23 32
r20 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=2.035
r21 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=2.405
+ $X2=0.265 $Y2=2.775
r22 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=2
r23 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=1.82
r24 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.405
r25 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.035
r26 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r27 7 13 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=0.99
+ $X2=0.225 $Y2=1.13
r28 7 9 19.5504 $w=2.78e-07 $l=4.75e-07 $layer=LI1_cond $X=0.225 $Y=0.99
+ $X2=0.225 $Y2=0.515
r29 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r30 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r31 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%VPWR 1 2 9 16 18 22 24 29 38 44
r39 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 39 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 38 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 36 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r47 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 30 38 17.8809 $w=1.7e-07 $l=6.18e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.232 $Y2=3.33
r49 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 29 43 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.612 $Y2=3.33
r51 29 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 24 38 17.8809 $w=1.7e-07 $l=6.17e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.232 $Y2=3.33
r55 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 22 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.55 $Y=2.135
+ $X2=3.55 $Y2=2.815
r59 16 43 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.612 $Y2=3.33
r60 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=2.815
r61 12 15 3.3587 $w=1.233e-06 $l=3.4e-07 $layer=LI1_cond $X=1.232 $Y=2.49
+ $X2=1.232 $Y2=2.83
r62 9 12 3.3587 $w=1.233e-06 $l=3.4e-07 $layer=LI1_cond $X=1.232 $Y=2.15
+ $X2=1.232 $Y2=2.49
r63 7 38 3.84952 $w=1.235e-06 $l=8.5e-08 $layer=LI1_cond $X=1.232 $Y=3.245
+ $X2=1.232 $Y2=3.33
r64 7 15 4.0996 $w=1.233e-06 $l=4.15e-07 $layer=LI1_cond $X=1.232 $Y=3.245
+ $X2=1.232 $Y2=2.83
r65 2 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.96 $X2=3.55 $Y2=2.815
r66 2 18 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.96 $X2=3.55 $Y2=2.135
r67 1 15 266.667 $w=1.7e-07 $l=1.27031e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=1.235 $Y2=2.83
r68 1 12 266.667 $w=1.7e-07 $l=1.37717e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=1.685 $Y2=2.49
r69 1 12 266.667 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.735 $Y2=2.49
r70 1 9 266.667 $w=1.7e-07 $l=7.79744e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=1.235 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r40 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 30 39 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.055
+ $Y2=0
r45 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.6
+ $Y2=0
r46 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r50 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r52 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r53 22 39 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.055
+ $Y2=0
r54 22 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.64
+ $Y2=0
r55 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r58 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r59 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r61 11 39 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r62 11 13 24.0657 $w=3.38e-07 $l=7.1e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.795
r63 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r64 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.515
r65 2 13 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.695 $X2=3.055 $Y2=0.795
r66 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O22A_1%A_299_139# 1 2 3 10 14 15 16 17 20
r39 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.56 $Y=1.13
+ $X2=3.56 $Y2=0.795
r40 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=1.215
+ $X2=3.56 $Y2=1.13
r41 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.395 $Y=1.215
+ $X2=2.705 $Y2=1.215
r42 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.62 $Y=1.13
+ $X2=2.705 $Y2=1.215
r43 14 23 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.62 $Y=0.935 $X2=2.62
+ $Y2=0.845
r44 14 15 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.62 $Y=0.935
+ $X2=2.62 $Y2=1.13
r45 10 23 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.845
+ $X2=2.62 $Y2=0.845
r46 10 12 55.1465 $w=1.78e-07 $l=8.95e-07 $layer=LI1_cond $X=2.535 $Y=0.845
+ $X2=1.64 $Y2=0.845
r47 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.65 $X2=3.56 $Y2=0.795
r48 2 23 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.695 $X2=2.54 $Y2=0.845
r49 1 12 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.695 $X2=1.64 $Y2=0.845
.ends


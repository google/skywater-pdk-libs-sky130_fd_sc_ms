* File: sky130_fd_sc_ms__dfrtn_1.pxi.spice
* Created: Fri Aug 28 17:22:18 2020
* 
x_PM_SKY130_FD_SC_MS__DFRTN_1%D N_D_c_232_n N_D_c_239_n N_D_M1030_g N_D_M1028_g
+ N_D_c_234_n N_D_c_235_n D D D N_D_c_236_n N_D_c_237_n
+ PM_SKY130_FD_SC_MS__DFRTN_1%D
x_PM_SKY130_FD_SC_MS__DFRTN_1%CLK_N N_CLK_N_c_270_n N_CLK_N_M1017_g
+ N_CLK_N_c_266_n N_CLK_N_M1013_g N_CLK_N_c_267_n N_CLK_N_c_268_n CLK_N
+ PM_SKY130_FD_SC_MS__DFRTN_1%CLK_N
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_510_74# N_A_510_74#_M1011_d N_A_510_74#_M1003_d
+ N_A_510_74#_M1006_g N_A_510_74#_c_334_n N_A_510_74#_M1014_g
+ N_A_510_74#_M1001_g N_A_510_74#_c_315_n N_A_510_74#_c_316_n
+ N_A_510_74#_c_317_n N_A_510_74#_M1022_g N_A_510_74#_c_318_n
+ N_A_510_74#_c_395_p N_A_510_74#_c_319_n N_A_510_74#_c_320_n
+ N_A_510_74#_c_321_n N_A_510_74#_c_322_n N_A_510_74#_c_323_n
+ N_A_510_74#_c_324_n N_A_510_74#_c_344_p N_A_510_74#_c_345_p
+ N_A_510_74#_c_325_n N_A_510_74#_c_326_n N_A_510_74#_c_327_n
+ N_A_510_74#_c_328_n N_A_510_74#_c_371_p N_A_510_74#_c_372_p
+ N_A_510_74#_c_329_n N_A_510_74#_c_330_n N_A_510_74#_c_338_n
+ N_A_510_74#_c_331_n N_A_510_74#_c_368_p N_A_510_74#_c_404_p
+ N_A_510_74#_c_332_n N_A_510_74#_c_333_n PM_SKY130_FD_SC_MS__DFRTN_1%A_510_74#
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_856_294# N_A_856_294#_M1020_d
+ N_A_856_294#_M1000_d N_A_856_294#_M1005_g N_A_856_294#_M1016_g
+ N_A_856_294#_c_502_n N_A_856_294#_c_503_n N_A_856_294#_c_504_n
+ N_A_856_294#_c_510_n N_A_856_294#_c_505_n N_A_856_294#_c_506_n
+ N_A_856_294#_c_507_n N_A_856_294#_c_540_p N_A_856_294#_c_541_p
+ N_A_856_294#_c_508_n PM_SKY130_FD_SC_MS__DFRTN_1%A_856_294#
x_PM_SKY130_FD_SC_MS__DFRTN_1%RESET_B N_RESET_B_M1024_g N_RESET_B_M1031_g
+ N_RESET_B_c_608_n N_RESET_B_c_609_n N_RESET_B_M1009_g N_RESET_B_M1018_g
+ N_RESET_B_M1010_g N_RESET_B_M1015_g N_RESET_B_c_596_n N_RESET_B_c_597_n
+ N_RESET_B_c_598_n N_RESET_B_c_599_n N_RESET_B_c_600_n N_RESET_B_c_601_n
+ RESET_B N_RESET_B_c_602_n N_RESET_B_c_603_n N_RESET_B_c_604_n
+ N_RESET_B_c_605_n N_RESET_B_c_606_n PM_SKY130_FD_SC_MS__DFRTN_1%RESET_B
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_714_119# N_A_714_119#_M1006_d
+ N_A_714_119#_M1012_d N_A_714_119#_M1018_d N_A_714_119#_M1020_g
+ N_A_714_119#_M1000_g N_A_714_119#_c_809_n N_A_714_119#_c_810_n
+ N_A_714_119#_c_826_n N_A_714_119#_c_811_n N_A_714_119#_c_818_n
+ N_A_714_119#_c_819_n N_A_714_119#_c_820_n N_A_714_119#_c_821_n
+ N_A_714_119#_c_812_n N_A_714_119#_c_813_n
+ PM_SKY130_FD_SC_MS__DFRTN_1%A_714_119#
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_300_347# N_A_300_347#_M1013_s
+ N_A_300_347#_M1017_s N_A_300_347#_c_914_n N_A_300_347#_M1011_g
+ N_A_300_347#_c_928_n N_A_300_347#_M1003_g N_A_300_347#_c_915_n
+ N_A_300_347#_c_916_n N_A_300_347#_c_917_n N_A_300_347#_c_929_n
+ N_A_300_347#_c_918_n N_A_300_347#_M1012_g N_A_300_347#_M1019_g
+ N_A_300_347#_c_920_n N_A_300_347#_M1007_g N_A_300_347#_c_932_n
+ N_A_300_347#_M1029_g N_A_300_347#_c_922_n N_A_300_347#_c_933_n
+ N_A_300_347#_c_944_n N_A_300_347#_c_947_n N_A_300_347#_c_948_n
+ N_A_300_347#_c_949_n N_A_300_347#_c_934_n N_A_300_347#_c_923_n
+ N_A_300_347#_c_936_n N_A_300_347#_c_937_n N_A_300_347#_c_924_n
+ N_A_300_347#_c_925_n N_A_300_347#_c_926_n N_A_300_347#_c_927_n
+ PM_SKY130_FD_SC_MS__DFRTN_1%A_300_347#
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_1598_93# N_A_1598_93#_M1004_d
+ N_A_1598_93#_M1015_d N_A_1598_93#_M1002_g N_A_1598_93#_M1008_g
+ N_A_1598_93#_c_1111_n N_A_1598_93#_c_1112_n N_A_1598_93#_c_1113_n
+ N_A_1598_93#_c_1114_n N_A_1598_93#_c_1107_n N_A_1598_93#_c_1116_n
+ N_A_1598_93#_c_1108_n PM_SKY130_FD_SC_MS__DFRTN_1%A_1598_93#
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_1266_119# N_A_1266_119#_M1007_d
+ N_A_1266_119#_M1001_d N_A_1266_119#_c_1194_n N_A_1266_119#_M1004_g
+ N_A_1266_119#_c_1195_n N_A_1266_119#_M1023_g N_A_1266_119#_c_1196_n
+ N_A_1266_119#_c_1206_n N_A_1266_119#_c_1207_n N_A_1266_119#_M1025_g
+ N_A_1266_119#_c_1197_n N_A_1266_119#_M1021_g N_A_1266_119#_c_1198_n
+ N_A_1266_119#_c_1215_n N_A_1266_119#_c_1208_n N_A_1266_119#_c_1199_n
+ N_A_1266_119#_c_1200_n N_A_1266_119#_c_1201_n N_A_1266_119#_c_1210_n
+ N_A_1266_119#_c_1223_n N_A_1266_119#_c_1202_n N_A_1266_119#_c_1203_n
+ PM_SKY130_FD_SC_MS__DFRTN_1%A_1266_119#
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_1934_94# N_A_1934_94#_M1021_s
+ N_A_1934_94#_M1025_s N_A_1934_94#_M1026_g N_A_1934_94#_M1027_g
+ N_A_1934_94#_c_1333_n N_A_1934_94#_c_1334_n N_A_1934_94#_c_1326_n
+ N_A_1934_94#_c_1327_n N_A_1934_94#_c_1328_n N_A_1934_94#_c_1329_n
+ N_A_1934_94#_c_1330_n N_A_1934_94#_c_1331_n
+ PM_SKY130_FD_SC_MS__DFRTN_1%A_1934_94#
x_PM_SKY130_FD_SC_MS__DFRTN_1%VPWR N_VPWR_M1030_s N_VPWR_M1031_d N_VPWR_M1017_d
+ N_VPWR_M1005_d N_VPWR_M1000_s N_VPWR_M1008_d N_VPWR_M1023_d N_VPWR_M1025_d
+ N_VPWR_c_1388_n N_VPWR_c_1389_n N_VPWR_c_1390_n N_VPWR_c_1391_n
+ N_VPWR_c_1392_n N_VPWR_c_1393_n N_VPWR_c_1394_n N_VPWR_c_1395_n
+ N_VPWR_c_1396_n N_VPWR_c_1397_n N_VPWR_c_1398_n N_VPWR_c_1399_n
+ N_VPWR_c_1400_n N_VPWR_c_1401_n VPWR N_VPWR_c_1402_n N_VPWR_c_1403_n
+ N_VPWR_c_1404_n N_VPWR_c_1405_n N_VPWR_c_1406_n N_VPWR_c_1387_n
+ N_VPWR_c_1408_n N_VPWR_c_1409_n N_VPWR_c_1410_n N_VPWR_c_1411_n
+ N_VPWR_c_1412_n PM_SKY130_FD_SC_MS__DFRTN_1%VPWR
x_PM_SKY130_FD_SC_MS__DFRTN_1%A_33_74# N_A_33_74#_M1028_s N_A_33_74#_M1006_s
+ N_A_33_74#_M1030_d N_A_33_74#_M1012_s N_A_33_74#_c_1515_n N_A_33_74#_c_1519_n
+ N_A_33_74#_c_1520_n N_A_33_74#_c_1516_n N_A_33_74#_c_1522_n
+ N_A_33_74#_c_1523_n N_A_33_74#_c_1524_n N_A_33_74#_c_1517_n
+ N_A_33_74#_c_1525_n N_A_33_74#_c_1526_n PM_SKY130_FD_SC_MS__DFRTN_1%A_33_74#
x_PM_SKY130_FD_SC_MS__DFRTN_1%Q N_Q_M1027_d N_Q_M1026_d N_Q_c_1601_n
+ N_Q_c_1602_n Q Q Q Q N_Q_c_1603_n PM_SKY130_FD_SC_MS__DFRTN_1%Q
x_PM_SKY130_FD_SC_MS__DFRTN_1%VGND N_VGND_M1024_d N_VGND_M1013_d N_VGND_M1009_d
+ N_VGND_M1002_d N_VGND_M1021_d N_VGND_c_1631_n N_VGND_c_1632_n N_VGND_c_1633_n
+ N_VGND_c_1634_n N_VGND_c_1635_n N_VGND_c_1636_n N_VGND_c_1637_n VGND
+ N_VGND_c_1638_n N_VGND_c_1639_n N_VGND_c_1640_n N_VGND_c_1641_n
+ N_VGND_c_1642_n N_VGND_c_1643_n N_VGND_c_1644_n N_VGND_c_1645_n
+ N_VGND_c_1646_n N_VGND_c_1647_n PM_SKY130_FD_SC_MS__DFRTN_1%VGND
cc_1 VNB N_D_c_232_n 0.0019217f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.92
cc_2 VNB N_D_M1028_g 0.027501f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_3 VNB N_D_c_234_n 0.0345854f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_4 VNB N_D_c_235_n 0.0229747f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_5 VNB N_D_c_236_n 0.0384952f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_6 VNB N_D_c_237_n 0.00478024f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_7 VNB N_CLK_N_c_266_n 0.0217863f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_8 VNB N_CLK_N_c_267_n 0.0399853f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.96
cc_9 VNB N_CLK_N_c_268_n 0.0137811f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_10 VNB CLK_N 0.00565793f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_11 VNB N_A_510_74#_M1006_g 0.023435f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_12 VNB N_A_510_74#_M1001_g 0.0165317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_510_74#_c_315_n 0.0171734f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_14 VNB N_A_510_74#_c_316_n 0.0191633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_510_74#_c_317_n 0.0231425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_510_74#_c_318_n 0.00558672f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_17 VNB N_A_510_74#_c_319_n 0.00979101f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=2.035
cc_18 VNB N_A_510_74#_c_320_n 0.00333238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_510_74#_c_321_n 0.00555068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_510_74#_c_322_n 0.062945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_510_74#_c_323_n 0.0166425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_510_74#_c_324_n 0.00103032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_510_74#_c_325_n 0.00384221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_510_74#_c_326_n 0.0193653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_510_74#_c_327_n 0.00260538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_510_74#_c_328_n 0.00739636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_510_74#_c_329_n 0.00166696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_510_74#_c_330_n 0.0294493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_510_74#_c_331_n 6.24913e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_510_74#_c_332_n 0.00628108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_510_74#_c_333_n 0.0169284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_856_294#_M1016_g 0.0305572f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_33 VNB N_A_856_294#_c_502_n 0.0155687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_856_294#_c_503_n 0.00201458f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_35 VNB N_A_856_294#_c_504_n 0.00112198f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_A_856_294#_c_505_n 0.00267139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_856_294#_c_506_n 0.0181271f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_38 VNB N_A_856_294#_c_507_n 0.00163478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_856_294#_c_508_n 0.0021497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_M1024_g 0.050311f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.07
cc_41 VNB N_RESET_B_M1009_g 0.0413741f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_42 VNB N_RESET_B_M1010_g 0.034399f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_43 VNB N_RESET_B_c_596_n 0.0114201f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_44 VNB N_RESET_B_c_597_n 0.00226973f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_45 VNB N_RESET_B_c_598_n 0.013881f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.125
cc_46 VNB N_RESET_B_c_599_n 5.71827e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_600_n 6.54175e-19 $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=2.035
cc_48 VNB N_RESET_B_c_601_n 0.00357755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_RESET_B_c_602_n 0.0287856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_603_n 0.0157912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_RESET_B_c_604_n 0.00223158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_c_605_n 0.0154637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_RESET_B_c_606_n 0.00570331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_714_119#_M1020_g 0.0201455f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.96
cc_55 VNB N_A_714_119#_c_809_n 0.0216047f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_56 VNB N_A_714_119#_c_810_n 0.00936918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_714_119#_c_811_n 0.00546417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_714_119#_c_812_n 0.00306892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_714_119#_c_813_n 0.00111181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_300_347#_c_914_n 0.0181086f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.96
cc_61 VNB N_A_300_347#_c_915_n 0.0502825f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_62 VNB N_A_300_347#_c_916_n 0.0684595f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_63 VNB N_A_300_347#_c_917_n 0.012382f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.995
cc_64 VNB N_A_300_347#_c_918_n 0.0516615f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_65 VNB N_A_300_347#_M1019_g 0.0385923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_300_347#_c_920_n 0.149745f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_67 VNB N_A_300_347#_M1007_g 0.030044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_300_347#_c_922_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_300_347#_c_923_n 0.00454971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_300_347#_c_924_n 0.00266304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_300_347#_c_925_n 0.00102467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_300_347#_c_926_n 0.00265148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_300_347#_c_927_n 0.018162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1598_93#_M1002_g 0.0473326f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_75 VNB N_A_1598_93#_c_1107_n 0.0107986f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_76 VNB N_A_1598_93#_c_1108_n 0.0121095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1266_119#_c_1194_n 0.0202606f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=0.96
cc_78 VNB N_A_1266_119#_c_1195_n 0.00226217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1266_119#_c_1196_n 0.0586053f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.465
cc_80 VNB N_A_1266_119#_c_1197_n 0.0219742f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_81 VNB N_A_1266_119#_c_1198_n 0.00948676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1266_119#_c_1199_n 0.00100139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1266_119#_c_1200_n 0.0107396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1266_119#_c_1201_n 0.0235899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1266_119#_c_1202_n 5.53899e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1266_119#_c_1203_n 0.024655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1934_94#_M1026_g 6.28484e-19 $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_88 VNB N_A_1934_94#_c_1326_n 0.00180273f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_89 VNB N_A_1934_94#_c_1327_n 2.65185e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1934_94#_c_1328_n 0.0106069f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_91 VNB N_A_1934_94#_c_1329_n 0.0403233f $X=-0.19 $Y=-0.245 $X2=0.237
+ $Y2=1.125
cc_92 VNB N_A_1934_94#_c_1330_n 0.00429191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1934_94#_c_1331_n 0.0213736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VPWR_c_1387_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_33_74#_c_1515_n 0.0122181f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_96 VNB N_A_33_74#_c_1516_n 0.015603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_33_74#_c_1517_n 0.0216357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_Q_c_1601_n 0.0243417f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_99 VNB N_Q_c_1602_n 0.00719696f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_100 VNB N_Q_c_1603_n 0.0236298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1631_n 0.0122824f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_102 VNB N_VGND_c_1632_n 0.00958887f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_103 VNB N_VGND_c_1633_n 0.0079779f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_104 VNB N_VGND_c_1634_n 0.0246564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1635_n 0.017712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1636_n 0.0309922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1637_n 0.00384695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1638_n 0.0226942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1639_n 0.0661307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1640_n 0.0716605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1641_n 0.0470737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1642_n 0.0198148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1643_n 0.610492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1644_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1645_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1646_n 0.00846329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1647_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VPB N_D_c_232_n 0.0175641f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.92
cc_119 VPB N_D_c_239_n 0.0220466f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.07
cc_120 VPB N_D_M1030_g 0.050484f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_121 VPB N_D_c_237_n 0.0217648f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_122 VPB N_CLK_N_c_270_n 0.0172106f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.63
cc_123 VPB N_CLK_N_c_267_n 0.0227968f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.96
cc_124 VPB N_CLK_N_c_268_n 0.00356384f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_125 VPB N_A_510_74#_c_334_n 0.00498296f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_126 VPB N_A_510_74#_M1014_g 0.0182608f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_127 VPB N_A_510_74#_M1001_g 0.036977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_510_74#_c_318_n 0.0172149f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_129 VPB N_A_510_74#_c_338_n 0.00134652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_510_74#_c_331_n 3.9332e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_856_294#_M1005_g 0.0361583f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_132 VPB N_A_856_294#_c_510_n 0.00689908f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_133 VPB N_A_856_294#_c_505_n 0.00151059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_856_294#_c_506_n 0.0120152f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_135 VPB N_A_856_294#_c_508_n 0.00238414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_M1031_g 0.0699098f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_137 VPB N_RESET_B_c_608_n 0.295722f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_138 VPB N_RESET_B_c_609_n 0.0138441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_RESET_B_M1018_g 0.0570425f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_140 VPB N_RESET_B_M1015_g 0.0509916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_RESET_B_c_596_n 0.0135354f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_142 VPB N_RESET_B_c_597_n 0.00395013f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_143 VPB N_RESET_B_c_598_n 0.00673887f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.125
cc_144 VPB N_RESET_B_c_599_n 5.68911e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_RESET_B_c_600_n 6.35107e-19 $X=-0.19 $Y=1.66 $X2=0.237 $Y2=2.035
cc_146 VPB N_RESET_B_c_601_n 0.00257552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_602_n 0.00607708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_c_603_n 0.0106707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_604_n 0.00127854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_605_n 0.0112707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_606_n 0.00331027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_714_119#_M1000_g 0.0287765f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_153 VPB N_A_714_119#_c_809_n 0.017529f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_154 VPB N_A_714_119#_c_810_n 0.00603589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_714_119#_c_811_n 0.00326143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_714_119#_c_818_n 0.0159486f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_157 VPB N_A_714_119#_c_819_n 0.00562343f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_158 VPB N_A_714_119#_c_820_n 0.00976667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_714_119#_c_821_n 0.0137564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_714_119#_c_812_n 0.00435853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_300_347#_c_928_n 0.0187075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_300_347#_c_929_n 0.0373826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_300_347#_c_918_n 0.0366414f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_164 VPB N_A_300_347#_M1012_g 0.0350994f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_165 VPB N_A_300_347#_c_932_n 0.0198187f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.665
cc_166 VPB N_A_300_347#_c_933_n 0.0317515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_300_347#_c_934_n 0.00237373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_300_347#_c_923_n 0.0168815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_300_347#_c_936_n 0.00232654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_300_347#_c_937_n 0.0462021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_300_347#_c_926_n 0.00280482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_300_347#_c_927_n 0.0167017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_1598_93#_M1002_g 0.01871f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_174 VPB N_A_1598_93#_M1008_g 0.0246517f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_175 VPB N_A_1598_93#_c_1111_n 0.00706063f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_176 VPB N_A_1598_93#_c_1112_n 0.0299411f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_177 VPB N_A_1598_93#_c_1113_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_178 VPB N_A_1598_93#_c_1114_n 0.00960971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_1598_93#_c_1107_n 0.00471733f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_180 VPB N_A_1598_93#_c_1116_n 0.00400474f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_181 VPB N_A_1266_119#_c_1195_n 0.023609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1266_119#_M1023_g 0.0438211f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=0.96
cc_183 VPB N_A_1266_119#_c_1206_n 0.0584058f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_184 VPB N_A_1266_119#_c_1207_n 0.0199894f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_185 VPB N_A_1266_119#_c_1208_n 0.00674641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1266_119#_c_1200_n 0.0132627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1266_119#_c_1210_n 8.88119e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1266_119#_c_1202_n 5.52803e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1934_94#_M1026_g 0.0309281f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_190 VPB N_A_1934_94#_c_1333_n 0.00267961f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_191 VPB N_A_1934_94#_c_1334_n 0.00737227f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_192 VPB N_A_1934_94#_c_1327_n 0.00591066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1388_n 0.0117348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1389_n 0.0298144f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_195 VPB N_VPWR_c_1390_n 0.00952052f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_196 VPB N_VPWR_c_1391_n 0.0150793f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=2.035
cc_197 VPB N_VPWR_c_1392_n 0.0160325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1393_n 0.0188116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1394_n 0.012578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1395_n 0.00904539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1396_n 0.0160669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1397_n 0.00975786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1398_n 0.0620036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1399_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1400_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1401_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1402_n 0.0165238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1403_n 0.0186862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1404_n 0.0619539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1405_n 0.0209223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1406_n 0.0197908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1387_n 0.100413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1408_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1409_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1410_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1411_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1412_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_33_74#_c_1515_n 0.00638129f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_219 VPB N_A_33_74#_c_1519_n 0.00347606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_33_74#_c_1520_n 0.020238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_33_74#_c_1516_n 0.00162035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_33_74#_c_1522_n 0.00104047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_33_74#_c_1523_n 0.00464675f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_224 VPB N_A_33_74#_c_1524_n 0.00709844f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.125
cc_225 VPB N_A_33_74#_c_1525_n 0.00693612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_33_74#_c_1526_n 0.00332765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB Q 0.00916683f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_228 VPB Q 0.0415238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_Q_c_1603_n 0.00763418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 N_D_M1028_g N_RESET_B_M1024_g 0.0435282f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_231 N_D_c_236_n N_RESET_B_M1024_g 0.00520474f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_232 N_D_c_232_n N_RESET_B_M1031_g 0.00462577f $X=0.36 $Y=1.92 $X2=0 $Y2=0
cc_233 N_D_c_239_n N_RESET_B_M1031_g 0.0171858f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_234 N_D_M1030_g N_RESET_B_c_609_n 0.0171858f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_235 N_D_c_236_n N_RESET_B_c_602_n 0.00877288f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_236 N_D_c_239_n N_VPWR_c_1389_n 0.00199186f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_237 N_D_M1030_g N_VPWR_c_1389_n 0.013284f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_238 N_D_c_237_n N_VPWR_c_1389_n 0.0140568f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_239 N_D_M1030_g N_VPWR_c_1402_n 0.00460063f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_240 N_D_M1030_g N_VPWR_c_1387_n 0.00908665f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_241 N_D_c_239_n N_A_33_74#_c_1515_n 0.00493555f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_242 N_D_M1030_g N_A_33_74#_c_1515_n 0.00297569f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_243 N_D_M1028_g N_A_33_74#_c_1515_n 0.00857134f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_244 N_D_c_234_n N_A_33_74#_c_1515_n 0.00517676f $X=0.352 $Y=1.11 $X2=0 $Y2=0
cc_245 N_D_c_236_n N_A_33_74#_c_1515_n 0.00665742f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_246 N_D_c_237_n N_A_33_74#_c_1515_n 0.0866708f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_247 N_D_M1030_g N_A_33_74#_c_1519_n 0.00403937f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_248 N_D_M1028_g N_A_33_74#_c_1517_n 0.0152419f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_249 N_D_c_234_n N_A_33_74#_c_1517_n 0.0040449f $X=0.352 $Y=1.11 $X2=0 $Y2=0
cc_250 N_D_c_237_n N_A_33_74#_c_1517_n 0.0188861f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_251 N_D_M1030_g N_A_33_74#_c_1525_n 0.013859f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_252 N_D_M1028_g N_VGND_c_1636_n 0.00291649f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_253 N_D_M1028_g N_VGND_c_1643_n 0.00362587f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_254 N_CLK_N_c_267_n N_RESET_B_M1024_g 0.00489911f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_255 CLK_N N_RESET_B_M1024_g 0.00149212f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_256 N_CLK_N_c_270_n N_RESET_B_c_608_n 0.0121828f $X=1.915 $Y=1.66 $X2=0 $Y2=0
cc_257 N_CLK_N_c_270_n N_RESET_B_c_596_n 0.00382256f $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_258 N_CLK_N_c_267_n N_RESET_B_c_596_n 0.0129154f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_259 N_CLK_N_c_268_n N_RESET_B_c_596_n 0.00347556f $X=1.915 $Y=1.435 $X2=0
+ $Y2=0
cc_260 CLK_N N_RESET_B_c_596_n 0.00897634f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_261 N_CLK_N_c_267_n N_RESET_B_c_597_n 8.07459e-19 $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_262 CLK_N N_RESET_B_c_597_n 7.30635e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_263 N_CLK_N_c_270_n N_RESET_B_c_602_n 2.43058e-19 $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_264 N_CLK_N_c_267_n N_RESET_B_c_602_n 0.0192274f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_265 N_CLK_N_c_270_n N_RESET_B_c_606_n 0.00138451f $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_266 N_CLK_N_c_267_n N_RESET_B_c_606_n 0.00365613f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_267 CLK_N N_RESET_B_c_606_n 0.0172783f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_268 N_CLK_N_c_266_n N_A_300_347#_c_914_n 0.0196269f $X=1.93 $Y=1.21 $X2=0
+ $Y2=0
cc_269 N_CLK_N_c_270_n N_A_300_347#_c_928_n 0.0334377f $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_270 N_CLK_N_c_268_n N_A_300_347#_c_918_n 0.0238835f $X=1.915 $Y=1.435 $X2=0
+ $Y2=0
cc_271 CLK_N N_A_300_347#_c_918_n 2.91382e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_272 N_CLK_N_c_270_n N_A_300_347#_c_944_n 0.010947f $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_273 N_CLK_N_c_267_n N_A_300_347#_c_944_n 0.00569548f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_274 CLK_N N_A_300_347#_c_944_n 0.00932989f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_275 N_CLK_N_c_266_n N_A_300_347#_c_947_n 0.00555768f $X=1.93 $Y=1.21 $X2=0
+ $Y2=0
cc_276 N_CLK_N_c_266_n N_A_300_347#_c_948_n 0.0121467f $X=1.93 $Y=1.21 $X2=0
+ $Y2=0
cc_277 N_CLK_N_c_266_n N_A_300_347#_c_949_n 3.9078e-19 $X=1.93 $Y=1.21 $X2=0
+ $Y2=0
cc_278 N_CLK_N_c_267_n N_A_300_347#_c_949_n 0.00437066f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_279 CLK_N N_A_300_347#_c_949_n 0.020061f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_280 N_CLK_N_c_270_n N_A_300_347#_c_934_n 0.00449677f $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_281 N_CLK_N_c_268_n N_A_300_347#_c_924_n 0.00449677f $X=1.915 $Y=1.435 $X2=0
+ $Y2=0
cc_282 N_CLK_N_c_266_n N_A_300_347#_c_925_n 0.00449677f $X=1.93 $Y=1.21 $X2=0
+ $Y2=0
cc_283 CLK_N N_A_300_347#_c_925_n 0.0173205f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_284 N_CLK_N_c_270_n N_VPWR_c_1390_n 0.00581454f $X=1.915 $Y=1.66 $X2=0 $Y2=0
cc_285 N_CLK_N_c_270_n N_VPWR_c_1391_n 0.00329659f $X=1.915 $Y=1.66 $X2=0 $Y2=0
cc_286 N_CLK_N_c_270_n N_VPWR_c_1387_n 0.00112709f $X=1.915 $Y=1.66 $X2=0 $Y2=0
cc_287 N_CLK_N_c_270_n N_A_33_74#_c_1520_n 0.0174663f $X=1.915 $Y=1.66 $X2=0
+ $Y2=0
cc_288 N_CLK_N_c_267_n N_A_33_74#_c_1520_n 0.00321633f $X=1.825 $Y=1.435 $X2=0
+ $Y2=0
cc_289 CLK_N N_A_33_74#_c_1520_n 7.01254e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_290 N_CLK_N_c_266_n N_VGND_c_1631_n 0.00311242f $X=1.93 $Y=1.21 $X2=0 $Y2=0
cc_291 N_CLK_N_c_266_n N_VGND_c_1632_n 0.00378344f $X=1.93 $Y=1.21 $X2=0 $Y2=0
cc_292 N_CLK_N_c_266_n N_VGND_c_1638_n 0.00451627f $X=1.93 $Y=1.21 $X2=0 $Y2=0
cc_293 N_CLK_N_c_266_n N_VGND_c_1643_n 0.0045447f $X=1.93 $Y=1.21 $X2=0 $Y2=0
cc_294 N_A_510_74#_c_334_n N_A_856_294#_M1005_g 0.0497452f $X=4.01 $Y=2.11 $X2=0
+ $Y2=0
cc_295 N_A_510_74#_c_318_n N_A_856_294#_M1005_g 0.0116006f $X=4.01 $Y=2.02 $X2=0
+ $Y2=0
cc_296 N_A_510_74#_c_322_n N_A_856_294#_M1016_g 0.00376909f $X=3.62 $Y=1.41
+ $X2=0 $Y2=0
cc_297 N_A_510_74#_c_324_n N_A_856_294#_M1016_g 0.00692821f $X=4.38 $Y=0.79
+ $X2=0 $Y2=0
cc_298 N_A_510_74#_c_344_p N_A_856_294#_M1016_g 0.00707231f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_299 N_A_510_74#_c_345_p N_A_856_294#_M1016_g 0.00117472f $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_300 N_A_510_74#_c_344_p N_A_856_294#_c_502_n 0.072849f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_301 N_A_510_74#_c_344_p N_A_856_294#_c_503_n 0.0109977f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_302 N_A_510_74#_c_345_p N_A_856_294#_c_503_n 0.00135883f $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_303 N_A_510_74#_c_326_n N_A_856_294#_c_504_n 0.0206843f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_304 N_A_510_74#_M1001_g N_A_856_294#_c_510_n 9.54046e-19 $X=6.81 $Y=2.46
+ $X2=0 $Y2=0
cc_305 N_A_510_74#_c_322_n N_A_856_294#_c_505_n 0.00113532f $X=3.62 $Y=1.41
+ $X2=0 $Y2=0
cc_306 N_A_510_74#_c_345_p N_A_856_294#_c_505_n 0.0041441f $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_307 N_A_510_74#_c_322_n N_A_856_294#_c_506_n 0.0214458f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_A_510_74#_c_345_p N_A_856_294#_c_506_n 7.42944e-19 $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_309 N_A_510_74#_c_322_n N_A_856_294#_c_507_n 5.57305e-19 $X=3.62 $Y=1.41
+ $X2=0 $Y2=0
cc_310 N_A_510_74#_M1001_g N_A_856_294#_c_508_n 0.0024704f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_311 N_A_510_74#_M1014_g N_RESET_B_c_608_n 0.0102218f $X=4.01 $Y=2.495 $X2=0
+ $Y2=0
cc_312 N_A_510_74#_c_324_n N_RESET_B_M1009_g 0.00125222f $X=4.38 $Y=0.79 $X2=0
+ $Y2=0
cc_313 N_A_510_74#_c_344_p N_RESET_B_M1009_g 0.0113546f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_314 N_A_510_74#_c_325_n N_RESET_B_M1009_g 0.00405244f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_315 N_A_510_74#_M1003_d N_RESET_B_c_596_n 5.99887e-19 $X=2.59 $Y=1.735 $X2=0
+ $Y2=0
cc_316 N_A_510_74#_c_334_n N_RESET_B_c_596_n 7.80952e-19 $X=4.01 $Y=2.11 $X2=0
+ $Y2=0
cc_317 N_A_510_74#_c_318_n N_RESET_B_c_596_n 0.00102117f $X=4.01 $Y=2.02 $X2=0
+ $Y2=0
cc_318 N_A_510_74#_c_321_n N_RESET_B_c_596_n 0.0101687f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_510_74#_c_322_n N_RESET_B_c_596_n 0.00602217f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_320 N_A_510_74#_c_338_n N_RESET_B_c_596_n 0.00536125f $X=2.73 $Y=1.915 $X2=0
+ $Y2=0
cc_321 N_A_510_74#_c_331_n N_RESET_B_c_596_n 0.0258163f $X=2.752 $Y=1.745 $X2=0
+ $Y2=0
cc_322 N_A_510_74#_c_368_p N_RESET_B_c_596_n 5.77133e-19 $X=2.792 $Y=1.09 $X2=0
+ $Y2=0
cc_323 N_A_510_74#_M1001_g N_RESET_B_c_598_n 0.00221676f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_324 N_A_510_74#_c_316_n N_RESET_B_c_598_n 0.00405791f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_325 N_A_510_74#_c_371_p N_RESET_B_c_598_n 0.00155657f $X=6.535 $Y=1.21 $X2=0
+ $Y2=0
cc_326 N_A_510_74#_c_372_p N_RESET_B_c_598_n 0.0169144f $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_327 N_A_510_74#_c_330_n N_RESET_B_c_598_n 0.011489f $X=7.255 $Y=1.29 $X2=0
+ $Y2=0
cc_328 N_A_510_74#_c_332_n N_RESET_B_c_598_n 0.00501712f $X=6.75 $Y=1.29 $X2=0
+ $Y2=0
cc_329 N_A_510_74#_c_321_n N_A_714_119#_M1006_d 0.00405707f $X=3.62 $Y=1.41
+ $X2=-0.19 $Y2=-0.245
cc_330 N_A_510_74#_c_325_n N_A_714_119#_M1020_g 0.00745398f $X=5.61 $Y=0.79
+ $X2=0 $Y2=0
cc_331 N_A_510_74#_c_326_n N_A_714_119#_M1020_g 0.00330666f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_332 N_A_510_74#_M1006_g N_A_714_119#_c_826_n 0.00188226f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_333 N_A_510_74#_c_321_n N_A_714_119#_c_826_n 0.0756934f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_334 N_A_510_74#_c_323_n N_A_714_119#_c_826_n 0.0171642f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_335 N_A_510_74#_c_318_n N_A_714_119#_c_811_n 0.0132003f $X=4.01 $Y=2.02 $X2=0
+ $Y2=0
cc_336 N_A_510_74#_c_322_n N_A_714_119#_c_811_n 0.0142202f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_337 N_A_510_74#_c_334_n N_A_714_119#_c_818_n 0.00184165f $X=4.01 $Y=2.11
+ $X2=0 $Y2=0
cc_338 N_A_510_74#_M1014_g N_A_714_119#_c_818_n 0.00290452f $X=4.01 $Y=2.495
+ $X2=0 $Y2=0
cc_339 N_A_510_74#_c_334_n N_A_714_119#_c_819_n 0.00151956f $X=4.01 $Y=2.11
+ $X2=0 $Y2=0
cc_340 N_A_510_74#_M1014_g N_A_714_119#_c_819_n 0.0167327f $X=4.01 $Y=2.495
+ $X2=0 $Y2=0
cc_341 N_A_510_74#_c_321_n N_A_714_119#_c_819_n 0.001505f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_342 N_A_510_74#_c_322_n N_A_714_119#_c_819_n 0.004295f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_343 N_A_510_74#_c_322_n N_A_714_119#_c_813_n 5.85608e-19 $X=3.62 $Y=1.41
+ $X2=0 $Y2=0
cc_344 N_A_510_74#_c_320_n N_A_300_347#_c_914_n 0.00175296f $X=2.94 $Y=0.36
+ $X2=0 $Y2=0
cc_345 N_A_510_74#_c_331_n N_A_300_347#_c_914_n 8.38974e-19 $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_346 N_A_510_74#_c_338_n N_A_300_347#_c_928_n 0.00356981f $X=2.73 $Y=1.915
+ $X2=0 $Y2=0
cc_347 N_A_510_74#_c_331_n N_A_300_347#_c_928_n 6.09784e-19 $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_348 N_A_510_74#_M1006_g N_A_300_347#_c_915_n 0.0135287f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_349 N_A_510_74#_c_395_p N_A_300_347#_c_915_n 0.0117407f $X=2.73 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_510_74#_c_319_n N_A_300_347#_c_915_n 0.0130864f $X=3.535 $Y=0.36
+ $X2=0 $Y2=0
cc_351 N_A_510_74#_c_320_n N_A_300_347#_c_915_n 0.00276418f $X=2.94 $Y=0.36
+ $X2=0 $Y2=0
cc_352 N_A_510_74#_c_321_n N_A_300_347#_c_915_n 7.68901e-19 $X=3.62 $Y=1.41
+ $X2=0 $Y2=0
cc_353 N_A_510_74#_c_331_n N_A_300_347#_c_915_n 0.00249267f $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_354 N_A_510_74#_c_368_p N_A_300_347#_c_915_n 0.00318247f $X=2.792 $Y=1.09
+ $X2=0 $Y2=0
cc_355 N_A_510_74#_M1006_g N_A_300_347#_c_916_n 0.00902735f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_356 N_A_510_74#_c_319_n N_A_300_347#_c_916_n 0.00670492f $X=3.535 $Y=0.36
+ $X2=0 $Y2=0
cc_357 N_A_510_74#_c_323_n N_A_300_347#_c_916_n 0.0072068f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_358 N_A_510_74#_c_404_p N_A_300_347#_c_916_n 0.0036181f $X=3.62 $Y=0.36 $X2=0
+ $Y2=0
cc_359 N_A_510_74#_c_318_n N_A_300_347#_c_929_n 0.0154492f $X=4.01 $Y=2.02 $X2=0
+ $Y2=0
cc_360 N_A_510_74#_c_321_n N_A_300_347#_c_929_n 0.0021958f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_361 N_A_510_74#_c_322_n N_A_300_347#_c_929_n 0.0162271f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_362 N_A_510_74#_c_322_n N_A_300_347#_c_918_n 0.0135287f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_363 N_A_510_74#_c_338_n N_A_300_347#_c_918_n 0.00568969f $X=2.73 $Y=1.915
+ $X2=0 $Y2=0
cc_364 N_A_510_74#_c_331_n N_A_300_347#_c_918_n 0.0298156f $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_365 N_A_510_74#_c_368_p N_A_300_347#_c_918_n 0.0010507f $X=2.792 $Y=1.09
+ $X2=0 $Y2=0
cc_366 N_A_510_74#_c_334_n N_A_300_347#_M1012_g 0.0154492f $X=4.01 $Y=2.11 $X2=0
+ $Y2=0
cc_367 N_A_510_74#_M1006_g N_A_300_347#_M1019_g 0.009038f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_368 N_A_510_74#_c_321_n N_A_300_347#_M1019_g 0.00208822f $X=3.62 $Y=1.41
+ $X2=0 $Y2=0
cc_369 N_A_510_74#_c_323_n N_A_300_347#_M1019_g 0.0191653f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_370 N_A_510_74#_c_324_n N_A_300_347#_M1019_g 0.00212663f $X=4.38 $Y=0.79
+ $X2=0 $Y2=0
cc_371 N_A_510_74#_c_323_n N_A_300_347#_c_920_n 0.00435896f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_372 N_A_510_74#_c_344_p N_A_300_347#_c_920_n 0.00966127f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_373 N_A_510_74#_c_326_n N_A_300_347#_c_920_n 0.00676815f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_374 N_A_510_74#_c_327_n N_A_300_347#_c_920_n 0.0041995f $X=5.695 $Y=0.34
+ $X2=0 $Y2=0
cc_375 N_A_510_74#_c_315_n N_A_300_347#_M1007_g 0.00954257f $X=6.9 $Y=1.29 $X2=0
+ $Y2=0
cc_376 N_A_510_74#_c_325_n N_A_300_347#_M1007_g 8.97611e-19 $X=5.61 $Y=0.79
+ $X2=0 $Y2=0
cc_377 N_A_510_74#_c_326_n N_A_300_347#_M1007_g 0.0169375f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_378 N_A_510_74#_c_328_n N_A_300_347#_M1007_g 0.0152469f $X=6.45 $Y=1.125
+ $X2=0 $Y2=0
cc_379 N_A_510_74#_c_372_p N_A_300_347#_M1007_g 8.5704e-19 $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_380 N_A_510_74#_M1001_g N_A_300_347#_c_933_n 0.0081292f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_381 N_A_510_74#_c_395_p N_A_300_347#_c_948_n 0.0163074f $X=2.73 $Y=0.56 $X2=0
+ $Y2=0
cc_382 N_A_510_74#_c_331_n N_A_300_347#_c_934_n 0.00686016f $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_383 N_A_510_74#_M1001_g N_A_300_347#_c_923_n 0.017003f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_384 N_A_510_74#_c_316_n N_A_300_347#_c_923_n 0.00107089f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_385 N_A_510_74#_c_371_p N_A_300_347#_c_923_n 8.672e-19 $X=6.535 $Y=1.21 $X2=0
+ $Y2=0
cc_386 N_A_510_74#_c_372_p N_A_300_347#_c_923_n 0.0348735f $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_387 N_A_510_74#_c_329_n N_A_300_347#_c_923_n 0.00717074f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_388 N_A_510_74#_c_330_n N_A_300_347#_c_923_n 0.00892364f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_389 N_A_510_74#_c_332_n N_A_300_347#_c_923_n 0.00691585f $X=6.75 $Y=1.29
+ $X2=0 $Y2=0
cc_390 N_A_510_74#_c_333_n N_A_300_347#_c_923_n 6.09268e-19 $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_391 N_A_510_74#_M1001_g N_A_300_347#_c_936_n 0.00257707f $X=6.81 $Y=2.46
+ $X2=0 $Y2=0
cc_392 N_A_510_74#_M1001_g N_A_300_347#_c_937_n 0.0194681f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_393 N_A_510_74#_c_316_n N_A_300_347#_c_937_n 0.00873909f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_394 N_A_510_74#_c_333_n N_A_300_347#_c_937_n 0.00582183f $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_395 N_A_510_74#_c_331_n N_A_300_347#_c_924_n 0.0263792f $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_396 N_A_510_74#_c_331_n N_A_300_347#_c_925_n 0.00877966f $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_397 N_A_510_74#_c_368_p N_A_300_347#_c_925_n 0.00611922f $X=2.792 $Y=1.09
+ $X2=0 $Y2=0
cc_398 N_A_510_74#_M1001_g N_A_300_347#_c_926_n 0.00134673f $X=6.81 $Y=2.46
+ $X2=0 $Y2=0
cc_399 N_A_510_74#_c_371_p N_A_300_347#_c_926_n 0.00994746f $X=6.535 $Y=1.21
+ $X2=0 $Y2=0
cc_400 N_A_510_74#_M1001_g N_A_300_347#_c_927_n 0.021585f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_401 N_A_510_74#_c_371_p N_A_300_347#_c_927_n 0.00106755f $X=6.535 $Y=1.21
+ $X2=0 $Y2=0
cc_402 N_A_510_74#_c_317_n N_A_1598_93#_M1002_g 0.0413341f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_403 N_A_510_74#_c_333_n N_A_1598_93#_M1002_g 0.00246675f $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_404 N_A_510_74#_c_328_n N_A_1266_119#_M1007_d 0.0153989f $X=6.45 $Y=1.125
+ $X2=-0.19 $Y2=-0.245
cc_405 N_A_510_74#_c_371_p N_A_1266_119#_M1007_d 0.00269935f $X=6.535 $Y=1.21
+ $X2=-0.19 $Y2=-0.245
cc_406 N_A_510_74#_c_332_n N_A_1266_119#_M1007_d 0.0025788f $X=6.75 $Y=1.29
+ $X2=-0.19 $Y2=-0.245
cc_407 N_A_510_74#_c_315_n N_A_1266_119#_c_1215_n 0.0198469f $X=6.9 $Y=1.29
+ $X2=0 $Y2=0
cc_408 N_A_510_74#_c_317_n N_A_1266_119#_c_1215_n 0.0148493f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_409 N_A_510_74#_c_328_n N_A_1266_119#_c_1215_n 0.0266855f $X=6.45 $Y=1.125
+ $X2=0 $Y2=0
cc_410 N_A_510_74#_c_332_n N_A_1266_119#_c_1215_n 0.0553581f $X=6.75 $Y=1.29
+ $X2=0 $Y2=0
cc_411 N_A_510_74#_M1001_g N_A_1266_119#_c_1208_n 0.00568969f $X=6.81 $Y=2.46
+ $X2=0 $Y2=0
cc_412 N_A_510_74#_c_317_n N_A_1266_119#_c_1199_n 0.00779099f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_413 N_A_510_74#_c_329_n N_A_1266_119#_c_1200_n 0.0080525f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_414 N_A_510_74#_c_333_n N_A_1266_119#_c_1200_n 6.25344e-19 $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_415 N_A_510_74#_c_316_n N_A_1266_119#_c_1223_n 0.00534427f $X=7.6 $Y=1.2
+ $X2=0 $Y2=0
cc_416 N_A_510_74#_c_329_n N_A_1266_119#_c_1223_n 0.00890259f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_417 N_A_510_74#_M1001_g N_VPWR_c_1398_n 0.00522773f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_418 N_A_510_74#_M1014_g N_VPWR_c_1387_n 0.00113998f $X=4.01 $Y=2.495 $X2=0
+ $Y2=0
cc_419 N_A_510_74#_M1001_g N_VPWR_c_1387_n 0.00991118f $X=6.81 $Y=2.46 $X2=0
+ $Y2=0
cc_420 N_A_510_74#_M1003_d N_A_33_74#_c_1520_n 0.00670029f $X=2.59 $Y=1.735
+ $X2=0 $Y2=0
cc_421 N_A_510_74#_c_338_n N_A_33_74#_c_1520_n 0.0247906f $X=2.73 $Y=1.915 $X2=0
+ $Y2=0
cc_422 N_A_510_74#_M1006_g N_A_33_74#_c_1516_n 0.00510675f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_423 N_A_510_74#_c_318_n N_A_33_74#_c_1516_n 6.4404e-19 $X=4.01 $Y=2.02 $X2=0
+ $Y2=0
cc_424 N_A_510_74#_c_395_p N_A_33_74#_c_1516_n 0.0339533f $X=2.73 $Y=0.56 $X2=0
+ $Y2=0
cc_425 N_A_510_74#_c_319_n N_A_33_74#_c_1516_n 0.0196918f $X=3.535 $Y=0.36 $X2=0
+ $Y2=0
cc_426 N_A_510_74#_c_321_n N_A_33_74#_c_1516_n 0.0609976f $X=3.62 $Y=1.41 $X2=0
+ $Y2=0
cc_427 N_A_510_74#_c_368_p N_A_33_74#_c_1522_n 0.0339533f $X=2.792 $Y=1.09 $X2=0
+ $Y2=0
cc_428 N_A_510_74#_c_331_n N_A_33_74#_c_1523_n 0.0339533f $X=2.752 $Y=1.745
+ $X2=0 $Y2=0
cc_429 N_A_510_74#_c_344_p N_VGND_M1009_d 0.0158358f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_430 N_A_510_74#_c_325_n N_VGND_M1009_d 0.00465623f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_431 N_A_510_74#_c_320_n N_VGND_c_1632_n 0.0100832f $X=2.94 $Y=0.36 $X2=0
+ $Y2=0
cc_432 N_A_510_74#_c_323_n N_VGND_c_1633_n 0.00810195f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_433 N_A_510_74#_c_324_n N_VGND_c_1633_n 0.00427355f $X=4.38 $Y=0.79 $X2=0
+ $Y2=0
cc_434 N_A_510_74#_c_344_p N_VGND_c_1633_n 0.0259789f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_435 N_A_510_74#_c_325_n N_VGND_c_1633_n 0.015351f $X=5.61 $Y=0.79 $X2=0 $Y2=0
cc_436 N_A_510_74#_c_327_n N_VGND_c_1633_n 0.0150385f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_437 N_A_510_74#_c_317_n N_VGND_c_1634_n 0.00102171f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_438 N_A_510_74#_c_319_n N_VGND_c_1639_n 0.0384101f $X=3.535 $Y=0.36 $X2=0
+ $Y2=0
cc_439 N_A_510_74#_c_320_n N_VGND_c_1639_n 0.0211124f $X=2.94 $Y=0.36 $X2=0
+ $Y2=0
cc_440 N_A_510_74#_c_323_n N_VGND_c_1639_n 0.0496716f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_441 N_A_510_74#_c_404_p N_VGND_c_1639_n 0.0115893f $X=3.62 $Y=0.36 $X2=0
+ $Y2=0
cc_442 N_A_510_74#_c_317_n N_VGND_c_1640_n 0.00332223f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_443 N_A_510_74#_c_326_n N_VGND_c_1640_n 0.0548435f $X=6.365 $Y=0.34 $X2=0
+ $Y2=0
cc_444 N_A_510_74#_c_327_n N_VGND_c_1640_n 0.0116199f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_445 N_A_510_74#_c_317_n N_VGND_c_1643_n 0.00477801f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_446 N_A_510_74#_c_319_n N_VGND_c_1643_n 0.0199841f $X=3.535 $Y=0.36 $X2=0
+ $Y2=0
cc_447 N_A_510_74#_c_320_n N_VGND_c_1643_n 0.0114232f $X=2.94 $Y=0.36 $X2=0
+ $Y2=0
cc_448 N_A_510_74#_c_323_n N_VGND_c_1643_n 0.025617f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_449 N_A_510_74#_c_344_p N_VGND_c_1643_n 0.0237285f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_450 N_A_510_74#_c_326_n N_VGND_c_1643_n 0.0291469f $X=6.365 $Y=0.34 $X2=0
+ $Y2=0
cc_451 N_A_510_74#_c_327_n N_VGND_c_1643_n 0.00583764f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_452 N_A_510_74#_c_404_p N_VGND_c_1643_n 0.00583135f $X=3.62 $Y=0.36 $X2=0
+ $Y2=0
cc_453 N_A_510_74#_c_345_p A_850_119# 0.00155242f $X=4.465 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_454 N_A_510_74#_c_344_p A_922_119# 0.00179164f $X=5.525 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_455 N_A_856_294#_M1005_g N_RESET_B_c_608_n 0.0108881f $X=4.4 $Y=2.495 $X2=0
+ $Y2=0
cc_456 N_A_856_294#_M1016_g N_RESET_B_M1009_g 0.0419483f $X=4.535 $Y=0.805 $X2=0
+ $Y2=0
cc_457 N_A_856_294#_c_502_n N_RESET_B_M1009_g 0.0119822f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_458 N_A_856_294#_c_507_n N_RESET_B_M1009_g 5.70855e-19 $X=4.445 $Y=1.47 $X2=0
+ $Y2=0
cc_459 N_A_856_294#_M1005_g N_RESET_B_M1018_g 0.0245463f $X=4.4 $Y=2.495 $X2=0
+ $Y2=0
cc_460 N_A_856_294#_c_502_n N_RESET_B_c_596_n 0.00880086f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_461 N_A_856_294#_c_505_n N_RESET_B_c_596_n 0.0277148f $X=4.445 $Y=1.635 $X2=0
+ $Y2=0
cc_462 N_A_856_294#_c_506_n N_RESET_B_c_596_n 0.0013891f $X=4.445 $Y=1.635 $X2=0
+ $Y2=0
cc_463 N_A_856_294#_c_502_n N_RESET_B_c_598_n 0.014851f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_464 N_A_856_294#_c_540_p N_RESET_B_c_598_n 0.00468242f $X=6.03 $Y=1.215 $X2=0
+ $Y2=0
cc_465 N_A_856_294#_c_541_p N_RESET_B_c_598_n 0.00919057f $X=6.11 $Y=2.135 $X2=0
+ $Y2=0
cc_466 N_A_856_294#_c_508_n N_RESET_B_c_598_n 0.0226321f $X=6.282 $Y=1.97 $X2=0
+ $Y2=0
cc_467 N_A_856_294#_c_502_n N_RESET_B_c_599_n 0.00289579f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_468 N_A_856_294#_c_505_n N_RESET_B_c_599_n 5.41012e-19 $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_469 N_A_856_294#_c_502_n N_RESET_B_c_603_n 0.0041539f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_470 N_A_856_294#_c_505_n N_RESET_B_c_603_n 0.00108349f $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_471 N_A_856_294#_c_506_n N_RESET_B_c_603_n 0.0419483f $X=4.445 $Y=1.635 $X2=0
+ $Y2=0
cc_472 N_A_856_294#_c_502_n N_RESET_B_c_604_n 0.0227858f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_473 N_A_856_294#_c_505_n N_RESET_B_c_604_n 0.0186562f $X=4.445 $Y=1.635 $X2=0
+ $Y2=0
cc_474 N_A_856_294#_c_506_n N_RESET_B_c_604_n 0.00112856f $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_475 N_A_856_294#_c_502_n N_A_714_119#_M1020_g 0.0134843f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_476 N_A_856_294#_c_504_n N_A_714_119#_M1020_g 0.011387f $X=6.03 $Y=0.76 $X2=0
+ $Y2=0
cc_477 N_A_856_294#_c_540_p N_A_714_119#_M1020_g 3.84191e-19 $X=6.03 $Y=1.215
+ $X2=0 $Y2=0
cc_478 N_A_856_294#_c_508_n N_A_714_119#_M1020_g 0.00824116f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_479 N_A_856_294#_c_510_n N_A_714_119#_M1000_g 4.94098e-19 $X=6.11 $Y=2.815
+ $X2=0 $Y2=0
cc_480 N_A_856_294#_c_541_p N_A_714_119#_M1000_g 0.00819794f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_481 N_A_856_294#_c_508_n N_A_714_119#_M1000_g 0.00561622f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_482 N_A_856_294#_c_502_n N_A_714_119#_c_809_n 0.00228823f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_483 N_A_856_294#_c_508_n N_A_714_119#_c_810_n 0.00997795f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_484 N_A_856_294#_M1016_g N_A_714_119#_c_826_n 2.5148e-19 $X=4.535 $Y=0.805
+ $X2=0 $Y2=0
cc_485 N_A_856_294#_M1005_g N_A_714_119#_c_811_n 0.00140573f $X=4.4 $Y=2.495
+ $X2=0 $Y2=0
cc_486 N_A_856_294#_M1016_g N_A_714_119#_c_811_n 0.00105532f $X=4.535 $Y=0.805
+ $X2=0 $Y2=0
cc_487 N_A_856_294#_c_503_n N_A_714_119#_c_811_n 0.00816185f $X=4.61 $Y=1.215
+ $X2=0 $Y2=0
cc_488 N_A_856_294#_c_505_n N_A_714_119#_c_811_n 0.0175333f $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_489 N_A_856_294#_c_506_n N_A_714_119#_c_811_n 0.0011032f $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_490 N_A_856_294#_c_507_n N_A_714_119#_c_811_n 0.00697204f $X=4.445 $Y=1.47
+ $X2=0 $Y2=0
cc_491 N_A_856_294#_M1005_g N_A_714_119#_c_818_n 0.017034f $X=4.4 $Y=2.495 $X2=0
+ $Y2=0
cc_492 N_A_856_294#_c_505_n N_A_714_119#_c_818_n 0.018171f $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_493 N_A_856_294#_c_506_n N_A_714_119#_c_818_n 9.78234e-19 $X=4.445 $Y=1.635
+ $X2=0 $Y2=0
cc_494 N_A_856_294#_M1005_g N_A_714_119#_c_819_n 0.00217523f $X=4.4 $Y=2.495
+ $X2=0 $Y2=0
cc_495 N_A_856_294#_M1005_g N_A_714_119#_c_820_n 7.08937e-19 $X=4.4 $Y=2.495
+ $X2=0 $Y2=0
cc_496 N_A_856_294#_c_541_p N_A_714_119#_c_821_n 0.0103534f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_497 N_A_856_294#_c_502_n N_A_714_119#_c_812_n 0.0234898f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_498 N_A_856_294#_c_508_n N_A_714_119#_c_812_n 0.0399257f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_499 N_A_856_294#_M1016_g N_A_714_119#_c_813_n 5.79331e-19 $X=4.535 $Y=0.805
+ $X2=0 $Y2=0
cc_500 N_A_856_294#_M1016_g N_A_300_347#_M1019_g 0.0424852f $X=4.535 $Y=0.805
+ $X2=0 $Y2=0
cc_501 N_A_856_294#_c_503_n N_A_300_347#_M1019_g 4.71906e-19 $X=4.61 $Y=1.215
+ $X2=0 $Y2=0
cc_502 N_A_856_294#_M1016_g N_A_300_347#_c_920_n 0.00998561f $X=4.535 $Y=0.805
+ $X2=0 $Y2=0
cc_503 N_A_856_294#_c_504_n N_A_300_347#_M1007_g 0.00547135f $X=6.03 $Y=0.76
+ $X2=0 $Y2=0
cc_504 N_A_856_294#_c_540_p N_A_300_347#_M1007_g 0.00198105f $X=6.03 $Y=1.215
+ $X2=0 $Y2=0
cc_505 N_A_856_294#_c_508_n N_A_300_347#_M1007_g 0.00421803f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_506 N_A_856_294#_c_541_p N_A_300_347#_c_923_n 0.0128981f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_507 N_A_856_294#_c_541_p N_A_300_347#_c_926_n 0.0229541f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_508 N_A_856_294#_c_508_n N_A_300_347#_c_926_n 0.0236964f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_509 N_A_856_294#_c_541_p N_A_300_347#_c_927_n 0.00343033f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_510 N_A_856_294#_M1005_g N_VPWR_c_1392_n 0.00396188f $X=4.4 $Y=2.495 $X2=0
+ $Y2=0
cc_511 N_A_856_294#_c_510_n N_VPWR_c_1394_n 0.0241513f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_512 N_A_856_294#_c_510_n N_VPWR_c_1398_n 0.0315916f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_513 N_A_856_294#_M1005_g N_VPWR_c_1387_n 0.00113998f $X=4.4 $Y=2.495 $X2=0
+ $Y2=0
cc_514 N_A_856_294#_c_510_n N_VPWR_c_1387_n 0.0261488f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_515 N_A_856_294#_c_502_n N_VGND_M1009_d 0.00417413f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_516 N_A_856_294#_M1016_g N_VGND_c_1643_n 9.07931e-19 $X=4.535 $Y=0.805 $X2=0
+ $Y2=0
cc_517 N_RESET_B_c_598_n N_A_714_119#_c_809_n 0.00272004f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_599_n N_A_714_119#_c_809_n 0.00140145f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_519 N_RESET_B_c_603_n N_A_714_119#_c_809_n 0.0214999f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_520 N_RESET_B_c_604_n N_A_714_119#_c_809_n 0.00169603f $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_521 N_RESET_B_c_598_n N_A_714_119#_c_810_n 0.00619558f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_596_n N_A_714_119#_c_811_n 0.0244744f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_523 N_RESET_B_M1018_g N_A_714_119#_c_818_n 0.0149606f $X=4.91 $Y=2.495 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_596_n N_A_714_119#_c_818_n 0.0198957f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_525 N_RESET_B_c_599_n N_A_714_119#_c_818_n 0.00176425f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_604_n N_A_714_119#_c_818_n 0.017712f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_527 N_RESET_B_c_608_n N_A_714_119#_c_819_n 0.0049782f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_528 N_RESET_B_c_596_n N_A_714_119#_c_819_n 0.00779596f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_RESET_B_M1018_g N_A_714_119#_c_820_n 0.0092892f $X=4.91 $Y=2.495 $X2=0
+ $Y2=0
cc_530 N_RESET_B_M1018_g N_A_714_119#_c_821_n 0.00433193f $X=4.91 $Y=2.495 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_598_n N_A_714_119#_c_821_n 0.0084368f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_532 N_RESET_B_c_599_n N_A_714_119#_c_821_n 0.00133381f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_603_n N_A_714_119#_c_821_n 0.00325305f $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_534 N_RESET_B_M1018_g N_A_714_119#_c_812_n 0.00674835f $X=4.91 $Y=2.495 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_598_n N_A_714_119#_c_812_n 0.0166072f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_536 N_RESET_B_c_599_n N_A_714_119#_c_812_n 0.00259167f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_RESET_B_c_603_n N_A_714_119#_c_812_n 5.08278e-19 $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_604_n N_A_714_119#_c_812_n 0.0191898f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_539 N_RESET_B_c_596_n N_A_714_119#_c_813_n 0.00233951f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_RESET_B_c_596_n N_A_300_347#_M1017_s 0.00243377f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_RESET_B_c_608_n N_A_300_347#_c_928_n 0.0121828f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_596_n N_A_300_347#_c_928_n 0.00356343f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_RESET_B_c_596_n N_A_300_347#_c_929_n 0.00533875f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_RESET_B_c_596_n N_A_300_347#_c_918_n 0.0164105f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_545 N_RESET_B_c_608_n N_A_300_347#_M1012_g 0.01074f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_596_n N_A_300_347#_M1019_g 0.00362894f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_RESET_B_M1009_g N_A_300_347#_c_920_n 0.00999433f $X=4.895 $Y=0.805
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_598_n N_A_300_347#_c_933_n 2.3419e-19 $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_549 N_RESET_B_M1031_g N_A_300_347#_c_944_n 0.00570626f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_596_n N_A_300_347#_c_944_n 0.0248592f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_596_n N_A_300_347#_c_948_n 0.0077618f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_552 N_RESET_B_M1024_g N_A_300_347#_c_949_n 0.00558603f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_596_n N_A_300_347#_c_949_n 0.00353251f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_RESET_B_c_596_n N_A_300_347#_c_934_n 0.0279904f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_598_n N_A_300_347#_c_923_n 0.0603286f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_598_n N_A_300_347#_c_937_n 0.00727375f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_RESET_B_c_596_n N_A_300_347#_c_924_n 0.00384355f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_598_n N_A_300_347#_c_926_n 0.0194318f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_598_n N_A_300_347#_c_927_n 0.00169661f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_560 N_RESET_B_M1010_g N_A_1598_93#_M1002_g 0.0206165f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_561 N_RESET_B_M1015_g N_A_1598_93#_M1002_g 0.0068596f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_598_n N_A_1598_93#_M1002_g 0.00903792f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_600_n N_A_1598_93#_M1002_g 0.00140024f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_601_n N_A_1598_93#_M1002_g 0.00248623f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_605_n N_A_1598_93#_M1002_g 0.0174849f $X=8.545 $Y=1.63 $X2=0
+ $Y2=0
cc_566 N_RESET_B_M1015_g N_A_1598_93#_M1008_g 0.0159607f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_567 N_RESET_B_M1015_g N_A_1598_93#_c_1111_n 0.0180187f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_598_n N_A_1598_93#_c_1111_n 0.00534563f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_600_n N_A_1598_93#_c_1111_n 0.00307024f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_570 N_RESET_B_c_601_n N_A_1598_93#_c_1111_n 0.0292669f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_605_n N_A_1598_93#_c_1111_n 0.00342754f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_572 N_RESET_B_M1015_g N_A_1598_93#_c_1112_n 0.0213501f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_601_n N_A_1598_93#_c_1112_n 2.32727e-19 $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_574 N_RESET_B_M1015_g N_A_1598_93#_c_1113_n 0.0125991f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_575 N_RESET_B_M1015_g N_A_1598_93#_c_1107_n 2.15799e-19 $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_576 N_RESET_B_c_605_n N_A_1598_93#_c_1107_n 0.00106075f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_577 N_RESET_B_M1015_g N_A_1598_93#_c_1116_n 0.00567658f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_601_n N_A_1598_93#_c_1116_n 0.00239474f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_579 N_RESET_B_M1010_g N_A_1598_93#_c_1108_n 0.00117144f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_580 N_RESET_B_M1010_g N_A_1266_119#_c_1194_n 0.0535388f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_581 N_RESET_B_M1015_g N_A_1266_119#_c_1195_n 0.0442479f $X=8.62 $Y=2.75 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_598_n N_A_1266_119#_c_1200_n 0.0245011f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_600_n N_A_1266_119#_c_1200_n 0.00232289f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_601_n N_A_1266_119#_c_1200_n 0.0115131f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_585 N_RESET_B_M1010_g N_A_1266_119#_c_1201_n 0.0144298f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_586 N_RESET_B_c_598_n N_A_1266_119#_c_1201_n 0.0108617f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_600_n N_A_1266_119#_c_1201_n 0.0025054f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_601_n N_A_1266_119#_c_1201_n 0.0302597f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_605_n N_A_1266_119#_c_1201_n 0.0041539f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_590 N_RESET_B_M1010_g N_A_1266_119#_c_1202_n 0.00109666f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_600_n N_A_1266_119#_c_1202_n 0.00111187f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_592 N_RESET_B_c_601_n N_A_1266_119#_c_1202_n 0.0199249f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_605_n N_A_1266_119#_c_1202_n 4.14158e-19 $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_601_n N_A_1266_119#_c_1203_n 0.0011399f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_595 N_RESET_B_c_605_n N_A_1266_119#_c_1203_n 0.0207482f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_596 N_RESET_B_c_596_n N_VPWR_M1017_d 0.00118222f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1031_g N_VPWR_c_1389_n 5.11614e-19 $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_598 N_RESET_B_c_609_n N_VPWR_c_1389_n 0.00183649f $X=1.04 $Y=3.15 $X2=0 $Y2=0
cc_599 N_RESET_B_M1031_g N_VPWR_c_1390_n 0.00383385f $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_600 N_RESET_B_c_608_n N_VPWR_c_1390_n 0.0216652f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_601 N_RESET_B_c_608_n N_VPWR_c_1391_n 0.0249582f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_602 N_RESET_B_c_608_n N_VPWR_c_1392_n 0.0222942f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_603 N_RESET_B_M1018_g N_VPWR_c_1392_n 0.0101094f $X=4.91 $Y=2.495 $X2=0 $Y2=0
cc_604 N_RESET_B_c_608_n N_VPWR_c_1393_n 0.00690969f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_605 N_RESET_B_M1018_g N_VPWR_c_1394_n 0.00890396f $X=4.91 $Y=2.495 $X2=0
+ $Y2=0
cc_606 N_RESET_B_M1015_g N_VPWR_c_1395_n 0.00733882f $X=8.62 $Y=2.75 $X2=0 $Y2=0
cc_607 N_RESET_B_c_609_n N_VPWR_c_1402_n 0.00736275f $X=1.04 $Y=3.15 $X2=0 $Y2=0
cc_608 N_RESET_B_c_608_n N_VPWR_c_1403_n 0.0230851f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_609 N_RESET_B_c_608_n N_VPWR_c_1404_n 0.0670325f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_610 N_RESET_B_M1015_g N_VPWR_c_1405_n 0.005209f $X=8.62 $Y=2.75 $X2=0 $Y2=0
cc_611 N_RESET_B_c_608_n N_VPWR_c_1387_n 0.12854f $X=4.82 $Y=3.15 $X2=0 $Y2=0
cc_612 N_RESET_B_c_609_n N_VPWR_c_1387_n 0.0121254f $X=1.04 $Y=3.15 $X2=0 $Y2=0
cc_613 N_RESET_B_M1015_g N_VPWR_c_1387_n 0.00983503f $X=8.62 $Y=2.75 $X2=0 $Y2=0
cc_614 N_RESET_B_M1024_g N_A_33_74#_c_1515_n 0.0120626f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_615 N_RESET_B_M1031_g N_A_33_74#_c_1515_n 0.00946659f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_597_n N_A_33_74#_c_1515_n 0.00111707f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_617 N_RESET_B_c_602_n N_A_33_74#_c_1515_n 0.00281219f $X=0.965 $Y=1.515 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_606_n N_A_33_74#_c_1515_n 0.0317711f $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_619 N_RESET_B_M1031_g N_A_33_74#_c_1519_n 0.0144943f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_620 N_RESET_B_M1031_g N_A_33_74#_c_1520_n 0.0175722f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_608_n N_A_33_74#_c_1520_n 0.0208063f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_596_n N_A_33_74#_c_1520_n 0.0183296f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_597_n N_A_33_74#_c_1520_n 0.00783911f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_624 N_RESET_B_c_602_n N_A_33_74#_c_1520_n 4.48841e-19 $X=0.965 $Y=1.515 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_606_n N_A_33_74#_c_1520_n 0.0127944f $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_626 N_RESET_B_c_596_n N_A_33_74#_c_1516_n 0.0272381f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_596_n N_A_33_74#_c_1522_n 0.00386488f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_628 N_RESET_B_c_608_n N_A_33_74#_c_1524_n 0.00508475f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_629 N_RESET_B_M1024_g N_A_33_74#_c_1517_n 0.00390091f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_630 N_RESET_B_M1031_g N_A_33_74#_c_1525_n 0.00402616f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_602_n N_A_33_74#_c_1525_n 0.00194221f $X=0.965 $Y=1.515 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_606_n N_A_33_74#_c_1525_n 4.07355e-19 $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_608_n N_A_33_74#_c_1526_n 0.00130391f $X=4.82 $Y=3.15 $X2=0
+ $Y2=0
cc_634 N_RESET_B_M1024_g N_VGND_c_1631_n 0.00587764f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_602_n N_VGND_c_1631_n 0.00152642f $X=0.965 $Y=1.515 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_606_n N_VGND_c_1631_n 0.0076285f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_637 N_RESET_B_M1009_g N_VGND_c_1633_n 0.00412761f $X=4.895 $Y=0.805 $X2=0
+ $Y2=0
cc_638 N_RESET_B_M1010_g N_VGND_c_1634_n 0.0103576f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_639 N_RESET_B_M1024_g N_VGND_c_1636_n 0.00461464f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_640 N_RESET_B_M1010_g N_VGND_c_1641_n 0.0035863f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_641 N_RESET_B_M1024_g N_VGND_c_1643_n 0.00913041f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_642 N_RESET_B_M1009_g N_VGND_c_1643_n 9.39239e-19 $X=4.895 $Y=0.805 $X2=0
+ $Y2=0
cc_643 N_RESET_B_M1010_g N_VGND_c_1643_n 0.00401353f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_644 N_A_714_119#_c_811_n N_A_300_347#_c_929_n 0.00199243f $X=3.965 $Y=2.02
+ $X2=0 $Y2=0
cc_645 N_A_714_119#_c_819_n N_A_300_347#_M1012_g 0.00899443f $X=4.055 $Y=2.105
+ $X2=0 $Y2=0
cc_646 N_A_714_119#_c_826_n N_A_300_347#_M1019_g 0.00380092f $X=3.96 $Y=0.855
+ $X2=0 $Y2=0
cc_647 N_A_714_119#_c_811_n N_A_300_347#_M1019_g 0.0022166f $X=3.965 $Y=2.02
+ $X2=0 $Y2=0
cc_648 N_A_714_119#_c_813_n N_A_300_347#_M1019_g 0.0033507f $X=4 $Y=1.075 $X2=0
+ $Y2=0
cc_649 N_A_714_119#_M1020_g N_A_300_347#_c_920_n 0.00882199f $X=5.815 $Y=0.965
+ $X2=0 $Y2=0
cc_650 N_A_714_119#_M1020_g N_A_300_347#_M1007_g 0.0106687f $X=5.815 $Y=0.965
+ $X2=0 $Y2=0
cc_651 N_A_714_119#_c_810_n N_A_300_347#_c_926_n 4.20447e-19 $X=5.855 $Y=1.635
+ $X2=0 $Y2=0
cc_652 N_A_714_119#_c_810_n N_A_300_347#_c_927_n 0.0214083f $X=5.855 $Y=1.635
+ $X2=0 $Y2=0
cc_653 N_A_714_119#_c_821_n N_VPWR_M1000_s 0.00508213f $X=5.53 $Y=2.02 $X2=0
+ $Y2=0
cc_654 N_A_714_119#_c_812_n N_VPWR_M1000_s 0.00133211f $X=5.53 $Y=1.635 $X2=0
+ $Y2=0
cc_655 N_A_714_119#_c_818_n N_VPWR_c_1392_n 0.0220954f $X=4.99 $Y=2.105 $X2=0
+ $Y2=0
cc_656 N_A_714_119#_c_819_n N_VPWR_c_1392_n 0.013467f $X=4.055 $Y=2.105 $X2=0
+ $Y2=0
cc_657 N_A_714_119#_c_820_n N_VPWR_c_1392_n 0.0265512f $X=5.135 $Y=2.495 $X2=0
+ $Y2=0
cc_658 N_A_714_119#_c_820_n N_VPWR_c_1393_n 0.00544596f $X=5.135 $Y=2.495 $X2=0
+ $Y2=0
cc_659 N_A_714_119#_M1000_g N_VPWR_c_1394_n 0.0166809f $X=5.88 $Y=2.46 $X2=0
+ $Y2=0
cc_660 N_A_714_119#_c_809_n N_VPWR_c_1394_n 0.00202602f $X=5.74 $Y=1.635 $X2=0
+ $Y2=0
cc_661 N_A_714_119#_c_820_n N_VPWR_c_1394_n 0.0264407f $X=5.135 $Y=2.495 $X2=0
+ $Y2=0
cc_662 N_A_714_119#_c_821_n N_VPWR_c_1394_n 0.0166816f $X=5.53 $Y=2.02 $X2=0
+ $Y2=0
cc_663 N_A_714_119#_M1000_g N_VPWR_c_1398_n 0.00460063f $X=5.88 $Y=2.46 $X2=0
+ $Y2=0
cc_664 N_A_714_119#_c_819_n N_VPWR_c_1404_n 0.00712978f $X=4.055 $Y=2.105 $X2=0
+ $Y2=0
cc_665 N_A_714_119#_M1000_g N_VPWR_c_1387_n 0.00913687f $X=5.88 $Y=2.46 $X2=0
+ $Y2=0
cc_666 N_A_714_119#_c_819_n N_VPWR_c_1387_n 0.0112276f $X=4.055 $Y=2.105 $X2=0
+ $Y2=0
cc_667 N_A_714_119#_c_820_n N_VPWR_c_1387_n 0.00925037f $X=5.135 $Y=2.495 $X2=0
+ $Y2=0
cc_668 N_A_714_119#_c_811_n N_A_33_74#_c_1516_n 0.0050068f $X=3.965 $Y=2.02
+ $X2=0 $Y2=0
cc_669 N_A_714_119#_c_811_n N_A_33_74#_c_1522_n 0.00701119f $X=3.965 $Y=2.02
+ $X2=0 $Y2=0
cc_670 N_A_714_119#_c_819_n N_A_33_74#_c_1523_n 0.00730611f $X=4.055 $Y=2.105
+ $X2=0 $Y2=0
cc_671 N_A_714_119#_c_819_n N_A_33_74#_c_1526_n 0.00859596f $X=4.055 $Y=2.105
+ $X2=0 $Y2=0
cc_672 N_A_300_347#_c_937_n N_A_1598_93#_M1002_g 0.0139896f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_673 N_A_300_347#_c_933_n N_A_1598_93#_M1008_g 0.0373867f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_674 N_A_300_347#_c_933_n N_A_1598_93#_c_1112_n 0.0139896f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_675 N_A_300_347#_c_923_n N_A_1266_119#_c_1215_n 0.00277079f $X=7.31 $Y=1.715
+ $X2=0 $Y2=0
cc_676 N_A_300_347#_c_933_n N_A_1266_119#_c_1208_n 9.05598e-19 $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_677 N_A_300_347#_c_936_n N_A_1266_119#_c_1208_n 0.0103637f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_678 N_A_300_347#_c_932_n N_A_1266_119#_c_1200_n 0.00364552f $X=7.66 $Y=2.455
+ $X2=0 $Y2=0
cc_679 N_A_300_347#_c_933_n N_A_1266_119#_c_1200_n 0.00468398f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_680 N_A_300_347#_c_923_n N_A_1266_119#_c_1200_n 0.01265f $X=7.31 $Y=1.715
+ $X2=0 $Y2=0
cc_681 N_A_300_347#_c_936_n N_A_1266_119#_c_1200_n 0.0415019f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_682 N_A_300_347#_c_937_n N_A_1266_119#_c_1200_n 0.0057575f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_683 N_A_300_347#_c_932_n N_A_1266_119#_c_1210_n 0.0176328f $X=7.66 $Y=2.455
+ $X2=0 $Y2=0
cc_684 N_A_300_347#_c_933_n N_A_1266_119#_c_1210_n 0.00139404f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_685 N_A_300_347#_c_936_n N_A_1266_119#_c_1210_n 0.010457f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_686 N_A_300_347#_c_944_n N_VPWR_M1017_d 0.00570078f $X=2.145 $Y=1.915 $X2=0
+ $Y2=0
cc_687 N_A_300_347#_c_934_n N_VPWR_M1017_d 0.00100198f $X=2.27 $Y=1.82 $X2=0
+ $Y2=0
cc_688 N_A_300_347#_c_928_n N_VPWR_c_1391_n 0.00499467f $X=2.5 $Y=1.66 $X2=0
+ $Y2=0
cc_689 N_A_300_347#_c_932_n N_VPWR_c_1395_n 0.00170129f $X=7.66 $Y=2.455 $X2=0
+ $Y2=0
cc_690 N_A_300_347#_c_932_n N_VPWR_c_1398_n 0.00386291f $X=7.66 $Y=2.455 $X2=0
+ $Y2=0
cc_691 N_A_300_347#_c_928_n N_VPWR_c_1387_n 0.00112709f $X=2.5 $Y=1.66 $X2=0
+ $Y2=0
cc_692 N_A_300_347#_M1012_g N_VPWR_c_1387_n 0.00113998f $X=3.56 $Y=2.495 $X2=0
+ $Y2=0
cc_693 N_A_300_347#_c_932_n N_VPWR_c_1387_n 0.00487503f $X=7.66 $Y=2.455 $X2=0
+ $Y2=0
cc_694 N_A_300_347#_M1017_s N_A_33_74#_c_1520_n 0.0075606f $X=1.5 $Y=1.735 $X2=0
+ $Y2=0
cc_695 N_A_300_347#_c_928_n N_A_33_74#_c_1520_n 0.0191482f $X=2.5 $Y=1.66 $X2=0
+ $Y2=0
cc_696 N_A_300_347#_c_918_n N_A_33_74#_c_1520_n 0.00759259f $X=3.08 $Y=1.86
+ $X2=0 $Y2=0
cc_697 N_A_300_347#_c_944_n N_A_33_74#_c_1520_n 0.0520912f $X=2.145 $Y=1.915
+ $X2=0 $Y2=0
cc_698 N_A_300_347#_c_924_n N_A_33_74#_c_1520_n 0.00111175f $X=2.42 $Y=1.41
+ $X2=0 $Y2=0
cc_699 N_A_300_347#_c_915_n N_A_33_74#_c_1516_n 0.0115859f $X=3.005 $Y=1.21
+ $X2=0 $Y2=0
cc_700 N_A_300_347#_c_929_n N_A_33_74#_c_1516_n 0.00896882f $X=3.47 $Y=1.86
+ $X2=0 $Y2=0
cc_701 N_A_300_347#_c_929_n N_A_33_74#_c_1522_n 0.0142446f $X=3.47 $Y=1.86 $X2=0
+ $Y2=0
cc_702 N_A_300_347#_M1012_g N_A_33_74#_c_1522_n 0.00687826f $X=3.56 $Y=2.495
+ $X2=0 $Y2=0
cc_703 N_A_300_347#_c_928_n N_A_33_74#_c_1523_n 0.00319711f $X=2.5 $Y=1.66 $X2=0
+ $Y2=0
cc_704 N_A_300_347#_c_928_n N_A_33_74#_c_1524_n 0.007817f $X=2.5 $Y=1.66 $X2=0
+ $Y2=0
cc_705 N_A_300_347#_M1012_g N_A_33_74#_c_1526_n 0.00338156f $X=3.56 $Y=2.495
+ $X2=0 $Y2=0
cc_706 N_A_300_347#_c_948_n N_VGND_M1013_d 0.00507268f $X=2.145 $Y=0.91 $X2=0
+ $Y2=0
cc_707 N_A_300_347#_c_925_n N_VGND_M1013_d 0.00125792f $X=2.325 $Y=1.22 $X2=0
+ $Y2=0
cc_708 N_A_300_347#_c_947_n N_VGND_c_1631_n 0.0219699f $X=1.695 $Y=0.56 $X2=0
+ $Y2=0
cc_709 N_A_300_347#_c_914_n N_VGND_c_1632_n 0.00328045f $X=2.475 $Y=1.21 $X2=0
+ $Y2=0
cc_710 N_A_300_347#_c_917_n N_VGND_c_1632_n 0.00213439f $X=3.08 $Y=0.18 $X2=0
+ $Y2=0
cc_711 N_A_300_347#_c_918_n N_VGND_c_1632_n 3.48011e-19 $X=3.08 $Y=1.86 $X2=0
+ $Y2=0
cc_712 N_A_300_347#_c_948_n N_VGND_c_1632_n 0.0239919f $X=2.145 $Y=0.91 $X2=0
+ $Y2=0
cc_713 N_A_300_347#_c_920_n N_VGND_c_1633_n 0.0251635f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_714 N_A_300_347#_c_947_n N_VGND_c_1638_n 0.0111284f $X=1.695 $Y=0.56 $X2=0
+ $Y2=0
cc_715 N_A_300_347#_c_914_n N_VGND_c_1639_n 0.00461464f $X=2.475 $Y=1.21 $X2=0
+ $Y2=0
cc_716 N_A_300_347#_c_917_n N_VGND_c_1639_n 0.0527072f $X=3.08 $Y=0.18 $X2=0
+ $Y2=0
cc_717 N_A_300_347#_c_920_n N_VGND_c_1640_n 0.0230598f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_718 N_A_300_347#_c_914_n N_VGND_c_1643_n 0.00683632f $X=2.475 $Y=1.21 $X2=0
+ $Y2=0
cc_719 N_A_300_347#_c_916_n N_VGND_c_1643_n 0.0239744f $X=4.1 $Y=0.18 $X2=0
+ $Y2=0
cc_720 N_A_300_347#_c_917_n N_VGND_c_1643_n 0.00600144f $X=3.08 $Y=0.18 $X2=0
+ $Y2=0
cc_721 N_A_300_347#_c_920_n N_VGND_c_1643_n 0.0470713f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_722 N_A_300_347#_c_922_n N_VGND_c_1643_n 0.00370846f $X=4.175 $Y=0.18 $X2=0
+ $Y2=0
cc_723 N_A_300_347#_c_947_n N_VGND_c_1643_n 0.0118586f $X=1.695 $Y=0.56 $X2=0
+ $Y2=0
cc_724 N_A_300_347#_c_948_n N_VGND_c_1643_n 0.0102384f $X=2.145 $Y=0.91 $X2=0
+ $Y2=0
cc_725 N_A_1598_93#_c_1107_n N_A_1266_119#_c_1194_n 0.0048734f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_726 N_A_1598_93#_c_1108_n N_A_1266_119#_c_1194_n 0.00750942f $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_727 N_A_1598_93#_c_1114_n N_A_1266_119#_c_1195_n 0.00514416f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_728 N_A_1598_93#_c_1116_n N_A_1266_119#_c_1195_n 0.00291268f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_729 N_A_1598_93#_c_1113_n N_A_1266_119#_M1023_g 0.0131468f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_730 N_A_1598_93#_c_1114_n N_A_1266_119#_M1023_g 0.0076155f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_731 N_A_1598_93#_c_1116_n N_A_1266_119#_M1023_g 0.015254f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_732 N_A_1598_93#_c_1114_n N_A_1266_119#_c_1196_n 6.15368e-19 $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_733 N_A_1598_93#_c_1107_n N_A_1266_119#_c_1196_n 0.0128412f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_734 N_A_1598_93#_c_1108_n N_A_1266_119#_c_1196_n 8.36802e-19 $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_735 N_A_1598_93#_c_1114_n N_A_1266_119#_c_1206_n 0.0109475f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_736 N_A_1598_93#_c_1107_n N_A_1266_119#_c_1206_n 0.00680794f $X=9.475
+ $Y=1.965 $X2=0 $Y2=0
cc_737 N_A_1598_93#_c_1114_n N_A_1266_119#_c_1207_n 3.91389e-19 $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_738 N_A_1598_93#_c_1107_n N_A_1266_119#_c_1197_n 7.21124e-19 $X=9.475
+ $Y=1.965 $X2=0 $Y2=0
cc_739 N_A_1598_93#_c_1108_n N_A_1266_119#_c_1197_n 7.36949e-19 $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_740 N_A_1598_93#_c_1108_n N_A_1266_119#_c_1198_n 0.0071021f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_741 N_A_1598_93#_M1002_g N_A_1266_119#_c_1215_n 0.00369318f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_742 N_A_1598_93#_M1002_g N_A_1266_119#_c_1199_n 0.00375809f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_743 N_A_1598_93#_M1002_g N_A_1266_119#_c_1200_n 0.0212281f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_744 N_A_1598_93#_c_1111_n N_A_1266_119#_c_1200_n 0.0293641f $X=8.68 $Y=2.15
+ $X2=0 $Y2=0
cc_745 N_A_1598_93#_M1002_g N_A_1266_119#_c_1201_n 0.0157592f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_746 N_A_1598_93#_c_1111_n N_A_1266_119#_c_1201_n 0.0023008f $X=8.68 $Y=2.15
+ $X2=0 $Y2=0
cc_747 N_A_1598_93#_c_1116_n N_A_1266_119#_c_1201_n 0.00676946f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_748 N_A_1598_93#_M1008_g N_A_1266_119#_c_1210_n 0.00189255f $X=8.08 $Y=2.75
+ $X2=0 $Y2=0
cc_749 N_A_1598_93#_c_1114_n N_A_1266_119#_c_1202_n 0.0128235f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_750 N_A_1598_93#_c_1107_n N_A_1266_119#_c_1202_n 0.0502151f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_751 N_A_1598_93#_c_1116_n N_A_1266_119#_c_1202_n 0.0110236f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_752 N_A_1598_93#_c_1108_n N_A_1266_119#_c_1202_n 0.0121056f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_753 N_A_1598_93#_c_1107_n N_A_1266_119#_c_1203_n 0.0103445f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_754 N_A_1598_93#_c_1113_n N_A_1934_94#_c_1333_n 0.00532392f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_755 N_A_1598_93#_c_1116_n N_A_1934_94#_c_1333_n 9.63229e-19 $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_756 N_A_1598_93#_c_1107_n N_A_1934_94#_c_1326_n 0.0270211f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_757 N_A_1598_93#_c_1108_n N_A_1934_94#_c_1326_n 0.0315201f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_758 N_A_1598_93#_c_1114_n N_A_1934_94#_c_1327_n 0.0140451f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_759 N_A_1598_93#_c_1107_n N_A_1934_94#_c_1327_n 0.0238206f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_760 N_A_1598_93#_c_1107_n N_A_1934_94#_c_1330_n 0.0278717f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_761 N_A_1598_93#_M1008_g N_VPWR_c_1395_n 0.012757f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_762 N_A_1598_93#_c_1111_n N_VPWR_c_1395_n 0.0266609f $X=8.68 $Y=2.15 $X2=0
+ $Y2=0
cc_763 N_A_1598_93#_c_1112_n N_VPWR_c_1395_n 0.00346833f $X=8.155 $Y=2.17 $X2=0
+ $Y2=0
cc_764 N_A_1598_93#_c_1113_n N_VPWR_c_1395_n 0.030414f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_765 N_A_1598_93#_c_1113_n N_VPWR_c_1396_n 0.0165069f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_766 N_A_1598_93#_c_1114_n N_VPWR_c_1396_n 0.0121819f $X=9.39 $Y=2.05 $X2=0
+ $Y2=0
cc_767 N_A_1598_93#_M1008_g N_VPWR_c_1398_n 0.00460063f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_768 N_A_1598_93#_c_1113_n N_VPWR_c_1405_n 0.0144623f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_769 N_A_1598_93#_M1008_g N_VPWR_c_1387_n 0.00908371f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_770 N_A_1598_93#_c_1113_n N_VPWR_c_1387_n 0.0118344f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_771 N_A_1598_93#_M1002_g N_VGND_c_1634_n 0.00889071f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_772 N_A_1598_93#_c_1108_n N_VGND_c_1634_n 0.0110474f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_773 N_A_1598_93#_M1002_g N_VGND_c_1640_n 0.0035863f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_774 N_A_1598_93#_c_1108_n N_VGND_c_1641_n 0.0112924f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_775 N_A_1598_93#_M1002_g N_VGND_c_1643_n 0.00401353f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_776 N_A_1598_93#_c_1108_n N_VGND_c_1643_n 0.0158807f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_777 N_A_1266_119#_c_1206_n N_A_1934_94#_M1026_g 0.0160315f $X=9.95 $Y=1.97
+ $X2=0 $Y2=0
cc_778 N_A_1266_119#_M1023_g N_A_1934_94#_c_1333_n 0.00440747f $X=9.07 $Y=2.75
+ $X2=0 $Y2=0
cc_779 N_A_1266_119#_c_1206_n N_A_1934_94#_c_1333_n 0.00292339f $X=9.95 $Y=1.97
+ $X2=0 $Y2=0
cc_780 N_A_1266_119#_c_1207_n N_A_1934_94#_c_1333_n 0.00196172f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_781 N_A_1266_119#_c_1207_n N_A_1934_94#_c_1334_n 0.00942028f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_782 N_A_1266_119#_c_1194_n N_A_1934_94#_c_1326_n 0.00140435f $X=8.995
+ $Y=1.125 $X2=0 $Y2=0
cc_783 N_A_1266_119#_c_1196_n N_A_1934_94#_c_1326_n 0.0161335f $X=9.955 $Y=1.2
+ $X2=0 $Y2=0
cc_784 N_A_1266_119#_c_1197_n N_A_1934_94#_c_1326_n 0.010444f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_785 N_A_1266_119#_M1023_g N_A_1934_94#_c_1327_n 0.00438224f $X=9.07 $Y=2.75
+ $X2=0 $Y2=0
cc_786 N_A_1266_119#_c_1206_n N_A_1934_94#_c_1327_n 0.0163005f $X=9.95 $Y=1.97
+ $X2=0 $Y2=0
cc_787 N_A_1266_119#_c_1207_n N_A_1934_94#_c_1327_n 0.00477196f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_788 N_A_1266_119#_c_1196_n N_A_1934_94#_c_1328_n 0.00434645f $X=9.955 $Y=1.2
+ $X2=0 $Y2=0
cc_789 N_A_1266_119#_c_1206_n N_A_1934_94#_c_1328_n 0.00435182f $X=9.95 $Y=1.97
+ $X2=0 $Y2=0
cc_790 N_A_1266_119#_c_1197_n N_A_1934_94#_c_1331_n 0.0160558f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_791 N_A_1266_119#_c_1200_n N_VPWR_c_1395_n 8.41106e-19 $X=7.815 $Y=2.535
+ $X2=0 $Y2=0
cc_792 N_A_1266_119#_c_1210_n N_VPWR_c_1395_n 0.0157085f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_793 N_A_1266_119#_M1023_g N_VPWR_c_1396_n 0.00609057f $X=9.07 $Y=2.75 $X2=0
+ $Y2=0
cc_794 N_A_1266_119#_c_1206_n N_VPWR_c_1396_n 0.00128121f $X=9.95 $Y=1.97 $X2=0
+ $Y2=0
cc_795 N_A_1266_119#_c_1207_n N_VPWR_c_1396_n 0.00378352f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_796 N_A_1266_119#_c_1207_n N_VPWR_c_1397_n 0.0042237f $X=10.04 $Y=2.045 $X2=0
+ $Y2=0
cc_797 N_A_1266_119#_c_1208_n N_VPWR_c_1398_n 0.0149856f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_798 N_A_1266_119#_c_1210_n N_VPWR_c_1398_n 0.00880705f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_799 N_A_1266_119#_c_1207_n N_VPWR_c_1400_n 0.005209f $X=10.04 $Y=2.045 $X2=0
+ $Y2=0
cc_800 N_A_1266_119#_M1023_g N_VPWR_c_1405_n 0.005209f $X=9.07 $Y=2.75 $X2=0
+ $Y2=0
cc_801 N_A_1266_119#_M1023_g N_VPWR_c_1387_n 0.00987509f $X=9.07 $Y=2.75 $X2=0
+ $Y2=0
cc_802 N_A_1266_119#_c_1207_n N_VPWR_c_1387_n 0.00987336f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_803 N_A_1266_119#_c_1208_n N_VPWR_c_1387_n 0.0186508f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_804 N_A_1266_119#_c_1210_n N_VPWR_c_1387_n 0.0135253f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_805 N_A_1266_119#_c_1210_n A_1550_508# 0.00328986f $X=7.435 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_806 N_A_1266_119#_c_1196_n N_Q_c_1601_n 2.48707e-19 $X=9.955 $Y=1.2 $X2=0
+ $Y2=0
cc_807 N_A_1266_119#_c_1206_n Q 4.96875e-19 $X=9.95 $Y=1.97 $X2=0 $Y2=0
cc_808 N_A_1266_119#_c_1207_n Q 4.96875e-19 $X=10.04 $Y=2.045 $X2=0 $Y2=0
cc_809 N_A_1266_119#_c_1194_n N_VGND_c_1634_n 0.00147671f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_810 N_A_1266_119#_c_1215_n N_VGND_c_1634_n 0.0196844f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_811 N_A_1266_119#_c_1201_n N_VGND_c_1634_n 0.0254301f $X=8.92 $Y=1.21 $X2=0
+ $Y2=0
cc_812 N_A_1266_119#_c_1197_n N_VGND_c_1635_n 0.0072589f $X=10.03 $Y=1.125 $X2=0
+ $Y2=0
cc_813 N_A_1266_119#_c_1215_n N_VGND_c_1640_n 0.0212446f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_814 N_A_1266_119#_c_1194_n N_VGND_c_1641_n 0.00414396f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_815 N_A_1266_119#_c_1197_n N_VGND_c_1641_n 0.00486718f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_816 N_A_1266_119#_c_1194_n N_VGND_c_1643_n 0.00477801f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_817 N_A_1266_119#_c_1197_n N_VGND_c_1643_n 0.00514438f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_818 N_A_1266_119#_c_1215_n N_VGND_c_1643_n 0.0353228f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_819 N_A_1266_119#_c_1215_n A_1550_119# 0.00494929f $X=7.73 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_820 N_A_1266_119#_c_1199_n A_1550_119# 6.55526e-19 $X=7.815 $Y=1.125
+ $X2=-0.19 $Y2=-0.245
cc_821 N_A_1934_94#_c_1334_n N_VPWR_c_1396_n 0.034692f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_822 N_A_1934_94#_M1026_g N_VPWR_c_1397_n 0.00385682f $X=10.545 $Y=2.4 $X2=0
+ $Y2=0
cc_823 N_A_1934_94#_c_1327_n N_VPWR_c_1397_n 0.0341417f $X=9.815 $Y=2.27 $X2=0
+ $Y2=0
cc_824 N_A_1934_94#_c_1328_n N_VPWR_c_1397_n 0.0104191f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_825 N_A_1934_94#_c_1329_n N_VPWR_c_1397_n 0.00162988f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_826 N_A_1934_94#_c_1334_n N_VPWR_c_1400_n 0.0145471f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_827 N_A_1934_94#_M1026_g N_VPWR_c_1406_n 0.005209f $X=10.545 $Y=2.4 $X2=0
+ $Y2=0
cc_828 N_A_1934_94#_M1026_g N_VPWR_c_1387_n 0.00986694f $X=10.545 $Y=2.4 $X2=0
+ $Y2=0
cc_829 N_A_1934_94#_c_1334_n N_VPWR_c_1387_n 0.0119735f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_830 N_A_1934_94#_c_1331_n N_Q_c_1601_n 0.00640271f $X=10.48 $Y=1.32 $X2=0
+ $Y2=0
cc_831 N_A_1934_94#_c_1326_n N_Q_c_1602_n 5.13862e-19 $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_832 N_A_1934_94#_c_1328_n N_Q_c_1602_n 0.00188005f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_833 N_A_1934_94#_c_1331_n N_Q_c_1602_n 0.00241276f $X=10.48 $Y=1.32 $X2=0
+ $Y2=0
cc_834 N_A_1934_94#_M1026_g Q 0.00475543f $X=10.545 $Y=2.4 $X2=0 $Y2=0
cc_835 N_A_1934_94#_c_1327_n Q 0.00727657f $X=9.815 $Y=2.27 $X2=0 $Y2=0
cc_836 N_A_1934_94#_c_1328_n Q 7.18422e-19 $X=10.48 $Y=1.485 $X2=0 $Y2=0
cc_837 N_A_1934_94#_c_1329_n Q 3.0165e-19 $X=10.48 $Y=1.485 $X2=0 $Y2=0
cc_838 N_A_1934_94#_M1026_g Q 0.0144587f $X=10.545 $Y=2.4 $X2=0 $Y2=0
cc_839 N_A_1934_94#_M1026_g N_Q_c_1603_n 0.0042683f $X=10.545 $Y=2.4 $X2=0 $Y2=0
cc_840 N_A_1934_94#_c_1328_n N_Q_c_1603_n 0.0262114f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_841 N_A_1934_94#_c_1329_n N_Q_c_1603_n 0.00769124f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_842 N_A_1934_94#_c_1331_n N_Q_c_1603_n 0.0040915f $X=10.48 $Y=1.32 $X2=0
+ $Y2=0
cc_843 N_A_1934_94#_c_1326_n N_VGND_c_1635_n 0.024751f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_844 N_A_1934_94#_c_1328_n N_VGND_c_1635_n 0.0194281f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_845 N_A_1934_94#_c_1329_n N_VGND_c_1635_n 0.00216466f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_846 N_A_1934_94#_c_1331_n N_VGND_c_1635_n 0.00292117f $X=10.48 $Y=1.32 $X2=0
+ $Y2=0
cc_847 N_A_1934_94#_c_1326_n N_VGND_c_1641_n 0.00541117f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_848 N_A_1934_94#_c_1331_n N_VGND_c_1642_n 0.00485341f $X=10.48 $Y=1.32 $X2=0
+ $Y2=0
cc_849 N_A_1934_94#_c_1326_n N_VGND_c_1643_n 0.00809617f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_850 N_A_1934_94#_c_1331_n N_VGND_c_1643_n 0.00514438f $X=10.48 $Y=1.32 $X2=0
+ $Y2=0
cc_851 N_VPWR_c_1389_n N_A_33_74#_c_1519_n 0.0165069f $X=0.275 $Y=2.75 $X2=0
+ $Y2=0
cc_852 N_VPWR_c_1390_n N_A_33_74#_c_1519_n 0.016253f $X=1.18 $Y=2.75 $X2=0 $Y2=0
cc_853 N_VPWR_c_1402_n N_A_33_74#_c_1519_n 0.0109793f $X=1.06 $Y=3.33 $X2=0
+ $Y2=0
cc_854 N_VPWR_c_1387_n N_A_33_74#_c_1519_n 0.00901959f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_855 N_VPWR_M1017_d N_A_33_74#_c_1520_n 0.00629868f $X=2.005 $Y=1.735 $X2=0
+ $Y2=0
cc_856 N_VPWR_c_1390_n N_A_33_74#_c_1520_n 0.0259654f $X=1.18 $Y=2.75 $X2=0
+ $Y2=0
cc_857 N_VPWR_c_1391_n N_A_33_74#_c_1520_n 0.0239372f $X=2.21 $Y=2.635 $X2=0
+ $Y2=0
cc_858 N_VPWR_c_1404_n N_A_33_74#_c_1524_n 0.00504459f $X=4.49 $Y=3.33 $X2=0
+ $Y2=0
cc_859 N_VPWR_c_1387_n N_A_33_74#_c_1524_n 0.00713738f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_860 N_VPWR_c_1397_n Q 0.0293476f $X=10.315 $Y=2.265 $X2=0 $Y2=0
cc_861 N_VPWR_c_1406_n Q 0.0154414f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_862 N_VPWR_c_1387_n Q 0.0127129f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_863 N_A_33_74#_c_1517_n A_120_74# 0.00489958f $X=0.625 $Y=0.57 $X2=-0.19
+ $Y2=-0.245
cc_864 N_A_33_74#_c_1515_n N_VGND_c_1631_n 9.26454e-19 $X=0.625 $Y=2.18 $X2=0
+ $Y2=0
cc_865 N_A_33_74#_c_1517_n N_VGND_c_1631_n 0.0120498f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_866 N_A_33_74#_c_1517_n N_VGND_c_1636_n 0.0239076f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_867 N_A_33_74#_c_1517_n N_VGND_c_1643_n 0.0198316f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_868 N_Q_c_1601_n N_VGND_c_1635_n 0.0261897f $X=10.755 $Y=0.605 $X2=0 $Y2=0
cc_869 N_Q_c_1601_n N_VGND_c_1642_n 0.0118258f $X=10.755 $Y=0.605 $X2=0 $Y2=0
cc_870 N_Q_c_1601_n N_VGND_c_1643_n 0.0126447f $X=10.755 $Y=0.605 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__sdfrbp_1.pxi.spice
* Created: Wed Sep  2 12:30:12 2020
* 
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_27_74# N_A_27_74#_M1038_s N_A_27_74#_M1018_s
+ N_A_27_74#_c_289_n N_A_27_74#_M1023_g N_A_27_74#_M1030_g N_A_27_74#_c_290_n
+ N_A_27_74#_c_291_n N_A_27_74#_c_292_n N_A_27_74#_c_293_n N_A_27_74#_c_297_n
+ N_A_27_74#_c_294_n N_A_27_74#_c_298_n N_A_27_74#_c_299_n N_A_27_74#_c_300_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_27_74#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%SCE N_SCE_M1038_g N_SCE_M1018_g N_SCE_M1017_g
+ N_SCE_M1032_g N_SCE_c_369_n N_SCE_c_370_n N_SCE_c_371_n N_SCE_c_372_n
+ N_SCE_c_373_n N_SCE_c_374_n SCE SCE SCE N_SCE_c_375_n N_SCE_c_376_n
+ N_SCE_c_377_n N_SCE_c_378_n SCE N_SCE_c_379_n PM_SKY130_FD_SC_MS__SDFRBP_1%SCE
x_PM_SKY130_FD_SC_MS__SDFRBP_1%D N_D_M1002_g N_D_M1027_g D N_D_c_456_n
+ N_D_c_457_n N_D_c_458_n PM_SKY130_FD_SC_MS__SDFRBP_1%D
x_PM_SKY130_FD_SC_MS__SDFRBP_1%SCD N_SCD_c_496_n N_SCD_M1022_g N_SCD_c_500_n
+ N_SCD_M1001_g N_SCD_c_498_n SCD SCD PM_SKY130_FD_SC_MS__SDFRBP_1%SCD
x_PM_SKY130_FD_SC_MS__SDFRBP_1%CLK N_CLK_c_539_n N_CLK_M1013_g N_CLK_M1025_g
+ N_CLK_c_540_n N_CLK_c_541_n CLK N_CLK_c_542_n N_CLK_c_543_n N_CLK_c_544_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%CLK
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_1037_119# N_A_1037_119#_M1014_d
+ N_A_1037_119#_M1035_d N_A_1037_119#_M1019_g N_A_1037_119#_c_600_n
+ N_A_1037_119#_M1036_g N_A_1037_119#_c_602_n N_A_1037_119#_M1029_g
+ N_A_1037_119#_c_603_n N_A_1037_119#_c_604_n N_A_1037_119#_M1033_g
+ N_A_1037_119#_c_605_n N_A_1037_119#_c_606_n N_A_1037_119#_c_607_n
+ N_A_1037_119#_c_608_n N_A_1037_119#_c_609_n N_A_1037_119#_c_610_n
+ N_A_1037_119#_c_611_n N_A_1037_119#_c_639_p N_A_1037_119#_c_637_p
+ N_A_1037_119#_c_662_p N_A_1037_119#_c_612_n N_A_1037_119#_c_613_n
+ N_A_1037_119#_c_733_p N_A_1037_119#_c_614_n N_A_1037_119#_c_624_n
+ N_A_1037_119#_c_615_n N_A_1037_119#_c_616_n N_A_1037_119#_c_617_n
+ N_A_1037_119#_c_618_n N_A_1037_119#_c_619_n N_A_1037_119#_c_627_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_1037_119#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_1369_93# N_A_1369_93#_M1041_d
+ N_A_1369_93#_M1007_d N_A_1369_93#_M1004_g N_A_1369_93#_M1006_g
+ N_A_1369_93#_c_812_n N_A_1369_93#_c_813_n N_A_1369_93#_c_814_n
+ N_A_1369_93#_c_815_n N_A_1369_93#_c_836_n N_A_1369_93#_c_816_n
+ N_A_1369_93#_c_817_n N_A_1369_93#_c_818_n N_A_1369_93#_c_819_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_1369_93#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%RESET_B N_RESET_B_M1028_g N_RESET_B_c_913_n
+ N_RESET_B_M1011_g N_RESET_B_c_914_n N_RESET_B_c_915_n N_RESET_B_M1034_g
+ N_RESET_B_M1040_g N_RESET_B_c_917_n N_RESET_B_M1009_g N_RESET_B_M1020_g
+ N_RESET_B_c_919_n N_RESET_B_c_927_n N_RESET_B_c_920_n N_RESET_B_c_928_n
+ N_RESET_B_c_921_n N_RESET_B_c_929_n N_RESET_B_c_930_n N_RESET_B_c_931_n
+ N_RESET_B_c_932_n N_RESET_B_c_933_n N_RESET_B_c_934_n RESET_B
+ N_RESET_B_c_936_n N_RESET_B_c_937_n N_RESET_B_c_938_n N_RESET_B_c_939_n
+ N_RESET_B_c_940_n N_RESET_B_c_941_n N_RESET_B_c_922_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%RESET_B
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_1235_119# N_A_1235_119#_M1031_d
+ N_A_1235_119#_M1019_d N_A_1235_119#_M1040_d N_A_1235_119#_M1041_g
+ N_A_1235_119#_M1007_g N_A_1235_119#_c_1158_n N_A_1235_119#_c_1165_n
+ N_A_1235_119#_c_1159_n N_A_1235_119#_c_1189_n N_A_1235_119#_c_1160_n
+ N_A_1235_119#_c_1161_n N_A_1235_119#_c_1162_n N_A_1235_119#_c_1168_n
+ N_A_1235_119#_c_1163_n PM_SKY130_FD_SC_MS__SDFRBP_1%A_1235_119#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_819_119# N_A_819_119#_M1013_s
+ N_A_819_119#_M1025_s N_A_819_119#_M1035_g N_A_819_119#_M1014_g
+ N_A_819_119#_c_1268_n N_A_819_119#_c_1269_n N_A_819_119#_c_1270_n
+ N_A_819_119#_c_1271_n N_A_819_119#_c_1272_n N_A_819_119#_c_1283_n
+ N_A_819_119#_c_1284_n N_A_819_119#_c_1273_n N_A_819_119#_M1031_g
+ N_A_819_119#_M1024_g N_A_819_119#_c_1286_n N_A_819_119#_M1015_g
+ N_A_819_119#_c_1274_n N_A_819_119#_c_1275_n N_A_819_119#_M1016_g
+ N_A_819_119#_c_1277_n N_A_819_119#_c_1290_n N_A_819_119#_c_1296_n
+ N_A_819_119#_c_1299_n N_A_819_119#_c_1278_n N_A_819_119#_c_1291_n
+ N_A_819_119#_c_1305_n N_A_819_119#_c_1308_n N_A_819_119#_c_1279_n
+ N_A_819_119#_c_1280_n N_A_819_119#_c_1281_n N_A_819_119#_c_1294_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_819_119#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_2008_48# N_A_2008_48#_M1012_d
+ N_A_2008_48#_M1020_d N_A_2008_48#_M1005_g N_A_2008_48#_c_1459_n
+ N_A_2008_48#_M1039_g N_A_2008_48#_c_1460_n N_A_2008_48#_c_1468_n
+ N_A_2008_48#_c_1469_n N_A_2008_48#_c_1470_n N_A_2008_48#_c_1471_n
+ N_A_2008_48#_c_1461_n N_A_2008_48#_c_1472_n N_A_2008_48#_c_1462_n
+ N_A_2008_48#_c_1463_n N_A_2008_48#_c_1474_n N_A_2008_48#_c_1464_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_2008_48#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_1747_74# N_A_1747_74#_M1029_d
+ N_A_1747_74#_M1015_d N_A_1747_74#_c_1590_n N_A_1747_74#_M1012_g
+ N_A_1747_74#_c_1591_n N_A_1747_74#_c_1592_n N_A_1747_74#_M1021_g
+ N_A_1747_74#_M1026_g N_A_1747_74#_c_1593_n N_A_1747_74#_M1010_g
+ N_A_1747_74#_c_1594_n N_A_1747_74#_c_1595_n N_A_1747_74#_M1008_g
+ N_A_1747_74#_M1003_g N_A_1747_74#_c_1606_n N_A_1747_74#_c_1607_n
+ N_A_1747_74#_c_1597_n N_A_1747_74#_c_1615_n N_A_1747_74#_c_1619_n
+ N_A_1747_74#_c_1609_n N_A_1747_74#_c_1610_n N_A_1747_74#_c_1598_n
+ N_A_1747_74#_c_1599_n N_A_1747_74#_c_1600_n N_A_1747_74#_c_1601_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_1747_74#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_2513_424# N_A_2513_424#_M1003_s
+ N_A_2513_424#_M1008_s N_A_2513_424#_M1037_g N_A_2513_424#_M1000_g
+ N_A_2513_424#_c_1762_n N_A_2513_424#_c_1767_n N_A_2513_424#_c_1763_n
+ N_A_2513_424#_c_1764_n N_A_2513_424#_c_1765_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_2513_424#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%VPWR N_VPWR_M1018_d N_VPWR_M1001_d N_VPWR_M1025_d
+ N_VPWR_M1006_d N_VPWR_M1007_s N_VPWR_M1039_d N_VPWR_M1021_d N_VPWR_M1008_d
+ N_VPWR_c_1811_n N_VPWR_c_1812_n N_VPWR_c_1813_n N_VPWR_c_1814_n
+ N_VPWR_c_1815_n N_VPWR_c_1816_n N_VPWR_c_1817_n N_VPWR_c_1930_n
+ N_VPWR_c_1818_n N_VPWR_c_1819_n N_VPWR_c_1820_n N_VPWR_c_1821_n
+ N_VPWR_c_1822_n N_VPWR_c_1823_n N_VPWR_c_1824_n N_VPWR_c_1825_n VPWR
+ N_VPWR_c_1826_n N_VPWR_c_1827_n N_VPWR_c_1828_n N_VPWR_c_1829_n
+ N_VPWR_c_1830_n N_VPWR_c_1831_n N_VPWR_c_1810_n N_VPWR_c_1833_n
+ N_VPWR_c_1834_n N_VPWR_c_1835_n N_VPWR_c_1836_n N_VPWR_c_1837_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%VPWR
x_PM_SKY130_FD_SC_MS__SDFRBP_1%A_413_90# N_A_413_90#_M1002_d N_A_413_90#_M1031_s
+ N_A_413_90#_M1027_d N_A_413_90#_M1011_d N_A_413_90#_M1019_s
+ N_A_413_90#_c_2006_n N_A_413_90#_c_1991_n N_A_413_90#_c_1992_n
+ N_A_413_90#_c_1999_n N_A_413_90#_c_2000_n N_A_413_90#_c_1993_n
+ N_A_413_90#_c_2001_n N_A_413_90#_c_2002_n N_A_413_90#_c_1994_n
+ N_A_413_90#_c_1995_n N_A_413_90#_c_1996_n N_A_413_90#_c_2004_n
+ N_A_413_90#_c_1997_n N_A_413_90#_c_2005_n
+ PM_SKY130_FD_SC_MS__SDFRBP_1%A_413_90#
x_PM_SKY130_FD_SC_MS__SDFRBP_1%Q_N N_Q_N_M1010_d N_Q_N_M1026_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_MS__SDFRBP_1%Q_N
x_PM_SKY130_FD_SC_MS__SDFRBP_1%Q N_Q_M1037_d N_Q_M1000_d Q Q Q Q Q Q Q
+ N_Q_c_2160_n PM_SKY130_FD_SC_MS__SDFRBP_1%Q
x_PM_SKY130_FD_SC_MS__SDFRBP_1%VGND N_VGND_M1038_d N_VGND_M1028_d N_VGND_M1013_d
+ N_VGND_M1034_d N_VGND_M1005_d N_VGND_M1010_s N_VGND_M1003_d N_VGND_c_2179_n
+ N_VGND_c_2180_n N_VGND_c_2181_n N_VGND_c_2182_n N_VGND_c_2183_n
+ N_VGND_c_2184_n N_VGND_c_2185_n N_VGND_c_2186_n N_VGND_c_2187_n VGND
+ N_VGND_c_2188_n N_VGND_c_2189_n N_VGND_c_2190_n N_VGND_c_2191_n
+ N_VGND_c_2192_n N_VGND_c_2193_n N_VGND_c_2194_n N_VGND_c_2195_n
+ N_VGND_c_2196_n N_VGND_c_2197_n N_VGND_c_2198_n N_VGND_c_2199_n
+ N_VGND_c_2200_n PM_SKY130_FD_SC_MS__SDFRBP_1%VGND
x_PM_SKY130_FD_SC_MS__SDFRBP_1%noxref_25 N_noxref_25_M1023_s N_noxref_25_M1022_d
+ N_noxref_25_c_2317_n N_noxref_25_c_2318_n N_noxref_25_c_2319_n
+ N_noxref_25_c_2320_n PM_SKY130_FD_SC_MS__SDFRBP_1%noxref_25
cc_1 VNB N_A_27_74#_c_289_n 0.0213036f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_2 VNB N_A_27_74#_c_290_n 0.0280153f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_3 VNB N_A_27_74#_c_291_n 0.0167958f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_4 VNB N_A_27_74#_c_292_n 0.0201543f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_5 VNB N_A_27_74#_c_293_n 0.0460387f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_6 VNB N_A_27_74#_c_294_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.145
cc_7 VNB N_SCE_M1038_g 0.0718805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_369_n 0.00457743f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_9 VNB N_SCE_c_370_n 0.0146141f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_10 VNB N_SCE_c_371_n 0.00965144f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.145
cc_11 VNB N_SCE_c_372_n 0.0119481f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_12 VNB N_SCE_c_373_n 0.00486821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_374_n 0.0284582f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.135
cc_14 VNB N_SCE_c_375_n 0.0181262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_c_376_n 0.0212613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_c_377_n 0.00874037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_SCE_c_378_n 0.00943038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_c_379_n 0.001771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_M1027_g 0.0241855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_D_c_456_n 0.0346496f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_21 VNB N_D_c_457_n 0.0056581f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_22 VNB N_D_c_458_n 0.0173597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCD_c_496_n 0.0263396f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_24 VNB N_SCD_M1022_g 0.0268436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_SCD_c_498_n 0.00366688f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_26 VNB SCD 0.00359665f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.16
cc_27 VNB N_CLK_c_539_n 0.0224328f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_28 VNB N_CLK_c_540_n 0.00141289f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_29 VNB N_CLK_c_541_n 0.0208908f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.98
cc_30 VNB N_CLK_c_542_n 0.0321028f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_31 VNB N_CLK_c_543_n 0.0216785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_CLK_c_544_n 0.0152241f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.135
cc_33 VNB N_A_1037_119#_c_600_n 0.00999582f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_34 VNB N_A_1037_119#_M1036_g 0.0409203f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_35 VNB N_A_1037_119#_c_602_n 0.0165132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1037_119#_c_603_n 0.0213887f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.145
cc_37 VNB N_A_1037_119#_c_604_n 0.007535f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_38 VNB N_A_1037_119#_c_605_n 0.00402601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1037_119#_c_606_n 0.00279065f $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.512
cc_40 VNB N_A_1037_119#_c_607_n 9.17021e-19 $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.465
cc_41 VNB N_A_1037_119#_c_608_n 0.0376244f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_42 VNB N_A_1037_119#_c_609_n 0.00219004f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_43 VNB N_A_1037_119#_c_610_n 0.00216636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1037_119#_c_611_n 0.00427035f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.98
cc_45 VNB N_A_1037_119#_c_612_n 0.00867477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1037_119#_c_613_n 0.00224459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1037_119#_c_614_n 0.00269633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1037_119#_c_615_n 5.95258e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1037_119#_c_616_n 0.00830295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1037_119#_c_617_n 0.0326227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1037_119#_c_618_n 0.00544115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1037_119#_c_619_n 0.010383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1369_93#_M1004_g 0.0329059f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_54 VNB N_A_1369_93#_c_812_n 0.00499007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1369_93#_c_813_n 0.0240804f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_56 VNB N_A_1369_93#_c_814_n 0.00402144f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.145
cc_57 VNB N_A_1369_93#_c_815_n 6.59562e-19 $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_58 VNB N_A_1369_93#_c_816_n 0.00177944f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.145
cc_59 VNB N_A_1369_93#_c_817_n 0.00845443f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.512
cc_60 VNB N_A_1369_93#_c_818_n 0.00273128f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.512
cc_61 VNB N_A_1369_93#_c_819_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_62 VNB N_RESET_B_M1028_g 0.015554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_RESET_B_c_913_n 0.0265591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_c_914_n 0.280456f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_65 VNB N_RESET_B_c_915_n 0.012806f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_66 VNB N_RESET_B_M1034_g 0.0247097f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_67 VNB N_RESET_B_c_917_n 0.0201149f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_68 VNB N_RESET_B_M1009_g 0.0341606f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.135
cc_69 VNB N_RESET_B_c_919_n 0.0133529f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_70 VNB N_RESET_B_c_920_n 0.0317695f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_71 VNB N_RESET_B_c_921_n 0.0234009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_RESET_B_c_922_n 0.0158526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1235_119#_M1041_g 0.0263955f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_74 VNB N_A_1235_119#_c_1158_n 6.70206e-19 $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_75 VNB N_A_1235_119#_c_1159_n 0.0107155f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.145
cc_76 VNB N_A_1235_119#_c_1160_n 5.52581e-19 $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.465
cc_77 VNB N_A_1235_119#_c_1161_n 0.00253125f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_78 VNB N_A_1235_119#_c_1162_n 0.00399797f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_79 VNB N_A_1235_119#_c_1163_n 0.0424031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_819_119#_c_1268_n 0.00908898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_819_119#_c_1269_n 0.00777684f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_82 VNB N_A_819_119#_c_1270_n 0.00404916f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_83 VNB N_A_819_119#_c_1271_n 0.0300812f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_84 VNB N_A_819_119#_c_1272_n 0.010326f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.145
cc_85 VNB N_A_819_119#_c_1273_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_86 VNB N_A_819_119#_c_1274_n 0.0212572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_819_119#_c_1275_n 0.0048066f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.135
cc_88 VNB N_A_819_119#_M1016_g 0.0521391f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_89 VNB N_A_819_119#_c_1277_n 0.00788042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_819_119#_c_1278_n 0.00164026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_819_119#_c_1279_n 0.00177279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_819_119#_c_1280_n 0.0177782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_819_119#_c_1281_n 0.0156093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2008_48#_M1005_g 0.0424527f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_95 VNB N_A_2008_48#_c_1459_n 0.0184816f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_96 VNB N_A_2008_48#_c_1460_n 0.00245359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2008_48#_c_1461_n 0.00907094f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.512
cc_98 VNB N_A_2008_48#_c_1462_n 6.5078e-19 $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.465
cc_99 VNB N_A_2008_48#_c_1463_n 0.00160142f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_100 VNB N_A_2008_48#_c_1464_n 0.00658078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1747_74#_c_1590_n 0.0180751f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.98
cc_102 VNB N_A_1747_74#_c_1591_n 0.031848f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.16
cc_103 VNB N_A_1747_74#_c_1592_n 0.0157622f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_104 VNB N_A_1747_74#_c_1593_n 0.0240396f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_105 VNB N_A_1747_74#_c_1594_n 0.0485708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1747_74#_c_1595_n 0.0663652f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=2.135
cc_107 VNB N_A_1747_74#_M1003_g 0.0405544f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_108 VNB N_A_1747_74#_c_1597_n 0.00927852f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.98
cc_109 VNB N_A_1747_74#_c_1598_n 0.00249714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1747_74#_c_1599_n 0.00130137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1747_74#_c_1600_n 0.0147798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1747_74#_c_1601_n 0.020816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2513_424#_M1037_g 0.0280908f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.66
cc_114 VNB N_A_2513_424#_M1000_g 0.00182328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2513_424#_c_1762_n 0.0126466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2513_424#_c_1763_n 0.00835153f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=2.135
cc_117 VNB N_A_2513_424#_c_1764_n 0.0333398f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.135
cc_118 VNB N_A_2513_424#_c_1765_n 4.48326e-19 $X=-0.19 $Y=-0.245 $X2=0.2
+ $Y2=2.512
cc_119 VNB N_VPWR_c_1810_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_413_90#_c_1991_n 0.0242946f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.145
cc_121 VNB N_A_413_90#_c_1992_n 0.00670543f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_122 VNB N_A_413_90#_c_1993_n 0.00242544f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_123 VNB N_A_413_90#_c_1994_n 0.00586596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_413_90#_c_1995_n 0.00197652f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=2.135
cc_125 VNB N_A_413_90#_c_1996_n 0.0057856f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_126 VNB N_A_413_90#_c_1997_n 0.00377909f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=2.16
cc_127 VNB Q_N 0.0123064f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_128 VNB Q 0.0267037f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_129 VNB Q 0.0127641f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.16
cc_130 VNB N_Q_c_2160_n 0.0251085f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=2.16
cc_131 VNB N_VGND_c_2179_n 0.0135998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2180_n 0.0137162f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.512
cc_133 VNB N_VGND_c_2181_n 0.0126266f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.512
cc_134 VNB N_VGND_c_2182_n 0.0079764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2183_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_136 VNB N_VGND_c_2184_n 0.0363017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2185_n 0.0097163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2186_n 0.0218665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2187_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2188_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2189_n 0.0628724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2190_n 0.0567011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2191_n 0.0609299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2192_n 0.0284194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2193_n 0.0193554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2194_n 0.728438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2195_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2196_n 0.00406166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2197_n 0.00631189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2198_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2199_n 0.0153005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2200_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_noxref_25_c_2317_n 0.00380385f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.66
cc_154 VNB N_noxref_25_c_2318_n 0.0295571f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_155 VNB N_noxref_25_c_2319_n 0.00398497f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_156 VNB N_noxref_25_c_2320_n 0.00452409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VPB N_A_27_74#_M1030_g 0.0223046f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_158 VPB N_A_27_74#_c_291_n 0.0237442f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_159 VPB N_A_27_74#_c_297_n 0.0219674f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=2.135
cc_160 VPB N_A_27_74#_c_298_n 0.0641672f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.512
cc_161 VPB N_A_27_74#_c_299_n 0.00655372f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_162 VPB N_A_27_74#_c_300_n 0.0279846f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_163 VPB N_SCE_M1018_g 0.0487569f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_164 VPB N_SCE_M1017_g 0.0353741f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_165 VPB N_SCE_c_369_n 0.0130807f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.31
cc_166 VPB N_SCE_c_373_n 0.00304854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SCE_c_375_n 0.0215244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_SCE_c_376_n 0.0217946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_SCE_c_379_n 0.00321268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_D_M1027_g 0.0518086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_SCD_c_500_n 0.0182479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_SCD_c_498_n 0.0465251f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.66
cc_173 VPB SCD 0.00459774f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.16
cc_174 VPB N_CLK_M1025_g 0.0256722f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.66
cc_175 VPB N_CLK_c_540_n 0.00356962f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_176 VPB N_CLK_c_543_n 0.0122193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1037_119#_M1019_g 0.0347523f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.66
cc_178 VPB N_A_1037_119#_c_600_n 0.0150583f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_179 VPB N_A_1037_119#_M1033_g 0.0267134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1037_119#_c_610_n 0.00192327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1037_119#_c_624_n 0.00533583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1037_119#_c_615_n 0.0026077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1037_119#_c_619_n 0.0208366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1037_119#_c_627_n 0.0351933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1369_93#_M1006_g 0.0464726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1369_93#_c_812_n 0.0022112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1369_93#_c_813_n 0.0200789f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.31
cc_188 VPB N_A_1369_93#_c_818_n 0.00419195f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.512
cc_189 VPB N_RESET_B_c_913_n 0.00966093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_M1011_g 0.0290245f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.66
cc_191 VPB N_RESET_B_M1040_g 0.0235919f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_192 VPB N_RESET_B_c_917_n 0.0118326f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_193 VPB N_RESET_B_c_927_n 0.0224929f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.135
cc_194 VPB N_RESET_B_c_928_n 0.0153435f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=2.16
cc_195 VPB N_RESET_B_c_929_n 0.0117494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_RESET_B_c_930_n 0.0277936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_931_n 0.0206518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_c_932_n 0.00360243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_RESET_B_c_933_n 0.0138334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_c_934_n 0.00662848f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB RESET_B 0.00207862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_RESET_B_c_936_n 0.0433488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_937_n 0.00263108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_938_n 0.0370056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_939_n 0.00182623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_940_n 0.0307002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_941_n 0.0048181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_RESET_B_c_922_n 0.00104493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1235_119#_M1007_g 0.0229573f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_210 VPB N_A_1235_119#_c_1165_n 0.00275976f $X=-0.19 $Y=1.66 $X2=1.23
+ $Y2=1.145
cc_211 VPB N_A_1235_119#_c_1159_n 0.012127f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_212 VPB N_A_1235_119#_c_1160_n 0.0125372f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_213 VPB N_A_1235_119#_c_1168_n 0.00176819f $X=-0.19 $Y=1.66 $X2=2.53
+ $Y2=2.135
cc_214 VPB N_A_1235_119#_c_1163_n 0.0168224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_819_119#_c_1270_n 0.0732417f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.31
cc_216 VPB N_A_819_119#_c_1283_n 0.0542667f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_217 VPB N_A_819_119#_c_1284_n 0.0106469f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_218 VPB N_A_819_119#_M1024_g 0.0384094f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_219 VPB N_A_819_119#_c_1286_n 0.179819f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.512
cc_220 VPB N_A_819_119#_M1015_g 0.0301782f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_221 VPB N_A_819_119#_c_1274_n 0.0205647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_819_119#_c_1275_n 0.00335889f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.135
cc_223 VPB N_A_819_119#_c_1290_n 0.00898883f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=2.16
cc_224 VPB N_A_819_119#_c_1291_n 0.00248311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_819_119#_c_1279_n 9.43952e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_819_119#_c_1280_n 0.0153562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_819_119#_c_1294_n 0.0165206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_2008_48#_c_1459_n 0.0363084f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_229 VPB N_A_2008_48#_M1039_g 0.0373974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_2008_48#_c_1460_n 0.00554437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2008_48#_c_1468_n 0.00200572f $X=-0.19 $Y=1.66 $X2=0.365
+ $Y2=1.145
cc_232 VPB N_A_2008_48#_c_1469_n 0.00187906f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_233 VPB N_A_2008_48#_c_1470_n 0.00270297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_2008_48#_c_1471_n 0.00272239f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_235 VPB N_A_2008_48#_c_1472_n 0.00849573f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.512
cc_236 VPB N_A_2008_48#_c_1462_n 0.00102188f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_237 VPB N_A_2008_48#_c_1474_n 0.00510534f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_238 VPB N_A_1747_74#_M1026_g 0.0263466f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_239 VPB N_A_1747_74#_c_1594_n 0.0251829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1747_74#_c_1595_n 0.00896715f $X=-0.19 $Y=1.66 $X2=2.365
+ $Y2=2.135
cc_241 VPB N_A_1747_74#_M1008_g 0.0469089f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_242 VPB N_A_1747_74#_c_1606_n 0.0264704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1747_74#_c_1607_n 0.0348437f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_244 VPB N_A_1747_74#_c_1597_n 0.00103641f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_245 VPB N_A_1747_74#_c_1609_n 0.00518853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1747_74#_c_1610_n 0.00295628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1747_74#_c_1599_n 0.00536586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_2513_424#_M1000_g 0.0295193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_2513_424#_c_1767_n 0.00663366f $X=-0.19 $Y=1.66 $X2=1.23
+ $Y2=1.145
cc_250 VPB N_VPWR_c_1811_n 0.00637601f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_251 VPB N_VPWR_c_1812_n 0.00661417f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_252 VPB N_VPWR_c_1813_n 0.00151893f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_253 VPB N_VPWR_c_1814_n 0.0138079f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_254 VPB N_VPWR_c_1815_n 0.0149001f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=2.16
cc_255 VPB N_VPWR_c_1816_n 0.0169489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1817_n 0.0142621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1818_n 0.0141394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1819_n 0.0338628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1820_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1821_n 0.033442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1822_n 0.00485379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1823_n 0.0562135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1824_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1825_n 5.14268e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1826_n 0.0456433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1827_n 0.0221228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1828_n 0.0505955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1829_n 0.020722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1830_n 0.0342915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1831_n 0.0189057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1810_n 0.128454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1833_n 0.00670471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1834_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1835_n 0.0066101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1836_n 0.00853483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1837_n 0.00535984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_413_90#_c_1992_n 0.00761494f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_278 VPB N_A_413_90#_c_1999_n 0.0115072f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_279 VPB N_A_413_90#_c_2000_n 0.00521527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_413_90#_c_2001_n 0.00664887f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_281 VPB N_A_413_90#_c_2002_n 0.00184105f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_282 VPB N_A_413_90#_c_1996_n 0.00541266f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_283 VPB N_A_413_90#_c_2004_n 0.00223406f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_284 VPB N_A_413_90#_c_2005_n 0.0123661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB Q_N 0.0163642f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_286 VPB Q 0.0100967f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_287 VPB Q 0.0417413f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.512
cc_288 VPB N_Q_c_2160_n 0.00779848f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=2.16
cc_289 N_A_27_74#_c_290_n N_SCE_M1038_g 0.00834942f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_291_n N_SCE_M1038_g 0.017345f $X=0.2 $Y=2.05 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_292_n N_SCE_M1038_g 0.0301676f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_293_n N_SCE_M1038_g 0.00651386f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_297_n N_SCE_M1018_g 0.0132272f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_298_n N_SCE_M1018_g 0.0182817f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_297_n N_SCE_M1017_g 0.0163411f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_298_n N_SCE_M1017_g 7.71431e-19 $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_298_n N_SCE_c_369_n 0.0185427f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_297_n N_SCE_c_372_n 0.0226621f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_299_n N_SCE_c_372_n 0.00221846f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_300_n N_SCE_c_372_n 3.5076e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_299_n N_SCE_c_373_n 0.0245971f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_300_n N_SCE_c_373_n 9.36187e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_299_n N_SCE_c_374_n 3.27278e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_300_n N_SCE_c_374_n 0.0181552f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_292_n N_SCE_c_375_n 0.00418009f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_292_n N_SCE_c_376_n 3.70854e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_293_n N_SCE_c_376_n 0.0219044f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_297_n N_SCE_c_376_n 0.00313888f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_291_n N_SCE_c_378_n 0.0195247f $X=0.2 $Y=2.05 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_292_n N_SCE_c_378_n 0.0626128f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_293_n N_SCE_c_378_n 0.00563186f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_298_n N_SCE_c_378_n 0.0467278f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_297_n N_SCE_c_379_n 0.0467278f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_299_n N_SCE_c_379_n 0.00165158f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_315 N_A_27_74#_M1030_g N_D_M1027_g 0.0149489f $X=2.485 $Y=2.64 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_297_n N_D_M1027_g 0.017008f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_299_n N_D_M1027_g 0.00136754f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_300_n N_D_M1027_g 0.0213178f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_292_n N_D_c_456_n 2.658e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_293_n N_D_c_456_n 0.0150607f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_289_n N_D_c_457_n 0.00525376f $X=1.485 $Y=0.98 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_292_n N_D_c_457_n 0.0286966f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_293_n N_D_c_457_n 7.30413e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_289_n N_D_c_458_n 0.0223399f $X=1.485 $Y=0.98 $X2=0 $Y2=0
cc_325 N_A_27_74#_M1030_g N_SCD_c_500_n 0.02946f $X=2.485 $Y=2.64 $X2=0 $Y2=0
cc_326 N_A_27_74#_M1030_g N_SCD_c_498_n 0.00353217f $X=2.485 $Y=2.64 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_299_n N_SCD_c_498_n 0.00371252f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_300_n N_SCD_c_498_n 0.0205599f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_299_n SCD 0.0195516f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_300_n SCD 3.48225e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_297_n N_VPWR_c_1811_n 0.0227172f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_332 N_A_27_74#_c_298_n N_VPWR_c_1811_n 0.0251436f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_M1030_g N_VPWR_c_1812_n 0.00125706f $X=2.485 $Y=2.64 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_298_n N_VPWR_c_1819_n 0.0408473f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_M1030_g N_VPWR_c_1826_n 0.00520371f $X=2.485 $Y=2.64 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_M1030_g N_VPWR_c_1810_n 0.00517166f $X=2.485 $Y=2.64 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_c_298_n N_VPWR_c_1810_n 0.0344402f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_M1030_g N_A_413_90#_c_2006_n 0.00998656f $X=2.485 $Y=2.64
+ $X2=0 $Y2=0
cc_339 N_A_27_74#_c_299_n N_A_413_90#_c_2006_n 0.0182477f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_300_n N_A_413_90#_c_2006_n 4.28484e-19 $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_M1030_g N_A_413_90#_c_2004_n 0.0106872f $X=2.485 $Y=2.64 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_297_n N_A_413_90#_c_2004_n 0.0181873f $X=2.365 $Y=2.135
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_c_299_n N_A_413_90#_c_2004_n 0.00362443f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_289_n N_VGND_c_2179_n 0.00108896f $X=1.485 $Y=0.98 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_290_n N_VGND_c_2179_n 0.0179429f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_346 N_A_27_74#_c_292_n N_VGND_c_2179_n 0.0288081f $X=1.23 $Y=1.145 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_290_n N_VGND_c_2188_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_348 N_A_27_74#_c_289_n N_VGND_c_2189_n 8.05596e-19 $X=1.485 $Y=0.98 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_290_n N_VGND_c_2194_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_289_n N_noxref_25_c_2317_n 9.72985e-19 $X=1.485 $Y=0.98
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_c_292_n N_noxref_25_c_2317_n 0.0201381f $X=1.23 $Y=1.145 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_293_n N_noxref_25_c_2317_n 0.00573089f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_353 N_A_27_74#_c_289_n N_noxref_25_c_2318_n 0.0139744f $X=1.485 $Y=0.98 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_292_n N_noxref_25_c_2318_n 0.00121356f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_355 N_A_27_74#_c_293_n N_noxref_25_c_2318_n 0.00100866f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_356 N_SCE_c_372_n N_D_M1027_g 0.0147488f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_357 N_SCE_c_373_n N_D_M1027_g 3.07837e-19 $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_358 N_SCE_c_376_n N_D_M1027_g 0.0821376f $X=1.615 $Y=1.715 $X2=0 $Y2=0
cc_359 N_SCE_c_379_n N_D_M1027_g 0.00533998f $X=1.795 $Y=1.685 $X2=0 $Y2=0
cc_360 N_SCE_c_371_n N_D_c_456_n 0.00877867f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_361 N_SCE_c_373_n N_D_c_456_n 0.00122493f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_362 N_SCE_c_374_n N_D_c_456_n 0.0213592f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_363 N_SCE_c_379_n N_D_c_456_n 0.00402499f $X=1.795 $Y=1.685 $X2=0 $Y2=0
cc_364 N_SCE_c_370_n N_D_c_457_n 2.24037e-19 $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_365 N_SCE_c_371_n N_D_c_457_n 0.00102769f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_366 N_SCE_c_373_n N_D_c_457_n 0.00246469f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_367 N_SCE_c_376_n N_D_c_457_n 9.21361e-19 $X=1.615 $Y=1.715 $X2=0 $Y2=0
cc_368 N_SCE_c_378_n N_D_c_457_n 0.0411265f $X=1.6 $Y=1.685 $X2=0 $Y2=0
cc_369 N_SCE_c_370_n N_D_c_458_n 0.00971463f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_370 N_SCE_c_373_n N_SCD_c_496_n 0.00685255f $X=2.5 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_371 N_SCE_c_377_n N_SCD_c_496_n 0.02052f $X=2.5 $Y=1.26 $X2=-0.19 $Y2=-0.245
cc_372 N_SCE_c_370_n N_SCD_M1022_g 0.0460512f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_373 N_SCE_c_377_n N_SCD_M1022_g 0.00782258f $X=2.5 $Y=1.26 $X2=0 $Y2=0
cc_374 N_SCE_c_373_n SCD 0.0148322f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_375 N_SCE_M1018_g N_VPWR_c_1811_n 0.0034688f $X=1.115 $Y=2.64 $X2=0 $Y2=0
cc_376 N_SCE_M1017_g N_VPWR_c_1811_n 0.0154602f $X=1.615 $Y=2.64 $X2=0 $Y2=0
cc_377 N_SCE_M1018_g N_VPWR_c_1819_n 0.00519929f $X=1.115 $Y=2.64 $X2=0 $Y2=0
cc_378 N_SCE_M1017_g N_VPWR_c_1826_n 0.00460063f $X=1.615 $Y=2.64 $X2=0 $Y2=0
cc_379 N_SCE_M1018_g N_VPWR_c_1810_n 0.00983675f $X=1.115 $Y=2.64 $X2=0 $Y2=0
cc_380 N_SCE_M1017_g N_VPWR_c_1810_n 0.00908371f $X=1.615 $Y=2.64 $X2=0 $Y2=0
cc_381 N_SCE_c_370_n N_A_413_90#_c_1991_n 0.00445896f $X=2.62 $Y=0.98 $X2=0
+ $Y2=0
cc_382 N_SCE_c_371_n N_A_413_90#_c_1991_n 0.00379357f $X=2.62 $Y=1.105 $X2=0
+ $Y2=0
cc_383 N_SCE_c_373_n N_A_413_90#_c_1991_n 0.00928826f $X=2.5 $Y=1.425 $X2=0
+ $Y2=0
cc_384 N_SCE_M1017_g N_A_413_90#_c_2004_n 0.00172668f $X=1.615 $Y=2.64 $X2=0
+ $Y2=0
cc_385 N_SCE_c_370_n N_A_413_90#_c_1997_n 0.00712912f $X=2.62 $Y=0.98 $X2=0
+ $Y2=0
cc_386 N_SCE_c_371_n N_A_413_90#_c_1997_n 0.004963f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_387 N_SCE_c_372_n N_A_413_90#_c_1997_n 0.00539971f $X=2.395 $Y=1.575 $X2=0
+ $Y2=0
cc_388 N_SCE_c_373_n N_A_413_90#_c_1997_n 0.016626f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_389 N_SCE_c_374_n N_A_413_90#_c_1997_n 0.00253045f $X=2.5 $Y=1.425 $X2=0
+ $Y2=0
cc_390 N_SCE_M1038_g N_VGND_c_2179_n 0.0141679f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_391 N_SCE_M1038_g N_VGND_c_2188_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_392 N_SCE_c_370_n N_VGND_c_2189_n 7.35405e-19 $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_393 N_SCE_M1038_g N_VGND_c_2194_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_394 N_SCE_M1038_g N_noxref_25_c_2317_n 7.01965e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_395 N_SCE_c_370_n N_noxref_25_c_2318_n 0.00865752f $X=2.62 $Y=0.98 $X2=0
+ $Y2=0
cc_396 N_SCE_M1038_g N_noxref_25_c_2319_n 6.37214e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_397 N_SCE_c_370_n N_noxref_25_c_2320_n 0.00130896f $X=2.62 $Y=0.98 $X2=0
+ $Y2=0
cc_398 N_D_M1027_g N_VPWR_c_1811_n 0.00217652f $X=2.035 $Y=2.64 $X2=0 $Y2=0
cc_399 N_D_M1027_g N_VPWR_c_1826_n 0.00520371f $X=2.035 $Y=2.64 $X2=0 $Y2=0
cc_400 N_D_M1027_g N_VPWR_c_1810_n 0.00982921f $X=2.035 $Y=2.64 $X2=0 $Y2=0
cc_401 N_D_M1027_g N_A_413_90#_c_2004_n 0.0123942f $X=2.035 $Y=2.64 $X2=0 $Y2=0
cc_402 N_D_c_456_n N_A_413_90#_c_1997_n 9.2104e-19 $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_403 N_D_c_457_n N_A_413_90#_c_1997_n 0.0209433f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_404 N_D_c_458_n N_A_413_90#_c_1997_n 0.00597193f $X=1.947 $Y=0.98 $X2=0 $Y2=0
cc_405 N_D_c_458_n N_VGND_c_2189_n 8.05596e-19 $X=1.947 $Y=0.98 $X2=0 $Y2=0
cc_406 N_D_c_456_n N_noxref_25_c_2318_n 0.0014811f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_407 N_D_c_457_n N_noxref_25_c_2318_n 0.0171941f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_408 N_D_c_458_n N_noxref_25_c_2318_n 0.0105212f $X=1.947 $Y=0.98 $X2=0 $Y2=0
cc_409 N_D_c_457_n noxref_26 0.00381079f $X=1.935 $Y=1.145 $X2=-0.19 $Y2=-0.245
cc_410 N_SCD_M1022_g N_RESET_B_M1028_g 0.015105f $X=3.01 $Y=0.695 $X2=0 $Y2=0
cc_411 N_SCD_c_496_n N_RESET_B_c_913_n 0.0207196f $X=3.01 $Y=1.255 $X2=0 $Y2=0
cc_412 N_SCD_M1022_g N_RESET_B_c_913_n 0.0106209f $X=3.01 $Y=0.695 $X2=0 $Y2=0
cc_413 SCD N_RESET_B_c_913_n 0.00399618f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_414 N_SCD_c_500_n N_RESET_B_M1011_g 0.0112676f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_415 N_SCD_c_498_n N_RESET_B_c_927_n 0.0319872f $X=3.04 $Y=1.945 $X2=0 $Y2=0
cc_416 N_SCD_c_500_n N_VPWR_c_1812_n 0.0102474f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_417 N_SCD_c_500_n N_VPWR_c_1826_n 0.00460063f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_418 N_SCD_c_500_n N_VPWR_c_1810_n 0.00444149f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_419 N_SCD_c_500_n N_A_413_90#_c_2006_n 0.0143512f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_420 N_SCD_c_498_n N_A_413_90#_c_2006_n 0.00193785f $X=3.04 $Y=1.945 $X2=0
+ $Y2=0
cc_421 SCD N_A_413_90#_c_2006_n 0.0184669f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_422 N_SCD_c_496_n N_A_413_90#_c_1991_n 0.00322121f $X=3.01 $Y=1.255 $X2=0
+ $Y2=0
cc_423 N_SCD_M1022_g N_A_413_90#_c_1991_n 0.0124958f $X=3.01 $Y=0.695 $X2=0
+ $Y2=0
cc_424 SCD N_A_413_90#_c_1991_n 0.0149668f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_425 N_SCD_c_496_n N_A_413_90#_c_1992_n 7.13262e-19 $X=3.01 $Y=1.255 $X2=0
+ $Y2=0
cc_426 N_SCD_M1022_g N_A_413_90#_c_1992_n 0.00203777f $X=3.01 $Y=0.695 $X2=0
+ $Y2=0
cc_427 N_SCD_c_498_n N_A_413_90#_c_1992_n 0.00317611f $X=3.04 $Y=1.945 $X2=0
+ $Y2=0
cc_428 SCD N_A_413_90#_c_1992_n 0.0514814f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_429 N_SCD_c_500_n N_A_413_90#_c_2004_n 0.00161343f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_430 N_SCD_M1022_g N_A_413_90#_c_1997_n 0.00135115f $X=3.01 $Y=0.695 $X2=0
+ $Y2=0
cc_431 N_SCD_c_500_n N_A_413_90#_c_2005_n 0.00188054f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_432 N_SCD_M1022_g N_VGND_c_2189_n 7.30329e-19 $X=3.01 $Y=0.695 $X2=0 $Y2=0
cc_433 N_SCD_M1022_g N_noxref_25_c_2318_n 0.00674254f $X=3.01 $Y=0.695 $X2=0
+ $Y2=0
cc_434 N_SCD_M1022_g N_noxref_25_c_2320_n 0.00799117f $X=3.01 $Y=0.695 $X2=0
+ $Y2=0
cc_435 N_CLK_c_544_n N_A_1037_119#_c_605_n 9.44493e-19 $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_CLK_M1025_g N_A_1037_119#_c_615_n 6.37706e-19 $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_437 N_CLK_c_541_n N_RESET_B_c_913_n 0.00133682f $X=4.395 $Y=1.477 $X2=0 $Y2=0
cc_438 N_CLK_c_542_n N_RESET_B_c_913_n 0.0212633f $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_439 N_CLK_c_544_n N_RESET_B_c_914_n 0.00999579f $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_440 N_CLK_c_540_n N_RESET_B_c_931_n 0.00190567f $X=4.56 $Y=1.61 $X2=0 $Y2=0
cc_441 N_CLK_c_541_n N_RESET_B_c_931_n 0.0052925f $X=4.395 $Y=1.477 $X2=0 $Y2=0
cc_442 N_CLK_M1025_g N_RESET_B_c_932_n 3.38591e-19 $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_443 N_CLK_c_541_n N_RESET_B_c_932_n 0.00434753f $X=4.395 $Y=1.477 $X2=0 $Y2=0
cc_444 N_CLK_M1025_g N_RESET_B_c_936_n 0.00527527f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_445 N_CLK_c_541_n N_RESET_B_c_936_n 0.00193077f $X=4.395 $Y=1.477 $X2=0 $Y2=0
cc_446 N_CLK_c_542_n N_RESET_B_c_936_n 0.0213386f $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_447 N_CLK_c_539_n N_RESET_B_c_937_n 3.35172e-19 $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_448 N_CLK_M1025_g N_RESET_B_c_937_n 0.00104729f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_449 N_CLK_c_541_n N_RESET_B_c_937_n 0.0296391f $X=4.395 $Y=1.477 $X2=0 $Y2=0
cc_450 N_CLK_c_542_n N_RESET_B_c_937_n 3.80123e-19 $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_451 N_CLK_c_541_n N_A_819_119#_M1013_s 0.00228945f $X=4.395 $Y=1.477
+ $X2=-0.19 $Y2=-0.245
cc_452 N_CLK_c_540_n N_A_819_119#_c_1296_n 0.0133012f $X=4.56 $Y=1.61 $X2=0
+ $Y2=0
cc_453 N_CLK_c_543_n N_A_819_119#_c_1296_n 0.00256125f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_454 N_CLK_c_544_n N_A_819_119#_c_1296_n 0.00731194f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_455 N_CLK_M1025_g N_A_819_119#_c_1299_n 0.0115718f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_456 N_CLK_c_540_n N_A_819_119#_c_1299_n 0.00404952f $X=4.56 $Y=1.61 $X2=0
+ $Y2=0
cc_457 N_CLK_c_540_n N_A_819_119#_c_1278_n 0.0147007f $X=4.56 $Y=1.61 $X2=0
+ $Y2=0
cc_458 N_CLK_c_543_n N_A_819_119#_c_1278_n 2.59598e-19 $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_459 N_CLK_c_544_n N_A_819_119#_c_1278_n 0.0043748f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_460 N_CLK_M1025_g N_A_819_119#_c_1291_n 0.00252678f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_461 N_CLK_c_539_n N_A_819_119#_c_1305_n 9.80044e-19 $X=4.395 $Y=1.51 $X2=0
+ $Y2=0
cc_462 N_CLK_c_541_n N_A_819_119#_c_1305_n 0.0133012f $X=4.395 $Y=1.477 $X2=0
+ $Y2=0
cc_463 N_CLK_c_544_n N_A_819_119#_c_1305_n 0.00627595f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_464 N_CLK_c_539_n N_A_819_119#_c_1308_n 3.66762e-19 $X=4.395 $Y=1.51 $X2=0
+ $Y2=0
cc_465 N_CLK_M1025_g N_A_819_119#_c_1308_n 0.0043986f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_466 N_CLK_c_540_n N_A_819_119#_c_1308_n 0.0116041f $X=4.56 $Y=1.61 $X2=0
+ $Y2=0
cc_467 N_CLK_c_541_n N_A_819_119#_c_1308_n 0.0027896f $X=4.395 $Y=1.477 $X2=0
+ $Y2=0
cc_468 N_CLK_c_543_n N_A_819_119#_c_1308_n 0.0038904f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_469 N_CLK_c_540_n N_A_819_119#_c_1279_n 0.0273204f $X=4.56 $Y=1.61 $X2=0
+ $Y2=0
cc_470 N_CLK_c_543_n N_A_819_119#_c_1279_n 0.00249677f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_471 N_CLK_c_540_n N_A_819_119#_c_1280_n 2.99534e-19 $X=4.56 $Y=1.61 $X2=0
+ $Y2=0
cc_472 N_CLK_c_543_n N_A_819_119#_c_1280_n 0.0252665f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_473 N_CLK_c_544_n N_A_819_119#_c_1281_n 0.0203845f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_474 N_CLK_M1025_g N_A_819_119#_c_1294_n 0.0455485f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_475 N_CLK_M1025_g N_VPWR_c_1813_n 0.017461f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_476 N_CLK_M1025_g N_VPWR_c_1821_n 0.00401239f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_477 N_CLK_M1025_g N_VPWR_c_1810_n 0.00589267f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_478 N_CLK_c_541_n N_A_413_90#_c_1992_n 0.0380255f $X=4.395 $Y=1.477 $X2=0
+ $Y2=0
cc_479 N_CLK_c_542_n N_A_413_90#_c_1992_n 0.0018935f $X=3.94 $Y=1.445 $X2=0
+ $Y2=0
cc_480 N_CLK_M1025_g N_A_413_90#_c_1999_n 0.0166738f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_481 N_CLK_M1025_g N_A_413_90#_c_2005_n 0.0128449f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_482 N_CLK_c_541_n N_VGND_c_2180_n 0.00368956f $X=4.395 $Y=1.477 $X2=0 $Y2=0
cc_483 N_CLK_c_542_n N_VGND_c_2180_n 7.67353e-19 $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_484 N_CLK_c_544_n N_VGND_c_2180_n 0.00353997f $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_485 N_CLK_c_544_n N_VGND_c_2181_n 0.00423158f $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_486 N_CLK_c_544_n N_VGND_c_2194_n 9.39239e-19 $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_487 N_A_1037_119#_c_612_n N_A_1369_93#_M1041_d 0.00176461f $X=8.78 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_488 N_A_1037_119#_M1036_g N_A_1369_93#_M1004_g 0.0307978f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_489 N_A_1037_119#_c_608_n N_A_1369_93#_M1004_g 0.0037178f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_490 N_A_1037_119#_c_611_n N_A_1369_93#_M1004_g 0.00314912f $X=7.1 $Y=0.595
+ $X2=0 $Y2=0
cc_491 N_A_1037_119#_M1019_g N_A_1369_93#_M1006_g 0.00360575f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_492 N_A_1037_119#_c_619_n N_A_1369_93#_M1006_g 0.00126194f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_493 N_A_1037_119#_c_600_n N_A_1369_93#_c_813_n 0.0307978f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_494 N_A_1037_119#_c_637_p N_A_1369_93#_c_813_n 4.26127e-19 $X=7.185 $Y=0.68
+ $X2=0 $Y2=0
cc_495 N_A_1037_119#_c_619_n N_A_1369_93#_c_813_n 6.28976e-19 $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_496 N_A_1037_119#_c_639_p N_A_1369_93#_c_814_n 0.0588266f $X=7.94 $Y=0.68
+ $X2=0 $Y2=0
cc_497 N_A_1037_119#_c_612_n N_A_1369_93#_c_814_n 0.0034413f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_498 N_A_1037_119#_c_637_p N_A_1369_93#_c_815_n 0.0111231f $X=7.185 $Y=0.68
+ $X2=0 $Y2=0
cc_499 N_A_1037_119#_c_602_n N_A_1369_93#_c_836_n 0.0041679f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_500 N_A_1037_119#_c_612_n N_A_1369_93#_c_836_n 0.0158584f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_501 N_A_1037_119#_c_604_n N_A_1369_93#_c_816_n 0.00444121f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_502 N_A_1037_119#_c_614_n N_A_1369_93#_c_816_n 0.00425045f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_503 N_A_1037_119#_c_604_n N_A_1369_93#_c_817_n 0.010636f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_504 N_A_1037_119#_c_614_n N_A_1369_93#_c_817_n 0.00854237f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_505 N_A_1037_119#_c_616_n N_A_1369_93#_c_817_n 0.011663f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_506 N_A_1037_119#_c_618_n N_A_1369_93#_c_817_n 0.00620138f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_507 N_A_1037_119#_c_624_n N_A_1369_93#_c_818_n 0.00513903f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_508 N_A_1037_119#_c_618_n N_A_1369_93#_c_818_n 0.0132001f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_509 N_A_1037_119#_c_602_n N_A_1369_93#_c_819_n 0.00251445f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_510 N_A_1037_119#_c_604_n N_A_1369_93#_c_819_n 8.10451e-19 $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_511 N_A_1037_119#_c_614_n N_A_1369_93#_c_819_n 9.81795e-19 $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_512 N_A_1037_119#_c_616_n N_A_1369_93#_c_819_n 0.00881609f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_513 N_A_1037_119#_M1036_g N_RESET_B_c_914_n 0.00882199f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_514 N_A_1037_119#_c_608_n N_RESET_B_c_914_n 0.034331f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_515 N_A_1037_119#_c_609_n N_RESET_B_c_914_n 0.00593026f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_516 N_A_1037_119#_c_608_n N_RESET_B_M1034_g 0.00421573f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_517 N_A_1037_119#_c_611_n N_RESET_B_M1034_g 0.00457302f $X=7.1 $Y=0.595 $X2=0
+ $Y2=0
cc_518 N_A_1037_119#_c_639_p N_RESET_B_M1034_g 0.0130455f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_519 N_A_1037_119#_c_662_p N_RESET_B_M1034_g 0.00387243f $X=8.025 $Y=0.595
+ $X2=0 $Y2=0
cc_520 N_A_1037_119#_c_639_p N_RESET_B_c_920_n 0.0013334f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_521 N_A_1037_119#_M1019_g N_RESET_B_c_931_n 0.00468421f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_522 N_A_1037_119#_c_600_n N_RESET_B_c_931_n 0.00384754f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_523 N_A_1037_119#_c_610_n N_RESET_B_c_931_n 0.0160518f $X=6.055 $Y=1.74 $X2=0
+ $Y2=0
cc_524 N_A_1037_119#_c_615_n N_RESET_B_c_931_n 0.0354867f $X=5.387 $Y=1.74 $X2=0
+ $Y2=0
cc_525 N_A_1037_119#_c_619_n N_RESET_B_c_931_n 0.0038641f $X=6.055 $Y=1.65 $X2=0
+ $Y2=0
cc_526 N_A_1037_119#_c_624_n N_RESET_B_c_933_n 0.0136948f $X=9.67 $Y=2.065 $X2=0
+ $Y2=0
cc_527 N_A_1037_119#_c_618_n N_RESET_B_c_933_n 0.0078678f $X=9.63 $Y=1.46 $X2=0
+ $Y2=0
cc_528 N_A_1037_119#_c_627_n N_RESET_B_c_933_n 0.00532527f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_529 N_A_1037_119#_c_602_n N_A_1235_119#_M1041_g 0.0262081f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_530 N_A_1037_119#_c_612_n N_A_1235_119#_M1041_g 0.0116741f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_531 N_A_1037_119#_c_600_n N_A_1235_119#_c_1158_n 4.04038e-19 $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_532 N_A_1037_119#_M1036_g N_A_1235_119#_c_1158_n 0.0145691f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_533 N_A_1037_119#_c_608_n N_A_1235_119#_c_1158_n 0.0426901f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_534 N_A_1037_119#_M1019_g N_A_1235_119#_c_1165_n 0.00506299f $X=6.115
+ $Y=2.525 $X2=0 $Y2=0
cc_535 N_A_1037_119#_c_600_n N_A_1235_119#_c_1165_n 8.9028e-19 $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_536 N_A_1037_119#_M1019_g N_A_1235_119#_c_1159_n 3.99449e-19 $X=6.115
+ $Y=2.525 $X2=0 $Y2=0
cc_537 N_A_1037_119#_M1036_g N_A_1235_119#_c_1159_n 0.00803125f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_538 N_A_1037_119#_c_604_n N_A_1235_119#_c_1163_n 0.00328288f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_539 N_A_1037_119#_c_606_n N_A_819_119#_c_1268_n 3.06294e-19 $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_540 N_A_1037_119#_c_607_n N_A_819_119#_c_1268_n 0.00650486f $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_541 N_A_1037_119#_c_606_n N_A_819_119#_c_1269_n 0.00182325f $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_542 N_A_1037_119#_c_607_n N_A_819_119#_c_1269_n 0.00842158f $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_543 N_A_1037_119#_M1019_g N_A_819_119#_c_1270_n 0.0253232f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_544 N_A_1037_119#_c_607_n N_A_819_119#_c_1270_n 6.92436e-19 $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_545 N_A_1037_119#_c_610_n N_A_819_119#_c_1270_n 0.00878462f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_546 N_A_1037_119#_c_615_n N_A_819_119#_c_1270_n 0.0184173f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_547 N_A_1037_119#_c_619_n N_A_819_119#_c_1270_n 0.0213783f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_548 N_A_1037_119#_c_608_n N_A_819_119#_c_1271_n 0.00108386f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_549 N_A_1037_119#_c_610_n N_A_819_119#_c_1271_n 0.00463817f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_550 N_A_1037_119#_c_619_n N_A_819_119#_c_1271_n 0.0102445f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_551 N_A_1037_119#_c_606_n N_A_819_119#_c_1272_n 0.00828721f $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_552 N_A_1037_119#_c_608_n N_A_819_119#_c_1272_n 0.00621399f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_553 N_A_1037_119#_M1019_g N_A_819_119#_c_1283_n 0.0123549f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_554 N_A_1037_119#_M1036_g N_A_819_119#_c_1273_n 0.0190129f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_555 N_A_1037_119#_c_605_n N_A_819_119#_c_1273_n 0.00410301f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_556 N_A_1037_119#_c_608_n N_A_819_119#_c_1273_n 0.00192639f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_557 N_A_1037_119#_M1019_g N_A_819_119#_M1024_g 0.0162604f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_558 N_A_1037_119#_c_600_n N_A_819_119#_M1024_g 0.00374845f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_559 N_A_1037_119#_M1033_g N_A_819_119#_M1015_g 0.00862099f $X=9.77 $Y=2.655
+ $X2=0 $Y2=0
cc_560 N_A_1037_119#_c_624_n N_A_819_119#_M1015_g 0.00164955f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_561 N_A_1037_119#_c_627_n N_A_819_119#_M1015_g 0.0045203f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_562 N_A_1037_119#_c_614_n N_A_819_119#_c_1274_n 3.3013e-19 $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_563 N_A_1037_119#_c_624_n N_A_819_119#_c_1274_n 0.00813875f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_564 N_A_1037_119#_c_617_n N_A_819_119#_c_1274_n 0.0126321f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_565 N_A_1037_119#_c_618_n N_A_819_119#_c_1274_n 0.0175647f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_566 N_A_1037_119#_c_627_n N_A_819_119#_c_1274_n 0.0191393f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_567 N_A_1037_119#_c_603_n N_A_819_119#_c_1275_n 0.0126321f $X=9.105 $Y=1.16
+ $X2=0 $Y2=0
cc_568 N_A_1037_119#_c_614_n N_A_819_119#_M1016_g 0.00266955f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_569 N_A_1037_119#_c_617_n N_A_819_119#_M1016_g 0.0176907f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_570 N_A_1037_119#_c_618_n N_A_819_119#_M1016_g 0.00700032f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_571 N_A_1037_119#_c_607_n N_A_819_119#_c_1277_n 0.00706417f $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_572 N_A_1037_119#_c_615_n N_A_819_119#_c_1299_n 0.00840728f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_573 N_A_1037_119#_c_607_n N_A_819_119#_c_1278_n 0.00560834f $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_574 N_A_1037_119#_c_615_n N_A_819_119#_c_1291_n 0.00717919f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_575 N_A_1037_119#_c_615_n N_A_819_119#_c_1308_n 0.004494f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_576 N_A_1037_119#_c_606_n N_A_819_119#_c_1279_n 0.00212908f $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_577 N_A_1037_119#_c_607_n N_A_819_119#_c_1279_n 0.00964804f $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_578 N_A_1037_119#_c_615_n N_A_819_119#_c_1279_n 0.020036f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_579 N_A_1037_119#_c_606_n N_A_819_119#_c_1280_n 0.0035545f $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_580 N_A_1037_119#_c_615_n N_A_819_119#_c_1280_n 0.00591228f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_581 N_A_1037_119#_c_605_n N_A_819_119#_c_1281_n 0.0105193f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_582 N_A_1037_119#_c_606_n N_A_819_119#_c_1281_n 0.00190426f $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_583 N_A_1037_119#_c_607_n N_A_819_119#_c_1281_n 0.00104006f $X=5.502 $Y=1.575
+ $X2=0 $Y2=0
cc_584 N_A_1037_119#_c_615_n N_A_819_119#_c_1294_n 0.00611642f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_585 N_A_1037_119#_c_618_n N_A_2008_48#_M1005_g 2.03511e-19 $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_586 N_A_1037_119#_c_624_n N_A_2008_48#_c_1459_n 0.0016211f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_587 N_A_1037_119#_c_627_n N_A_2008_48#_c_1459_n 0.0346924f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_588 N_A_1037_119#_M1033_g N_A_2008_48#_M1039_g 0.0346924f $X=9.77 $Y=2.655
+ $X2=0 $Y2=0
cc_589 N_A_1037_119#_c_612_n N_A_1747_74#_M1029_d 0.0019485f $X=8.78 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_590 N_A_1037_119#_c_733_p N_A_1747_74#_M1029_d 0.0100293f $X=8.865 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_591 N_A_1037_119#_c_616_n N_A_1747_74#_M1029_d 0.00256528f $X=9.27 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_592 N_A_1037_119#_M1033_g N_A_1747_74#_c_1615_n 0.00188718f $X=9.77 $Y=2.655
+ $X2=0 $Y2=0
cc_593 N_A_1037_119#_c_624_n N_A_1747_74#_c_1615_n 0.0330459f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_594 N_A_1037_119#_c_618_n N_A_1747_74#_c_1615_n 0.0143899f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_595 N_A_1037_119#_c_627_n N_A_1747_74#_c_1615_n 0.00236589f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_596 N_A_1037_119#_c_602_n N_A_1747_74#_c_1619_n 7.45707e-19 $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_597 N_A_1037_119#_c_612_n N_A_1747_74#_c_1619_n 0.00160036f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_598 N_A_1037_119#_c_733_p N_A_1747_74#_c_1619_n 0.0234496f $X=8.865 $Y=0.905
+ $X2=0 $Y2=0
cc_599 N_A_1037_119#_c_616_n N_A_1747_74#_c_1619_n 0.0221981f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_600 N_A_1037_119#_c_617_n N_A_1747_74#_c_1619_n 0.00683469f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_601 N_A_1037_119#_c_618_n N_A_1747_74#_c_1619_n 0.00536065f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_602 N_A_1037_119#_M1033_g N_A_1747_74#_c_1609_n 0.0151069f $X=9.77 $Y=2.655
+ $X2=0 $Y2=0
cc_603 N_A_1037_119#_c_624_n N_A_1747_74#_c_1609_n 0.0168861f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_604 N_A_1037_119#_c_627_n N_A_1747_74#_c_1609_n 0.00125859f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_605 N_A_1037_119#_c_733_p N_A_1747_74#_c_1598_n 0.00463964f $X=8.865 $Y=0.905
+ $X2=0 $Y2=0
cc_606 N_A_1037_119#_c_616_n N_A_1747_74#_c_1598_n 0.00785017f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_607 N_A_1037_119#_c_617_n N_A_1747_74#_c_1598_n 2.98286e-19 $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_608 N_A_1037_119#_c_624_n N_A_1747_74#_c_1599_n 0.0483469f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_609 N_A_1037_119#_c_618_n N_A_1747_74#_c_1599_n 0.0109876f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_610 N_A_1037_119#_c_627_n N_A_1747_74#_c_1599_n 0.00418902f $X=9.77 $Y=2.065
+ $X2=0 $Y2=0
cc_611 N_A_1037_119#_c_614_n N_A_1747_74#_c_1600_n 0.015348f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_612 N_A_1037_119#_c_616_n N_A_1747_74#_c_1600_n 0.00613506f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_613 N_A_1037_119#_c_617_n N_A_1747_74#_c_1600_n 0.00101813f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_614 N_A_1037_119#_c_618_n N_A_1747_74#_c_1600_n 0.0202102f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_615 N_A_1037_119#_M1033_g N_VPWR_c_1828_n 0.00463536f $X=9.77 $Y=2.655 $X2=0
+ $Y2=0
cc_616 N_A_1037_119#_M1019_g N_VPWR_c_1810_n 0.00112709f $X=6.115 $Y=2.525 $X2=0
+ $Y2=0
cc_617 N_A_1037_119#_M1033_g N_VPWR_c_1810_n 0.00619157f $X=9.77 $Y=2.655 $X2=0
+ $Y2=0
cc_618 N_A_1037_119#_M1035_d N_A_413_90#_c_1999_n 0.00612038f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_619 N_A_1037_119#_c_610_n N_A_413_90#_c_1999_n 0.00140057f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_620 N_A_1037_119#_c_615_n N_A_413_90#_c_1999_n 0.0302568f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_621 N_A_1037_119#_M1019_g N_A_413_90#_c_2000_n 0.00209388f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_622 N_A_1037_119#_c_610_n N_A_413_90#_c_2000_n 0.00102338f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_623 N_A_1037_119#_c_615_n N_A_413_90#_c_2000_n 0.00230268f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_624 N_A_1037_119#_c_605_n N_A_413_90#_c_1993_n 0.0208662f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_625 N_A_1037_119#_c_608_n N_A_413_90#_c_1993_n 0.0133345f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_626 N_A_1037_119#_M1019_g N_A_413_90#_c_2001_n 0.0158867f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_627 N_A_1037_119#_c_600_n N_A_413_90#_c_2001_n 0.00272338f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_628 N_A_1037_119#_c_610_n N_A_413_90#_c_2001_n 0.0118264f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_629 N_A_1037_119#_c_619_n N_A_413_90#_c_2001_n 0.001604f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_630 N_A_1037_119#_c_610_n N_A_413_90#_c_2002_n 0.0126264f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_631 N_A_1037_119#_c_615_n N_A_413_90#_c_2002_n 0.0143123f $X=5.387 $Y=1.74
+ $X2=0 $Y2=0
cc_632 N_A_1037_119#_c_619_n N_A_413_90#_c_2002_n 0.0018949f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_633 N_A_1037_119#_M1036_g N_A_413_90#_c_1994_n 0.00502428f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_634 N_A_1037_119#_c_608_n N_A_413_90#_c_1994_n 0.00422476f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_635 N_A_1037_119#_c_610_n N_A_413_90#_c_1994_n 0.00885768f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_636 N_A_1037_119#_c_619_n N_A_413_90#_c_1994_n 0.0064095f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_637 N_A_1037_119#_c_605_n N_A_413_90#_c_1995_n 4.34295e-19 $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_638 N_A_1037_119#_c_606_n N_A_413_90#_c_1995_n 0.0125704f $X=5.502 $Y=1.275
+ $X2=0 $Y2=0
cc_639 N_A_1037_119#_c_610_n N_A_413_90#_c_1995_n 0.0100819f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_640 N_A_1037_119#_c_619_n N_A_413_90#_c_1995_n 6.82307e-19 $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_641 N_A_1037_119#_M1019_g N_A_413_90#_c_1996_n 0.00381322f $X=6.115 $Y=2.525
+ $X2=0 $Y2=0
cc_642 N_A_1037_119#_c_600_n N_A_413_90#_c_1996_n 0.0116858f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_643 N_A_1037_119#_M1036_g N_A_413_90#_c_1996_n 0.0087802f $X=6.53 $Y=0.805
+ $X2=0 $Y2=0
cc_644 N_A_1037_119#_c_610_n N_A_413_90#_c_1996_n 0.0256541f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_645 N_A_1037_119#_c_619_n N_A_413_90#_c_1996_n 0.0020471f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_646 N_A_1037_119#_c_639_p N_VGND_M1034_d 0.0173685f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_647 N_A_1037_119#_c_662_p N_VGND_M1034_d 0.00302969f $X=8.025 $Y=0.595 $X2=0
+ $Y2=0
cc_648 N_A_1037_119#_c_613_n N_VGND_M1034_d 6.57704e-19 $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_649 N_A_1037_119#_c_605_n N_VGND_c_2181_n 0.0152912f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_650 N_A_1037_119#_c_609_n N_VGND_c_2181_n 0.0144411f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_651 N_A_1037_119#_c_608_n N_VGND_c_2182_n 0.0113026f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_652 N_A_1037_119#_c_639_p N_VGND_c_2182_n 0.0246763f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_653 N_A_1037_119#_c_613_n N_VGND_c_2182_n 0.0148567f $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_654 N_A_1037_119#_c_608_n N_VGND_c_2190_n 0.114006f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_655 N_A_1037_119#_c_609_n N_VGND_c_2190_n 0.0170431f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_656 N_A_1037_119#_c_639_p N_VGND_c_2190_n 0.0038254f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_657 N_A_1037_119#_c_602_n N_VGND_c_2191_n 0.00278271f $X=8.66 $Y=1.085 $X2=0
+ $Y2=0
cc_658 N_A_1037_119#_c_639_p N_VGND_c_2191_n 0.00323133f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_659 N_A_1037_119#_c_612_n N_VGND_c_2191_n 0.0543743f $X=8.78 $Y=0.34 $X2=0
+ $Y2=0
cc_660 N_A_1037_119#_c_613_n N_VGND_c_2191_n 0.0119262f $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_661 N_A_1037_119#_c_602_n N_VGND_c_2194_n 0.00358525f $X=8.66 $Y=1.085 $X2=0
+ $Y2=0
cc_662 N_A_1037_119#_c_608_n N_VGND_c_2194_n 0.0593877f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_1037_119#_c_609_n N_VGND_c_2194_n 0.00857552f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_664 N_A_1037_119#_c_639_p N_VGND_c_2194_n 0.0132173f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_665 N_A_1037_119#_c_612_n N_VGND_c_2194_n 0.0304188f $X=8.78 $Y=0.34 $X2=0
+ $Y2=0
cc_666 N_A_1037_119#_c_613_n N_VGND_c_2194_n 0.00656035f $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_667 N_A_1037_119#_c_637_p A_1399_119# 0.00131685f $X=7.185 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_668 N_A_1369_93#_M1004_g N_RESET_B_c_914_n 0.00882199f $X=6.92 $Y=0.805 $X2=0
+ $Y2=0
cc_669 N_A_1369_93#_c_815_n N_RESET_B_c_914_n 3.3965e-19 $X=7.235 $Y=1.02 $X2=0
+ $Y2=0
cc_670 N_A_1369_93#_M1004_g N_RESET_B_M1034_g 0.0377196f $X=6.92 $Y=0.805 $X2=0
+ $Y2=0
cc_671 N_A_1369_93#_c_814_n N_RESET_B_M1034_g 0.00787198f $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_672 N_A_1369_93#_c_815_n N_RESET_B_M1034_g 0.00122241f $X=7.235 $Y=1.02 $X2=0
+ $Y2=0
cc_673 N_A_1369_93#_M1004_g N_RESET_B_c_917_n 0.00306867f $X=6.92 $Y=0.805 $X2=0
+ $Y2=0
cc_674 N_A_1369_93#_M1006_g N_RESET_B_c_917_n 0.00439725f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_675 N_A_1369_93#_c_812_n N_RESET_B_c_917_n 0.0015409f $X=7.125 $Y=1.615 $X2=0
+ $Y2=0
cc_676 N_A_1369_93#_c_813_n N_RESET_B_c_917_n 0.0175447f $X=7.125 $Y=1.615 $X2=0
+ $Y2=0
cc_677 N_A_1369_93#_c_812_n N_RESET_B_c_920_n 0.00368383f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_678 N_A_1369_93#_c_813_n N_RESET_B_c_920_n 0.00405967f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_679 N_A_1369_93#_c_814_n N_RESET_B_c_920_n 0.0142771f $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_680 N_A_1369_93#_M1006_g N_RESET_B_c_928_n 0.0211295f $X=6.955 $Y=2.525 $X2=0
+ $Y2=0
cc_681 N_A_1369_93#_M1006_g N_RESET_B_c_931_n 0.0115372f $X=6.955 $Y=2.525 $X2=0
+ $Y2=0
cc_682 N_A_1369_93#_c_812_n N_RESET_B_c_931_n 0.00661774f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_683 N_A_1369_93#_c_813_n N_RESET_B_c_931_n 0.00189194f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_684 N_A_1369_93#_M1007_d N_RESET_B_c_933_n 0.00242247f $X=8.635 $Y=1.735
+ $X2=0 $Y2=0
cc_685 N_A_1369_93#_c_817_n N_RESET_B_c_933_n 0.00655969f $X=8.81 $Y=1.415 $X2=0
+ $Y2=0
cc_686 N_A_1369_93#_c_818_n N_RESET_B_c_933_n 0.0248508f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_687 N_A_1369_93#_c_814_n N_A_1235_119#_M1041_g 0.0108107f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_688 N_A_1369_93#_c_836_n N_A_1235_119#_M1041_g 0.00970467f $X=8.445 $Y=0.81
+ $X2=0 $Y2=0
cc_689 N_A_1369_93#_c_816_n N_A_1235_119#_M1041_g 0.0031265f $X=8.525 $Y=1.245
+ $X2=0 $Y2=0
cc_690 N_A_1369_93#_c_819_n N_A_1235_119#_M1041_g 0.0021525f $X=8.445 $Y=1.02
+ $X2=0 $Y2=0
cc_691 N_A_1369_93#_M1004_g N_A_1235_119#_c_1158_n 0.00671859f $X=6.92 $Y=0.805
+ $X2=0 $Y2=0
cc_692 N_A_1369_93#_M1004_g N_A_1235_119#_c_1159_n 0.00664117f $X=6.92 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_A_1369_93#_M1006_g N_A_1235_119#_c_1159_n 0.00837363f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_694 N_A_1369_93#_c_812_n N_A_1235_119#_c_1159_n 0.0504904f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_695 N_A_1369_93#_c_815_n N_A_1235_119#_c_1159_n 0.00751148f $X=7.235 $Y=1.02
+ $X2=0 $Y2=0
cc_696 N_A_1369_93#_M1006_g N_A_1235_119#_c_1189_n 0.011764f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_697 N_A_1369_93#_c_812_n N_A_1235_119#_c_1189_n 0.00251284f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_698 N_A_1369_93#_c_813_n N_A_1235_119#_c_1189_n 0.00224896f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_699 N_A_1369_93#_M1006_g N_A_1235_119#_c_1160_n 0.00479487f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_700 N_A_1369_93#_c_812_n N_A_1235_119#_c_1160_n 0.0170914f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_701 N_A_1369_93#_c_813_n N_A_1235_119#_c_1160_n 0.00155061f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_702 N_A_1369_93#_c_812_n N_A_1235_119#_c_1161_n 0.0228386f $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_703 N_A_1369_93#_c_813_n N_A_1235_119#_c_1161_n 7.19249e-19 $X=7.125 $Y=1.615
+ $X2=0 $Y2=0
cc_704 N_A_1369_93#_c_814_n N_A_1235_119#_c_1161_n 0.0135117f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_705 N_A_1369_93#_c_814_n N_A_1235_119#_c_1162_n 0.0516286f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_706 N_A_1369_93#_c_817_n N_A_1235_119#_c_1162_n 0.0120015f $X=8.81 $Y=1.415
+ $X2=0 $Y2=0
cc_707 N_A_1369_93#_c_818_n N_A_1235_119#_c_1162_n 0.00540759f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_708 N_A_1369_93#_M1006_g N_A_1235_119#_c_1168_n 0.00107811f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_709 N_A_1369_93#_c_814_n N_A_1235_119#_c_1163_n 0.00505406f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_710 N_A_1369_93#_c_817_n N_A_1235_119#_c_1163_n 0.0121855f $X=8.81 $Y=1.415
+ $X2=0 $Y2=0
cc_711 N_A_1369_93#_c_818_n N_A_1235_119#_c_1163_n 0.00825581f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_712 N_A_1369_93#_c_819_n N_A_1235_119#_c_1163_n 0.00275569f $X=8.445 $Y=1.02
+ $X2=0 $Y2=0
cc_713 N_A_1369_93#_M1006_g N_A_819_119#_M1024_g 0.0402741f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_714 N_A_1369_93#_M1006_g N_A_819_119#_c_1286_n 0.0120603f $X=6.955 $Y=2.525
+ $X2=0 $Y2=0
cc_715 N_A_1369_93#_c_818_n N_A_819_119#_c_1286_n 0.00262042f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_716 N_A_1369_93#_c_818_n N_A_819_119#_M1015_g 0.0145988f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_717 N_A_1369_93#_c_818_n N_A_819_119#_c_1275_n 0.00507363f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_718 N_A_1369_93#_c_818_n N_A_1747_74#_c_1615_n 0.0261048f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_719 N_A_1369_93#_c_818_n N_A_1747_74#_c_1610_n 0.0128087f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_720 N_A_1369_93#_M1006_g N_VPWR_c_1814_n 0.00393159f $X=6.955 $Y=2.525 $X2=0
+ $Y2=0
cc_721 N_A_1369_93#_c_814_n N_VPWR_c_1815_n 2.9437e-19 $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_722 N_A_1369_93#_c_817_n N_VPWR_c_1815_n 0.00213947f $X=8.81 $Y=1.415 $X2=0
+ $Y2=0
cc_723 N_A_1369_93#_c_818_n N_VPWR_c_1815_n 0.0357016f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_724 N_A_1369_93#_c_819_n N_VPWR_c_1815_n 0.00582847f $X=8.445 $Y=1.02 $X2=0
+ $Y2=0
cc_725 N_A_1369_93#_c_818_n N_VPWR_c_1828_n 0.0056446f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_726 N_A_1369_93#_M1006_g N_VPWR_c_1810_n 0.00112709f $X=6.955 $Y=2.525 $X2=0
+ $Y2=0
cc_727 N_A_1369_93#_c_818_n N_VPWR_c_1810_n 0.00682683f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_728 N_A_1369_93#_c_814_n N_VGND_M1034_d 0.0074698f $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_729 N_A_1369_93#_c_815_n A_1399_119# 0.00134092f $X=7.235 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_730 N_RESET_B_c_920_n N_A_1235_119#_M1041_g 0.0050753f $X=7.605 $Y=1.165
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_933_n N_A_1235_119#_M1007_g 0.00808965f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_RESET_B_M1034_g N_A_1235_119#_c_1158_n 8.68322e-19 $X=7.31 $Y=0.805
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_931_n N_A_1235_119#_c_1165_n 0.00851067f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_931_n N_A_1235_119#_c_1159_n 0.025309f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_931_n N_A_1235_119#_c_1189_n 0.0198099f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_RESET_B_M1040_g N_A_1235_119#_c_1160_n 0.0206938f $X=7.555 $Y=2.525
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_917_n N_A_1235_119#_c_1160_n 0.0101718f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_928_n N_A_1235_119#_c_1160_n 0.0173189f $X=7.465 $Y=2 $X2=0
+ $Y2=0
cc_739 N_RESET_B_c_931_n N_A_1235_119#_c_1160_n 0.0311602f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_934_n N_A_1235_119#_c_1160_n 0.00470341f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_939_n N_A_1235_119#_c_1160_n 0.0355881f $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_917_n N_A_1235_119#_c_1161_n 0.00434972f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_920_n N_A_1235_119#_c_1161_n 0.00295398f $X=7.605 $Y=1.165
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_917_n N_A_1235_119#_c_1162_n 0.00921867f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_745 N_RESET_B_c_931_n N_A_1235_119#_c_1162_n 0.00551265f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_933_n N_A_1235_119#_c_1162_n 0.00588285f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_934_n N_A_1235_119#_c_1162_n 0.0026603f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_938_n N_A_1235_119#_c_1162_n 0.00668769f $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_939_n N_A_1235_119#_c_1162_n 0.0134428f $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_917_n N_A_1235_119#_c_1163_n 0.0179208f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_933_n N_A_1235_119#_c_1163_n 0.00394795f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_934_n N_A_1235_119#_c_1163_n 7.15345e-19 $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_938_n N_A_1235_119#_c_1163_n 0.00483051f $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_939_n N_A_1235_119#_c_1163_n 5.47888e-19 $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_755 N_RESET_B_c_931_n N_A_819_119#_M1025_s 0.00116494f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_931_n N_A_819_119#_c_1270_n 0.00219472f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_914_n N_A_819_119#_c_1273_n 0.00882199f $X=7.235 $Y=0.18
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_931_n N_A_819_119#_M1024_g 0.00317501f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1040_g N_A_819_119#_c_1286_n 0.0119874f $X=7.555 $Y=2.525
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_933_n N_A_819_119#_M1015_g 0.011734f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_761 N_RESET_B_c_933_n N_A_819_119#_c_1274_n 0.0043462f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_914_n N_A_819_119#_c_1296_n 0.00142396f $X=7.235 $Y=0.18
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_931_n N_A_819_119#_c_1299_n 0.0225786f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_932_n N_A_819_119#_c_1291_n 5.46046e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_937_n N_A_819_119#_c_1291_n 0.00346024f $X=3.95 $Y=1.985
+ $X2=0 $Y2=0
cc_766 N_RESET_B_M1028_g N_A_819_119#_c_1305_n 0.00401892f $X=3.485 $Y=0.65
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_914_n N_A_819_119#_c_1305_n 0.00440229f $X=7.235 $Y=0.18
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_919_n N_A_819_119#_c_1305_n 4.31847e-19 $X=3.487 $Y=1.145
+ $X2=0 $Y2=0
cc_769 N_RESET_B_M1011_g N_A_819_119#_c_1308_n 0.00277356f $X=3.595 $Y=2.64
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_931_n N_A_819_119#_c_1308_n 0.0114462f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_932_n N_A_819_119#_c_1308_n 0.0020276f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_936_n N_A_819_119#_c_1308_n 5.9362e-19 $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_937_n N_A_819_119#_c_1308_n 0.0142721f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_931_n N_A_819_119#_c_1279_n 0.00588539f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_931_n N_A_819_119#_c_1280_n 5.3491e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_914_n N_A_819_119#_c_1281_n 0.0103518f $X=7.235 $Y=0.18 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_931_n N_A_819_119#_c_1294_n 0.00385098f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_778 N_RESET_B_M1009_g N_A_2008_48#_M1005_g 0.0358144f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_922_n N_A_2008_48#_M1005_g 0.00188557f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_780 N_RESET_B_c_921_n N_A_2008_48#_c_1459_n 0.0030428f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_933_n N_A_2008_48#_c_1459_n 0.00247648f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_782 RESET_B N_A_2008_48#_c_1459_n 7.14482e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_783 N_RESET_B_c_941_n N_A_2008_48#_c_1459_n 0.00169359f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_784 N_RESET_B_c_922_n N_A_2008_48#_c_1459_n 0.0249721f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_785 N_RESET_B_c_929_n N_A_2008_48#_M1039_g 0.00373821f $X=10.81 $Y=2.22 $X2=0
+ $Y2=0
cc_786 N_RESET_B_c_930_n N_A_2008_48#_M1039_g 0.0149506f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_787 N_RESET_B_c_933_n N_A_2008_48#_M1039_g 0.00762753f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_940_n N_A_2008_48#_M1039_g 6.88508e-19 $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_789 N_RESET_B_c_929_n N_A_2008_48#_c_1460_n 0.00199769f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_930_n N_A_2008_48#_c_1460_n 0.00241136f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_933_n N_A_2008_48#_c_1460_n 0.0174665f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_792 RESET_B N_A_2008_48#_c_1460_n 0.00269473f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_793 N_RESET_B_c_940_n N_A_2008_48#_c_1460_n 4.38169e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_941_n N_A_2008_48#_c_1460_n 0.0344591f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_795 N_RESET_B_c_922_n N_A_2008_48#_c_1460_n 2.34208e-19 $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_796 N_RESET_B_c_930_n N_A_2008_48#_c_1468_n 0.00995223f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_933_n N_A_2008_48#_c_1468_n 0.00560031f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_798 RESET_B N_A_2008_48#_c_1468_n 0.00309934f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_799 N_RESET_B_c_941_n N_A_2008_48#_c_1468_n 0.00989058f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_930_n N_A_2008_48#_c_1470_n 0.00721892f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_801 N_RESET_B_c_929_n N_A_2008_48#_c_1471_n 0.0015825f $X=10.81 $Y=2.22 $X2=0
+ $Y2=0
cc_802 N_RESET_B_c_930_n N_A_2008_48#_c_1471_n 5.62382e-19 $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_803 RESET_B N_A_2008_48#_c_1471_n 0.00125949f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_804 N_RESET_B_c_940_n N_A_2008_48#_c_1471_n 0.00110518f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_805 N_RESET_B_c_941_n N_A_2008_48#_c_1471_n 0.0258608f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_940_n N_A_2008_48#_c_1462_n 8.24141e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_807 N_RESET_B_c_941_n N_A_2008_48#_c_1462_n 0.00968802f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_808 N_RESET_B_c_922_n N_A_2008_48#_c_1462_n 0.00111902f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_930_n N_A_2008_48#_c_1474_n 0.00362988f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_810 RESET_B N_A_2008_48#_c_1474_n 7.29139e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_811 N_RESET_B_c_940_n N_A_2008_48#_c_1474_n 8.21335e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_812 N_RESET_B_c_941_n N_A_2008_48#_c_1474_n 0.0169044f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_813 N_RESET_B_M1009_g N_A_2008_48#_c_1464_n 0.00108873f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_814 N_RESET_B_c_933_n N_A_1747_74#_M1015_d 0.00138561f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_815 N_RESET_B_M1009_g N_A_1747_74#_c_1590_n 0.0481778f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_816 N_RESET_B_c_921_n N_A_1747_74#_c_1591_n 0.00304958f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_817 N_RESET_B_c_940_n N_A_1747_74#_c_1591_n 0.00202705f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_818 N_RESET_B_M1009_g N_A_1747_74#_c_1592_n 0.00503338f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_819 N_RESET_B_c_921_n N_A_1747_74#_c_1595_n 0.0113835f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_820 N_RESET_B_c_940_n N_A_1747_74#_c_1595_n 0.0205072f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_821 N_RESET_B_c_922_n N_A_1747_74#_c_1595_n 0.00965718f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_822 N_RESET_B_c_929_n N_A_1747_74#_c_1606_n 0.00655145f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_823 N_RESET_B_c_941_n N_A_1747_74#_c_1606_n 8.64724e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_824 N_RESET_B_c_930_n N_A_1747_74#_c_1607_n 0.0189805f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_825 N_RESET_B_c_933_n N_A_1747_74#_c_1615_n 0.0211312f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_826 N_RESET_B_c_930_n N_A_1747_74#_c_1609_n 7.97616e-19 $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_827 N_RESET_B_c_933_n N_A_1747_74#_c_1609_n 0.0153789f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_828 N_RESET_B_c_933_n N_A_1747_74#_c_1599_n 0.0224891f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_829 N_RESET_B_c_922_n N_A_1747_74#_c_1599_n 9.47605e-19 $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_830 N_RESET_B_M1009_g N_A_1747_74#_c_1601_n 0.0173454f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_831 N_RESET_B_c_921_n N_A_1747_74#_c_1601_n 0.0168092f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_832 N_RESET_B_c_933_n N_A_1747_74#_c_1601_n 0.0108974f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_833 RESET_B N_A_1747_74#_c_1601_n 0.00277891f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_834 N_RESET_B_c_940_n N_A_1747_74#_c_1601_n 0.00194273f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_835 N_RESET_B_c_941_n N_A_1747_74#_c_1601_n 0.0211796f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_836 N_RESET_B_c_922_n N_A_1747_74#_c_1601_n 0.00355179f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_837 N_RESET_B_c_931_n N_VPWR_M1025_d 3.376e-19 $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_838 N_RESET_B_c_933_n N_VPWR_M1007_s 0.00248619f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_839 N_RESET_B_M1011_g N_VPWR_c_1812_n 0.00502238f $X=3.595 $Y=2.64 $X2=0
+ $Y2=0
cc_840 N_RESET_B_M1040_g N_VPWR_c_1814_n 0.00391542f $X=7.555 $Y=2.525 $X2=0
+ $Y2=0
cc_841 N_RESET_B_c_931_n N_VPWR_c_1814_n 6.82537e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_842 N_RESET_B_M1040_g N_VPWR_c_1815_n 0.00605413f $X=7.555 $Y=2.525 $X2=0
+ $Y2=0
cc_843 N_RESET_B_c_917_n N_VPWR_c_1815_n 0.00159571f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_844 N_RESET_B_c_933_n N_VPWR_c_1815_n 0.025533f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_845 N_RESET_B_c_934_n N_VPWR_c_1815_n 0.00264729f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_846 N_RESET_B_c_938_n N_VPWR_c_1815_n 0.00113137f $X=7.86 $Y=1.985 $X2=0
+ $Y2=0
cc_847 N_RESET_B_c_939_n N_VPWR_c_1815_n 0.0204823f $X=7.86 $Y=1.985 $X2=0 $Y2=0
cc_848 N_RESET_B_c_930_n N_VPWR_c_1816_n 0.00483774f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_849 N_RESET_B_c_933_n N_VPWR_c_1816_n 0.00113818f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_850 N_RESET_B_M1011_g N_VPWR_c_1821_n 0.00474321f $X=3.595 $Y=2.64 $X2=0
+ $Y2=0
cc_851 N_RESET_B_c_930_n N_VPWR_c_1829_n 0.00586114f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_852 N_RESET_B_M1011_g N_VPWR_c_1810_n 0.0049737f $X=3.595 $Y=2.64 $X2=0 $Y2=0
cc_853 N_RESET_B_M1040_g N_VPWR_c_1810_n 0.00112709f $X=7.555 $Y=2.525 $X2=0
+ $Y2=0
cc_854 N_RESET_B_c_930_n N_VPWR_c_1810_n 0.00619157f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_855 N_RESET_B_c_927_n N_A_413_90#_c_2006_n 0.00109147f $X=3.415 $Y=1.82 $X2=0
+ $Y2=0
cc_856 N_RESET_B_M1028_g N_A_413_90#_c_1991_n 0.00805057f $X=3.485 $Y=0.65 $X2=0
+ $Y2=0
cc_857 N_RESET_B_c_919_n N_A_413_90#_c_1991_n 0.00814139f $X=3.487 $Y=1.145
+ $X2=0 $Y2=0
cc_858 N_RESET_B_c_913_n N_A_413_90#_c_1992_n 0.0197229f $X=3.49 $Y=1.82 $X2=0
+ $Y2=0
cc_859 N_RESET_B_M1011_g N_A_413_90#_c_1992_n 0.00921141f $X=3.595 $Y=2.64 $X2=0
+ $Y2=0
cc_860 N_RESET_B_c_919_n N_A_413_90#_c_1992_n 0.00216416f $X=3.487 $Y=1.145
+ $X2=0 $Y2=0
cc_861 N_RESET_B_c_927_n N_A_413_90#_c_1992_n 0.0138017f $X=3.415 $Y=1.82 $X2=0
+ $Y2=0
cc_862 N_RESET_B_c_932_n N_A_413_90#_c_1992_n 0.00108246f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_863 N_RESET_B_c_937_n N_A_413_90#_c_1992_n 0.0228178f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_864 N_RESET_B_c_931_n N_A_413_90#_c_1999_n 0.016634f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_865 N_RESET_B_c_932_n N_A_413_90#_c_1999_n 0.00665688f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_866 N_RESET_B_c_936_n N_A_413_90#_c_1999_n 0.00191895f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_867 N_RESET_B_c_937_n N_A_413_90#_c_1999_n 0.0064556f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_868 N_RESET_B_c_931_n N_A_413_90#_c_2000_n 0.00166662f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_869 N_RESET_B_c_931_n N_A_413_90#_c_2001_n 0.0199643f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_870 N_RESET_B_c_931_n N_A_413_90#_c_2002_n 0.0117838f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_871 N_RESET_B_c_931_n N_A_413_90#_c_1996_n 0.0113119f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_872 N_RESET_B_M1011_g N_A_413_90#_c_2005_n 0.0225344f $X=3.595 $Y=2.64 $X2=0
+ $Y2=0
cc_873 N_RESET_B_c_932_n N_A_413_90#_c_2005_n 0.00122942f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_874 N_RESET_B_c_936_n N_A_413_90#_c_2005_n 0.00741283f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_875 N_RESET_B_c_937_n N_A_413_90#_c_2005_n 0.0158802f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_876 N_RESET_B_M1028_g N_VGND_c_2180_n 0.00438348f $X=3.485 $Y=0.65 $X2=0
+ $Y2=0
cc_877 N_RESET_B_c_914_n N_VGND_c_2180_n 0.021597f $X=7.235 $Y=0.18 $X2=0 $Y2=0
cc_878 N_RESET_B_c_914_n N_VGND_c_2181_n 0.0252774f $X=7.235 $Y=0.18 $X2=0 $Y2=0
cc_879 N_RESET_B_c_914_n N_VGND_c_2182_n 0.00986746f $X=7.235 $Y=0.18 $X2=0
+ $Y2=0
cc_880 N_RESET_B_M1009_g N_VGND_c_2183_n 0.0110663f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_881 N_RESET_B_c_914_n N_VGND_c_2186_n 0.0250888f $X=7.235 $Y=0.18 $X2=0 $Y2=0
cc_882 N_RESET_B_c_915_n N_VGND_c_2189_n 0.00583607f $X=3.56 $Y=0.18 $X2=0 $Y2=0
cc_883 N_RESET_B_c_914_n N_VGND_c_2190_n 0.0526108f $X=7.235 $Y=0.18 $X2=0 $Y2=0
cc_884 N_RESET_B_M1009_g N_VGND_c_2192_n 0.00383152f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_885 N_RESET_B_c_914_n N_VGND_c_2194_n 0.0925762f $X=7.235 $Y=0.18 $X2=0 $Y2=0
cc_886 N_RESET_B_c_915_n N_VGND_c_2194_n 0.0113334f $X=3.56 $Y=0.18 $X2=0 $Y2=0
cc_887 N_RESET_B_M1009_g N_VGND_c_2194_n 0.0075694f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_888 N_RESET_B_M1028_g N_noxref_25_c_2320_n 0.00320551f $X=3.485 $Y=0.65 $X2=0
+ $Y2=0
cc_889 N_A_1235_119#_c_1165_n N_A_819_119#_c_1283_n 0.00357117f $X=6.675
+ $Y=2.585 $X2=0 $Y2=0
cc_890 N_A_1235_119#_c_1158_n N_A_819_119#_c_1273_n 0.00402473f $X=6.675 $Y=0.76
+ $X2=0 $Y2=0
cc_891 N_A_1235_119#_c_1165_n N_A_819_119#_M1024_g 0.0142007f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_892 N_A_1235_119#_c_1159_n N_A_819_119#_M1024_g 0.00208145f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_893 N_A_1235_119#_M1007_g N_A_819_119#_c_1286_n 0.0123711f $X=8.545 $Y=2.235
+ $X2=0 $Y2=0
cc_894 N_A_1235_119#_c_1189_n N_A_819_119#_c_1286_n 0.00152355f $X=7.405
+ $Y=2.405 $X2=0 $Y2=0
cc_895 N_A_1235_119#_c_1160_n N_A_819_119#_c_1286_n 0.00646428f $X=7.49 $Y=2.32
+ $X2=0 $Y2=0
cc_896 N_A_1235_119#_c_1168_n N_A_819_119#_c_1286_n 0.00202544f $X=6.76 $Y=2.537
+ $X2=0 $Y2=0
cc_897 N_A_1235_119#_M1007_g N_A_819_119#_M1015_g 0.0080851f $X=8.545 $Y=2.235
+ $X2=0 $Y2=0
cc_898 N_A_1235_119#_c_1163_n N_A_819_119#_c_1275_n 0.0080851f $X=8.23 $Y=1.42
+ $X2=0 $Y2=0
cc_899 N_A_1235_119#_c_1189_n N_VPWR_M1006_d 0.00711651f $X=7.405 $Y=2.405 $X2=0
+ $Y2=0
cc_900 N_A_1235_119#_c_1189_n N_VPWR_c_1814_n 0.0233006f $X=7.405 $Y=2.405 $X2=0
+ $Y2=0
cc_901 N_A_1235_119#_c_1160_n N_VPWR_c_1814_n 0.00393012f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_902 N_A_1235_119#_c_1168_n N_VPWR_c_1814_n 0.00129738f $X=6.76 $Y=2.537 $X2=0
+ $Y2=0
cc_903 N_A_1235_119#_M1007_g N_VPWR_c_1815_n 0.0174235f $X=8.545 $Y=2.235 $X2=0
+ $Y2=0
cc_904 N_A_1235_119#_c_1160_n N_VPWR_c_1815_n 0.0313212f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_905 N_A_1235_119#_c_1162_n N_VPWR_c_1815_n 0.00271335f $X=8.105 $Y=1.41 $X2=0
+ $Y2=0
cc_906 N_A_1235_119#_c_1163_n N_VPWR_c_1815_n 0.00636177f $X=8.23 $Y=1.42 $X2=0
+ $Y2=0
cc_907 N_A_1235_119#_c_1165_n N_VPWR_c_1823_n 0.010458f $X=6.675 $Y=2.585 $X2=0
+ $Y2=0
cc_908 N_A_1235_119#_c_1168_n N_VPWR_c_1823_n 0.00389335f $X=6.76 $Y=2.537 $X2=0
+ $Y2=0
cc_909 N_A_1235_119#_c_1160_n N_VPWR_c_1827_n 0.00728415f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_910 N_A_1235_119#_M1007_g N_VPWR_c_1810_n 9.455e-19 $X=8.545 $Y=2.235 $X2=0
+ $Y2=0
cc_911 N_A_1235_119#_c_1165_n N_VPWR_c_1810_n 0.0131156f $X=6.675 $Y=2.585 $X2=0
+ $Y2=0
cc_912 N_A_1235_119#_c_1189_n N_VPWR_c_1810_n 0.00795073f $X=7.405 $Y=2.405
+ $X2=0 $Y2=0
cc_913 N_A_1235_119#_c_1160_n N_VPWR_c_1810_n 0.0151926f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_914 N_A_1235_119#_c_1168_n N_VPWR_c_1810_n 0.00470184f $X=6.76 $Y=2.537 $X2=0
+ $Y2=0
cc_915 N_A_1235_119#_c_1165_n N_A_413_90#_c_2000_n 0.01209f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_916 N_A_1235_119#_c_1165_n N_A_413_90#_c_2001_n 0.0210346f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_917 N_A_1235_119#_c_1159_n N_A_413_90#_c_2001_n 0.0137765f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_918 N_A_1235_119#_c_1158_n N_A_413_90#_c_1994_n 0.0239547f $X=6.675 $Y=0.76
+ $X2=0 $Y2=0
cc_919 N_A_1235_119#_c_1159_n N_A_413_90#_c_1994_n 0.0136236f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_920 N_A_1235_119#_c_1159_n N_A_413_90#_c_1996_n 0.0586249f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_921 N_A_1235_119#_M1041_g N_VGND_c_2182_n 0.00117551f $X=8.23 $Y=0.69 $X2=0
+ $Y2=0
cc_922 N_A_1235_119#_M1041_g N_VGND_c_2191_n 0.00278271f $X=8.23 $Y=0.69 $X2=0
+ $Y2=0
cc_923 N_A_1235_119#_M1041_g N_VGND_c_2194_n 0.00358525f $X=8.23 $Y=0.69 $X2=0
+ $Y2=0
cc_924 N_A_1235_119#_c_1158_n A_1321_119# 0.00165713f $X=6.675 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_925 N_A_1235_119#_c_1159_n A_1321_119# 9.96634e-19 $X=6.76 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_926 N_A_819_119#_M1016_g N_A_2008_48#_M1005_g 0.0422064f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_927 N_A_819_119#_c_1274_n N_A_2008_48#_c_1459_n 0.0427595f $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_928 N_A_819_119#_M1015_g N_A_1747_74#_c_1615_n 2.54907e-19 $X=8.995 $Y=2.235
+ $X2=0 $Y2=0
cc_929 N_A_819_119#_c_1274_n N_A_1747_74#_c_1615_n 0.00468179f $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_930 N_A_819_119#_M1016_g N_A_1747_74#_c_1619_n 0.0150881f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_931 N_A_819_119#_M1015_g N_A_1747_74#_c_1610_n 0.00218567f $X=8.995 $Y=2.235
+ $X2=0 $Y2=0
cc_932 N_A_819_119#_M1016_g N_A_1747_74#_c_1598_n 0.00884302f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_933 N_A_819_119#_M1016_g N_A_1747_74#_c_1599_n 0.0014557f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_934 N_A_819_119#_c_1274_n N_A_1747_74#_c_1600_n 4.03784e-19 $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_935 N_A_819_119#_M1016_g N_A_1747_74#_c_1600_n 0.0141061f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_936 N_A_819_119#_c_1299_n N_VPWR_M1025_d 0.00325331f $X=4.815 $Y=2.03 $X2=0
+ $Y2=0
cc_937 N_A_819_119#_c_1270_n N_VPWR_c_1813_n 0.00211235f $X=5.605 $Y=3.075 $X2=0
+ $Y2=0
cc_938 N_A_819_119#_c_1284_n N_VPWR_c_1813_n 7.02368e-19 $X=5.68 $Y=3.15 $X2=0
+ $Y2=0
cc_939 N_A_819_119#_c_1294_n N_VPWR_c_1813_n 0.0105232f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_940 N_A_819_119#_M1024_g N_VPWR_c_1814_n 0.00617223f $X=6.565 $Y=2.525 $X2=0
+ $Y2=0
cc_941 N_A_819_119#_c_1286_n N_VPWR_c_1814_n 0.0253641f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_942 N_A_819_119#_c_1286_n N_VPWR_c_1815_n 0.0210786f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_943 N_A_819_119#_M1015_g N_VPWR_c_1815_n 0.00681114f $X=8.995 $Y=2.235 $X2=0
+ $Y2=0
cc_944 N_A_819_119#_c_1284_n N_VPWR_c_1823_n 0.0448726f $X=5.68 $Y=3.15 $X2=0
+ $Y2=0
cc_945 N_A_819_119#_c_1294_n N_VPWR_c_1823_n 0.00401239f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_946 N_A_819_119#_c_1286_n N_VPWR_c_1827_n 0.0250026f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_947 N_A_819_119#_c_1286_n N_VPWR_c_1828_n 0.0193431f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_948 N_A_819_119#_c_1283_n N_VPWR_c_1810_n 0.0234229f $X=6.475 $Y=3.15 $X2=0
+ $Y2=0
cc_949 N_A_819_119#_c_1284_n N_VPWR_c_1810_n 0.00588524f $X=5.68 $Y=3.15 $X2=0
+ $Y2=0
cc_950 N_A_819_119#_c_1286_n N_VPWR_c_1810_n 0.0674076f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_951 N_A_819_119#_c_1290_n N_VPWR_c_1810_n 0.00500367f $X=6.565 $Y=3.15 $X2=0
+ $Y2=0
cc_952 N_A_819_119#_c_1294_n N_VPWR_c_1810_n 0.00500915f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_953 N_A_819_119#_c_1305_n N_A_413_90#_c_1991_n 0.00323663f $X=4.49 $Y=0.802
+ $X2=0 $Y2=0
cc_954 N_A_819_119#_M1025_s N_A_413_90#_c_1999_n 0.00770925f $X=4.275 $Y=1.935
+ $X2=0 $Y2=0
cc_955 N_A_819_119#_c_1270_n N_A_413_90#_c_1999_n 0.0134859f $X=5.605 $Y=3.075
+ $X2=0 $Y2=0
cc_956 N_A_819_119#_c_1299_n N_A_413_90#_c_1999_n 0.0110961f $X=4.815 $Y=2.03
+ $X2=0 $Y2=0
cc_957 N_A_819_119#_c_1308_n N_A_413_90#_c_1999_n 0.0137082f $X=4.46 $Y=2.03
+ $X2=0 $Y2=0
cc_958 N_A_819_119#_c_1279_n N_A_413_90#_c_1999_n 0.00140597f $X=5.13 $Y=1.61
+ $X2=0 $Y2=0
cc_959 N_A_819_119#_c_1294_n N_A_413_90#_c_1999_n 0.0160652f $X=5.13 $Y=1.86
+ $X2=0 $Y2=0
cc_960 N_A_819_119#_c_1270_n N_A_413_90#_c_2000_n 0.0076682f $X=5.605 $Y=3.075
+ $X2=0 $Y2=0
cc_961 N_A_819_119#_c_1283_n N_A_413_90#_c_2000_n 0.00412947f $X=6.475 $Y=3.15
+ $X2=0 $Y2=0
cc_962 N_A_819_119#_c_1271_n N_A_413_90#_c_1993_n 0.00406792f $X=6.025 $Y=1.165
+ $X2=0 $Y2=0
cc_963 N_A_819_119#_c_1273_n N_A_413_90#_c_1993_n 0.00350442f $X=6.1 $Y=1.09
+ $X2=0 $Y2=0
cc_964 N_A_819_119#_M1024_g N_A_413_90#_c_2001_n 0.0023028f $X=6.565 $Y=2.525
+ $X2=0 $Y2=0
cc_965 N_A_819_119#_c_1270_n N_A_413_90#_c_2002_n 0.0012967f $X=5.605 $Y=3.075
+ $X2=0 $Y2=0
cc_966 N_A_819_119#_c_1271_n N_A_413_90#_c_1994_n 0.00971137f $X=6.025 $Y=1.165
+ $X2=0 $Y2=0
cc_967 N_A_819_119#_c_1271_n N_A_413_90#_c_1995_n 0.00629199f $X=6.025 $Y=1.165
+ $X2=0 $Y2=0
cc_968 N_A_819_119#_c_1269_n N_A_413_90#_c_1996_n 0.00572173f $X=5.605 $Y=1.41
+ $X2=0 $Y2=0
cc_969 N_A_819_119#_c_1296_n N_VGND_M1013_d 0.00857319f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_970 N_A_819_119#_c_1278_n N_VGND_M1013_d 0.005277f $X=4.9 $Y=1.445 $X2=0
+ $Y2=0
cc_971 N_A_819_119#_c_1305_n N_VGND_c_2180_n 0.00723274f $X=4.49 $Y=0.802 $X2=0
+ $Y2=0
cc_972 N_A_819_119#_c_1296_n N_VGND_c_2181_n 0.0255675f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_973 N_A_819_119#_c_1281_n N_VGND_c_2181_n 0.0016944f $X=5.13 $Y=1.41 $X2=0
+ $Y2=0
cc_974 N_A_819_119#_M1016_g N_VGND_c_2183_n 0.00177088f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_975 N_A_819_119#_c_1305_n N_VGND_c_2186_n 0.00480704f $X=4.49 $Y=0.802 $X2=0
+ $Y2=0
cc_976 N_A_819_119#_M1016_g N_VGND_c_2191_n 0.00358451f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_977 N_A_819_119#_M1016_g N_VGND_c_2194_n 0.00569641f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_978 N_A_819_119#_c_1296_n N_VGND_c_2194_n 0.00593113f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_979 N_A_819_119#_c_1305_n N_VGND_c_2194_n 0.00701863f $X=4.49 $Y=0.802 $X2=0
+ $Y2=0
cc_980 N_A_819_119#_c_1281_n N_VGND_c_2194_n 8.47775e-19 $X=5.13 $Y=1.41 $X2=0
+ $Y2=0
cc_981 N_A_2008_48#_c_1463_n N_A_1747_74#_c_1590_n 0.0023753f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_982 N_A_2008_48#_c_1464_n N_A_1747_74#_c_1590_n 0.00741302f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_983 N_A_2008_48#_c_1461_n N_A_1747_74#_c_1591_n 0.00406259f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_984 N_A_2008_48#_c_1463_n N_A_1747_74#_c_1591_n 0.00385495f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_985 N_A_2008_48#_c_1464_n N_A_1747_74#_c_1591_n 0.00768727f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_986 N_A_2008_48#_c_1471_n N_A_1747_74#_M1026_g 6.65497e-19 $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_987 N_A_2008_48#_c_1472_n N_A_1747_74#_M1026_g 0.00349104f $X=11.675 $Y=1.715
+ $X2=0 $Y2=0
cc_988 N_A_2008_48#_c_1463_n N_A_1747_74#_c_1593_n 0.00507794f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_989 N_A_2008_48#_c_1464_n N_A_1747_74#_c_1593_n 0.00413357f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_990 N_A_2008_48#_c_1461_n N_A_1747_74#_c_1595_n 0.00447579f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_991 N_A_2008_48#_c_1472_n N_A_1747_74#_c_1595_n 0.0175993f $X=11.675 $Y=1.715
+ $X2=0 $Y2=0
cc_992 N_A_2008_48#_c_1462_n N_A_1747_74#_c_1595_n 0.00406088f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_993 N_A_2008_48#_c_1463_n N_A_1747_74#_c_1595_n 0.0258377f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_994 N_A_2008_48#_c_1471_n N_A_1747_74#_c_1606_n 0.0105602f $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_995 N_A_2008_48#_c_1472_n N_A_1747_74#_c_1606_n 0.00280977f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_996 N_A_2008_48#_c_1462_n N_A_1747_74#_c_1606_n 0.00167941f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_997 N_A_2008_48#_c_1470_n N_A_1747_74#_c_1607_n 0.00645245f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_998 N_A_2008_48#_c_1471_n N_A_1747_74#_c_1607_n 0.00434752f $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_999 N_A_2008_48#_c_1474_n N_A_1747_74#_c_1607_n 0.0142091f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1000 N_A_2008_48#_M1005_g N_A_1747_74#_c_1619_n 0.00100268f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1001 N_A_2008_48#_M1039_g N_A_1747_74#_c_1609_n 0.00925232f $X=10.16 $Y=2.655
+ $X2=0 $Y2=0
cc_1002 N_A_2008_48#_c_1469_n N_A_1747_74#_c_1609_n 0.00364064f $X=10.525
+ $Y=2.405 $X2=0 $Y2=0
cc_1003 N_A_2008_48#_M1005_g N_A_1747_74#_c_1598_n 0.00151652f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1004 N_A_2008_48#_M1005_g N_A_1747_74#_c_1599_n 0.00175137f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1005 N_A_2008_48#_c_1459_n N_A_1747_74#_c_1599_n 0.0146343f $X=10.16 $Y=1.98
+ $X2=0 $Y2=0
cc_1006 N_A_2008_48#_M1039_g N_A_1747_74#_c_1599_n 0.00699016f $X=10.16 $Y=2.655
+ $X2=0 $Y2=0
cc_1007 N_A_2008_48#_c_1460_n N_A_1747_74#_c_1599_n 0.0472741f $X=10.36 $Y=1.815
+ $X2=0 $Y2=0
cc_1008 N_A_2008_48#_c_1469_n N_A_1747_74#_c_1599_n 0.00843626f $X=10.525
+ $Y=2.405 $X2=0 $Y2=0
cc_1009 N_A_2008_48#_M1005_g N_A_1747_74#_c_1600_n 0.00782885f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1010 N_A_2008_48#_M1005_g N_A_1747_74#_c_1601_n 0.0151836f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1011 N_A_2008_48#_c_1459_n N_A_1747_74#_c_1601_n 0.00516648f $X=10.16 $Y=1.98
+ $X2=0 $Y2=0
cc_1012 N_A_2008_48#_c_1460_n N_A_1747_74#_c_1601_n 0.0174506f $X=10.36 $Y=1.815
+ $X2=0 $Y2=0
cc_1013 N_A_2008_48#_c_1461_n N_A_1747_74#_c_1601_n 0.00792529f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_1014 N_A_2008_48#_c_1472_n N_A_1747_74#_c_1601_n 0.00127707f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_1015 N_A_2008_48#_c_1462_n N_A_1747_74#_c_1601_n 0.0125719f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_1016 N_A_2008_48#_c_1463_n N_A_1747_74#_c_1601_n 0.0245935f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1017 N_A_2008_48#_c_1464_n N_A_1747_74#_c_1601_n 0.017591f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_1018 N_A_2008_48#_c_1468_n N_VPWR_M1039_d 0.00127931f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1019 N_A_2008_48#_c_1469_n N_VPWR_M1039_d 0.00292266f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1020 N_A_2008_48#_c_1474_n N_VPWR_M1021_d 5.96727e-19 $X=11.13 $Y=2.405 $X2=0
+ $Y2=0
cc_1021 N_A_2008_48#_c_1459_n N_VPWR_c_1816_n 6.36779e-19 $X=10.16 $Y=1.98 $X2=0
+ $Y2=0
cc_1022 N_A_2008_48#_M1039_g N_VPWR_c_1816_n 0.0052036f $X=10.16 $Y=2.655 $X2=0
+ $Y2=0
cc_1023 N_A_2008_48#_c_1468_n N_VPWR_c_1816_n 0.00943806f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1024 N_A_2008_48#_c_1469_n N_VPWR_c_1816_n 0.0186301f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1025 N_A_2008_48#_c_1470_n N_VPWR_c_1816_n 0.00796567f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1026 N_A_2008_48#_c_1470_n N_VPWR_c_1930_n 0.00796754f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1027 N_A_2008_48#_c_1471_n N_VPWR_c_1930_n 0.0240111f $X=11.32 $Y=2.32 $X2=0
+ $Y2=0
cc_1028 N_A_2008_48#_c_1472_n N_VPWR_c_1930_n 0.0184768f $X=11.675 $Y=1.715
+ $X2=0 $Y2=0
cc_1029 N_A_2008_48#_c_1474_n N_VPWR_c_1930_n 0.0135228f $X=11.13 $Y=2.405 $X2=0
+ $Y2=0
cc_1030 N_A_2008_48#_c_1470_n N_VPWR_c_1825_n 0.00744121f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1031 N_A_2008_48#_c_1474_n N_VPWR_c_1825_n 9.81877e-19 $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1032 N_A_2008_48#_M1039_g N_VPWR_c_1828_n 0.00591817f $X=10.16 $Y=2.655 $X2=0
+ $Y2=0
cc_1033 N_A_2008_48#_c_1470_n N_VPWR_c_1829_n 0.0102777f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1034 N_A_2008_48#_M1039_g N_VPWR_c_1810_n 0.00619157f $X=10.16 $Y=2.655 $X2=0
+ $Y2=0
cc_1035 N_A_2008_48#_c_1468_n N_VPWR_c_1810_n 0.00699598f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1036 N_A_2008_48#_c_1469_n N_VPWR_c_1810_n 0.00241369f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1037 N_A_2008_48#_c_1470_n N_VPWR_c_1810_n 0.0112587f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1038 N_A_2008_48#_c_1474_n N_VPWR_c_1810_n 0.00666881f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1039 N_A_2008_48#_c_1471_n Q_N 0.00449177f $X=11.32 $Y=2.32 $X2=0 $Y2=0
cc_1040 N_A_2008_48#_c_1472_n Q_N 0.0138803f $X=11.675 $Y=1.715 $X2=0 $Y2=0
cc_1041 N_A_2008_48#_c_1463_n Q_N 0.0510002f $X=11.76 $Y=1.63 $X2=0 $Y2=0
cc_1042 N_A_2008_48#_c_1461_n N_VGND_M1010_s 0.00795702f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1043 N_A_2008_48#_c_1463_n N_VGND_M1010_s 0.00751007f $X=11.76 $Y=1.63 $X2=0
+ $Y2=0
cc_1044 N_A_2008_48#_M1005_g N_VGND_c_2183_n 0.0106684f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1045 N_A_2008_48#_c_1464_n N_VGND_c_2183_n 0.0133829f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1046 N_A_2008_48#_M1005_g N_VGND_c_2191_n 0.00383152f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1047 N_A_2008_48#_c_1461_n N_VGND_c_2192_n 0.00463151f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1048 N_A_2008_48#_c_1464_n N_VGND_c_2192_n 0.0140232f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1049 N_A_2008_48#_M1005_g N_VGND_c_2194_n 0.0075694f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1050 N_A_2008_48#_c_1461_n N_VGND_c_2194_n 0.00869887f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1051 N_A_2008_48#_c_1464_n N_VGND_c_2194_n 0.0117897f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1052 N_A_2008_48#_c_1461_n N_VGND_c_2199_n 0.0253659f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1053 N_A_2008_48#_c_1464_n N_VGND_c_2199_n 0.00410713f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1054 N_A_1747_74#_M1003_g N_A_2513_424#_M1037_g 0.0206457f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1055 N_A_1747_74#_c_1597_n N_A_2513_424#_M1000_g 0.0170449f $X=12.915 $Y=1.52
+ $X2=0 $Y2=0
cc_1056 N_A_1747_74#_c_1593_n N_A_2513_424#_c_1762_n 0.00194375f $X=11.965
+ $Y=1.235 $X2=0 $Y2=0
cc_1057 N_A_1747_74#_M1003_g N_A_2513_424#_c_1762_n 0.0144342f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1058 N_A_1747_74#_c_1594_n N_A_2513_424#_c_1767_n 0.00619956f $X=12.825
+ $Y=1.52 $X2=0 $Y2=0
cc_1059 N_A_1747_74#_M1008_g N_A_2513_424#_c_1767_n 0.0285135f $X=12.915 $Y=2.54
+ $X2=0 $Y2=0
cc_1060 N_A_1747_74#_c_1597_n N_A_2513_424#_c_1767_n 0.00107618f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1061 N_A_1747_74#_M1003_g N_A_2513_424#_c_1763_n 0.00833371f $X=12.93
+ $Y=0.645 $X2=0 $Y2=0
cc_1062 N_A_1747_74#_c_1597_n N_A_2513_424#_c_1763_n 0.0134747f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1063 N_A_1747_74#_M1003_g N_A_2513_424#_c_1764_n 0.0214527f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1064 N_A_1747_74#_c_1594_n N_A_2513_424#_c_1765_n 0.0160204f $X=12.825
+ $Y=1.52 $X2=0 $Y2=0
cc_1065 N_A_1747_74#_c_1595_n N_A_2513_424#_c_1765_n 2.29508e-19 $X=12.04
+ $Y=1.52 $X2=0 $Y2=0
cc_1066 N_A_1747_74#_M1003_g N_A_2513_424#_c_1765_n 0.00105416f $X=12.93
+ $Y=0.645 $X2=0 $Y2=0
cc_1067 N_A_1747_74#_c_1597_n N_A_2513_424#_c_1765_n 7.76856e-19 $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1068 N_A_1747_74#_M1026_g N_VPWR_c_1817_n 0.00730664f $X=11.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1069 N_A_1747_74#_c_1595_n N_VPWR_c_1930_n 9.58405e-19 $X=12.04 $Y=1.52 $X2=0
+ $Y2=0
cc_1070 N_A_1747_74#_c_1606_n N_VPWR_c_1930_n 0.00300744f $X=11.29 $Y=2.22 $X2=0
+ $Y2=0
cc_1071 N_A_1747_74#_c_1607_n N_VPWR_c_1930_n 0.00229229f $X=11.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1072 N_A_1747_74#_M1008_g N_VPWR_c_1818_n 0.00646597f $X=12.915 $Y=2.54 $X2=0
+ $Y2=0
cc_1073 N_A_1747_74#_c_1607_n N_VPWR_c_1825_n 0.00599998f $X=11.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1074 N_A_1747_74#_c_1609_n N_VPWR_c_1828_n 0.0143964f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1075 N_A_1747_74#_c_1610_n N_VPWR_c_1828_n 0.00507318f $X=9.325 $Y=2.59 $X2=0
+ $Y2=0
cc_1076 N_A_1747_74#_c_1607_n N_VPWR_c_1829_n 0.00586114f $X=11.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1077 N_A_1747_74#_M1026_g N_VPWR_c_1830_n 0.00553757f $X=11.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1078 N_A_1747_74#_M1008_g N_VPWR_c_1830_n 0.005209f $X=12.915 $Y=2.54 $X2=0
+ $Y2=0
cc_1079 N_A_1747_74#_M1026_g N_VPWR_c_1810_n 0.0109825f $X=11.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1080 N_A_1747_74#_M1008_g N_VPWR_c_1810_n 0.00987912f $X=12.915 $Y=2.54 $X2=0
+ $Y2=0
cc_1081 N_A_1747_74#_c_1607_n N_VPWR_c_1810_n 0.00619157f $X=11.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1082 N_A_1747_74#_c_1609_n N_VPWR_c_1810_n 0.023561f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1083 N_A_1747_74#_c_1610_n N_VPWR_c_1810_n 0.00697584f $X=9.325 $Y=2.59 $X2=0
+ $Y2=0
cc_1084 N_A_1747_74#_c_1609_n A_1972_489# 0.00160657f $X=9.925 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_1085 N_A_1747_74#_M1026_g Q_N 0.00522079f $X=11.925 $Y=2.4 $X2=0 $Y2=0
cc_1086 N_A_1747_74#_c_1593_n Q_N 0.0192064f $X=11.965 $Y=1.235 $X2=0 $Y2=0
cc_1087 N_A_1747_74#_c_1594_n Q_N 0.0259435f $X=12.825 $Y=1.52 $X2=0 $Y2=0
cc_1088 N_A_1747_74#_c_1595_n Q_N 0.00977739f $X=12.04 $Y=1.52 $X2=0 $Y2=0
cc_1089 N_A_1747_74#_M1008_g Q_N 0.00389012f $X=12.915 $Y=2.54 $X2=0 $Y2=0
cc_1090 N_A_1747_74#_M1003_g Q_N 0.00438444f $X=12.93 $Y=0.645 $X2=0 $Y2=0
cc_1091 N_A_1747_74#_c_1590_n N_VGND_c_2183_n 0.00170773f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1092 N_A_1747_74#_c_1619_n N_VGND_c_2183_n 0.0133993f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1093 N_A_1747_74#_c_1598_n N_VGND_c_2183_n 8.97539e-19 $X=9.69 $Y=1.005 $X2=0
+ $Y2=0
cc_1094 N_A_1747_74#_c_1601_n N_VGND_c_2183_n 0.0179642f $X=11.26 $Y=1.27 $X2=0
+ $Y2=0
cc_1095 N_A_1747_74#_c_1593_n N_VGND_c_2184_n 0.00434272f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1096 N_A_1747_74#_M1003_g N_VGND_c_2184_n 0.00461464f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1097 N_A_1747_74#_M1003_g N_VGND_c_2185_n 0.0103391f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1098 N_A_1747_74#_c_1619_n N_VGND_c_2191_n 0.0207002f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1099 N_A_1747_74#_c_1590_n N_VGND_c_2192_n 0.00434272f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1100 N_A_1747_74#_c_1590_n N_VGND_c_2194_n 0.00825669f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1101 N_A_1747_74#_c_1593_n N_VGND_c_2194_n 0.0083017f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1102 N_A_1747_74#_M1003_g N_VGND_c_2194_n 0.00914946f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1103 N_A_1747_74#_c_1619_n N_VGND_c_2194_n 0.0219224f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1104 N_A_1747_74#_c_1590_n N_VGND_c_2199_n 0.00289541f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1105 N_A_1747_74#_c_1593_n N_VGND_c_2199_n 0.00583402f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1106 N_A_2513_424#_M1000_g N_VPWR_c_1818_n 0.00378136f $X=13.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1107 N_A_2513_424#_c_1767_n N_VPWR_c_1818_n 0.0508632f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1108 N_A_2513_424#_c_1763_n N_VPWR_c_1818_n 0.0222736f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1109 N_A_2513_424#_c_1764_n N_VPWR_c_1818_n 0.00251384f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1110 N_A_2513_424#_c_1767_n N_VPWR_c_1830_n 0.012541f $X=12.69 $Y=2.265 $X2=0
+ $Y2=0
cc_1111 N_A_2513_424#_M1000_g N_VPWR_c_1831_n 0.00553757f $X=13.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1112 N_A_2513_424#_M1000_g N_VPWR_c_1810_n 0.0109239f $X=13.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1113 N_A_2513_424#_c_1767_n N_VPWR_c_1810_n 0.0103123f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1114 N_A_2513_424#_c_1762_n Q_N 0.0571733f $X=12.715 $Y=0.645 $X2=0 $Y2=0
cc_1115 N_A_2513_424#_c_1767_n Q_N 0.0895803f $X=12.69 $Y=2.265 $X2=0 $Y2=0
cc_1116 N_A_2513_424#_c_1765_n Q_N 0.0215198f $X=12.712 $Y=1.465 $X2=0 $Y2=0
cc_1117 N_A_2513_424#_M1037_g Q 0.00811057f $X=13.42 $Y=0.74 $X2=0 $Y2=0
cc_1118 N_A_2513_424#_M1037_g Q 0.00301691f $X=13.42 $Y=0.74 $X2=0 $Y2=0
cc_1119 N_A_2513_424#_c_1763_n Q 0.00111755f $X=13.38 $Y=1.465 $X2=0 $Y2=0
cc_1120 N_A_2513_424#_c_1764_n Q 0.00234039f $X=13.38 $Y=1.465 $X2=0 $Y2=0
cc_1121 N_A_2513_424#_M1000_g Q 0.00201151f $X=13.435 $Y=2.4 $X2=0 $Y2=0
cc_1122 N_A_2513_424#_M1037_g N_Q_c_2160_n 0.0040915f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1123 N_A_2513_424#_M1000_g N_Q_c_2160_n 0.00503704f $X=13.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1124 N_A_2513_424#_c_1763_n N_Q_c_2160_n 0.0250949f $X=13.38 $Y=1.465 $X2=0
+ $Y2=0
cc_1125 N_A_2513_424#_c_1764_n N_Q_c_2160_n 0.00791816f $X=13.38 $Y=1.465 $X2=0
+ $Y2=0
cc_1126 N_A_2513_424#_c_1762_n N_VGND_c_2184_n 0.00778672f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1127 N_A_2513_424#_M1037_g N_VGND_c_2185_n 0.00330159f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1128 N_A_2513_424#_c_1762_n N_VGND_c_2185_n 0.035427f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1129 N_A_2513_424#_c_1763_n N_VGND_c_2185_n 0.0145561f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1130 N_A_2513_424#_c_1764_n N_VGND_c_2185_n 0.00172388f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1131 N_A_2513_424#_M1037_g N_VGND_c_2193_n 0.00434272f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1132 N_A_2513_424#_M1037_g N_VGND_c_2194_n 0.00824587f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1133 N_A_2513_424#_c_1762_n N_VGND_c_2194_n 0.00976756f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1134 N_VPWR_M1001_d N_A_413_90#_c_2006_n 0.0103023f $X=3.115 $Y=2.32 $X2=0
+ $Y2=0
cc_1135 N_VPWR_c_1812_n N_A_413_90#_c_2006_n 0.0236174f $X=3.265 $Y=2.815 $X2=0
+ $Y2=0
cc_1136 N_VPWR_c_1810_n N_A_413_90#_c_2006_n 0.023363f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1137 N_VPWR_M1025_d N_A_413_90#_c_1999_n 0.00371121f $X=4.735 $Y=1.935 $X2=0
+ $Y2=0
cc_1138 N_VPWR_c_1813_n N_A_413_90#_c_1999_n 0.016342f $X=4.87 $Y=2.88 $X2=0
+ $Y2=0
cc_1139 N_VPWR_c_1821_n N_A_413_90#_c_1999_n 0.010522f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1140 N_VPWR_c_1823_n N_A_413_90#_c_1999_n 0.00976707f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_1141 N_VPWR_c_1810_n N_A_413_90#_c_1999_n 0.0371338f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1142 N_VPWR_c_1823_n N_A_413_90#_c_2000_n 0.0056737f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_1143 N_VPWR_c_1810_n N_A_413_90#_c_2000_n 0.00686828f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1144 N_VPWR_c_1811_n N_A_413_90#_c_2004_n 0.0180221f $X=1.39 $Y=2.475 $X2=0
+ $Y2=0
cc_1145 N_VPWR_c_1812_n N_A_413_90#_c_2004_n 0.00657142f $X=3.265 $Y=2.815 $X2=0
+ $Y2=0
cc_1146 N_VPWR_c_1826_n N_A_413_90#_c_2004_n 0.0155867f $X=3.085 $Y=3.33 $X2=0
+ $Y2=0
cc_1147 N_VPWR_c_1810_n N_A_413_90#_c_2004_n 0.0119322f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1148 N_VPWR_M1001_d N_A_413_90#_c_2005_n 0.00106248f $X=3.115 $Y=2.32 $X2=0
+ $Y2=0
cc_1149 N_VPWR_c_1812_n N_A_413_90#_c_2005_n 0.0213403f $X=3.265 $Y=2.815 $X2=0
+ $Y2=0
cc_1150 N_VPWR_c_1821_n N_A_413_90#_c_2005_n 0.0176368f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1151 N_VPWR_c_1810_n N_A_413_90#_c_2005_n 0.0196785f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1152 N_VPWR_c_1817_n Q_N 0.0378068f $X=11.592 $Y=3.245 $X2=0 $Y2=0
cc_1153 N_VPWR_c_1830_n Q_N 0.0146357f $X=13.045 $Y=3.33 $X2=0 $Y2=0
cc_1154 N_VPWR_c_1810_n Q_N 0.0121141f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1155 N_VPWR_c_1818_n Q 0.00249537f $X=13.21 $Y=1.985 $X2=0 $Y2=0
cc_1156 N_VPWR_c_1831_n Q 0.0124046f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1157 N_VPWR_c_1810_n Q 0.0102675f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1158 N_A_413_90#_c_2006_n A_515_464# 0.0121424f $X=3.445 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_1159 N_A_413_90#_c_1991_n N_noxref_25_c_2318_n 0.0146432f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1160 N_A_413_90#_c_1997_n N_noxref_25_c_2318_n 0.0224658f $X=2.435 $Y=0.76
+ $X2=0 $Y2=0
cc_1161 N_A_413_90#_c_1991_n N_noxref_25_c_2320_n 0.0222684f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1162 N_A_413_90#_c_1997_n N_noxref_25_c_2320_n 0.00518589f $X=2.435 $Y=0.76
+ $X2=0 $Y2=0
cc_1163 Q_N N_VGND_c_2184_n 0.0145639f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1164 Q_N N_VGND_c_2194_n 0.0119984f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1165 Q_N N_VGND_c_2199_n 0.00297405f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1166 Q N_VGND_c_2185_n 0.0297276f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1167 Q N_VGND_c_2193_n 0.0161257f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1168 Q N_VGND_c_2194_n 0.013291f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1169 N_VGND_c_2179_n N_noxref_25_c_2317_n 0.0253895f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1170 N_VGND_c_2189_n N_noxref_25_c_2318_n 0.109804f $X=3.56 $Y=0 $X2=0 $Y2=0
cc_1171 N_VGND_c_2194_n N_noxref_25_c_2318_n 0.0641003f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1172 N_VGND_c_2179_n N_noxref_25_c_2319_n 0.0121617f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1173 N_VGND_c_2189_n N_noxref_25_c_2319_n 0.0176516f $X=3.56 $Y=0 $X2=0 $Y2=0
cc_1174 N_VGND_c_2194_n N_noxref_25_c_2319_n 0.00966868f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1175 N_VGND_c_2180_n N_noxref_25_c_2320_n 0.027964f $X=3.7 $Y=0.585 $X2=0
+ $Y2=0
cc_1176 N_VGND_c_2189_n N_noxref_25_c_2320_n 0.0229596f $X=3.56 $Y=0 $X2=0 $Y2=0
cc_1177 N_VGND_c_2194_n N_noxref_25_c_2320_n 0.0126481f $X=13.68 $Y=0 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o2111a_2.pex.spice
* Created: Fri Aug 28 17:51:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2111A_2%A1 5 7 9 10 11 15
c24 11 0 1.15392e-19 $X=0.72 $Y=1.295
c25 7 0 1.31769e-19 $X=0.7 $Y=1.22
r26 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r27 11 16 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r28 10 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r29 7 15 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.7 $Y=1.22
+ $X2=0.685 $Y2=1.385
r30 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.7
+ $Y2=0.74
r31 3 15 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.685 $Y=1.55
+ $X2=0.685 $Y2=1.385
r32 3 5 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.685 $Y=1.55
+ $X2=0.685 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%A2 3 7 8 11 13
c31 13 0 1.15392e-19 $X=1.18 $Y=1.22
c32 8 0 1.73321e-19 $X=1.2 $Y=1.295
r33 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.385
+ $X2=1.18 $Y2=1.55
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.385
+ $X2=1.18 $Y2=1.22
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.385 $X2=1.18 $Y2=1.385
r36 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=1.295 $X2=1.18
+ $Y2=1.385
r37 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.27 $Y=0.74 $X2=1.27
+ $Y2=1.22
r38 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.105 $Y=2.34
+ $X2=1.105 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%B1 3 7 8 11 13
c37 13 0 4.15525e-20 $X=1.75 $Y=1.22
r38 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.385
+ $X2=1.75 $Y2=1.55
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.385
+ $X2=1.75 $Y2=1.22
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.385 $X2=1.75 $Y2=1.385
r41 8 12 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=1.74 $Y=1.295 $X2=1.74
+ $Y2=1.385
r42 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.77 $Y=0.74 $X2=1.77
+ $Y2=1.22
r43 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.675 $Y=2.34
+ $X2=1.675 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%C1 3 7 9 12
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.515
+ $X2=2.32 $Y2=1.68
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.515
+ $X2=2.32 $Y2=1.35
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.515 $X2=2.32 $Y2=1.515
r45 9 13 8.57632 $w=4.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.32 $Y2=1.565
r46 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=2.34
+ $X2=2.315 $Y2=1.68
r47 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.23 $Y=0.74 $X2=2.23
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%D1 3 7 9 15 16
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.515 $X2=3.09 $Y2=1.515
r40 13 15 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.815 $Y=1.515
+ $X2=3.09 $Y2=1.515
r41 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.8 $Y=1.515
+ $X2=2.815 $Y2=1.515
r42 9 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.515
r43 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.68
+ $X2=2.815 $Y2=1.515
r44 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.815 $Y=1.68
+ $X2=2.815 $Y2=2.34
r45 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.35 $X2=2.8
+ $Y2=1.515
r46 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.8 $Y=1.35 $X2=2.8
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%A_239_368# 1 2 3 12 16 20 24 26 28 30 34 36
+ 40 42 43 44 45 49 57
r113 57 58 6.71517 $w=3.23e-07 $l=4.5e-08 $layer=POLY_cond $X=4.245 $Y=1.465
+ $X2=4.29 $Y2=1.465
r114 56 57 57.452 $w=3.23e-07 $l=3.85e-07 $layer=POLY_cond $X=3.86 $Y=1.465
+ $X2=4.245 $Y2=1.465
r115 55 56 9.69969 $w=3.23e-07 $l=6.5e-08 $layer=POLY_cond $X=3.795 $Y=1.465
+ $X2=3.86 $Y2=1.465
r116 53 55 17.161 $w=3.23e-07 $l=1.15e-07 $layer=POLY_cond $X=3.68 $Y=1.465
+ $X2=3.795 $Y2=1.465
r117 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.465 $X2=3.68 $Y2=1.465
r118 50 52 17.702 $w=2.55e-07 $l=3.7e-07 $layer=LI1_cond $X=3.68 $Y=1.095
+ $X2=3.68 $Y2=1.465
r119 44 52 9.25285 $w=2.55e-07 $l=2.0106e-07 $layer=LI1_cond $X=3.6 $Y=1.63
+ $X2=3.68 $Y2=1.465
r120 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.6 $Y=1.63 $X2=3.6
+ $Y2=1.95
r121 42 50 3.11056 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=1.095
+ $X2=3.68 $Y2=1.095
r122 42 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.515 $Y=1.095
+ $X2=3.18 $Y2=1.095
r123 38 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.015 $Y=1.01
+ $X2=3.18 $Y2=1.095
r124 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.015 $Y=1.01
+ $X2=3.015 $Y2=0.515
r125 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=2.035
+ $X2=2.54 $Y2=2.035
r126 36 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.515 $Y=2.035
+ $X2=3.6 $Y2=1.95
r127 36 37 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.515 $Y=2.035
+ $X2=2.705 $Y2=2.035
r128 32 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=2.12
+ $X2=2.54 $Y2=2.035
r129 32 34 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.54 $Y=2.12
+ $X2=2.54 $Y2=2.375
r130 31 47 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=1.45 $Y2=1.97
r131 30 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.035
+ $X2=2.54 $Y2=2.035
r132 30 31 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.375 $Y=2.035
+ $X2=1.615 $Y2=2.035
r133 26 47 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.45 $Y=2.12 $X2=1.45
+ $Y2=1.97
r134 26 28 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.45 $Y=2.12
+ $X2=1.45 $Y2=2.695
r135 22 58 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.29 $Y=1.3
+ $X2=4.29 $Y2=1.465
r136 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.29 $Y=1.3
+ $X2=4.29 $Y2=0.74
r137 18 57 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.63
+ $X2=4.245 $Y2=1.465
r138 18 20 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.245 $Y=1.63
+ $X2=4.245 $Y2=2.4
r139 14 56 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.86 $Y=1.3
+ $X2=3.86 $Y2=1.465
r140 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.86 $Y=1.3
+ $X2=3.86 $Y2=0.74
r141 10 55 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.63
+ $X2=3.795 $Y2=1.465
r142 10 12 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.795 $Y=1.63
+ $X2=3.795 $Y2=2.4
r143 3 49 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.84 $X2=2.54 $Y2=2.035
r144 3 34 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.405
+ $Y=1.84 $X2=2.54 $Y2=2.375
r145 2 47 400 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=1.84 $X2=1.45 $Y2=1.985
r146 2 28 400 $w=1.7e-07 $l=9.74192e-07 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=1.84 $X2=1.45 $Y2=2.695
r147 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.875
+ $Y=0.37 $X2=3.015 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%VPWR 1 2 3 4 15 21 25 27 29 34 35 37 38 39
+ 50 54 60 64
r58 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 58 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 58 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 55 60 14.7259 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.28 $Y2=3.33
r64 55 57 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 54 63 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.577 $Y2=3.33
r66 54 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 53 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 50 60 14.7259 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=3.28 $Y2=3.33
r70 50 52 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r74 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 39 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 39 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 37 48 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.95 $Y2=3.33
r81 36 52 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.95 $Y2=3.33
r83 34 42 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.295 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=3.33
+ $X2=0.46 $Y2=3.33
r85 33 45 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.46 $Y2=3.33
r87 29 32 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.52 $Y=1.985
+ $X2=4.52 $Y2=2.815
r88 27 63 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.577 $Y2=3.33
r89 27 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.52 $Y2=2.815
r90 23 60 3.15573 $w=8.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=3.33
r91 23 25 12.8468 $w=8.08e-07 $l=8.7e-07 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=2.375
r92 19 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r93 19 21 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.375
r94 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.46 $Y=1.985
+ $X2=0.46 $Y2=2.695
r95 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.46 $Y=3.245
+ $X2=0.46 $Y2=3.33
r96 13 18 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.46 $Y=3.245
+ $X2=0.46 $Y2=2.695
r97 4 32 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.84 $X2=4.52 $Y2=2.815
r98 4 29 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.84 $X2=4.52 $Y2=1.985
r99 3 25 150 $w=1.7e-07 $l=8.40982e-07 $layer=licon1_PDIFF $count=4 $X=2.905
+ $Y=1.84 $X2=3.52 $Y2=2.375
r100 2 21 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=1.765
+ $Y=1.84 $X2=1.95 $Y2=2.375
r101 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.84 $X2=0.46 $Y2=2.695
r102 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.84 $X2=0.46 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%X 1 2 9 11 15 16 17 28
r32 21 28 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=4.075 $Y=0.965
+ $X2=4.075 $Y2=0.925
r33 17 30 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=4.075 $Y=0.987
+ $X2=4.075 $Y2=1.13
r34 17 21 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=4.075 $Y=0.987
+ $X2=4.075 $Y2=0.965
r35 17 28 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=4.075 $Y=0.902
+ $X2=4.075 $Y2=0.925
r36 16 17 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=4.075 $Y=0.515
+ $X2=4.075 $Y2=0.902
r37 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.1 $Y=1.82 $X2=4.1
+ $Y2=1.13
r38 9 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=1.985
+ $X2=4.02 $Y2=1.82
r39 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.02 $Y=1.985
+ $X2=4.02 $Y2=2.815
r40 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.02 $Y2=2.815
r41 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.02 $Y2=1.985
r42 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.37 $X2=4.075 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%A_54_74# 1 2 7 9 11 13 15
r27 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=0.84
+ $X2=1.555 $Y2=0.925
r28 13 15 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.555 $Y=0.84
+ $X2=1.555 $Y2=0.515
r29 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0.925
+ $X2=0.415 $Y2=0.925
r30 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0.925
+ $X2=1.555 $Y2=0.925
r31 11 12 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.39 $Y=0.925
+ $X2=0.58 $Y2=0.925
r32 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=0.84 $X2=0.415
+ $Y2=0.925
r33 7 9 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.415 $Y=0.84
+ $X2=0.415 $Y2=0.515
r34 2 20 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=1.345
+ $Y=0.37 $X2=1.555 $Y2=0.925
r35 2 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.345
+ $Y=0.37 $X2=1.555 $Y2=0.515
r36 1 18 182 $w=1.7e-07 $l=6.5372e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.37 $X2=0.485 $Y2=0.925
r37 1 9 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.37 $X2=0.485 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111A_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r52 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r55 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r56 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.575
+ $Y2=0
r58 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=4.08
+ $Y2=0
r59 34 46 4.13553 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.61
+ $Y2=0
r60 34 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.08
+ $Y2=0
r61 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r62 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 30 40 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=0.985
+ $Y2=0
r64 30 32 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=1.22 $Y=0 $X2=3.12
+ $Y2=0
r65 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.575
+ $Y2=0
r66 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.12
+ $Y2=0
r67 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r68 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 24 40 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.985
+ $Y2=0
r70 24 26 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.72
+ $Y2=0
r71 22 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r72 22 41 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r73 18 46 3.11253 $w=2.65e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.552 $Y=0.085
+ $X2=4.61 $Y2=0
r74 18 20 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=4.552 $Y=0.085
+ $X2=4.552 $Y2=0.515
r75 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0
r76 14 16 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.63
r77 10 40 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0
r78 10 12 11.7063 $w=4.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0.545
r79 3 20 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.365
+ $Y=0.37 $X2=4.51 $Y2=0.515
r80 2 16 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.37 $X2=3.645 $Y2=0.63
r81 1 12 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.37 $X2=0.985 $Y2=0.545
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor3_1 A B C VGND VNB VPB VPWR X
X0 VGND C a_232_162# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_81_268# a_232_162# a_363_394# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_897_54# a_786_100# a_363_394# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 VGND a_897_54# a_1116_383# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_371_74# C a_81_268# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_897_54# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 a_1116_383# a_786_100# a_371_74# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X7 X a_81_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND B a_786_100# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_1116_383# a_786_100# a_363_394# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VPWR C a_232_162# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X11 a_371_74# B a_897_54# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X12 a_363_394# B a_897_54# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_897_54# a_786_100# a_371_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_81_268# a_232_162# a_371_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X15 VPWR a_897_54# a_1116_383# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 X a_81_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VPWR B a_786_100# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_363_394# B a_1116_383# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X19 a_897_54# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_363_394# C a_81_268# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X21 a_371_74# B a_1116_383# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_313_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_476_48# A2_N a_835_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VPWR A2_N a_476_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 VPWR a_313_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VGND a_313_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_313_392# a_476_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VGND a_313_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_476_48# a_313_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 a_313_392# a_476_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X9 VGND B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 X a_313_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 X a_313_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VPWR B1 a_41_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 X a_313_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_313_392# B2 a_41_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_476_48# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X18 a_835_94# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_27_74# a_476_48# a_313_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_41_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X21 X a_313_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_27_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_41_392# B2 a_313_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
.ends

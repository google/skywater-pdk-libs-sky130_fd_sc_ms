* File: sky130_fd_sc_ms__a21boi_1.pex.spice
* Created: Fri Aug 28 16:58:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21BOI_1%B1_N 1 3 5 7 9 10 11 12 18 19
r46 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=1.44 $X2=0.285 $Y2=1.44
r47 21 23 22.2462 $w=3.9e-07 $l=1.8e-07 $layer=POLY_cond $X=0.352 $Y=1.26
+ $X2=0.352 $Y2=1.44
r48 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=0.42 $X2=0.285 $Y2=0.42
r49 16 21 8.93446 $w=4.35e-07 $l=8.21584e-08 $layer=POLY_cond $X=0.337 $Y=1.185
+ $X2=0.352 $Y2=1.26
r50 16 18 97.8064 $w=4.35e-07 $l=7.65e-07 $layer=POLY_cond $X=0.337 $Y=1.185
+ $X2=0.337 $Y2=0.42
r51 12 24 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.285 $Y=1.295
+ $X2=0.285 $Y2=1.44
r52 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.285 $Y=0.925
+ $X2=0.285 $Y2=1.295
r53 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.285 $Y=0.555
+ $X2=0.285 $Y2=0.925
r54 10 19 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.285 $Y=0.555
+ $X2=0.285 $Y2=0.42
r55 7 9 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1 $Y=1.185 $X2=1
+ $Y2=0.835
r56 6 21 25.2441 $w=1.5e-07 $l=2.03e-07 $layer=POLY_cond $X=0.555 $Y=1.26
+ $X2=0.352 $Y2=1.26
r57 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=1.26
+ $X2=1 $Y2=1.185
r58 5 6 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.925 $Y=1.26
+ $X2=0.555 $Y2=1.26
r59 1 23 45.6156 $w=3.9e-07 $l=3.18575e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.352 $Y2=1.44
r60 1 3 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.495 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%A_29_424# 1 2 9 11 13 16 18 19 22 25 27 30
+ 33 34 38
r74 37 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.665 $Y=1.385
+ $X2=1.68 $Y2=1.385
r75 31 37 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.45 $Y=1.385
+ $X2=1.665 $Y2=1.385
r76 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.385 $X2=1.45 $Y2=1.385
r77 28 34 0.588983 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=0.95 $Y=1.385
+ $X2=0.847 $Y2=1.385
r78 28 30 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.95 $Y=1.385 $X2=1.45
+ $Y2=1.385
r79 26 34 8.03064 $w=1.87e-07 $l=1.73292e-07 $layer=LI1_cond $X=0.83 $Y=1.55
+ $X2=0.847 $Y2=1.385
r80 26 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.83 $Y=1.55
+ $X2=0.83 $Y2=1.775
r81 25 34 8.03064 $w=1.87e-07 $l=1.65e-07 $layer=LI1_cond $X=0.847 $Y=1.22
+ $X2=0.847 $Y2=1.385
r82 25 33 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=0.847 $Y=1.22
+ $X2=0.847 $Y2=1.05
r83 20 33 7.40596 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=0.885
+ $X2=0.785 $Y2=1.05
r84 20 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.785 $Y=0.885
+ $X2=0.785 $Y2=0.795
r85 18 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.745 $Y=1.86
+ $X2=0.83 $Y2=1.775
r86 18 19 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.745 $Y=1.86
+ $X2=0.435 $Y2=1.86
r87 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=1.945
+ $X2=0.435 $Y2=1.86
r88 14 16 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.27 $Y=1.945
+ $X2=0.27 $Y2=2.265
r89 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.22
+ $X2=1.68 $Y2=1.385
r90 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.68 $Y=1.22 $X2=1.68
+ $Y2=0.74
r91 7 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.55
+ $X2=1.665 $Y2=1.385
r92 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.665 $Y=1.55
+ $X2=1.665 $Y2=2.4
r93 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=2.12 $X2=0.27 $Y2=2.265
r94 1 22 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.56 $X2=0.785 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%A1 3 7 9 12 13
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.68
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.35
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r44 9 13 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=1.515
r45 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.11 $Y=0.74 $X2=2.11
+ $Y2=1.35
r46 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.115 $Y=2.4
+ $X2=2.115 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%A2 3 6 8 9 13 15
r29 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.385
+ $X2=2.67 $Y2=1.55
r30 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.385
+ $X2=2.67 $Y2=1.22
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.385 $X2=2.67 $Y2=1.385
r32 9 14 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.67 $Y2=1.365
r33 8 14 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.365 $X2=2.67
+ $Y2=1.365
r34 6 16 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.595 $Y=2.4
+ $X2=2.595 $Y2=1.55
r35 3 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.58 $Y=0.74 $X2=2.58
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r44 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 25 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.76 $Y2=3.33
r46 25 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.76 $Y2=3.33
r50 20 22 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 16 30 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.19 $Y=3.33 $X2=2.16
+ $Y2=3.33
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=3.33
+ $X2=2.355 $Y2=3.33
r55 15 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.52 $Y=3.33 $X2=3.12
+ $Y2=3.33
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.52 $Y=3.33
+ $X2=2.355 $Y2=3.33
r57 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=3.245
+ $X2=2.355 $Y2=3.33
r58 11 13 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.355 $Y=3.245
+ $X2=2.355 $Y2=2.485
r59 7 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r60 7 9 44.4843 $w=2.48e-07 $l=9.65e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.28
r61 2 13 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=2.205
+ $Y=1.84 $X2=2.355 $Y2=2.485
r62 1 9 300 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.12 $X2=0.72 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%Y 1 2 7 10 13 16 17 18 19 23
r49 31 33 6.29226 $w=3.49e-07 $l=1.8e-07 $layer=LI1_cond $X=1.305 $Y=1.805
+ $X2=1.305 $Y2=1.985
r50 19 29 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=1.305 $Y=2.775
+ $X2=1.305 $Y2=2.815
r51 18 19 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.305 $Y=2.405
+ $X2=1.305 $Y2=2.775
r52 18 23 6.94085 $w=4.38e-07 $l=2.65e-07 $layer=LI1_cond $X=1.305 $Y=2.405
+ $X2=1.305 $Y2=2.14
r53 17 23 3.4677 $w=4.4e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=2.035
+ $X2=1.305 $Y2=2.14
r54 17 33 1.74785 $w=3.49e-07 $l=5e-08 $layer=LI1_cond $X=1.305 $Y=2.035
+ $X2=1.305 $Y2=1.985
r55 15 16 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.882 $Y=1.01
+ $X2=1.882 $Y2=1.18
r56 13 15 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.935 $Y=0.515
+ $X2=1.935 $Y2=1.01
r57 10 16 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.79 $Y=1.72
+ $X2=1.79 $Y2=1.18
r58 8 31 4.95691 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.525 $Y=1.805
+ $X2=1.305 $Y2=1.805
r59 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.705 $Y=1.805
+ $X2=1.79 $Y2=1.72
r60 7 8 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.705 $Y=1.805
+ $X2=1.525 $Y2=1.805
r61 2 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=1.985
r62 2 29 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=2.815
r63 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.755
+ $Y=0.37 $X2=1.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%A_351_368# 1 2 9 13 16 18
r27 20 21 3.12451 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=2.145
+ $X2=2.82 $Y2=2.23
r28 18 20 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.82 $Y=1.985
+ $X2=2.82 $Y2=2.145
r29 13 21 6.6412 $w=2.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.837 $Y=2.4
+ $X2=2.837 $Y2=2.23
r30 10 16 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.02 $Y=2.145
+ $X2=1.872 $Y2=2.145
r31 9 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=2.145
+ $X2=2.82 $Y2=2.145
r32 9 10 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.655 $Y=2.145
+ $X2=2.02 $Y2=2.145
r33 2 18 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.84 $X2=2.82 $Y2=1.985
r34 2 13 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.685
+ $Y=1.84 $X2=2.82 $Y2=2.4
r35 1 16 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.755
+ $Y=1.84 $X2=1.89 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_1%VGND 1 2 8 11 15 17 22 29 30 33 36
r39 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.795
+ $Y2=0
r44 27 29 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=3.12
+ $Y2=0
r45 23 33 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.375
+ $Y2=0
r46 23 25 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.68
+ $Y2=0
r47 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.795
+ $Y2=0
r48 22 25 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=1.68
+ $Y2=0
r49 20 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r50 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 17 33 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.375
+ $Y2=0
r52 17 19 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.24
+ $Y2=0
r53 15 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r54 15 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r55 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0
r57 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0.515
r58 8 14 2.62105 $w=5.1e-07 $l=9e-08 $layer=LI1_cond $X=1.375 $Y=0.505 $X2=1.375
+ $Y2=0.595
r59 7 33 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0
r60 7 8 9.85006 $w=5.08e-07 $l=4.2e-07 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0.505
r61 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.655
+ $Y=0.37 $X2=2.795 $Y2=0.515
r62 1 14 91 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.56 $X2=1.465 $Y2=0.595
.ends


* File: sky130_fd_sc_ms__clkbuf_2.pxi.spice
* Created: Wed Sep  2 12:00:28 2020
* 
x_PM_SKY130_FD_SC_MS__CLKBUF_2%A_43_192# N_A_43_192#_M1002_d N_A_43_192#_M1003_d
+ N_A_43_192#_M1000_g N_A_43_192#_M1004_g N_A_43_192#_M1005_g
+ N_A_43_192#_M1001_g N_A_43_192#_c_48_n N_A_43_192#_c_49_n N_A_43_192#_c_61_p
+ N_A_43_192#_c_78_p N_A_43_192#_c_57_n N_A_43_192#_c_50_n N_A_43_192#_c_51_n
+ N_A_43_192#_c_52_n N_A_43_192#_c_59_n N_A_43_192#_c_53_n
+ PM_SKY130_FD_SC_MS__CLKBUF_2%A_43_192#
x_PM_SKY130_FD_SC_MS__CLKBUF_2%A N_A_M1003_g N_A_M1002_g N_A_c_124_n N_A_c_125_n
+ A A A N_A_c_126_n N_A_c_127_n PM_SKY130_FD_SC_MS__CLKBUF_2%A
x_PM_SKY130_FD_SC_MS__CLKBUF_2%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_c_162_n
+ N_VPWR_c_163_n N_VPWR_c_164_n VPWR N_VPWR_c_165_n N_VPWR_c_166_n
+ N_VPWR_c_161_n N_VPWR_c_168_n PM_SKY130_FD_SC_MS__CLKBUF_2%VPWR
x_PM_SKY130_FD_SC_MS__CLKBUF_2%X N_X_M1004_d N_X_M1000_d N_X_c_194_n N_X_c_192_n
+ X PM_SKY130_FD_SC_MS__CLKBUF_2%X
x_PM_SKY130_FD_SC_MS__CLKBUF_2%VGND N_VGND_M1004_s N_VGND_M1005_s N_VGND_c_220_n
+ N_VGND_c_221_n N_VGND_c_222_n VGND N_VGND_c_223_n N_VGND_c_224_n
+ N_VGND_c_225_n N_VGND_c_226_n PM_SKY130_FD_SC_MS__CLKBUF_2%VGND
cc_1 VNB N_A_43_192#_M1000_g 0.00166642f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A_43_192#_M1004_g 0.025695f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_A_43_192#_M1005_g 0.0206266f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.58
cc_4 VNB N_A_43_192#_M1001_g 0.00139804f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_5 VNB N_A_43_192#_c_48_n 0.00366521f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.125
cc_6 VNB N_A_43_192#_c_49_n 0.00120535f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=2.32
cc_7 VNB N_A_43_192#_c_50_n 0.0396899f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=2.32
cc_8 VNB N_A_43_192#_c_51_n 8.13082e-19 $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.63
cc_9 VNB N_A_43_192#_c_52_n 0.0254971f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=0.58
cc_10 VNB N_A_43_192#_c_53_n 0.125169f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.295
cc_11 VNB N_A_M1002_g 0.0299202f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.63
cc_12 VNB N_A_c_124_n 0.0231477f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.96
cc_13 VNB N_A_c_125_n 0.00993024f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_14 VNB N_A_c_126_n 0.016251f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_15 VNB N_A_c_127_n 0.00804942f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_16 VNB N_VPWR_c_161_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.125
cc_17 VNB N_X_c_192_n 0.00135547f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.96
cc_18 VNB X 0.00425977f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_19 VNB N_VGND_c_220_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.63
cc_20 VNB N_VGND_c_221_n 0.0326954f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_21 VNB N_VGND_c_222_n 0.012368f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_22 VNB N_VGND_c_223_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.58
cc_23 VNB N_VGND_c_224_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.125
cc_24 VNB N_VGND_c_225_n 0.138933f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=1.125
cc_25 VNB N_VGND_c_226_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.405
cc_26 VPB N_A_43_192#_M1000_g 0.0245517f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_27 VPB N_A_43_192#_M1001_g 0.0212867f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_28 VPB N_A_43_192#_c_49_n 0.00771408f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.32
cc_29 VPB N_A_43_192#_c_57_n 0.0217468f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=2.815
cc_30 VPB N_A_43_192#_c_50_n 0.025967f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=2.32
cc_31 VPB N_A_43_192#_c_59_n 0.00723806f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=2.405
cc_32 VPB N_A_M1003_g 0.025304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A_c_125_n 0.00626001f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_34 VPB N_A_c_127_n 0.002588f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_35 VPB N_VPWR_c_162_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.63
cc_36 VPB N_VPWR_c_163_n 0.0219477f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_37 VPB N_VPWR_c_164_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_38 VPB N_VPWR_c_165_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.58
cc_39 VPB N_VPWR_c_166_n 0.0182732f $X=-0.19 $Y=1.66 $X2=0.38 $Y2=1.125
cc_40 VPB N_VPWR_c_161_n 0.0499503f $X=-0.19 $Y=1.66 $X2=0.38 $Y2=1.125
cc_41 VPB N_VPWR_c_168_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=2.405
cc_42 VPB N_X_c_194_n 0.00377904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_X_c_192_n 8.13921e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.96
cc_44 N_A_43_192#_M1001_g N_A_M1003_g 0.0476457f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_45 N_A_43_192#_c_61_p N_A_M1003_g 0.0110395f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_46 N_A_43_192#_c_57_n N_A_M1003_g 8.73643e-19 $X=1.63 $Y=2.815 $X2=0 $Y2=0
cc_47 N_A_43_192#_c_50_n N_A_M1003_g 0.006356f $X=1.75 $Y=2.32 $X2=0 $Y2=0
cc_48 N_A_43_192#_M1005_g N_A_M1002_g 0.0145334f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_49 N_A_43_192#_c_50_n N_A_M1002_g 0.00514634f $X=1.75 $Y=2.32 $X2=0 $Y2=0
cc_50 N_A_43_192#_c_52_n N_A_M1002_g 0.00696419f $X=1.64 $Y=0.58 $X2=0 $Y2=0
cc_51 N_A_43_192#_c_53_n N_A_M1002_g 0.0020866f $X=0.945 $Y=1.295 $X2=0 $Y2=0
cc_52 N_A_43_192#_M1001_g N_A_c_124_n 0.0217016f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_53 N_A_43_192#_c_59_n N_A_c_125_n 0.00106699f $X=1.63 $Y=2.405 $X2=0 $Y2=0
cc_54 N_A_43_192#_c_50_n N_A_c_126_n 0.0164695f $X=1.75 $Y=2.32 $X2=0 $Y2=0
cc_55 N_A_43_192#_c_52_n N_A_c_126_n 0.00331415f $X=1.64 $Y=0.58 $X2=0 $Y2=0
cc_56 N_A_43_192#_c_53_n N_A_c_126_n 0.0217016f $X=0.945 $Y=1.295 $X2=0 $Y2=0
cc_57 N_A_43_192#_c_61_p N_A_c_127_n 0.0263694f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_58 N_A_43_192#_c_50_n N_A_c_127_n 0.0752414f $X=1.75 $Y=2.32 $X2=0 $Y2=0
cc_59 N_A_43_192#_c_52_n N_A_c_127_n 0.0012973f $X=1.64 $Y=0.58 $X2=0 $Y2=0
cc_60 N_A_43_192#_c_53_n N_A_c_127_n 0.00840431f $X=0.945 $Y=1.295 $X2=0 $Y2=0
cc_61 N_A_43_192#_c_49_n N_VPWR_M1000_s 0.0205644f $X=0.3 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_62 N_A_43_192#_c_78_p N_VPWR_M1000_s 0.00920379f $X=0.385 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_63 N_A_43_192#_c_61_p N_VPWR_M1001_s 0.00326225f $X=1.535 $Y=2.405 $X2=0
+ $Y2=0
cc_64 N_A_43_192#_M1000_g N_VPWR_c_163_n 0.0118211f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_65 N_A_43_192#_M1001_g N_VPWR_c_163_n 0.00125818f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A_43_192#_c_61_p N_VPWR_c_163_n 0.0021187f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_67 N_A_43_192#_c_78_p N_VPWR_c_163_n 0.0116597f $X=0.385 $Y=2.405 $X2=0 $Y2=0
cc_68 N_A_43_192#_M1000_g N_VPWR_c_164_n 0.00125818f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A_43_192#_M1001_g N_VPWR_c_164_n 0.0106899f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A_43_192#_c_61_p N_VPWR_c_164_n 0.0166513f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_71 N_A_43_192#_c_57_n N_VPWR_c_164_n 0.0112375f $X=1.63 $Y=2.815 $X2=0 $Y2=0
cc_72 N_A_43_192#_M1000_g N_VPWR_c_165_n 0.00460063f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_43_192#_M1001_g N_VPWR_c_165_n 0.00460063f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_74 N_A_43_192#_c_57_n N_VPWR_c_166_n 0.0132845f $X=1.63 $Y=2.815 $X2=0 $Y2=0
cc_75 N_A_43_192#_M1000_g N_VPWR_c_161_n 0.0046086f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A_43_192#_M1001_g N_VPWR_c_161_n 0.0046086f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_43_192#_c_61_p N_VPWR_c_161_n 0.0246034f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_78 N_A_43_192#_c_78_p N_VPWR_c_161_n 6.15054e-19 $X=0.385 $Y=2.405 $X2=0
+ $Y2=0
cc_79 N_A_43_192#_c_57_n N_VPWR_c_161_n 0.0110013f $X=1.63 $Y=2.815 $X2=0 $Y2=0
cc_80 N_A_43_192#_c_61_p N_X_M1000_d 0.00473092f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_81 N_A_43_192#_M1000_g N_X_c_194_n 0.0058762f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_82 N_A_43_192#_M1001_g N_X_c_194_n 0.00454626f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_43_192#_c_49_n N_X_c_194_n 0.0130972f $X=0.3 $Y=2.32 $X2=0 $Y2=0
cc_84 N_A_43_192#_c_61_p N_X_c_194_n 0.0165698f $X=1.535 $Y=2.405 $X2=0 $Y2=0
cc_85 N_A_43_192#_c_53_n N_X_c_194_n 0.00172428f $X=0.945 $Y=1.295 $X2=0 $Y2=0
cc_86 N_A_43_192#_M1000_g N_X_c_192_n 0.00111019f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_43_192#_M1004_g N_X_c_192_n 0.0025553f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_88 N_A_43_192#_M1005_g N_X_c_192_n 0.00452402f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_89 N_A_43_192#_M1001_g N_X_c_192_n 0.00377148f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_43_192#_c_48_n N_X_c_192_n 0.0478089f $X=0.38 $Y=1.125 $X2=0 $Y2=0
cc_91 N_A_43_192#_c_49_n N_X_c_192_n 0.00661604f $X=0.3 $Y=2.32 $X2=0 $Y2=0
cc_92 N_A_43_192#_c_53_n N_X_c_192_n 0.0283479f $X=0.945 $Y=1.295 $X2=0 $Y2=0
cc_93 N_A_43_192#_M1004_g X 0.00682464f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_94 N_A_43_192#_M1005_g X 0.0057329f $X=0.925 $Y=0.58 $X2=0 $Y2=0
cc_95 N_A_43_192#_c_53_n X 0.00250405f $X=0.945 $Y=1.295 $X2=0 $Y2=0
cc_96 N_A_43_192#_M1004_g N_VGND_c_221_n 0.00545557f $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_97 N_A_43_192#_c_48_n N_VGND_c_221_n 0.0128908f $X=0.38 $Y=1.125 $X2=0 $Y2=0
cc_98 N_A_43_192#_c_53_n N_VGND_c_221_n 0.00115565f $X=0.945 $Y=1.295 $X2=0
+ $Y2=0
cc_99 N_A_43_192#_M1005_g N_VGND_c_222_n 0.00337454f $X=0.925 $Y=0.58 $X2=0
+ $Y2=0
cc_100 N_A_43_192#_c_52_n N_VGND_c_222_n 0.0190076f $X=1.64 $Y=0.58 $X2=0 $Y2=0
cc_101 N_A_43_192#_M1004_g N_VGND_c_223_n 0.00434272f $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_102 N_A_43_192#_M1005_g N_VGND_c_223_n 0.00422942f $X=0.925 $Y=0.58 $X2=0
+ $Y2=0
cc_103 N_A_43_192#_c_52_n N_VGND_c_224_n 0.0156722f $X=1.64 $Y=0.58 $X2=0 $Y2=0
cc_104 N_A_43_192#_M1004_g N_VGND_c_225_n 0.00823942f $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_105 N_A_43_192#_M1005_g N_VGND_c_225_n 0.00784309f $X=0.925 $Y=0.58 $X2=0
+ $Y2=0
cc_106 N_A_43_192#_c_52_n N_VGND_c_225_n 0.0130167f $X=1.64 $Y=0.58 $X2=0 $Y2=0
cc_107 N_A_c_127_n N_VPWR_M1001_s 0.00224384f $X=1.41 $Y=1.175 $X2=0 $Y2=0
cc_108 N_A_M1003_g N_VPWR_c_164_n 0.0112285f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_M1003_g N_VPWR_c_166_n 0.00460063f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_M1003_g N_VPWR_c_161_n 0.00464669f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_M1003_g N_X_c_192_n 3.45524e-19 $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_c_126_n N_X_c_192_n 5.11958e-19 $X=1.41 $Y=1.175 $X2=0 $Y2=0
cc_113 N_A_c_127_n N_X_c_192_n 0.0670495f $X=1.41 $Y=1.175 $X2=0 $Y2=0
cc_114 N_A_M1002_g X 0.00106277f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_115 N_A_M1002_g N_VGND_c_222_n 0.0054557f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_116 N_A_c_126_n N_VGND_c_222_n 4.52883e-19 $X=1.41 $Y=1.175 $X2=0 $Y2=0
cc_117 N_A_c_127_n N_VGND_c_222_n 0.0179246f $X=1.41 $Y=1.175 $X2=0 $Y2=0
cc_118 N_A_M1002_g N_VGND_c_224_n 0.00434272f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_119 N_A_M1002_g N_VGND_c_225_n 0.00824429f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_120 X N_VGND_c_221_n 0.0165704f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_121 X N_VGND_c_222_n 0.018898f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_122 X N_VGND_c_223_n 0.0146803f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_123 X N_VGND_c_225_n 0.0121149f $X=0.635 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o41ai_1.pex.spice
* Created: Wed Sep  2 12:27:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O41AI_1%B1 1 3 6 8 9 10
c37 10 0 9.14826e-20 $X=0.24 $Y=1.295
c38 6 0 1.72297e-19 $X=0.725 $Y=2.4
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r40 10 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r41 8 13 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=0.635 $Y=1.385
+ $X2=0.27 $Y2=1.385
r42 8 9 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.635 $Y=1.385 $X2=0.725
+ $Y2=1.385
r43 4 9 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.725 $Y=1.55
+ $X2=0.725 $Y2=1.385
r44 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.725 $Y=1.55
+ $X2=0.725 $Y2=2.4
r45 1 9 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.71 $Y=1.22
+ $X2=0.725 $Y2=1.385
r46 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.71 $Y=1.22 $X2=0.71
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%A4 3 7 9 12 13
c46 13 0 5.13055e-20 $X=1.22 $Y=1.515
c47 12 0 4.0177e-20 $X=1.22 $Y=1.515
c48 3 0 8.61844e-20 $X=1.225 $Y=2.4
r49 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.515
+ $X2=1.22 $Y2=1.68
r50 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.515
+ $X2=1.22 $Y2=1.35
r51 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.515 $X2=1.22 $Y2=1.515
r52 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.515
r53 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.255 $Y=0.74
+ $X2=1.255 $Y2=1.35
r54 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.225 $Y=2.4
+ $X2=1.225 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%A3 3 7 9 10 11 12 19 20
r46 19 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.515
+ $X2=1.79 $Y2=1.68
r47 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.515
+ $X2=1.79 $Y2=1.35
r48 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.515 $X2=1.79 $Y2=1.515
r49 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.405
+ $X2=1.68 $Y2=2.775
r50 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.405
r51 9 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.79 $Y2=1.515
r52 9 23 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.68 $Y2=1.68
r53 9 10 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.68 $Y=1.715 $X2=1.68
+ $Y2=2.035
r54 9 23 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.715
+ $X2=1.68 $Y2=1.68
r55 7 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.84 $Y=0.74 $X2=1.84
+ $Y2=1.35
r56 3 22 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.715 $Y=2.4
+ $X2=1.715 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%A2 3 7 14 15 17 18 19 35 37
r43 27 37 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=2.17 $Y=2.045
+ $X2=2.17 $Y2=2.035
r44 18 19 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.17 $Y=2.405
+ $X2=2.17 $Y2=2.775
r45 17 37 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=2.17 $Y=1.997
+ $X2=2.17 $Y2=2.035
r46 17 35 4.73668 $w=2.48e-07 $l=7.7e-08 $layer=LI1_cond $X=2.17 $Y=1.997
+ $X2=2.17 $Y2=1.92
r47 17 18 14.8896 $w=2.48e-07 $l=3.23e-07 $layer=LI1_cond $X=2.17 $Y=2.082
+ $X2=2.17 $Y2=2.405
r48 17 27 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=2.17 $Y=2.082
+ $X2=2.17 $Y2=2.045
r49 15 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.515
+ $X2=2.36 $Y2=1.68
r50 15 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.515
+ $X2=2.36 $Y2=1.35
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.515 $X2=2.36 $Y2=1.515
r52 11 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.21 $Y=1.515
+ $X2=2.36 $Y2=1.515
r53 9 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.68 $X2=2.21
+ $Y2=1.515
r54 9 35 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.21 $Y=1.68 $X2=2.21
+ $Y2=1.92
r55 7 26 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.285 $Y=2.4
+ $X2=2.285 $Y2=1.68
r56 3 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.27 $Y=0.74 $X2=2.27
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%A1 3 7 9 12 13
r28 12 15 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.952 $Y=1.515
+ $X2=2.952 $Y2=1.68
r29 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.952 $Y=1.515
+ $X2=2.952 $Y2=1.35
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.515 $X2=2.975 $Y2=1.515
r31 9 13 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=3.022 $Y=1.665
+ $X2=3.022 $Y2=1.515
r32 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.855 $Y=2.4
+ $X2=2.855 $Y2=1.68
r33 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.84 $Y=0.74 $X2=2.84
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%VPWR 1 2 9 12 13 15 20 22 24 37
c35 20 0 8.61844e-20 $X=0.495 $Y=2.815
r36 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 25 33 6.74725 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=0.665 $Y=3.33
+ $X2=0.332 $Y2=3.33
r44 25 27 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.665 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 24 36 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r46 24 30 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 22 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 22 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 20 21 4.19009 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.39 $Y=2.815
+ $X2=0.39 $Y2=2.65
r50 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=3.12 $Y=2.115 $X2=3.12
+ $Y2=2.815
r51 13 36 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r52 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r53 12 33 2.89747 $w=5.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.39 $Y=3.245
+ $X2=0.332 $Y2=3.33
r54 11 20 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=0.39 $Y=2.925
+ $X2=0.39 $Y2=2.815
r55 11 12 6.959 $w=5.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.39 $Y=2.925 $X2=0.39
+ $Y2=3.245
r56 9 21 17.8227 $w=4.28e-07 $l=6.65e-07 $layer=LI1_cond $X=0.33 $Y=1.985
+ $X2=0.33 $Y2=2.65
r57 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.815
r58 2 15 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.115
r59 1 20 600 $w=1.7e-07 $l=1.14089e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.495 $Y2=2.815
r60 1 9 300 $w=1.7e-07 $l=3.85746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.455 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%Y 1 2 8 13 17 20 21 23 26
c42 13 0 1.72297e-19 $X=1 $Y=2.815
r43 23 30 15.8183 $w=6.48e-07 $l=4.55e-07 $layer=LI1_cond $X=0.45 $Y=0.555
+ $X2=0.45 $Y2=1.01
r44 23 26 0.736048 $w=6.48e-07 $l=4e-08 $layer=LI1_cond $X=0.45 $Y=0.555
+ $X2=0.45 $Y2=0.515
r45 20 22 1.00633 $w=4.48e-07 $l=5e-09 $layer=LI1_cond $X=0.94 $Y=2.115 $X2=0.94
+ $Y2=2.12
r46 20 21 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=2.115
+ $X2=0.94 $Y2=1.95
r47 15 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.69 $Y=1.435
+ $X2=0.8 $Y2=1.435
r48 13 22 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1 $Y=2.815 $X2=1
+ $Y2=2.12
r49 9 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.52 $X2=0.8
+ $Y2=1.435
r50 9 21 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.8 $Y=1.52 $X2=0.8
+ $Y2=1.95
r51 8 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.35 $X2=0.69
+ $Y2=1.435
r52 8 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.69 $Y=1.35 $X2=0.69
+ $Y2=1.01
r53 2 20 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=0.815
+ $Y=1.84 $X2=1 $Y2=2.115
r54 2 13 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=0.815
+ $Y=1.84 $X2=1 $Y2=2.815
r55 1 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.35
+ $Y=0.37 $X2=0.495 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%A_157_74# 1 2 3 12 14 15 18 20 24 26
r53 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.055 $Y=1.01
+ $X2=3.055 $Y2=0.515
r54 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=1.095
+ $X2=2.055 $Y2=1.095
r55 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.89 $Y=1.095
+ $X2=3.055 $Y2=1.01
r56 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.89 $Y=1.095
+ $X2=2.22 $Y2=1.095
r57 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.01
+ $X2=2.055 $Y2=1.095
r58 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.055 $Y=1.01
+ $X2=2.055 $Y2=0.515
r59 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=1.095
+ $X2=2.055 $Y2=1.095
r60 14 15 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.89 $Y=1.095
+ $X2=1.205 $Y2=1.095
r61 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.08 $Y=1.01
+ $X2=1.205 $Y2=1.095
r62 10 12 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.08 $Y=1.01
+ $X2=1.08 $Y2=0.515
r63 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.515
r64 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.37 $X2=2.055 $Y2=0.515
r65 1 12 91 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=2 $X=0.785
+ $Y=0.37 $X2=1.04 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r40 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r41 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r43 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r44 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r46 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r47 19 31 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.16
+ $Y2=0
r48 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.555
+ $Y2=0
r49 18 34 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=3.12
+ $Y2=0
r50 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.555
+ $Y2=0
r51 16 28 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.2
+ $Y2=0
r52 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.54
+ $Y2=0
r53 15 31 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=2.16
+ $Y2=0
r54 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.54
+ $Y2=0
r55 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=0.085
+ $X2=2.555 $Y2=0
r56 11 13 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.555 $Y=0.085
+ $X2=2.555 $Y2=0.595
r57 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.085 $X2=1.54
+ $Y2=0
r58 7 9 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.54 $Y=0.085 $X2=1.54
+ $Y2=0.595
r59 2 13 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.37 $X2=2.555 $Y2=0.595
r60 1 9 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=1.33
+ $Y=0.37 $X2=1.54 $Y2=0.595
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ms__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__nor4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.350000 9.475000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 7.555000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.920000 1.350000 5.155000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.413400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.920000 0.550000 1.930000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.373400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.570000 0.350000 1.820000 0.980000 ;
        RECT 1.570000 0.980000 2.830000 1.150000 ;
        RECT 2.025000 1.820000 3.305000 1.950000 ;
        RECT 2.025000 1.950000 5.635000 1.990000 ;
        RECT 2.025000 1.990000 2.355000 2.735000 ;
        RECT 2.500000 0.350000 2.830000 0.980000 ;
        RECT 2.500000 1.150000 2.830000 1.300000 ;
        RECT 2.500000 1.300000 3.750000 1.470000 ;
        RECT 2.975000 1.990000 5.635000 2.120000 ;
        RECT 2.975000 2.120000 3.305000 2.735000 ;
        RECT 3.500000 0.350000 3.750000 1.010000 ;
        RECT 3.500000 1.010000 9.465000 1.180000 ;
        RECT 3.500000 1.180000 3.750000 1.300000 ;
        RECT 4.905000 0.350000 5.235000 1.010000 ;
        RECT 5.405000 1.180000 5.635000 1.950000 ;
        RECT 6.250000 0.350000 6.580000 1.010000 ;
        RECT 7.250000 0.350000 7.580000 1.010000 ;
        RECT 8.275000 0.350000 8.525000 1.010000 ;
        RECT 9.215000 0.350000 9.465000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 10.080000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 10.270000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  2.100000  0.365000 3.245000 ;
      RECT 0.275000  0.420000  0.890000 0.750000 ;
      RECT 0.565000  2.100000  0.895000 2.980000 ;
      RECT 0.720000  0.750000  0.890000 1.320000 ;
      RECT 0.720000  1.320000  2.330000 1.650000 ;
      RECT 0.720000  1.650000  0.890000 2.100000 ;
      RECT 1.060000  0.085000  1.390000 1.130000 ;
      RECT 1.075000  2.100000  1.345000 3.245000 ;
      RECT 1.575000  1.820000  1.825000 2.905000 ;
      RECT 1.575000  2.905000  3.755000 3.075000 ;
      RECT 2.000000  0.085000  2.330000 0.790000 ;
      RECT 2.525000  2.160000  2.805000 2.905000 ;
      RECT 3.000000  0.085000  3.330000 1.130000 ;
      RECT 3.475000  2.320000  5.705000 2.460000 ;
      RECT 3.475000  2.460000  4.755000 2.490000 ;
      RECT 3.475000  2.490000  3.755000 2.905000 ;
      RECT 3.925000  2.660000  4.255000 2.905000 ;
      RECT 3.925000  2.905000  7.715000 3.075000 ;
      RECT 3.930000  0.085000  4.735000 0.840000 ;
      RECT 4.425000  2.290000  5.705000 2.320000 ;
      RECT 4.425000  2.490000  4.755000 2.720000 ;
      RECT 4.925000  2.630000  5.255000 2.905000 ;
      RECT 5.405000  0.085000  6.080000 0.840000 ;
      RECT 5.440000  2.460000  5.705000 2.540000 ;
      RECT 5.935000  1.950000  9.965000 2.120000 ;
      RECT 5.935000  2.120000  6.265000 2.735000 ;
      RECT 6.435000  2.290000  6.765000 2.905000 ;
      RECT 6.750000  0.085000  7.080000 0.805000 ;
      RECT 6.935000  2.120000  7.265000 2.735000 ;
      RECT 7.465000  2.290000  7.715000 2.905000 ;
      RECT 7.750000  0.085000  8.105000 0.805000 ;
      RECT 7.885000  2.120000  8.115000 2.980000 ;
      RECT 8.285000  2.290000  8.535000 3.245000 ;
      RECT 8.705000  0.085000  9.035000 0.805000 ;
      RECT 8.735000  2.120000  9.065000 2.980000 ;
      RECT 9.265000  2.290000  9.515000 3.245000 ;
      RECT 9.635000  0.085000  9.965000 1.130000 ;
      RECT 9.715000  1.820000  9.965000 1.950000 ;
      RECT 9.715000  2.120000  9.965000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_ms__nor4b_4
END LIBRARY

* File: sky130_fd_sc_ms__nor3_1.pxi.spice
* Created: Fri Aug 28 17:47:47 2020
* 
x_PM_SKY130_FD_SC_MS__NOR3_1%A N_A_M1001_g N_A_c_42_n N_A_M1003_g A A N_A_c_44_n
+ PM_SKY130_FD_SC_MS__NOR3_1%A
x_PM_SKY130_FD_SC_MS__NOR3_1%B N_B_M1005_g N_B_M1004_g B N_B_c_75_n
+ PM_SKY130_FD_SC_MS__NOR3_1%B
x_PM_SKY130_FD_SC_MS__NOR3_1%C N_C_M1000_g N_C_M1002_g C N_C_c_112_n N_C_c_113_n
+ PM_SKY130_FD_SC_MS__NOR3_1%C
x_PM_SKY130_FD_SC_MS__NOR3_1%VPWR N_VPWR_M1001_s N_VPWR_c_135_n N_VPWR_c_136_n
+ N_VPWR_c_137_n VPWR N_VPWR_c_138_n N_VPWR_c_134_n
+ PM_SKY130_FD_SC_MS__NOR3_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR3_1%Y N_Y_M1003_d N_Y_M1002_d N_Y_M1000_d N_Y_c_160_n
+ N_Y_c_161_n N_Y_c_162_n N_Y_c_163_n N_Y_c_164_n Y Y Y Y
+ PM_SKY130_FD_SC_MS__NOR3_1%Y
x_PM_SKY130_FD_SC_MS__NOR3_1%VGND N_VGND_M1003_s N_VGND_M1004_d N_VGND_c_211_n
+ N_VGND_c_212_n N_VGND_c_213_n N_VGND_c_214_n N_VGND_c_215_n VGND
+ N_VGND_c_216_n N_VGND_c_217_n N_VGND_c_218_n N_VGND_c_219_n
+ PM_SKY130_FD_SC_MS__NOR3_1%VGND
cc_1 VNB N_A_M1001_g 0.00559392f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A_c_42_n 0.0204394f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_3 VNB A 0.00896353f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_44_n 0.056984f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_5 VNB N_B_M1005_g 0.0015035f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_B_M1004_g 0.0218836f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_7 VNB B 0.00387716f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_B_c_75_n 0.0290066f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_9 VNB N_C_M1000_g 0.00198273f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_C_M1002_g 0.0310069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_C_c_112_n 0.0577187f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_12 VNB N_C_c_113_n 0.00431086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_134_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.232 $Y2=1.385
cc_14 VNB N_Y_c_160_n 0.00369654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_161_n 0.00168586f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_16 VNB N_Y_c_162_n 0.0160949f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_17 VNB N_Y_c_163_n 0.0227723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_164_n 0.00398282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_211_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_VGND_c_212_n 0.0158675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_213_n 0.0110726f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_22 VNB N_VGND_c_214_n 0.00568581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_215_n 0.00626527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_216_n 0.0150599f $X=-0.19 $Y=-0.245 $X2=0.232 $Y2=1.665
cc_25 VNB N_VGND_c_217_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_218_n 0.138456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_219_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A_M1001_g 0.0253567f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_29 VPB A 0.00799818f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_30 VPB N_B_M1005_g 0.023009f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_31 VPB B 0.00359542f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_32 VPB N_C_M1000_g 0.0304465f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_33 VPB N_C_c_113_n 0.00726331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_135_n 0.0140744f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_35 VPB N_VPWR_c_136_n 0.0395973f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_36 VPB N_VPWR_c_137_n 0.0063263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_138_n 0.0397956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_134_n 0.0513904f $X=-0.19 $Y=1.66 $X2=0.232 $Y2=1.385
cc_39 VPB N_Y_c_160_n 0.00221067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB Y 0.049735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 N_A_M1001_g N_B_M1005_g 0.0739843f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_42 N_A_c_42_n N_B_M1004_g 0.0113716f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_43 N_A_c_44_n N_B_M1004_g 0.0034836f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_44 N_A_c_44_n B 4.32487e-19 $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_45 N_A_c_44_n N_B_c_75_n 0.0204192f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_46 A N_VPWR_c_135_n 0.0223626f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A_c_44_n N_VPWR_c_135_n 0.00115632f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_48 N_A_M1001_g N_VPWR_c_136_n 0.0106922f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_49 N_A_M1001_g N_VPWR_c_137_n 0.00328578f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_50 N_A_M1001_g N_VPWR_c_138_n 0.00460063f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_51 N_A_M1001_g N_VPWR_c_134_n 0.00908371f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_52 N_A_M1001_g N_Y_c_160_n 0.0230441f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_53 N_A_c_42_n N_Y_c_160_n 0.00310315f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_54 A N_Y_c_160_n 0.0429724f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A_c_44_n N_Y_c_160_n 0.00817501f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_56 N_A_c_42_n N_Y_c_161_n 2.26494e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_57 N_A_c_42_n N_Y_c_164_n 0.00948239f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A_c_42_n N_VGND_c_212_n 0.00707603f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_59 A N_VGND_c_213_n 0.0221597f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_c_44_n N_VGND_c_213_n 0.00172545f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_61 N_A_c_42_n N_VGND_c_214_n 4.67172e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A_c_42_n N_VGND_c_215_n 0.00286134f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A_c_44_n N_VGND_c_215_n 9.43085e-19 $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_64 N_A_c_42_n N_VGND_c_216_n 0.00383152f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_65 N_A_c_42_n N_VGND_c_218_n 0.00757637f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_66 N_B_M1005_g N_C_M1000_g 0.0542681f $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_67 N_B_M1004_g N_C_M1002_g 0.0280261f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_68 B N_C_c_112_n 0.00409514f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B_c_75_n N_C_c_112_n 0.0209151f $X=0.96 $Y=1.465 $X2=0 $Y2=0
cc_70 B N_C_c_113_n 0.0388905f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_71 N_B_c_75_n N_C_c_113_n 2.3211e-19 $X=0.96 $Y=1.465 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_VPWR_c_136_n 5.45649e-19 $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_73 N_B_M1005_g N_VPWR_c_137_n 4.58619e-19 $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_74 N_B_M1005_g N_VPWR_c_138_n 0.00349978f $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_75 N_B_M1005_g N_VPWR_c_134_n 0.00429988f $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_76 N_B_M1005_g N_Y_c_160_n 0.00450827f $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_77 N_B_M1004_g N_Y_c_160_n 0.00356835f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_78 B N_Y_c_160_n 0.036899f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_79 N_B_c_75_n N_Y_c_160_n 0.0020371f $X=0.96 $Y=1.465 $X2=0 $Y2=0
cc_80 N_B_M1004_g N_Y_c_161_n 2.26494e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_81 N_B_M1004_g N_Y_c_162_n 0.0157822f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_82 B N_Y_c_162_n 0.0357518f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_83 N_B_c_75_n N_Y_c_162_n 0.00469027f $X=0.96 $Y=1.465 $X2=0 $Y2=0
cc_84 N_B_M1004_g N_Y_c_163_n 5.9203e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_85 N_B_c_75_n N_Y_c_164_n 4.44413e-19 $X=0.96 $Y=1.465 $X2=0 $Y2=0
cc_86 N_B_M1005_g Y 0.0457758f $X=0.915 $Y=2.4 $X2=0 $Y2=0
cc_87 B Y 0.0343349f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_88 N_B_c_75_n Y 5.33374e-19 $X=0.96 $Y=1.465 $X2=0 $Y2=0
cc_89 N_B_M1004_g N_VGND_c_212_n 4.66889e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_90 N_B_M1004_g N_VGND_c_214_n 0.00803107f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_VGND_c_216_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_92 N_B_M1004_g N_VGND_c_218_n 0.00757637f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_93 N_C_M1000_g N_VPWR_c_138_n 0.00349978f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_94 N_C_M1000_g N_VPWR_c_134_n 0.00433878f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_95 N_C_M1002_g N_Y_c_162_n 0.0193333f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_96 N_C_c_112_n N_Y_c_162_n 0.00305934f $X=1.65 $Y=1.465 $X2=0 $Y2=0
cc_97 N_C_c_113_n N_Y_c_162_n 0.0276802f $X=1.65 $Y=1.465 $X2=0 $Y2=0
cc_98 N_C_M1002_g N_Y_c_163_n 0.00889319f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_99 N_C_M1000_g Y 0.0414213f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_100 N_C_c_112_n Y 0.00152081f $X=1.65 $Y=1.465 $X2=0 $Y2=0
cc_101 N_C_c_113_n Y 0.026488f $X=1.65 $Y=1.465 $X2=0 $Y2=0
cc_102 N_C_M1002_g N_VGND_c_214_n 0.00503266f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_103 N_C_M1002_g N_VGND_c_217_n 0.00434272f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_104 N_C_M1002_g N_VGND_c_218_n 0.00824429f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_105 N_VPWR_c_137_n N_Y_c_160_n 0.0255419f $X=0.27 $Y=2.455 $X2=0 $Y2=0
cc_106 N_VPWR_c_138_n N_Y_c_160_n 0.00421728f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_107 N_VPWR_c_134_n N_Y_c_160_n 0.00350217f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_108 N_VPWR_c_138_n Y 0.0484359f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_109 N_VPWR_c_134_n Y 0.0394057f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_110 A_117_368# N_Y_c_160_n 0.00134035f $X=0.585 $Y=1.84 $X2=0.615 $Y2=1.95
cc_111 A_117_368# Y 0.0030224f $X=0.585 $Y=1.84 $X2=1.595 $Y2=2.32
cc_112 A_201_368# Y 0.00228446f $X=1.005 $Y=1.84 $X2=1.595 $Y2=2.32
cc_113 N_Y_c_162_n N_VGND_M1004_d 0.00253871f $X=1.475 $Y=1.005 $X2=0 $Y2=0
cc_114 N_Y_c_161_n N_VGND_c_212_n 0.0130608f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_115 N_Y_c_164_n N_VGND_c_213_n 0.0104845f $X=0.71 $Y=0.965 $X2=0 $Y2=0
cc_116 N_Y_c_161_n N_VGND_c_214_n 0.0130983f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_117 N_Y_c_162_n N_VGND_c_214_n 0.0215485f $X=1.475 $Y=1.005 $X2=0 $Y2=0
cc_118 N_Y_c_163_n N_VGND_c_214_n 0.0142986f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_119 N_Y_c_161_n N_VGND_c_216_n 0.00791198f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_120 N_Y_c_163_n N_VGND_c_217_n 0.0145639f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_121 N_Y_c_161_n N_VGND_c_218_n 0.00688042f $X=0.71 $Y=0.53 $X2=0 $Y2=0
cc_122 N_Y_c_163_n N_VGND_c_218_n 0.0119984f $X=1.64 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o21a_1.spice
* Created: Wed Sep  2 12:21:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21a_1.pex.spice"
.subckt sky130_fd_sc_ms__o21a_1  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_83_244#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_320_74#_M1002_d N_B1_M1002_g N_A_83_244#_M1002_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_320_74#_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_320_74#_M1001_d N_A1_M1001_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_83_244#_M1003_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.365857 AS=0.3136 PD=1.98286 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1000 N_A_83_244#_M1000_d N_B1_M1000_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=0.84
+ AD=0.142891 AS=0.274393 PD=1.20978 PS=1.48714 NRD=0 NRS=39.8531 M=1 R=4.66667
+ SA=90001 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1007 A_379_387# N_A2_M1007_g N_A_83_244#_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.170109 PD=1.39 PS=1.44022 NRD=27.5603 NRS=9.8303 M=1 R=5.55556
+ SA=90001.3 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_379_387# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.195 PD=2.56 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90001.8 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__o21a_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o22a_1.spice
* Created: Fri Aug 28 17:57:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o22a_1.pex.spice"
.subckt sky130_fd_sc_ms__o22a_1  VNB VPB B1 B2 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_83_260#_M1009_g N_X_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_83_260#_M1003_d N_B1_M1003_g N_A_299_139#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1024 AS=0.1705 PD=0.96 PS=1.85 NRD=3.744 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 N_A_299_139#_M1006_d N_B2_M1006_g N_A_83_260#_M1003_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=3.744 M=1 R=4.26667
+ SA=75000.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_299_139#_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.144737 AS=0.0896 PD=1.125 PS=0.92 NRD=15.936 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_299_139#_M1000_d N_A1_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.18205 AS=0.144737 PD=1.85 PS=1.125 NRD=0 NRS=14.052 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A_83_260#_M1002_g N_X_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.66566 AS=0.3136 PD=2.48302 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1005 A_401_392# N_B1_M1005_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.59434 PD=1.24 PS=2.21698 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_83_260#_M1007_d N_B2_M1007_g A_401_392# VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.12 PD=1.27 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90002
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1008 A_575_392# N_A2_M1008_g N_A_83_260#_M1007_d VPB PSHORT L=0.18 W=1 AD=0.18
+ AS=0.135 PD=1.36 PS=1.27 NRD=24.6053 NRS=0 M=1 R=5.55556 SA=90002.5 SB=90000.7
+ A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_575_392# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.18 PD=2.56 PS=1.36 NRD=0 NRS=24.6053 M=1 R=5.55556 SA=90003 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.81875 P=12.19
c_348 A_401_392# 0 1.51466e-19 $X=2.005 $Y=1.96
*
.include "sky130_fd_sc_ms__o22a_1.pxi.spice"
*
.ends
*
*

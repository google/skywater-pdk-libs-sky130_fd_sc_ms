* File: sky130_fd_sc_ms__buf_8.spice
* Created: Wed Sep  2 11:59:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__buf_8.pex.spice"
.subckt sky130_fd_sc_ms__buf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_A_27_74#_M1006_d N_A_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.12025 PD=2.05 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1015 N_A_27_74#_M1015_d N_A_M1015_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12025 PD=1.02 PS=1.065 NRD=0 NRS=7.296 M=1 R=4.93333 SA=75000.7
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1015_d N_A_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1000 N_X_M1000_d N_A_27_74#_M1000_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1000_d N_A_27_74#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1012_d N_A_27_74#_M1012_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.5
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1012_d N_A_27_74#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.9
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1016 N_X_M1016_d N_A_27_74#_M1016_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.5
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1017 N_X_M1016_d N_A_27_74#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.9
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1019 N_X_M1019_d N_A_27_74#_M1019_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1554 PD=1.025 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.5
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1019_d N_A_27_74#_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.2627 PD=1.025 PS=2.19 NRD=0.804 NRS=11.34 M=1 R=4.93333
+ SA=75004.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_74#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1001_d N_A_M1002_g N_A_27_74#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_74#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90004 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1003_d N_A_27_74#_M1004_g N_X_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.5
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_27_74#_M1005_g N_X_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1005_d N_A_27_74#_M1007_g N_X_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_74#_M1008_g N_X_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1008_d N_A_27_74#_M1010_g N_X_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.5
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1011 N_VPWR_M1011_d N_A_27_74#_M1011_g N_X_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1708 AS=0.1512 PD=1.425 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.9
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1011_d N_A_27_74#_M1014_g N_X_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1708 AS=0.1596 PD=1.425 PS=1.405 NRD=5.2599 NRS=1.7533 M=1 R=6.22222
+ SA=90004.4 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_27_74#_M1021_g N_X_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1596 PD=2.8 PS=1.405 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__buf_8.pxi.spice"
*
.ends
*
*

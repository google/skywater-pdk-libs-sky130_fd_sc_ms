* File: sky130_fd_sc_ms__or4bb_4.spice
* Created: Wed Sep  2 12:29:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4bb_4.pex.spice"
.subckt sky130_fd_sc_ms__or4bb_4  VNB VPB D_N C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_N_M1008_g N_A_27_94#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.137739 AS=0.1824 PD=1.08058 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1008_d N_A_193_277#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.159261 AS=0.1036 PD=1.24942 PS=1.02 NRD=12.156 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_193_277#_M1015_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19035 AS=0.1036 PD=1.37 PS=1.02 NRD=32.784 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1015_d N_A_193_277#_M1019_g N_X_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19035 AS=0.24235 PD=1.37 PS=1.395 NRD=32.784 NRS=0 M=1 R=4.93333
+ SA=75001.7 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_193_277#_M1020_g N_X_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13883 AS=0.24235 PD=1.17971 PS=1.395 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_A_681_368#_M1009_d N_C_N_M1009_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1719 AS=0.12007 PD=1.85 PS=1.02029 NRD=0 NRS=15.936 M=1 R=4.26667
+ SA=75003.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_193_277#_M1017_d N_A_27_94#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.53465 AS=0.327 PD=2.185 PS=3.11 NRD=0 NRS=62.736 M=1 R=4.93333
+ SA=75000.2 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_681_368#_M1021_g N_A_193_277#_M1017_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.18315 AS=0.53465 PD=1.235 PS=2.185 NRD=11.34 NRS=0 M=1
+ R=4.93333 SA=75001.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_193_277#_M1014_d N_B_M1014_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.17205 AS=0.18315 PD=1.205 PS=1.235 NRD=0 NRS=23.508 M=1 R=4.93333
+ SA=75002.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_193_277#_M1014_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.4625 AS=0.17205 PD=2.73 PS=1.205 NRD=0 NRS=30 M=1 R=4.93333 SA=75003.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_D_N_M1011_g N_A_27_94#_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.191226 AS=0.28 PD=1.40566 PS=2.56 NRD=17.7103 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90003 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_193_277#_M1003_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.214174 PD=1.39 PS=1.57434 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90000.7 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1003_d N_A_193_277#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2044 PD=1.39 PS=1.485 NRD=0 NRS=7.0329 M=1 R=6.22222 SA=90001.1
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1012_d N_A_193_277#_M1012_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.2044 PD=1.67 PS=1.485 NRD=6.1464 NRS=7.8997 M=1 R=6.22222
+ SA=90001.7 SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1013 N_X_M1012_d N_A_193_277#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.205298 PD=1.67 PS=1.55849 NRD=41.3306 NRS=0 M=1 R=6.22222
+ SA=90002.4 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1022 N_A_681_368#_M1022_d N_C_N_M1022_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.183302 PD=2.56 PS=1.39151 NRD=0 NRS=16.7253 M=1 R=5.55556
+ SA=90003 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_A_193_277#_M1006_d N_A_27_94#_M1006_g N_A_791_392#_M1006_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1010 N_A_193_277#_M1006_d N_A_27_94#_M1010_g N_A_791_392#_M1010_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1016 N_A_791_392#_M1010_s N_A_681_368#_M1016_g N_A_1063_392#_M1016_s VPB
+ PSHORT L=0.18 W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1
+ R=5.55556 SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1018 N_A_791_392#_M1018_d N_A_681_368#_M1018_g N_A_1063_392#_M1016_s VPB
+ PSHORT L=0.18 W=1 AD=0.28 AS=0.16 PD=2.56 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_1273_392#_M1000_d N_B_M1000_g N_A_1063_392#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1023 N_A_1273_392#_M1023_d N_B_M1023_g N_A_1063_392#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1002 N_A_1273_392#_M1023_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1004 N_A_1273_392#_M1004_d N_A_M1004_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.16 PD=2.56 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__or4bb_4.pxi.spice"
*
.ends
*
*

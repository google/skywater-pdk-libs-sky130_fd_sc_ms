# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfstp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.820000 1.585000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.990000 0.370000 14.345000 1.150000 ;
        RECT 13.995000 1.820000 14.755000 2.150000 ;
        RECT 13.995000 2.150000 14.275000 2.980000 ;
        RECT 14.175000 1.150000 14.345000 1.320000 ;
        RECT 14.175000 1.320000 14.755000 1.490000 ;
        RECT 14.325000 1.490000 14.755000 1.820000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.140000 2.780000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 1.410000 2.045000 1.580000 ;
        RECT 0.475000 1.580000 0.805000 2.140000 ;
        RECT 1.795000 1.250000 2.045000 1.410000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.205000 1.210000  7.555000 1.555000 ;
        RECT 11.445000 1.180000 11.875000 1.800000 ;
      LAYER mcon ;
        RECT  7.355000 1.210000  7.525000 1.380000 ;
        RECT 11.675000 1.210000 11.845000 1.380000 ;
      LAYER met1 ;
        RECT  7.295000 1.180000  7.585000 1.225000 ;
        RECT  7.295000 1.225000 11.905000 1.365000 ;
        RECT  7.295000 1.365000  7.585000 1.410000 ;
        RECT 11.615000 1.180000 11.905000 1.225000 ;
        RECT 11.615000 1.365000 11.905000 1.410000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.300000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.880000 0.085000 ;
        RECT  0.615000  0.085000  1.070000 0.680000 ;
        RECT  2.460000  0.085000  2.790000 0.740000 ;
        RECT  3.520000  0.085000  3.850000 1.010000 ;
        RECT  6.130000  0.085000  6.460000 0.360000 ;
        RECT  7.510000  0.085000  8.010000 0.680000 ;
        RECT  8.690000  0.085000  9.020000 0.715000 ;
        RECT 11.640000  0.085000 12.330000 0.600000 ;
        RECT 13.555000  0.085000 13.805000 1.150000 ;
        RECT 14.515000  0.085000 14.765000 1.150000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.880000 3.415000 ;
        RECT  0.565000 2.660000  0.895000 3.245000 ;
        RECT  2.560000 2.830000  2.890000 3.245000 ;
        RECT  3.545000 2.580000  3.875000 3.245000 ;
        RECT  6.095000 2.425000  6.345000 3.245000 ;
        RECT  7.535000 2.065000  7.705000 3.245000 ;
        RECT  8.435000 2.405000  8.685000 3.245000 ;
        RECT 11.080000 2.645000 11.330000 3.245000 ;
        RECT 12.510000 2.650000 12.840000 3.245000 ;
        RECT 13.540000 1.820000 13.825000 3.245000 ;
        RECT 14.445000 2.320000 14.775000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.350000  0.445000 0.900000 ;
      RECT  0.115000 0.900000  1.225000 1.230000 ;
      RECT  0.115000 1.230000  0.285000 2.310000 ;
      RECT  0.115000 2.310000  0.365000 2.320000 ;
      RECT  0.115000 2.320000  2.045000 2.490000 ;
      RECT  0.115000 2.490000  0.365000 2.980000 ;
      RECT  1.435000 2.660000  2.385000 2.910000 ;
      RECT  1.560000 0.350000  1.890000 0.910000 ;
      RECT  1.560000 0.910000  2.385000 1.080000 ;
      RECT  1.795000 1.830000  2.045000 2.320000 ;
      RECT  2.215000 1.080000  2.385000 2.490000 ;
      RECT  2.215000 2.490000  3.120000 2.660000 ;
      RECT  2.950000 2.240000  4.915000 2.410000 ;
      RECT  2.950000 2.410000  3.120000 2.490000 ;
      RECT  2.960000 0.350000  3.350000 1.010000 ;
      RECT  2.960000 1.010000  3.130000 1.820000 ;
      RECT  2.960000 1.820000  4.215000 2.070000 ;
      RECT  3.885000 1.350000  4.215000 1.820000 ;
      RECT  4.030000 0.255000  5.170000 0.425000 ;
      RECT  4.030000 0.425000  4.200000 1.130000 ;
      RECT  4.075000 2.580000  4.325000 2.895000 ;
      RECT  4.075000 2.895000  5.730000 3.065000 ;
      RECT  4.420000 0.595000  4.830000 0.845000 ;
      RECT  4.420000 0.845000  4.590000 1.900000 ;
      RECT  4.420000 1.900000  4.915000 2.070000 ;
      RECT  4.585000 2.070000  4.915000 2.240000 ;
      RECT  4.585000 2.410000  4.915000 2.725000 ;
      RECT  4.760000 1.015000  5.170000 1.185000 ;
      RECT  4.760000 1.185000  4.965000 1.730000 ;
      RECT  5.000000 0.425000  5.170000 1.015000 ;
      RECT  5.115000 2.265000  5.365000 2.725000 ;
      RECT  5.135000 1.375000  6.880000 1.545000 ;
      RECT  5.135000 1.545000  5.305000 2.265000 ;
      RECT  5.340000 0.385000  5.590000 1.375000 ;
      RECT  5.475000 1.715000  5.730000 2.045000 ;
      RECT  5.560000 2.045000  5.730000 2.085000 ;
      RECT  5.560000 2.085000  6.685000 2.255000 ;
      RECT  5.560000 2.255000  5.730000 2.895000 ;
      RECT  5.940000 1.715000  6.270000 1.745000 ;
      RECT  5.940000 1.745000  7.025000 1.915000 ;
      RECT  5.980000 0.530000  7.020000 0.700000 ;
      RECT  5.980000 0.700000  6.310000 1.205000 ;
      RECT  6.515000 2.255000  6.685000 2.905000 ;
      RECT  6.515000 2.905000  7.365000 3.075000 ;
      RECT  6.550000 0.870000  7.925000 1.040000 ;
      RECT  6.550000 1.040000  6.880000 1.375000 ;
      RECT  6.550000 1.545000  6.880000 1.570000 ;
      RECT  6.690000 0.350000  7.020000 0.530000 ;
      RECT  6.855000 1.915000  7.025000 2.735000 ;
      RECT  7.195000 1.725000 10.170000 1.805000 ;
      RECT  7.195000 1.805000  8.425000 1.895000 ;
      RECT  7.195000 1.895000  7.365000 2.905000 ;
      RECT  7.755000 1.040000  7.925000 1.225000 ;
      RECT  7.755000 1.225000  8.085000 1.555000 ;
      RECT  7.905000 2.065000  9.830000 2.145000 ;
      RECT  7.905000 2.145000  8.765000 2.235000 ;
      RECT  7.905000 2.235000  8.235000 2.755000 ;
      RECT  8.180000 0.350000  8.510000 0.885000 ;
      RECT  8.180000 0.885000 10.080000 1.055000 ;
      RECT  8.255000 1.475000 10.170000 1.725000 ;
      RECT  8.595000 1.975000  9.830000 2.065000 ;
      RECT  9.000000 2.315000  9.330000 2.905000 ;
      RECT  9.000000 2.905000 10.435000 3.075000 ;
      RECT  9.250000 0.255000 10.580000 0.425000 ;
      RECT  9.250000 0.425000  9.580000 0.715000 ;
      RECT  9.500000 2.145000  9.830000 2.735000 ;
      RECT  9.750000 0.595000 10.080000 0.885000 ;
      RECT 10.000000 1.805000 10.720000 2.135000 ;
      RECT 10.105000 2.305000 11.860000 2.475000 ;
      RECT 10.105000 2.475000 10.435000 2.905000 ;
      RECT 10.250000 0.425000 10.580000 0.810000 ;
      RECT 10.410000 0.810000 10.580000 1.400000 ;
      RECT 10.410000 1.400000 11.060000 1.570000 ;
      RECT 10.890000 1.570000 11.060000 1.970000 ;
      RECT 10.890000 1.970000 12.465000 2.140000 ;
      RECT 10.890000 2.140000 11.860000 2.305000 ;
      RECT 10.945000 0.790000 12.805000 0.960000 ;
      RECT 10.945000 0.960000 11.275000 1.230000 ;
      RECT 11.530000 2.475000 11.860000 2.980000 ;
      RECT 12.060000 2.310000 12.805000 2.480000 ;
      RECT 12.060000 2.480000 12.310000 2.980000 ;
      RECT 12.135000 1.130000 12.465000 1.970000 ;
      RECT 12.500000 0.350000 12.805000 0.790000 ;
      RECT 12.635000 0.960000 12.805000 2.310000 ;
      RECT 13.035000 0.470000 13.365000 1.320000 ;
      RECT 13.035000 1.320000 14.005000 1.650000 ;
      RECT 13.035000 1.650000 13.370000 2.980000 ;
  END
END sky130_fd_sc_ms__sdfstp_2

* File: sky130_fd_sc_ms__nand3b_4.pex.spice
* Created: Wed Sep  2 12:14:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND3B_4%A_N 3 5 7 8 10 12 13 20 21
c51 20 0 5.29186e-20 $X=0.93 $Y=1.515
r52 19 21 46.0284 $w=4.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.557
+ $X2=1.095 $Y2=1.557
r53 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.515 $X2=0.93 $Y2=1.515
r54 17 19 4.69045 $w=4.15e-07 $l=3.5e-08 $layer=POLY_cond $X=0.895 $Y=1.557
+ $X2=0.93 $Y2=1.557
r55 13 20 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.76 $Y=1.665
+ $X2=0.76 $Y2=1.515
r56 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=1.345 $Y=1.765
+ $X2=1.345 $Y2=2.26
r57 8 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.255 $Y=1.69
+ $X2=1.345 $Y2=1.765
r58 8 21 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.255 $Y=1.69
+ $X2=1.095 $Y2=1.69
r59 5 17 22.3416 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.895 $Y=1.765
+ $X2=0.895 $Y2=1.557
r60 5 7 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=0.895 $Y=1.765
+ $X2=0.895 $Y2=2.26
r61 1 17 12.0612 $w=4.15e-07 $l=9e-08 $layer=POLY_cond $X=0.805 $Y=1.557
+ $X2=0.895 $Y2=1.557
r62 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.805 $Y=1.35
+ $X2=0.805 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%C 1 3 4 5 6 8 9 11 14 18 20 22 24 25 26 27
+ 31
c78 5 0 2.71579e-20 $X=1.485 $Y=1.3
r79 41 43 15.279 $w=4.55e-07 $l=1.25e-07 $layer=POLY_cond $X=2.95 $Y=1.452
+ $X2=3.075 $Y2=1.452
r80 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.515 $X2=2.95 $Y2=1.515
r81 39 41 39.7253 $w=4.55e-07 $l=3.25e-07 $layer=POLY_cond $X=2.625 $Y=1.452
+ $X2=2.95 $Y2=1.452
r82 37 39 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=2.61 $Y=1.452
+ $X2=2.625 $Y2=1.452
r83 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r84 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.515 $X2=1.93 $Y2=1.515
r85 31 33 71.5055 $w=4.55e-07 $l=5.85e-07 $layer=POLY_cond $X=2.515 $Y=1.452
+ $X2=1.93 $Y2=1.452
r86 27 42 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.95 $Y2=1.565
r87 26 42 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.95 $Y2=1.565
r88 26 38 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.61
+ $Y2=1.565
r89 25 38 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.61 $Y2=1.565
r90 25 34 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.93 $Y2=1.565
r91 23 33 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=1.915 $Y=1.452
+ $X2=1.93 $Y2=1.452
r92 23 24 11.0167 $w=3.02e-07 $l=7.5e-08 $layer=POLY_cond $X=1.915 $Y=1.452
+ $X2=1.84 $Y2=1.452
r93 20 43 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=3.09 $Y=1.452
+ $X2=3.075 $Y2=1.452
r94 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.09 $Y=1.225
+ $X2=3.09 $Y2=0.78
r95 16 43 24.5593 $w=1.8e-07 $l=2.28e-07 $layer=POLY_cond $X=3.075 $Y=1.68
+ $X2=3.075 $Y2=1.452
r96 16 18 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.075 $Y=1.68
+ $X2=3.075 $Y2=2.4
r97 12 39 24.5593 $w=1.8e-07 $l=2.28e-07 $layer=POLY_cond $X=2.625 $Y=1.68
+ $X2=2.625 $Y2=1.452
r98 12 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.625 $Y=1.68
+ $X2=2.625 $Y2=2.4
r99 9 37 2.44463 $w=4.55e-07 $l=2e-08 $layer=POLY_cond $X=2.59 $Y=1.452 $X2=2.61
+ $Y2=1.452
r100 9 31 9.16737 $w=4.55e-07 $l=7.5e-08 $layer=POLY_cond $X=2.59 $Y=1.452
+ $X2=2.515 $Y2=1.452
r101 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.59 $Y=1.225
+ $X2=2.59 $Y2=0.78
r102 6 24 15.6242 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=1.84 $Y=1.225
+ $X2=1.84 $Y2=1.452
r103 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.84 $Y=1.225
+ $X2=1.84 $Y2=0.78
r104 4 24 11.0167 $w=3.02e-07 $l=1.85753e-07 $layer=POLY_cond $X=1.765 $Y=1.3
+ $X2=1.84 $Y2=1.452
r105 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.765 $Y=1.3
+ $X2=1.485 $Y2=1.3
r106 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.225
+ $X2=1.485 $Y2=1.3
r107 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.41 $Y=1.225
+ $X2=1.41 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%A_89_172# 1 2 9 11 13 16 18 20 21 23 25 26
+ 28 30 31 32 34 39 40 44 48 52 53 66
c127 52 0 1.74867e-19 $X=1.35 $Y=1.095
c128 26 0 2.37294e-19 $X=5.32 $Y=1.26
c129 18 0 3.1443e-19 $X=4.535 $Y=1.185
r130 57 59 9.37338 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.407
+ $X2=3.69 $Y2=1.407
r131 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.765
+ $Y=1.465 $X2=3.765 $Y2=1.465
r132 53 56 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.685 $Y2=1.465
r133 48 50 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.59 $Y=1.005
+ $X2=0.59 $Y2=1.095
r134 45 64 9.37338 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=4.445 $Y=1.407
+ $X2=4.52 $Y2=1.407
r135 44 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.445 $Y=1.465
+ $X2=3.77 $Y2=1.465
r136 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.445
+ $Y=1.465 $X2=4.445 $Y2=1.465
r137 41 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=1.095
+ $X2=1.35 $Y2=1.095
r138 40 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.095
+ $X2=3.685 $Y2=1.095
r139 40 41 141.246 $w=1.68e-07 $l=2.165e-06 $layer=LI1_cond $X=3.6 $Y=1.095
+ $X2=1.435 $Y2=1.095
r140 38 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=1.18
+ $X2=1.35 $Y2=1.095
r141 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.35 $Y=1.18
+ $X2=1.35 $Y2=1.95
r142 34 39 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.265 $Y=2.045
+ $X2=1.35 $Y2=1.95
r143 34 36 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.265 $Y=2.045
+ $X2=1.12 $Y2=2.045
r144 33 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=1.095
+ $X2=0.59 $Y2=1.095
r145 32 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=1.095
+ $X2=1.35 $Y2=1.095
r146 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.265 $Y=1.095
+ $X2=0.755 $Y2=1.095
r147 28 30 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.395 $Y=1.185
+ $X2=5.395 $Y2=0.74
r148 27 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.04 $Y=1.26
+ $X2=4.965 $Y2=1.26
r149 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.32 $Y=1.26
+ $X2=5.395 $Y2=1.185
r150 26 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.32 $Y=1.26
+ $X2=5.04 $Y2=1.26
r151 23 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=1.26
r152 23 25 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=0.74
r153 21 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.89 $Y=1.26
+ $X2=4.965 $Y2=1.26
r154 21 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.89 $Y=1.26
+ $X2=4.61 $Y2=1.26
r155 18 66 35.5547 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=4.535 $Y=1.407
+ $X2=4.61 $Y2=1.407
r156 18 64 1.87468 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=4.535 $Y=1.407
+ $X2=4.52 $Y2=1.407
r157 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=0.74
r158 14 64 24.0211 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=4.52 $Y=1.63
+ $X2=4.52 $Y2=1.407
r159 14 16 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.52 $Y=1.63
+ $X2=4.52 $Y2=2.4
r160 11 45 45.6171 $w=4.45e-07 $l=3.65e-07 $layer=POLY_cond $X=4.08 $Y=1.407
+ $X2=4.445 $Y2=1.407
r161 11 57 39.3682 $w=4.45e-07 $l=3.15e-07 $layer=POLY_cond $X=4.08 $Y=1.407
+ $X2=3.765 $Y2=1.407
r162 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.08 $Y=1.185
+ $X2=4.08 $Y2=0.74
r163 7 59 24.0211 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=3.69 $Y=1.63
+ $X2=3.69 $Y2=1.407
r164 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.69 $Y=1.63 $X2=3.69
+ $Y2=2.4
r165 2 36 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.84 $X2=1.12 $Y2=2.045
r166 1 48 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.445
+ $Y=0.86 $X2=0.59 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%B 1 3 4 5 8 10 12 15 19 23 25 26 27 39 40
c67 40 0 6.5646e-20 $X=6.965 $Y=1.485
c68 39 0 1.64144e-19 $X=6.965 $Y=1.485
c69 8 0 1.10856e-19 $X=5.895 $Y=0.74
r70 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.965
+ $Y=1.485 $X2=6.965 $Y2=1.485
r71 37 39 26.155 $w=3.87e-07 $l=2.1e-07 $layer=POLY_cond $X=6.755 $Y=1.522
+ $X2=6.965 $Y2=1.522
r72 36 37 53.5556 $w=3.87e-07 $l=4.3e-07 $layer=POLY_cond $X=6.325 $Y=1.522
+ $X2=6.755 $Y2=1.522
r73 34 36 47.3282 $w=3.87e-07 $l=3.8e-07 $layer=POLY_cond $X=5.945 $Y=1.522
+ $X2=6.325 $Y2=1.522
r74 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.945
+ $Y=1.485 $X2=5.945 $Y2=1.485
r75 32 34 4.35917 $w=3.87e-07 $l=3.5e-08 $layer=POLY_cond $X=5.91 $Y=1.522
+ $X2=5.945 $Y2=1.522
r76 31 32 1.86822 $w=3.87e-07 $l=1.5e-08 $layer=POLY_cond $X=5.895 $Y=1.522
+ $X2=5.91 $Y2=1.522
r77 27 40 0.127242 $w=4.68e-07 $l=5e-09 $layer=LI1_cond $X=6.96 $Y=1.415
+ $X2=6.965 $Y2=1.415
r78 26 27 12.2153 $w=4.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.415
+ $X2=6.96 $Y2=1.415
r79 25 26 12.2153 $w=4.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6 $Y=1.415 $X2=6.48
+ $Y2=1.415
r80 25 35 1.39967 $w=4.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6 $Y=1.415 $X2=5.945
+ $Y2=1.415
r81 21 39 27.4005 $w=3.87e-07 $l=3.04697e-07 $layer=POLY_cond $X=7.185 $Y=1.32
+ $X2=6.965 $Y2=1.522
r82 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.185 $Y=1.32
+ $X2=7.185 $Y2=0.74
r83 17 37 25.0561 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=6.755 $Y=1.32
+ $X2=6.755 $Y2=1.522
r84 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.755 $Y=1.32
+ $X2=6.755 $Y2=0.74
r85 13 36 25.0561 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=6.325 $Y=1.32
+ $X2=6.325 $Y2=1.522
r86 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.325 $Y=1.32
+ $X2=6.325 $Y2=0.74
r87 10 32 20.6767 $w=1.8e-07 $l=2.03e-07 $layer=POLY_cond $X=5.91 $Y=1.725
+ $X2=5.91 $Y2=1.522
r88 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.91 $Y=1.725
+ $X2=5.91 $Y2=2.4
r89 6 31 25.0561 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=5.895 $Y=1.32
+ $X2=5.895 $Y2=1.522
r90 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.895 $Y=1.32
+ $X2=5.895 $Y2=0.74
r91 4 31 38.0952 $w=3.87e-07 $l=2.0944e-07 $layer=POLY_cond $X=5.74 $Y=1.65
+ $X2=5.895 $Y2=1.522
r92 4 5 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.74 $Y=1.65 $X2=5.55
+ $Y2=1.65
r93 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.46 $Y=1.725
+ $X2=5.55 $Y2=1.65
r94 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.46 $Y=1.725 $X2=5.46
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%VPWR 1 2 3 4 5 16 18 22 24 26 33 48 54 56
+ 61 64 76 79
c69 76 0 1.64144e-19 $X=7.4 $Y=2.325
r70 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r71 76 78 0.461248 $w=1.058e-06 $l=4e-08 $layer=LI1_cond $X=7.4 $Y=2.787
+ $X2=7.44 $Y2=2.787
r72 74 76 9.74386 $w=1.058e-06 $l=8.45e-07 $layer=LI1_cond $X=6.555 $Y=2.787
+ $X2=7.4 $Y2=2.787
r73 72 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r74 71 74 0.864839 $w=1.058e-06 $l=7.5e-08 $layer=LI1_cond $X=6.48 $Y=2.787
+ $X2=6.555 $Y2=2.787
r75 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r76 69 71 3.97826 $w=1.058e-06 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=2.787
+ $X2=6.48 $Y2=2.787
r77 67 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r78 66 69 1.55671 $w=1.058e-06 $l=1.35e-07 $layer=LI1_cond $X=6 $Y=2.787
+ $X2=6.135 $Y2=2.787
r79 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r80 63 64 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=3.032
+ $X2=5.4 $Y2=3.032
r81 60 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r82 59 63 3.04883 $w=7.63e-07 $l=1.95e-07 $layer=LI1_cond $X=5.04 $Y=3.032
+ $X2=5.235 $Y2=3.032
r83 59 61 15.8294 $w=7.63e-07 $l=4.6e-07 $layer=LI1_cond $X=5.04 $Y=3.032
+ $X2=4.58 $Y2=3.032
r84 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r86 53 54 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=3.032
+ $X2=2.565 $Y2=3.032
r87 50 53 3.7524 $w=7.63e-07 $l=2.4e-07 $layer=LI1_cond $X=2.16 $Y=3.032 $X2=2.4
+ $Y2=3.032
r88 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r89 47 50 7.89568 $w=7.63e-07 $l=5.05e-07 $layer=LI1_cond $X=1.655 $Y=3.032
+ $X2=2.16 $Y2=3.032
r90 47 48 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=3.032
+ $X2=1.49 $Y2=3.032
r91 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 41 61 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=4.58
+ $Y2=3.33
r94 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 39 56 11.2236 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.382 $Y2=3.33
r96 39 41 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 37 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r98 37 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 36 54 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.565 $Y2=3.33
r100 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 33 56 11.2236 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.382 $Y2=3.33
r102 33 36 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 32 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 32 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 31 48 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=1.49 $Y2=3.33
r106 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 29 44 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r108 29 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 26 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 26 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r111 24 66 11.613 $w=1.058e-06 $l=5.57798e-07 $layer=LI1_cond $X=5.97 $Y=3.33
+ $X2=6 $Y2=2.787
r112 24 64 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.97 $Y=3.33
+ $X2=5.4 $Y2=3.33
r113 20 56 2.04857 $w=4.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.382 $Y=3.245
+ $X2=3.382 $Y2=3.33
r114 20 22 10.3902 $w=4.93e-07 $l=4.3e-07 $layer=LI1_cond $X=3.382 $Y=3.245
+ $X2=3.382 $Y2=2.815
r115 16 44 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r116 16 18 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.495
r117 5 76 200 $w=1.7e-07 $l=1.6245e-06 $layer=licon1_PDIFF $count=3 $X=6 $Y=1.84
+ $X2=7.4 $Y2=2.325
r118 5 74 200 $w=1.7e-07 $l=7.59737e-07 $layer=licon1_PDIFF $count=3 $X=6
+ $Y=1.84 $X2=6.555 $Y2=2.325
r119 5 69 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6
+ $Y=1.84 $X2=6.135 $Y2=2.815
r120 4 63 300 $w=1.7e-07 $l=1.249e-06 $layer=licon1_PDIFF $count=2 $X=4.61
+ $Y=1.84 $X2=5.235 $Y2=2.815
r121 3 22 600 $w=1.7e-07 $l=1.07715e-06 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.84 $X2=3.38 $Y2=2.815
r122 2 53 300 $w=1.7e-07 $l=1.37532e-06 $layer=licon1_PDIFF $count=2 $X=1.435
+ $Y=1.84 $X2=2.4 $Y2=2.815
r123 2 47 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.84 $X2=1.655 $Y2=2.815
r124 1 18 600 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%Y 1 2 3 4 5 20 21 24 30 32 34 35 36 37 41
c65 41 0 1.74292e-19 $X=5.04 $Y=1.13
c66 36 0 1.10856e-19 $X=5.04 $Y=1.295
c67 34 0 1.70138e-19 $X=5.04 $Y=1.98
r68 36 37 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.665
r69 36 41 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.13
r70 35 41 3.90668 $w=2.3e-07 $l=2.22486e-07 $layer=LI1_cond $X=5.135 $Y=0.95
+ $X2=5.04 $Y2=1.13
r71 33 37 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.04 $Y=1.82
+ $X2=5.04 $Y2=1.665
r72 33 34 2.55462 $w=2.3e-07 $l=1.6e-07 $layer=LI1_cond $X=5.04 $Y=1.82 $X2=5.04
+ $Y2=1.98
r73 28 34 3.89311 $w=3.2e-07 $l=1.15e-07 $layer=LI1_cond $X=5.155 $Y=1.98
+ $X2=5.04 $Y2=1.98
r74 28 30 19.0873 $w=3.18e-07 $l=5.3e-07 $layer=LI1_cond $X=5.155 $Y=1.98
+ $X2=5.685 $Y2=1.98
r75 24 35 3.19638 $w=3.3e-07 $l=2.17371e-07 $layer=LI1_cond $X=4.925 $Y=0.965
+ $X2=5.135 $Y2=0.95
r76 24 26 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=4.925 $Y=0.965
+ $X2=4.305 $Y2=0.965
r77 21 32 7.64885 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=3.91 $Y=1.98
+ $X2=3.75 $Y2=1.98
r78 21 23 13.8653 $w=3.18e-07 $l=3.85e-07 $layer=LI1_cond $X=3.91 $Y=1.98
+ $X2=4.295 $Y2=1.98
r79 20 34 3.89311 $w=3.2e-07 $l=1.15e-07 $layer=LI1_cond $X=4.925 $Y=1.98
+ $X2=5.04 $Y2=1.98
r80 20 23 22.6887 $w=3.18e-07 $l=6.3e-07 $layer=LI1_cond $X=4.925 $Y=1.98
+ $X2=4.295 $Y2=1.98
r81 18 32 52.5359 $w=1.88e-07 $l=9e-07 $layer=LI1_cond $X=2.85 $Y=2.045 $X2=3.75
+ $Y2=2.045
r82 5 30 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=5.55
+ $Y=1.84 $X2=5.685 $Y2=2.02
r83 4 23 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.78
+ $Y=1.84 $X2=4.295 $Y2=1.985
r84 3 18 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.84 $X2=2.85 $Y2=2.045
r85 2 35 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.37 $X2=5.18 $Y2=0.91
r86 1 26 182 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.37 $X2=4.305 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%VGND 1 2 3 12 15 22 23 24 30 42 43 47
c67 1 0 1.74867e-19 $X=0.88 $Y=0.41
r68 47 50 8.17727 $w=4.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.215 $Y=0
+ $X2=2.215 $Y2=0.335
r69 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r71 39 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=7.44
+ $Y2=0
r72 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r73 37 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r74 37 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r75 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r76 34 47 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.215
+ $Y2=0
r77 34 36 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=3.12
+ $Y2=0
r78 33 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r79 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r80 30 47 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=2.215
+ $Y2=0
r81 30 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=1.68
+ $Y2=0
r82 28 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r83 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r84 24 43 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=7.44
+ $Y2=0
r85 24 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r86 22 36 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.12
+ $Y2=0
r87 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.305
+ $Y2=0
r88 21 39 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.6
+ $Y2=0
r89 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.305
+ $Y2=0
r90 17 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r91 15 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.72
+ $Y2=0
r92 15 19 10.8563 $w=3.43e-07 $l=3.25e-07 $layer=LI1_cond $X=1.107 $Y=0
+ $X2=1.107 $Y2=0.325
r93 15 17 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.107 $Y=0 $X2=1.28
+ $Y2=0
r94 10 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0
r95 10 12 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0.615
r96 3 12 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.41 $X2=3.305 $Y2=0.615
r97 2 50 182 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.41 $X2=2.215 $Y2=0.335
r98 1 19 182 $w=1.7e-07 $l=2.64102e-07 $layer=licon1_NDIFF $count=1 $X=0.88
+ $Y=0.41 $X2=1.105 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%A_297_82# 1 2 3 4 14 16 17 18 20 21 22 23
+ 25 32 33 34 36 39 40 42
c125 39 0 2.57607e-20 $X=1.46 $Y=0.615
r126 42 44 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.805 $Y=0.615
+ $X2=2.805 $Y2=0.755
r127 38 40 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0.615
+ $X2=1.79 $Y2=0.615
r128 38 39 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0.615
+ $X2=1.46 $Y2=0.615
r129 35 36 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=7.33 $Y=1.01
+ $X2=7.33 $Y2=1.82
r130 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.245 $Y=1.905
+ $X2=7.33 $Y2=1.82
r131 33 34 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=7.245 $Y=1.905
+ $X2=6.23 $Y2=1.905
r132 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.145 $Y=1.99
+ $X2=6.23 $Y2=1.905
r133 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.145 $Y=1.99
+ $X2=6.145 $Y2=2.31
r134 27 30 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=6.11 $Y=0.925
+ $X2=6.97 $Y2=0.925
r135 25 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.245 $Y=0.925
+ $X2=7.33 $Y2=1.01
r136 25 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.245 $Y=0.925
+ $X2=6.97 $Y2=0.925
r137 23 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0.755
+ $X2=2.805 $Y2=0.755
r138 23 40 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.64 $Y=0.755
+ $X2=1.79 $Y2=0.755
r139 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.06 $Y=2.395
+ $X2=6.145 $Y2=2.31
r140 21 22 344.144 $w=1.68e-07 $l=5.275e-06 $layer=LI1_cond $X=6.06 $Y=2.395
+ $X2=0.785 $Y2=2.395
r141 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=2.31
+ $X2=0.785 $Y2=2.395
r142 19 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.7 $Y=2.12 $X2=0.7
+ $Y2=2.31
r143 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.7 $Y2=2.12
r144 17 18 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.255 $Y2=2.035
r145 16 39 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=0.255 $Y=0.665
+ $X2=1.46 $Y2=0.665
r146 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.95
+ $X2=0.255 $Y2=2.035
r147 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.255 $Y2=0.665
r148 13 14 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.17 $Y2=1.95
r149 4 30 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=6.83
+ $Y=0.37 $X2=6.97 $Y2=0.925
r150 3 27 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.37 $X2=6.11 $Y2=0.925
r151 2 42 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.41 $X2=2.805 $Y2=0.615
r152 1 38 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.41 $X2=1.625 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__NAND3B_4%A_744_74# 1 2 3 4 5 20 24 29 32
c35 32 0 1.71648e-19 $X=5.515 $Y=0.51
c36 29 0 1.40137e-19 $X=4.03 $Y=0.49
r37 31 32 6.52497 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0.51
+ $X2=5.515 $Y2=0.51
r38 27 29 6.95017 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=0.49
+ $X2=4.03 $Y2=0.49
r39 22 24 30.9719 $w=3.18e-07 $l=8.6e-07 $layer=LI1_cond $X=6.54 $Y=0.51 $X2=7.4
+ $Y2=0.51
r40 20 31 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=5.835 $Y=0.51
+ $X2=5.68 $Y2=0.51
r41 20 22 25.3898 $w=3.18e-07 $l=7.05e-07 $layer=LI1_cond $X=5.835 $Y=0.51
+ $X2=6.54 $Y2=0.51
r42 19 32 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=4.75 $Y=0.475
+ $X2=5.515 $Y2=0.475
r43 19 29 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.75 $Y=0.475
+ $X2=4.03 $Y2=0.475
r44 5 24 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=7.26 $Y=0.37
+ $X2=7.4 $Y2=0.55
r45 4 22 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.4 $Y=0.37
+ $X2=6.54 $Y2=0.55
r46 3 31 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.37 $X2=5.68 $Y2=0.55
r47 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.61
+ $Y=0.37 $X2=4.75 $Y2=0.515
r48 1 27 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.37 $X2=3.865 $Y2=0.53
.ends


* File: sky130_fd_sc_ms__nand3_2.spice
* Created: Fri Aug 28 17:43:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand3_2.pex.spice"
.subckt sky130_fd_sc_ms__nand3_2  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1000 N_A_27_74#_M1000_d N_C_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.1036 PD=2.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_C_M1010_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1007 N_A_283_74#_M1007_d N_B_M1007_g N_A_27_74#_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.176975 AS=0.1036 PD=1.375 PS=1.02 NRD=29.856 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 N_A_283_74#_M1007_d N_A_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.176975 AS=0.1036 PD=1.375 PS=1.02 NRD=29.856 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_283_74#_M1011_d N_A_M1011_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.179175 AS=0.1036 PD=1.375 PS=1.02 NRD=30.336 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1009 N_A_283_74#_M1011_d N_B_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.179175 AS=0.1998 PD=1.375 PS=2.02 NRD=30.336 NRS=0 M=1 R=4.93333
+ SA=75002.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90002.5
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1004_d N_C_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6 SB=90002.1
+ A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.154
+ AS=0.1792 PD=1.395 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90001.6
+ A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1003_d VPB PSHORT L=0.18 W=1.12 AD=0.1764
+ AS=0.154 PD=1.435 PS=1.395 NRD=7.0329 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1001_d N_A_M1006_g N_Y_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.1764
+ AS=0.1512 PD=1.435 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1006_s N_B_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__nand3_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__edfxtp_1.pex.spice
* Created: Wed Sep  2 12:08:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%D 3 7 11 12 17 18 20 22
c43 18 0 6.13878e-20 $X=0.52 $Y=1.145
c44 3 0 1.15294e-19 $X=0.495 $Y=2.75
r45 20 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.825
+ $X2=0.52 $Y2=1.99
r46 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.825 $X2=0.52 $Y2=1.825
r47 17 20 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.52 $Y=1.145
+ $X2=0.52 $Y2=1.825
r48 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.145 $X2=0.52 $Y2=1.145
r49 12 21 4.85239 $w=3.78e-07 $l=1.6e-07 $layer=LI1_cond $X=0.615 $Y=1.665
+ $X2=0.615 $Y2=1.825
r50 11 12 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.665
r51 11 18 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.145
r52 10 17 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.98
+ $X2=0.52 $Y2=1.145
r53 7 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.58 $Y=0.58 $X2=0.58
+ $Y2=0.98
r54 3 22 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=2.75
+ $X2=0.495 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_159_446# 1 2 9 12 15 19 22 26 27 28 29 30
+ 31 34 38 40 42 44 53
c124 53 0 1.98585e-19 $X=2.38 $Y=1.55
c125 44 0 1.9156e-19 $X=2.22 $Y=1.55
c126 42 0 1.34182e-19 $X=1.79 $Y=1.695
c127 31 0 1.15294e-19 $X=1.305 $Y=1.695
c128 28 0 1.9799e-19 $X=1.57 $Y=0.855
c129 19 0 6.13878e-20 $X=1.05 $Y=2.305
r130 45 53 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.22 $Y=1.55
+ $X2=2.38 $Y2=1.55
r131 44 47 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.22 $Y=1.55
+ $X2=2.22 $Y2=1.695
r132 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.55 $X2=2.22 $Y2=1.55
r133 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=1.695
+ $X2=1.79 $Y2=1.695
r134 40 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=1.695
+ $X2=2.22 $Y2=1.695
r135 40 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.055 $Y=1.695
+ $X2=1.875 $Y2=1.695
r136 36 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=1.78
+ $X2=1.79 $Y2=1.695
r137 36 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.79 $Y=1.78
+ $X2=1.79 $Y2=2.495
r138 32 34 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.695 $Y=0.77
+ $X2=1.695 $Y2=0.645
r139 30 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.695
+ $X2=1.79 $Y2=1.695
r140 30 31 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.705 $Y=1.695
+ $X2=1.305 $Y2=1.695
r141 28 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.57 $Y=0.855
+ $X2=1.695 $Y2=0.77
r142 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.57 $Y=0.855
+ $X2=1.305 $Y2=0.855
r143 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.505 $X2=1.14 $Y2=1.505
r144 24 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.61
+ $X2=1.305 $Y2=1.695
r145 24 26 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.14 $Y=1.61
+ $X2=1.14 $Y2=1.505
r146 23 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=0.94
+ $X2=1.305 $Y2=0.855
r147 23 26 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=1.14 $Y=0.94
+ $X2=1.14 $Y2=1.505
r148 21 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.14 $Y=1.845
+ $X2=1.14 $Y2=1.505
r149 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.845
+ $X2=1.14 $Y2=2.01
r150 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.385
+ $X2=2.38 $Y2=1.55
r151 13 15 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.38 $Y=1.385
+ $X2=2.38 $Y2=0.645
r152 12 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.05 $Y=2.23
+ $X2=1.05 $Y2=2.305
r153 12 22 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.05 $Y=2.23
+ $X2=1.05 $Y2=2.01
r154 7 19 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.885 $Y=2.305
+ $X2=1.05 $Y2=2.305
r155 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=0.885 $Y=2.38
+ $X2=0.885 $Y2=2.75
r156 2 38 600 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=2.18 $X2=1.79 $Y2=2.495
r157 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.435 $X2=1.735 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%DE 3 5 6 10 11 13 14 16 17 18 19 21 22 26
+ 29 31
c88 31 0 3.25741e-19 $X=1.68 $Y=1.44
c89 26 0 1.98585e-19 $X=1.68 $Y=1.295
c90 10 0 3.01092e-20 $X=1.74 $Y=1.955
r91 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.275
+ $X2=1.68 $Y2=1.44
r92 26 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.275 $X2=1.68 $Y2=1.275
r93 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.695 $Y=2.105
+ $X2=2.695 $Y2=2.39
r94 17 19 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.605 $Y=2.03
+ $X2=2.695 $Y2=2.105
r95 17 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.605 $Y=2.03
+ $X2=2.105 $Y2=2.03
r96 14 18 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.015 $Y=2.03
+ $X2=2.105 $Y2=2.03
r97 14 23 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.015 $Y=2.03
+ $X2=1.74 $Y2=2.03
r98 14 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.015 $Y=2.105
+ $X2=2.015 $Y2=2.5
r99 11 22 13.5877 $w=2.4e-07 $l=2.14243e-07 $layer=POLY_cond $X=1.95 $Y=0.95
+ $X2=1.77 $Y2=1.025
r100 11 13 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.95 $Y=0.95
+ $X2=1.95 $Y2=0.645
r101 10 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.74 $Y=1.955
+ $X2=1.74 $Y2=2.03
r102 10 31 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.74 $Y=1.955
+ $X2=1.74 $Y2=1.44
r103 7 22 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.68 $Y=1.1
+ $X2=1.77 $Y2=1.025
r104 7 29 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.68 $Y=1.1
+ $X2=1.68 $Y2=1.275
r105 5 22 12.1617 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.515 $Y=1.025
+ $X2=1.77 $Y2=1.025
r106 5 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.515 $Y=1.025 $X2=1.045
+ $Y2=1.025
r107 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.97 $Y=0.95
+ $X2=1.045 $Y2=1.025
r108 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.97 $Y=0.95 $X2=0.97
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_533_61# 1 2 9 13 15 17 18 19 22 26 29 33
+ 36 40 43 44 45 51 52 55 56 60 67
c197 44 0 2.65373e-20 $X=11.615 $Y=1.665
r198 55 58 76.7264 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=2.92 $Y=1.21
+ $X2=2.92 $Y2=1.715
r199 55 57 46.8261 $w=5.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.21
+ $X2=2.92 $Y2=1.045
r200 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.83
+ $Y=1.21 $X2=2.83 $Y2=1.21
r201 52 67 6.51792 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=11.765 $Y=1.665
+ $X2=11.765 $Y2=1.55
r202 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=1.665
+ $X2=11.76 $Y2=1.665
r203 48 56 13.983 $w=3.73e-07 $l=4.55e-07 $layer=LI1_cond $X=2.742 $Y=1.665
+ $X2=2.742 $Y2=1.21
r204 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r205 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r206 44 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=11.76 $Y2=1.665
r207 44 45 10.9282 $w=1.4e-07 $l=8.83e-06 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=2.785 $Y2=1.665
r208 42 67 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.76 $Y=0.81
+ $X2=11.76 $Y2=1.55
r209 40 42 10.9338 $w=3.53e-07 $l=2.4e-07 $layer=LI1_cond $X=11.667 $Y=0.57
+ $X2=11.667 $Y2=0.81
r210 36 43 4.2255 $w=2.85e-07 $l=1.32605e-07 $layer=LI1_cond $X=11.765 $Y=2.095
+ $X2=11.72 $Y2=2.207
r211 35 52 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=11.765 $Y=1.67
+ $X2=11.765 $Y2=1.665
r212 35 36 20.4078 $w=2.38e-07 $l=4.25e-07 $layer=LI1_cond $X=11.765 $Y=1.67
+ $X2=11.765 $Y2=2.095
r213 31 43 4.2255 $w=2.85e-07 $l=1.13e-07 $layer=LI1_cond $X=11.72 $Y=2.32
+ $X2=11.72 $Y2=2.207
r214 31 33 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.72 $Y=2.32
+ $X2=11.72 $Y2=2.435
r215 29 61 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.83 $Y=2.185
+ $X2=10.83 $Y2=2.35
r216 29 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.83 $Y=2.185
+ $X2=10.83 $Y2=2.02
r217 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.83
+ $Y=2.185 $X2=10.83 $Y2=2.185
r218 26 43 2.20607 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=11.555 $Y=2.207
+ $X2=11.72 $Y2=2.207
r219 26 28 37.1343 $w=2.23e-07 $l=7.25e-07 $layer=LI1_cond $X=11.555 $Y=2.207
+ $X2=10.83 $Y2=2.207
r220 24 60 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=10.89 $Y=1.015
+ $X2=10.89 $Y2=2.02
r221 22 61 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=10.785 $Y=2.72
+ $X2=10.785 $Y2=2.35
r222 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.815 $Y=0.94
+ $X2=10.89 $Y2=1.015
r223 18 19 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.815 $Y=0.94
+ $X2=10.375 $Y2=0.94
r224 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.3 $Y=0.865
+ $X2=10.375 $Y2=0.94
r225 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.3 $Y=0.865
+ $X2=10.3 $Y2=0.58
r226 13 58 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.085 $Y=2.39
+ $X2=3.085 $Y2=1.715
r227 9 57 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.74 $Y=0.645 $X2=2.74
+ $Y2=1.045
r228 2 33 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.585
+ $Y=2.29 $X2=11.72 $Y2=2.435
r229 1 40 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=11.48
+ $Y=0.37 $X2=11.62 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%CLK 3 4 8 10 13 15
c40 13 0 1.4577e-19 $X=3.615 $Y=1.385
r41 13 16 14.2284 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=3.632 $Y=1.385
+ $X2=3.632 $Y2=1.475
r42 13 15 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.632 $Y=1.385
+ $X2=3.632 $Y2=1.22
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.385 $X2=3.615 $Y2=1.385
r44 10 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.615 $Y=1.295
+ $X2=3.615 $Y2=1.385
r45 6 8 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.06 $Y=1.55 $X2=4.06
+ $Y2=2.32
r46 5 16 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.815 $Y=1.475
+ $X2=3.632 $Y2=1.475
r47 4 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.97 $Y=1.475
+ $X2=4.06 $Y2=1.55
r48 4 5 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=3.97 $Y=1.475
+ $X2=3.815 $Y2=1.475
r49 3 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.74 $Y=0.74 $X2=3.74
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_958_74# 1 2 9 11 13 16 19 23 25 26 27 32
+ 33 36 37 40 41 42 44 45 46 47 49 50 53 56 59 61 64 65 69 76
c217 69 0 2.65373e-20 $X=10.44 $Y=1.42
c218 56 0 2.80716e-20 $X=6.67 $Y=1.145
c219 53 0 1.61107e-19 $X=6.085 $Y=2.135
c220 40 0 1.62788e-19 $X=7.675 $Y=0.935
c221 11 0 1.96074e-19 $X=6.67 $Y=0.98
r222 69 80 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.44 $Y=1.42
+ $X2=10.44 $Y2=1.585
r223 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.44
+ $Y=1.42 $X2=10.44 $Y2=1.42
r224 65 68 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.44 $Y=1.29
+ $X2=10.44 $Y2=1.42
r225 64 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.36 $Y=1.385
+ $X2=9.36 $Y2=1.22
r226 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.36
+ $Y=1.385 $X2=9.36 $Y2=1.385
r227 61 63 4.29259 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.285 $Y=1.29
+ $X2=9.285 $Y2=1.385
r228 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.67
+ $Y=1.145 $X2=6.67 $Y2=1.145
r229 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=2.135 $X2=6.085 $Y2=2.135
r230 50 52 5.47436 $w=3.9e-07 $l=1.75e-07 $layer=LI1_cond $X=5.91 $Y=2.06
+ $X2=6.085 $Y2=2.06
r231 48 61 3.44395 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.46 $Y=1.29
+ $X2=9.285 $Y2=1.29
r232 47 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.275 $Y=1.29
+ $X2=10.44 $Y2=1.29
r233 47 48 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=10.275 $Y=1.29
+ $X2=9.46 $Y2=1.29
r234 45 61 12.2 $w=2.7e-07 $l=3.46627e-07 $layer=LI1_cond $X=9.11 $Y=1.02
+ $X2=9.285 $Y2=1.29
r235 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.11 $Y=1.02
+ $X2=8.44 $Y2=1.02
r236 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.355 $Y=0.935
+ $X2=8.44 $Y2=1.02
r237 43 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.355 $Y=0.425
+ $X2=8.355 $Y2=0.935
r238 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.27 $Y=0.34
+ $X2=8.355 $Y2=0.425
r239 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.27 $Y=0.34
+ $X2=7.76 $Y2=0.34
r240 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.675 $Y=0.425
+ $X2=7.76 $Y2=0.34
r241 39 40 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.675 $Y=0.425
+ $X2=7.675 $Y2=0.935
r242 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=1.02
+ $X2=7.675 $Y2=0.935
r243 37 59 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.59 $Y=1.02
+ $X2=6.96 $Y2=1.02
r244 36 59 6.09592 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=1.122
+ $X2=6.96 $Y2=1.122
r245 36 55 6.30002 $w=3.73e-07 $l=2.05e-07 $layer=LI1_cond $X=6.875 $Y=1.122
+ $X2=6.67 $Y2=1.122
r246 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.875 $Y=0.425
+ $X2=6.875 $Y2=0.935
r247 34 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=0.34
+ $X2=5.91 $Y2=0.34
r248 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.79 $Y=0.34
+ $X2=6.875 $Y2=0.425
r249 33 34 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.79 $Y=0.34
+ $X2=5.995 $Y2=0.34
r250 32 50 5.6248 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.91 $Y=1.82 $X2=5.91
+ $Y2=2.06
r251 31 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=0.425
+ $X2=5.91 $Y2=0.34
r252 31 32 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.91 $Y=0.425
+ $X2=5.91 $Y2=1.82
r253 27 50 3.08808 $w=3.9e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.825 $Y=1.98
+ $X2=5.91 $Y2=2.06
r254 27 29 6.84263 $w=3.18e-07 $l=1.9e-07 $layer=LI1_cond $X=5.825 $Y=1.98
+ $X2=5.635 $Y2=1.98
r255 25 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.825 $Y=0.34
+ $X2=5.91 $Y2=0.34
r256 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.825 $Y=0.34
+ $X2=5.095 $Y2=0.34
r257 21 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.93 $Y=0.425
+ $X2=5.095 $Y2=0.34
r258 21 23 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.93 $Y=0.425
+ $X2=4.93 $Y2=0.515
r259 19 80 441.185 $w=1.8e-07 $l=1.135e-06 $layer=POLY_cond $X=10.365 $Y=2.72
+ $X2=10.365 $Y2=1.585
r260 16 76 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.4 $Y=0.74 $X2=9.4
+ $Y2=1.22
r261 11 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=0.98
+ $X2=6.67 $Y2=1.145
r262 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.67 $Y=0.98
+ $X2=6.67 $Y2=0.66
r263 7 53 56.2646 $w=2.57e-07 $l=3.73497e-07 $layer=POLY_cond $X=6.385 $Y=2.3
+ $X2=6.085 $Y2=2.135
r264 7 9 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=6.385 $Y=2.3
+ $X2=6.385 $Y2=2.75
r265 2 29 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.84 $X2=5.635 $Y2=2.02
r266 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.79
+ $Y=0.37 $X2=4.93 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_763_74# 1 2 11 13 15 17 20 22 23 28 32 36
+ 42 45 46 50 51 53 56 57 59 60 65 66 70 72
c184 59 0 1.61107e-19 $X=6.875 $Y=2.165
c185 51 0 5.61815e-20 $X=4.735 $Y=1.635
r186 66 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.9 $Y=1.635
+ $X2=9.9 $Y2=1.8
r187 66 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.9 $Y=1.635
+ $X2=9.9 $Y2=1.47
r188 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.9
+ $Y=1.635 $X2=9.9 $Y2=1.635
r189 62 65 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=9.715 $Y=1.635
+ $X2=9.9 $Y2=1.635
r190 60 73 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=6.862 $Y=2.165
+ $X2=6.862 $Y2=2.33
r191 60 72 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=6.862 $Y=2.165
+ $X2=6.862 $Y2=2
r192 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.875
+ $Y=2.165 $X2=6.875 $Y2=2.165
r193 55 62 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.715 $Y=1.725
+ $X2=9.715 $Y2=1.635
r194 55 56 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=9.715 $Y=1.725
+ $X2=9.715 $Y2=2.41
r195 54 59 14.482 $w=2.78e-07 $l=4.10244e-07 $layer=LI1_cond $X=7.115 $Y=2.495
+ $X2=6.935 $Y2=2.165
r196 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.63 $Y=2.495
+ $X2=9.715 $Y2=2.41
r197 53 54 164.08 $w=1.68e-07 $l=2.515e-06 $layer=LI1_cond $X=9.63 $Y=2.495
+ $X2=7.115 $Y2=2.495
r198 51 70 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.735 $Y=1.635
+ $X2=4.735 $Y2=1.655
r199 51 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.635
+ $X2=4.735 $Y2=1.47
r200 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.735
+ $Y=1.635 $X2=4.735 $Y2=1.635
r201 48 50 8.03336 $w=6.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.285 $Y=1.805
+ $X2=4.735 $Y2=1.805
r202 46 48 2.94557 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=1.805
+ $X2=4.285 $Y2=1.805
r203 45 46 10.5816 $w=6.7e-07 $l=3.751e-07 $layer=LI1_cond $X=4.035 $Y=1.47
+ $X2=4.12 $Y2=1.805
r204 45 57 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.035 $Y=1.47
+ $X2=4.035 $Y2=1.01
r205 40 57 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0.845
+ $X2=3.955 $Y2=1.01
r206 40 42 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.955 $Y=0.845
+ $X2=3.955 $Y2=0.515
r207 36 75 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=9.91 $Y=0.58
+ $X2=9.91 $Y2=1.47
r208 32 76 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=9.83 $Y=2.46
+ $X2=9.83 $Y2=1.8
r209 28 73 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=6.835 $Y=2.75
+ $X2=6.835 $Y2=2.33
r210 24 72 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.76 $Y=1.73
+ $X2=6.76 $Y2=2
r211 23 39 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.78 $Y=1.655
+ $X2=5.705 $Y2=1.655
r212 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.685 $Y=1.655
+ $X2=6.76 $Y2=1.73
r213 22 23 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=6.685 $Y=1.655
+ $X2=5.78 $Y2=1.655
r214 18 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.705 $Y=1.58
+ $X2=5.705 $Y2=1.655
r215 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=5.705 $Y=1.58
+ $X2=5.705 $Y2=0.66
r216 15 39 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.41 $Y=1.655
+ $X2=5.705 $Y2=1.655
r217 15 17 179.411 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=5.41 $Y=1.73
+ $X2=5.41 $Y2=2.4
r218 14 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.655
+ $X2=4.735 $Y2=1.655
r219 13 15 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.32 $Y=1.655
+ $X2=5.41 $Y2=1.655
r220 13 14 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.32 $Y=1.655
+ $X2=4.9 $Y2=1.655
r221 11 69 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=4.715 $Y=0.74
+ $X2=4.715 $Y2=1.47
r222 2 48 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=4.15
+ $Y=1.76 $X2=4.285 $Y2=1.94
r223 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.815
+ $Y=0.37 $X2=3.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_1409_64# 1 2 9 13 17 21 23 24 25 29 31 36
+ 37 39 46 54
c102 46 0 2.74064e-19 $X=7.46 $Y=1.367
c103 13 0 1.96559e-19 $X=7.34 $Y=2.75
r104 47 48 18.6009 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=8.015 $Y=1.44
+ $X2=8.355 $Y2=1.44
r105 44 54 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=7.295 $Y=1.365
+ $X2=7.34 $Y2=1.365
r106 44 51 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.295 $Y=1.365
+ $X2=7.12 $Y2=1.365
r107 43 46 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=1.367
+ $X2=7.46 $Y2=1.367
r108 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.295
+ $Y=1.365 $X2=7.295 $Y2=1.365
r109 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.775
+ $Y=1.44 $X2=8.775 $Y2=1.44
r110 37 48 4.43115 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=1.44
+ $X2=8.355 $Y2=1.44
r111 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.44 $Y=1.44
+ $X2=8.775 $Y2=1.44
r112 35 48 2.32876 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.355 $Y=1.605
+ $X2=8.355 $Y2=1.44
r113 35 36 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.355 $Y=1.605
+ $X2=8.355 $Y2=2.07
r114 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.27 $Y=2.155
+ $X2=8.355 $Y2=2.07
r115 31 33 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.27 $Y=2.155
+ $X2=8.11 $Y2=2.155
r116 27 47 2.32876 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=1.275
+ $X2=8.015 $Y2=1.44
r117 27 29 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.015 $Y=1.275
+ $X2=8.015 $Y2=0.85
r118 25 47 5.36928 $w=2.23e-07 $l=1.18427e-07 $layer=LI1_cond $X=7.93 $Y=1.36
+ $X2=8.015 $Y2=1.44
r119 25 46 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=7.93 $Y=1.36
+ $X2=7.46 $Y2=1.36
r120 23 40 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.805 $Y=1.44
+ $X2=8.775 $Y2=1.44
r121 23 24 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.805 $Y=1.44
+ $X2=8.895 $Y2=1.44
r122 19 24 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=8.91 $Y=1.275
+ $X2=8.895 $Y2=1.44
r123 19 21 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=8.91 $Y=1.275
+ $X2=8.91 $Y2=0.74
r124 15 24 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.895 $Y=1.605
+ $X2=8.895 $Y2=1.44
r125 15 17 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=8.895 $Y=1.605
+ $X2=8.895 $Y2=2.46
r126 11 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.34 $Y=1.53
+ $X2=7.34 $Y2=1.365
r127 11 13 474.226 $w=1.8e-07 $l=1.22e-06 $layer=POLY_cond $X=7.34 $Y=1.53
+ $X2=7.34 $Y2=2.75
r128 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.12 $Y=1.2
+ $X2=7.12 $Y2=1.365
r129 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.12 $Y=1.2 $X2=7.12
+ $Y2=0.66
r130 2 33 600 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=7.975
+ $Y=2.025 $X2=8.11 $Y2=2.155
r131 1 29 182 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_NDIFF $count=1 $X=7.875
+ $Y=0.45 $X2=8.015 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_1156_90# 1 2 9 13 16 17 23 28 29 32 33 34
c97 9 0 2.85555e-19 $X=7.8 $Y=0.77
r98 33 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.865 $Y=1.7
+ $X2=7.865 $Y2=1.865
r99 33 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.865 $Y=1.7
+ $X2=7.865 $Y2=1.535
r100 32 34 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=7.865 $Y=1.722
+ $X2=7.7 $Y2=1.722
r101 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.865
+ $Y=1.7 $X2=7.865 $Y2=1.7
r102 28 29 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=6.595 $Y=2.75
+ $X2=6.595 $Y2=2.52
r103 24 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=1.715
+ $X2=6.5 $Y2=1.715
r104 23 26 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=1.715
+ $X2=6.5 $Y2=1.715
r105 23 34 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=6.585 $Y=1.715
+ $X2=7.7 $Y2=1.715
r106 20 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=1.8 $X2=6.5
+ $Y2=1.715
r107 20 29 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.5 $Y=1.8 $X2=6.5
+ $Y2=2.52
r108 17 19 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=6.335 $Y=0.68
+ $X2=6.39 $Y2=0.68
r109 16 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.25 $Y=1.63
+ $X2=6.25 $Y2=1.715
r110 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.25 $Y=0.765
+ $X2=6.335 $Y2=0.68
r111 15 16 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.25 $Y=0.765
+ $X2=6.25 $Y2=1.63
r112 13 38 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.885 $Y=2.445
+ $X2=7.885 $Y2=1.865
r113 9 37 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=7.8 $Y=0.77 $X2=7.8
+ $Y2=1.535
r114 2 28 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=6.475
+ $Y=2.54 $X2=6.61 $Y2=2.75
r115 1 19 182 $w=1.7e-07 $l=7.15821e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.45 $X2=6.39 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_1895_74# 1 2 9 13 15 17 19 22 24 27 29 30
+ 33 37 38 40 43 44 47
c128 30 0 1.36277e-19 $X=9.78 $Y=0.92
r129 50 51 27.9638 $w=4.1e-07 $l=7.5e-08 $layer=POLY_cond $X=11.38 $Y=1.26
+ $X2=11.38 $Y2=1.335
r130 44 50 12.2083 $w=4.1e-07 $l=9e-08 $layer=POLY_cond $X=11.38 $Y=1.17
+ $X2=11.38 $Y2=1.26
r131 44 49 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=11.38 $Y=1.17
+ $X2=11.38 $Y2=1.005
r132 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.34
+ $Y=1.17 $X2=11.34 $Y2=1.17
r133 41 47 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.945 $Y=1.17
+ $X2=10.86 $Y2=1.085
r134 41 43 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=10.945 $Y=1.17
+ $X2=11.34 $Y2=1.17
r135 39 47 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=10.86 $Y=1.335
+ $X2=10.86 $Y2=1.085
r136 39 40 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=1.335
+ $X2=10.86 $Y2=1.755
r137 38 46 16.9994 $w=2.36e-07 $l=3.49929e-07 $layer=LI1_cond $X=10.405 $Y=1.84
+ $X2=10.095 $Y2=1.925
r138 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.775 $Y=1.84
+ $X2=10.86 $Y2=1.755
r139 37 38 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.775 $Y=1.84
+ $X2=10.405 $Y2=1.84
r140 33 35 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=10.095 $Y=2.105
+ $X2=10.095 $Y2=2.835
r141 31 46 0.361987 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=10.095 $Y=2.095
+ $X2=10.095 $Y2=1.925
r142 31 33 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=10.095 $Y=2.095
+ $X2=10.095 $Y2=2.105
r143 29 47 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.775 $Y=0.92
+ $X2=10.86 $Y2=1.085
r144 29 30 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=10.775 $Y=0.92
+ $X2=9.78 $Y2=0.92
r145 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.615 $Y=0.835
+ $X2=9.78 $Y2=0.92
r146 25 27 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=9.615 $Y=0.835
+ $X2=9.615 $Y2=0.515
r147 20 24 18.8402 $w=1.65e-07 $l=8.7892e-08 $layer=POLY_cond $X=12.465 $Y=1.335
+ $X2=12.437 $Y2=1.26
r148 20 22 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=12.465 $Y=1.335
+ $X2=12.465 $Y2=2.4
r149 17 24 18.8402 $w=1.65e-07 $l=9.3675e-08 $layer=POLY_cond $X=12.395 $Y=1.185
+ $X2=12.437 $Y2=1.26
r150 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=12.395 $Y=1.185
+ $X2=12.395 $Y2=0.74
r151 16 50 26.4667 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=11.585 $Y=1.26
+ $X2=11.38 $Y2=1.26
r152 15 24 6.66866 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=12.32 $Y=1.26
+ $X2=12.437 $Y2=1.26
r153 15 16 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=12.32 $Y=1.26
+ $X2=11.585 $Y2=1.26
r154 13 51 495.605 $w=1.8e-07 $l=1.275e-06 $layer=POLY_cond $X=11.495 $Y=2.61
+ $X2=11.495 $Y2=1.335
r155 9 49 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=11.405 $Y=0.58
+ $X2=11.405 $Y2=1.005
r156 2 35 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=9.92
+ $Y=1.96 $X2=10.055 $Y2=2.835
r157 2 33 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.92
+ $Y=1.96 $X2=10.055 $Y2=2.105
r158 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.475
+ $Y=0.37 $X2=9.615 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%A_27_508# 1 2 3 4 5 6 20 23 25 28 29 30 32
+ 33 34 36 37 40 41 43 45 46 49 54 56 60 64
c172 64 0 1.4577e-19 $X=3.31 $Y=2.39
c173 43 0 5.61815e-20 $X=5.49 $Y=0.7
c174 34 0 3.01092e-20 $X=2.215 $Y=2.035
r175 64 65 0.189441 $w=3.22e-07 $l=5e-09 $layer=LI1_cond $X=3.287 $Y=2.39
+ $X2=3.287 $Y2=2.395
r176 58 60 5.98039 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=2.955 $Y=0.645
+ $X2=3.185 $Y2=0.645
r177 51 54 4.96245 $w=4.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.17 $Y=0.575
+ $X2=0.365 $Y2=0.575
r178 47 49 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=6.12 $Y=2.69 $X2=6.12
+ $Y2=2.75
r179 46 70 20.8849 $w=2.44e-07 $l=4.53211e-07 $layer=LI1_cond $X=5.61 $Y=2.605
+ $X2=5.215 $Y2=2.48
r180 45 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.995 $Y=2.605
+ $X2=6.12 $Y2=2.69
r181 45 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.995 $Y=2.605
+ $X2=5.61 $Y2=2.605
r182 41 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.49 $Y=1.565
+ $X2=5.215 $Y2=1.565
r183 41 43 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.49 $Y=1.48
+ $X2=5.49 $Y2=0.7
r184 40 70 2.85362 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.215 $Y=2.31
+ $X2=5.215 $Y2=2.48
r185 39 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=1.65
+ $X2=5.215 $Y2=1.565
r186 39 40 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.215 $Y=1.65
+ $X2=5.215 $Y2=2.31
r187 38 65 4.47834 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.475 $Y=2.395
+ $X2=3.287 $Y2=2.395
r188 37 70 5.3849 $w=2.44e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.13 $Y=2.395
+ $X2=5.215 $Y2=2.48
r189 37 38 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=5.13 $Y=2.395
+ $X2=3.475 $Y2=2.395
r190 35 60 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.185 $Y=0.875
+ $X2=3.185 $Y2=0.645
r191 35 36 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=3.185 $Y=0.875
+ $X2=3.185 $Y2=1.95
r192 33 64 13.4503 $w=3.22e-07 $l=4.38646e-07 $layer=LI1_cond $X=3.1 $Y=2.035
+ $X2=3.287 $Y2=2.39
r193 33 36 5.92483 $w=3.22e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.035
+ $X2=3.185 $Y2=1.95
r194 33 34 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.1 $Y=2.035
+ $X2=2.215 $Y2=2.035
r195 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=2.12
+ $X2=2.215 $Y2=2.035
r196 31 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.13 $Y=2.12
+ $X2=2.13 $Y2=2.905
r197 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.13 $Y2=2.905
r198 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.535 $Y2=2.99
r199 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=2.905
+ $X2=1.535 $Y2=2.99
r200 27 28 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.45 $Y=2.35
+ $X2=1.45 $Y2=2.905
r201 26 56 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.435 $Y=2.265
+ $X2=0.26 $Y2=2.265
r202 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.365 $Y=2.265
+ $X2=1.45 $Y2=2.35
r203 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.365 $Y=2.265
+ $X2=0.435 $Y2=2.265
r204 21 56 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.35
+ $X2=0.26 $Y2=2.265
r205 21 23 13.1708 $w=3.48e-07 $l=4e-07 $layer=LI1_cond $X=0.26 $Y=2.35 $X2=0.26
+ $Y2=2.75
r206 20 56 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.17 $Y=2.18
+ $X2=0.26 $Y2=2.265
r207 19 51 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=0.575
r208 19 20 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.18
r209 6 49 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=2.54 $X2=6.16 $Y2=2.75
r210 5 64 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=2.18 $X2=3.31 $Y2=2.39
r211 4 23 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
r212 3 43 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.45 $X2=5.49 $Y2=0.7
r213 2 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.435 $X2=2.955 $Y2=0.645
r214 1 54 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=0.22
+ $Y=0.37 $X2=0.365 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 53 55 60 61 63 64 66 67 69 70 71 89 93 102 109 115 118 121 125
r134 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r135 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r136 118 119 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r137 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r138 113 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r139 113 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r140 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r141 110 121 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=11.385 $Y=3.33
+ $X2=11.115 $Y2=3.33
r142 110 112 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=11.385 $Y=3.33
+ $X2=12.24 $Y2=3.33
r143 109 124 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=12.605 $Y=3.33
+ $X2=12.782 $Y2=3.33
r144 109 112 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.605 $Y=3.33
+ $X2=12.24 $Y2=3.33
r145 108 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r146 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r147 105 108 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r148 104 107 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r149 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r150 102 121 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=10.845 $Y=3.33
+ $X2=11.115 $Y2=3.33
r151 102 107 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=10.845 $Y=3.33
+ $X2=10.8 $Y2=3.33
r152 101 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r153 101 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 98 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.74 $Y=3.33
+ $X2=7.575 $Y2=3.33
r156 98 100 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.74 $Y=3.33
+ $X2=8.4 $Y2=3.33
r157 97 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r158 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r159 94 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.145 $Y2=3.33
r160 94 96 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.52 $Y2=3.33
r161 93 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=3.33
+ $X2=7.575 $Y2=3.33
r162 93 96 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=7.41 $Y=3.33
+ $X2=5.52 $Y2=3.33
r163 92 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r164 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r165 89 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=5.145 $Y2=3.33
r166 89 91 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=4.08 $Y2=3.33
r167 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r169 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r170 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r171 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r172 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r173 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r174 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r176 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r177 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r178 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 71 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r180 71 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r181 69 100 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.4 $Y2=3.33
r182 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.67 $Y2=3.33
r183 68 104 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.835 $Y=3.33
+ $X2=8.88 $Y2=3.33
r184 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.835 $Y=3.33
+ $X2=8.67 $Y2=3.33
r185 66 87 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=3.33 $X2=3.6
+ $Y2=3.33
r186 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.67 $Y=3.33
+ $X2=3.835 $Y2=3.33
r187 65 91 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4 $Y=3.33 $X2=4.08
+ $Y2=3.33
r188 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=3.33 $X2=3.835
+ $Y2=3.33
r189 63 81 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r190 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.51 $Y2=3.33
r191 62 84 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.51 $Y2=3.33
r193 60 74 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r194 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.07 $Y2=3.33
r195 59 78 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.2 $Y2=3.33
r196 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.07 $Y2=3.33
r197 55 58 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.73 $Y=1.985
+ $X2=12.73 $Y2=2.815
r198 53 124 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=12.73 $Y=3.245
+ $X2=12.782 $Y2=3.33
r199 53 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.73 $Y=3.245
+ $X2=12.73 $Y2=2.815
r200 49 121 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=11.115 $Y=3.245
+ $X2=11.115 $Y2=3.33
r201 49 51 12.293 $w=5.38e-07 $l=5.55e-07 $layer=LI1_cond $X=11.115 $Y=3.245
+ $X2=11.115 $Y2=2.69
r202 45 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.67 $Y=3.245
+ $X2=8.67 $Y2=3.33
r203 45 47 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.67 $Y=3.245
+ $X2=8.67 $Y2=2.835
r204 41 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=3.245
+ $X2=7.575 $Y2=3.33
r205 41 43 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.575 $Y=3.245
+ $X2=7.575 $Y2=2.835
r206 37 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=3.33
r207 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=2.815
r208 33 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=3.245
+ $X2=3.835 $Y2=3.33
r209 33 35 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.835 $Y=3.245
+ $X2=3.835 $Y2=2.735
r210 29 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=3.33
r211 29 31 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=2.455
r212 25 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r213 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.75
r214 8 58 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.555
+ $Y=1.84 $X2=12.69 $Y2=2.815
r215 8 55 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.555
+ $Y=1.84 $X2=12.69 $Y2=1.985
r216 7 51 600 $w=1.7e-07 $l=3.43402e-07 $layer=licon1_PDIFF $count=1 $X=10.875
+ $Y=2.51 $X2=11.14 $Y2=2.69
r217 6 47 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=1.96 $X2=8.67 $Y2=2.835
r218 5 43 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=7.43
+ $Y=2.54 $X2=7.575 $Y2=2.835
r219 4 39 600 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=5.06
+ $Y=1.84 $X2=5.185 $Y2=2.815
r220 3 35 600 $w=1.7e-07 $l=1.03797e-06 $layer=licon1_PDIFF $count=1 $X=3.705
+ $Y=1.76 $X2=3.835 $Y2=2.735
r221 2 31 600 $w=1.7e-07 $l=4.83322e-07 $layer=licon1_PDIFF $count=1 $X=2.105
+ $Y=2.18 $X2=2.47 $Y2=2.455
r222 1 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=2.54 $X2=1.11 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%Q 1 2 9 13 14 15 16 17 35 37
r28 23 37 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=12.24 $Y=1.715
+ $X2=12.24 $Y2=1.665
r29 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.24 $Y=2.405
+ $X2=12.24 $Y2=2.775
r30 15 16 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=12.24 $Y=1.985
+ $X2=12.24 $Y2=2.405
r31 14 37 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=12.24 $Y=1.647
+ $X2=12.24 $Y2=1.665
r32 14 35 3.8025 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=12.24 $Y=1.647
+ $X2=12.24 $Y2=1.55
r33 14 15 8.8354 $w=3.28e-07 $l=2.53e-07 $layer=LI1_cond $X=12.24 $Y=1.732
+ $X2=12.24 $Y2=1.985
r34 14 23 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=12.24 $Y=1.732
+ $X2=12.24 $Y2=1.715
r35 13 35 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=12.21 $Y=1.13
+ $X2=12.21 $Y2=1.55
r36 7 13 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.18 $Y=0.965
+ $X2=12.18 $Y2=1.13
r37 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=12.18 $Y=0.965
+ $X2=12.18 $Y2=0.515
r38 2 17 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=12.115
+ $Y=1.84 $X2=12.24 $Y2=2.815
r39 2 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=12.115
+ $Y=1.84 $X2=12.24 $Y2=1.985
r40 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.035
+ $Y=0.37 $X2=12.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXTP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 57 58 60 61 62 64 69 78 99 105 108 111 116 122 125
c148 43 0 1.96074e-19 $X=7.335 $Y=0.595
c149 1 0 1.9799e-19 $X=1.045 $Y=0.37
r150 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r151 120 122 8.97006 $w=7.48e-07 $l=3e-08 $layer=LI1_cond $X=11.28 $Y=0.29
+ $X2=11.31 $Y2=0.29
r152 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r153 118 120 1.43529 $w=7.48e-07 $l=9e-08 $layer=LI1_cond $X=11.19 $Y=0.29
+ $X2=11.28 $Y2=0.29
r154 115 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r155 114 118 6.21961 $w=7.48e-07 $l=3.9e-07 $layer=LI1_cond $X=10.8 $Y=0.29
+ $X2=11.19 $Y2=0.29
r156 114 116 15.6681 $w=7.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.8 $Y=0.29
+ $X2=10.35 $Y2=0.29
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r158 111 112 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r159 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r160 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r161 103 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r162 103 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.28 $Y2=0
r163 102 122 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=11.31 $Y2=0
r164 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r165 99 124 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.737 $Y2=0
r166 99 102 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.24 $Y2=0
r167 98 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r168 97 116 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=10.32 $Y=0 $X2=10.35
+ $Y2=0
r169 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r170 95 98 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r171 94 97 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r172 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r173 91 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r174 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r175 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r176 87 90 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r177 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r178 85 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r179 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r180 82 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=0
+ $X2=4.46 $Y2=0
r181 82 84 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=4.585 $Y=0
+ $X2=6.96 $Y2=0
r182 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r183 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r184 78 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.46 $Y2=0
r185 78 80 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.08 $Y2=0
r186 77 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r187 77 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.16 $Y2=0
r188 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r189 74 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0
+ $X2=2.165 $Y2=0
r190 74 76 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=3.12
+ $Y2=0
r191 73 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r192 73 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r193 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r194 70 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0
+ $X2=1.185 $Y2=0
r195 70 72 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.68
+ $Y2=0
r196 69 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.165
+ $Y2=0
r197 69 72 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.68
+ $Y2=0
r198 67 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r199 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r200 64 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0
+ $X2=1.185 $Y2=0
r201 64 66 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.72
+ $Y2=0
r202 62 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r203 62 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=4.56 $Y2=0
r204 60 90 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.4
+ $Y2=0
r205 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.735
+ $Y2=0
r206 59 94 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=8.86 $Y=0 $X2=8.88
+ $Y2=0
r207 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.86 $Y=0 $X2=8.735
+ $Y2=0
r208 57 84 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=6.96
+ $Y2=0
r209 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.295
+ $Y2=0
r210 56 87 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.44
+ $Y2=0
r211 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.295
+ $Y2=0
r212 54 76 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.12
+ $Y2=0
r213 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.525
+ $Y2=0
r214 53 80 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=4.08
+ $Y2=0
r215 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.525
+ $Y2=0
r216 49 124 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.737 $Y2=0
r217 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.68 $Y2=0.515
r218 45 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0
r219 45 47 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0.555
r220 41 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0
r221 41 43 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0.595
r222 37 111 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r223 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.515
r224 33 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0
r225 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.505
r226 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r227 29 31 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.645
r228 25 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r229 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.515
r230 8 51 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=12.47
+ $Y=0.37 $X2=12.68 $Y2=0.515
r231 7 118 91 $w=1.7e-07 $l=8.77596e-07 $layer=licon1_NDIFF $count=2 $X=10.375
+ $Y=0.37 $X2=11.19 $Y2=0.5
r232 6 47 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.55
+ $Y=0.37 $X2=8.695 $Y2=0.555
r233 5 43 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.45 $X2=7.335 $Y2=0.595
r234 4 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.36
+ $Y=0.37 $X2=4.5 $Y2=0.515
r235 3 35 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.37 $X2=3.525 $Y2=0.505
r236 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.435 $X2=2.165 $Y2=0.645
r237 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.515
.ends


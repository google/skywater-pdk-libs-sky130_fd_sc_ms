* File: sky130_fd_sc_ms__nor4bb_2.pex.spice
* Created: Fri Aug 28 17:50:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%C_N 3 7 9 10 17
r32 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.635 $X2=1.03 $Y2=1.635
r33 15 17 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=1.635
+ $X2=1.03 $Y2=1.635
r34 13 15 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=0.505 $Y=1.635
+ $X2=0.865 $Y2=1.635
r35 10 18 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.635
+ $X2=1.03 $Y2=1.635
r36 9 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.72 $Y=1.635 $X2=1.03
+ $Y2=1.635
r37 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=1.47
+ $X2=0.865 $Y2=1.635
r38 5 7 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.865 $Y=1.47
+ $X2=0.865 $Y2=0.69
r39 1 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.8
+ $X2=0.505 $Y2=1.635
r40 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.8 $X2=0.505
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%D_N 1 3 6 8 15
r35 13 15 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.635
+ $X2=1.825 $Y2=1.635
r36 10 13 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.48 $Y=1.635
+ $X2=1.66 $Y2=1.635
r37 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.635 $X2=1.66 $Y2=1.635
r38 4 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.8
+ $X2=1.825 $Y2=1.635
r39 4 6 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.825 $Y=1.8 $X2=1.825
+ $Y2=2.46
r40 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=1.47
+ $X2=1.48 $Y2=1.635
r41 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.48 $Y=1.47 $X2=1.48
+ $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%A_311_124# 1 2 9 13 17 21 23 29 35 39 40 47
+ 53
c73 17 0 1.04248e-19 $X=3.27 $Y=0.74
r74 53 54 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=3.27 $Y=1.515
+ $X2=3.285 $Y2=1.515
r75 50 51 0.748447 $w=3.22e-07 $l=5e-09 $layer=POLY_cond $X=2.835 $Y=1.515
+ $X2=2.84 $Y2=1.515
r76 47 50 13.1455 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.745 $Y=1.515
+ $X2=2.835 $Y2=1.515
r77 46 47 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=2.32 $Y=1.515
+ $X2=2.745 $Y2=1.515
r78 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.515 $X2=2.32 $Y2=1.515
r79 39 41 0.877092 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=2.105 $Y=2.135
+ $X2=2.105 $Y2=2.14
r80 39 40 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.135
+ $X2=2.105 $Y2=1.97
r81 36 53 40.4161 $w=3.22e-07 $l=2.7e-07 $layer=POLY_cond $X=3 $Y=1.515 $X2=3.27
+ $Y2=1.515
r82 36 51 23.9503 $w=3.22e-07 $l=1.6e-07 $layer=POLY_cond $X=3 $Y=1.515 $X2=2.84
+ $Y2=1.515
r83 35 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3 $Y=1.515
+ $X2=2.325 $Y2=1.515
r84 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.515 $X2=3 $Y2=1.515
r85 31 45 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.68
+ $X2=2.24 $Y2=1.515
r86 31 40 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.24 $Y=1.68
+ $X2=2.24 $Y2=1.97
r87 29 41 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.05 $Y=2.815
+ $X2=2.05 $Y2=2.14
r88 23 45 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.24 $Y=1.175
+ $X2=2.24 $Y2=1.515
r89 23 25 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.155 $Y=1.175
+ $X2=1.79 $Y2=1.175
r90 19 54 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.68
+ $X2=3.285 $Y2=1.515
r91 19 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.285 $Y=1.68
+ $X2=3.285 $Y2=2.4
r92 15 53 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.35
+ $X2=3.27 $Y2=1.515
r93 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.27 $Y=1.35
+ $X2=3.27 $Y2=0.74
r94 11 51 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.35
+ $X2=2.84 $Y2=1.515
r95 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.84 $Y=1.35
+ $X2=2.84 $Y2=0.74
r96 7 50 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.68
+ $X2=2.835 $Y2=1.515
r97 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.835 $Y=1.68
+ $X2=2.835 $Y2=2.4
r98 2 39 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.96 $X2=2.05 $Y2=2.135
r99 2 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.96 $X2=2.05 $Y2=2.815
r100 1 25 182 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.62 $X2=1.79 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%A_27_392# 1 2 9 13 17 21 27 29 31 32 35 38
+ 39 41 45 46 47 52 54 59
c135 21 0 3.67831e-20 $X=4.335 $Y=0.74
c136 17 0 1.11683e-19 $X=4.285 $Y=2.4
r137 59 60 7.48447 $w=3.22e-07 $l=5e-08 $layer=POLY_cond $X=4.285 $Y=1.515
+ $X2=4.335 $Y2=1.515
r138 58 59 56.882 $w=3.22e-07 $l=3.8e-07 $layer=POLY_cond $X=3.905 $Y=1.515
+ $X2=4.285 $Y2=1.515
r139 57 58 17.9627 $w=3.22e-07 $l=1.2e-07 $layer=POLY_cond $X=3.785 $Y=1.515
+ $X2=3.905 $Y2=1.515
r140 53 57 0.748447 $w=3.22e-07 $l=5e-09 $layer=POLY_cond $X=3.78 $Y=1.515
+ $X2=3.785 $Y2=1.515
r141 52 54 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.78 $Y=1.515
+ $X2=3.78 $Y2=1.35
r142 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.515 $X2=3.78 $Y2=1.515
r143 47 49 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.58 $Y=0.795
+ $X2=2.58 $Y2=1.095
r144 43 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.7 $Y=1.18 $X2=3.7
+ $Y2=1.35
r145 42 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=1.095
+ $X2=2.58 $Y2=1.095
r146 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=1.095
+ $X2=3.7 $Y2=1.18
r147 41 42 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.615 $Y=1.095
+ $X2=2.665 $Y2=1.095
r148 40 46 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0.795
+ $X2=0.65 $Y2=0.795
r149 39 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.795
+ $X2=2.58 $Y2=0.795
r150 39 40 109.604 $w=1.68e-07 $l=1.68e-06 $layer=LI1_cond $X=2.495 $Y=0.795
+ $X2=0.815 $Y2=0.795
r151 37 46 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.88
+ $X2=0.65 $Y2=0.795
r152 37 38 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.65 $Y=0.88
+ $X2=0.65 $Y2=1.13
r153 33 46 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.71
+ $X2=0.65 $Y2=0.795
r154 33 35 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.65 $Y=0.71
+ $X2=0.65 $Y2=0.525
r155 31 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.485 $Y=1.215
+ $X2=0.65 $Y2=1.13
r156 31 32 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.485 $Y=1.215
+ $X2=0.285 $Y2=1.215
r157 27 45 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=1.97
r158 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=2.815
r159 23 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.3
+ $X2=0.285 $Y2=1.215
r160 23 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.2 $Y=1.3 $X2=0.2
+ $Y2=1.97
r161 19 60 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.35
+ $X2=4.335 $Y2=1.515
r162 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.335 $Y=1.35
+ $X2=4.335 $Y2=0.74
r163 15 59 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.68
+ $X2=4.285 $Y2=1.515
r164 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.285 $Y=1.68
+ $X2=4.285 $Y2=2.4
r165 11 58 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=1.35
+ $X2=3.905 $Y2=1.515
r166 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.905 $Y=1.35
+ $X2=3.905 $Y2=0.74
r167 7 57 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.68
+ $X2=3.785 $Y2=1.515
r168 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.785 $Y=1.68
+ $X2=3.785 $Y2=2.4
r169 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r170 2 27 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.135
r171 1 35 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.505
+ $Y=0.37 $X2=0.65 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%B 3 7 11 13 15 21 22 30 34
c57 13 0 1.98445e-19 $X=5.745 $Y=1.77
c58 3 0 1.75889e-19 $X=4.835 $Y=0.74
r59 30 32 15.1075 $w=3.35e-07 $l=1.05e-07 $layer=POLY_cond $X=5.64 $Y=1.56
+ $X2=5.745 $Y2=1.56
r60 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.515 $X2=5.64 $Y2=1.515
r61 22 31 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.64
+ $Y2=1.565
r62 21 31 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.64 $Y2=1.565
r63 21 34 4.39439 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.405 $Y2=1.565
r64 19 27 34.5313 $w=3.35e-07 $l=2.4e-07 $layer=POLY_cond $X=5.025 $Y=1.56
+ $X2=5.265 $Y2=1.56
r65 19 25 27.3373 $w=3.35e-07 $l=1.9e-07 $layer=POLY_cond $X=5.025 $Y=1.56
+ $X2=4.835 $Y2=1.56
r66 18 34 15.3659 $w=2.83e-07 $l=3.8e-07 $layer=LI1_cond $X=5.025 $Y=1.492
+ $X2=5.405 $Y2=1.492
r67 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.025
+ $Y=1.515 $X2=5.025 $Y2=1.515
r68 13 32 17.2825 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.745 $Y=1.77
+ $X2=5.745 $Y2=1.56
r69 13 15 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=5.745 $Y=1.77
+ $X2=5.745 $Y2=2.4
r70 9 30 49.6388 $w=3.35e-07 $l=3.45e-07 $layer=POLY_cond $X=5.295 $Y=1.56
+ $X2=5.64 $Y2=1.56
r71 9 27 4.31642 $w=3.35e-07 $l=3e-08 $layer=POLY_cond $X=5.295 $Y=1.56
+ $X2=5.265 $Y2=1.56
r72 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.295 $Y=1.68
+ $X2=5.295 $Y2=2.4
r73 5 27 21.5811 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=1.56
r74 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=0.74
r75 1 25 21.5811 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.835 $Y=1.35
+ $X2=4.835 $Y2=1.56
r76 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.835 $Y=1.35
+ $X2=4.835 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%A 3 7 11 15 17 18 27
r47 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.815
+ $Y=1.515 $X2=6.815 $Y2=1.515
r48 25 27 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.705 $Y=1.515
+ $X2=6.815 $Y2=1.515
r49 24 25 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.695 $Y=1.515
+ $X2=6.705 $Y2=1.515
r50 23 24 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=6.245 $Y=1.515
+ $X2=6.695 $Y2=1.515
r51 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.23 $Y=1.515
+ $X2=6.245 $Y2=1.515
r52 18 28 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.815 $Y2=1.565
r53 17 28 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.815 $Y2=1.565
r54 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.705 $Y=1.35
+ $X2=6.705 $Y2=1.515
r55 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.705 $Y=1.35
+ $X2=6.705 $Y2=0.74
r56 9 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.68
+ $X2=6.695 $Y2=1.515
r57 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.695 $Y=1.68
+ $X2=6.695 $Y2=2.4
r58 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.68
+ $X2=6.245 $Y2=1.515
r59 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.245 $Y=1.68
+ $X2=6.245 $Y2=2.4
r60 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.35
+ $X2=6.23 $Y2=1.515
r61 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.23 $Y=1.35 $X2=6.23
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%VPWR 1 2 9 18 21 22 23 25 35 36 39
r59 40 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 39 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 39 40 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r63 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r64 32 33 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r65 30 39 17.0061 $w=1.7e-07 $l=5.5e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.165 $Y2=3.33
r66 30 32 279.556 $w=1.68e-07 $l=4.285e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=6 $Y2=3.33
r67 28 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 25 39 17.0061 $w=1.7e-07 $l=5.5e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.165 $Y2=3.33
r70 25 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 23 33 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 23 40 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 21 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=3.33 $X2=6
+ $Y2=3.33
r74 21 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=3.33
+ $X2=6.47 $Y2=3.33
r75 20 35 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.96 $Y2=3.33
r76 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.47 $Y2=3.33
r77 16 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=3.33
r78 16 18 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=2.455
r79 12 15 3.77091 $w=1.098e-06 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=2.475
+ $X2=1.165 $Y2=2.815
r80 9 12 3.77091 $w=1.098e-06 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=2.135
+ $X2=1.165 $Y2=2.475
r81 7 39 3.68071 $w=1.1e-06 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=3.245
+ $X2=1.165 $Y2=3.33
r82 7 15 4.76909 $w=1.098e-06 $l=4.3e-07 $layer=LI1_cond $X=1.165 $Y=3.245
+ $X2=1.165 $Y2=2.815
r83 2 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.335
+ $Y=1.84 $X2=6.47 $Y2=2.455
r84 1 15 266.667 $w=1.7e-07 $l=1.1038e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=1.165 $Y2=2.815
r85 1 12 266.667 $w=1.7e-07 $l=1.23596e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=1.6 $Y2=2.475
r86 1 12 266.667 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.475
r87 1 9 266.667 $w=1.7e-07 $l=6.51652e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=1.165 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%A_493_368# 1 2 3 12 16 17 18 19 20 27
c41 16 0 1.11683e-19 $X=3.395 $Y=2.99
r42 21 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=2.275
+ $X2=3.56 $Y2=2.275
r43 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=2.275
+ $X2=4.51 $Y2=2.275
r44 20 21 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.345 $Y=2.275
+ $X2=3.725 $Y2=2.275
r45 18 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=2.36 $X2=3.56
+ $Y2=2.275
r46 18 19 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.56 $Y=2.36
+ $X2=3.56 $Y2=2.905
r47 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=3.56 $Y2=2.905
r48 16 17 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=2.775 $Y2=2.99
r49 12 15 32.9269 $w=2.78e-07 $l=8e-07 $layer=LI1_cond $X=2.635 $Y=2.015
+ $X2=2.635 $Y2=2.815
r50 10 17 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.635 $Y=2.905
+ $X2=2.775 $Y2=2.99
r51 10 15 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.635 $Y=2.905
+ $X2=2.635 $Y2=2.815
r52 3 27 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=4.375
+ $Y=1.84 $X2=4.51 $Y2=2.275
r53 2 25 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=3.375
+ $Y=1.84 $X2=3.56 $Y2=2.355
r54 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.61 $Y2=2.815
r55 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.61 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%Y 1 2 3 4 5 18 20 23 25 26 30 32 36 39 44
+ 46 49 51 54 55
c114 49 0 1.04248e-19 $X=4.12 $Y=1.095
c115 46 0 1.75889e-19 $X=4.12 $Y=0.515
c116 18 0 3.67831e-20 $X=3.955 $Y=0.755
r117 51 55 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.285 $Y=1.665
+ $X2=4.56 $Y2=1.665
r118 51 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.2 $Y=1.665 $X2=4.2
+ $Y2=1.935
r119 46 48 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.12 $Y=0.515
+ $X2=4.12 $Y2=0.755
r120 39 41 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.055 $Y=0.675
+ $X2=3.055 $Y2=0.755
r121 34 36 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=6.45 $Y=1.01
+ $X2=6.45 $Y2=0.515
r122 33 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.215 $Y=1.095
+ $X2=5.09 $Y2=1.095
r123 32 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.325 $Y=1.095
+ $X2=6.45 $Y2=1.01
r124 32 33 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=6.325 $Y=1.095
+ $X2=5.215 $Y2=1.095
r125 28 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=1.01
+ $X2=5.09 $Y2=1.095
r126 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.09 $Y=1.01
+ $X2=5.09 $Y2=0.515
r127 27 49 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=1.095
+ $X2=4.12 $Y2=1.095
r128 26 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.965 $Y=1.095
+ $X2=5.09 $Y2=1.095
r129 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.965 $Y=1.095
+ $X2=4.285 $Y2=1.095
r130 25 51 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.2 $Y=1.55
+ $X2=4.2 $Y2=1.665
r131 24 49 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.2 $Y=1.18
+ $X2=4.12 $Y2=1.095
r132 24 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.2 $Y=1.18 $X2=4.2
+ $Y2=1.55
r133 23 49 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=1.01
+ $X2=4.12 $Y2=1.095
r134 22 48 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=0.84
+ $X2=4.12 $Y2=0.755
r135 22 23 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.12 $Y=0.84
+ $X2=4.12 $Y2=1.01
r136 21 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=1.935
+ $X2=3.1 $Y2=1.935
r137 20 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=1.935
+ $X2=4.2 $Y2=1.935
r138 20 21 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.115 $Y=1.935
+ $X2=3.225 $Y2=1.935
r139 19 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0.755
+ $X2=3.055 $Y2=0.755
r140 18 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0.755
+ $X2=4.12 $Y2=0.755
r141 18 19 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.955 $Y=0.755
+ $X2=3.22 $Y2=0.755
r142 5 44 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=1.84 $X2=3.06 $Y2=2.015
r143 4 36 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=6.305
+ $Y=0.37 $X2=6.49 $Y2=0.515
r144 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.515
r145 2 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.98
+ $Y=0.37 $X2=4.12 $Y2=0.515
r146 1 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%A_775_368# 1 2 9 11 12 15
r26 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.52 $Y=2.905
+ $X2=5.52 $Y2=2.455
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.355 $Y=2.99
+ $X2=5.52 $Y2=2.905
r28 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=5.355 $Y=2.99
+ $X2=4.175 $Y2=2.99
r29 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.035 $Y=2.905
+ $X2=4.175 $Y2=2.99
r30 7 9 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=4.035 $Y=2.905
+ $X2=4.035 $Y2=2.695
r31 2 15 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.385
+ $Y=1.84 $X2=5.52 $Y2=2.455
r32 1 9 600 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.84 $X2=4.06 $Y2=2.695
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%A_985_368# 1 2 3 10 12 14 18 20 22 24 29
c42 18 0 1.98445e-19 $X=6.02 $Y=2.43
r43 22 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=2.12 $X2=6.92
+ $Y2=2.035
r44 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.92 $Y=2.12
+ $X2=6.92 $Y2=2.815
r45 21 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.185 $Y=2.035
+ $X2=6.02 $Y2=2.035
r46 20 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.92 $Y2=2.035
r47 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.185 $Y2=2.035
r48 16 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=2.12 $X2=6.02
+ $Y2=2.035
r49 16 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.02 $Y=2.12 $X2=6.02
+ $Y2=2.43
r50 15 27 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=5.155 $Y=2.035
+ $X2=5.03 $Y2=1.97
r51 14 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=6.02 $Y2=2.035
r52 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=5.155 $Y2=2.035
r53 10 27 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=5.03 $Y=2.12 $X2=5.03
+ $Y2=1.97
r54 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=5.03 $Y=2.12 $X2=5.03
+ $Y2=2.57
r55 3 31 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.84 $X2=6.92 $Y2=2.035
r56 3 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.84 $X2=6.92 $Y2=2.815
r57 2 29 600 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.84 $X2=6.02 $Y2=2.035
r58 2 18 300 $w=1.7e-07 $l=6.76203e-07 $layer=licon1_PDIFF $count=2 $X=5.835
+ $Y=1.84 $X2=6.02 $Y2=2.43
r59 1 27 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.84 $X2=5.07 $Y2=1.985
r60 1 12 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=1.84 $X2=5.07 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_2%VGND 1 2 3 4 5 6 21 25 27 29 32 38 40 49 53
+ 58 63 76 79 83 92
r87 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 84 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r89 83 88 10.4851 $w=7.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.77 $Y=0 $X2=5.77
+ $Y2=0.675
r90 83 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r91 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r93 67 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r94 67 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r95 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r96 64 83 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=5.77
+ $Y2=0
r97 64 66 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.48
+ $Y2=0
r98 63 91 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r99 63 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r100 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r101 62 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r102 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r103 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=4.62
+ $Y2=0
r104 59 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=0
+ $X2=5.04 $Y2=0
r105 58 83 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.77
+ $Y2=0
r106 58 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.04
+ $Y2=0
r107 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r108 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 54 76 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=3.587 $Y2=0
r110 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=4.08 $Y2=0
r111 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.62
+ $Y2=0
r112 53 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.455 $Y=0
+ $X2=4.08 $Y2=0
r113 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r114 49 76 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.587
+ $Y2=0
r115 49 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.12
+ $Y2=0
r116 48 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r117 48 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r118 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r119 45 47 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=2.16 $Y2=0
r120 43 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r122 40 73 10.2521 $w=5.23e-07 $l=4.5e-07 $layer=LI1_cond $X=1.252 $Y=0
+ $X2=1.252 $Y2=0.45
r123 40 45 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=1.252 $Y=0
+ $X2=1.515 $Y2=0
r124 40 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 40 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r126 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r127 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r128 38 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r129 34 51 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=3.12
+ $Y2=0
r130 32 47 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.16
+ $Y2=0
r131 32 36 8.70931 $w=5.13e-07 $l=3.75e-07 $layer=LI1_cond $X=2.452 $Y=0
+ $X2=2.452 $Y2=0.375
r132 32 34 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=2.452 $Y=0 $X2=2.71
+ $Y2=0
r133 27 91 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r134 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r135 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=0.085
+ $X2=4.62 $Y2=0
r136 23 25 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=4.62 $Y=0.085
+ $X2=4.62 $Y2=0.675
r137 19 76 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.587 $Y=0.085
+ $X2=3.587 $Y2=0
r138 19 21 7.68295 $w=3.73e-07 $l=2.5e-07 $layer=LI1_cond $X=3.587 $Y=0.085
+ $X2=3.587 $Y2=0.335
r139 6 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.78
+ $Y=0.37 $X2=6.92 $Y2=0.515
r140 5 88 91 $w=1.7e-07 $l=8.13326e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=6.015 $Y2=0.675
r141 4 25 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.37 $X2=4.62 $Y2=0.675
r142 3 21 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=3.345
+ $Y=0.37 $X2=3.585 $Y2=0.335
r143 2 36 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.23 $X2=2.45 $Y2=0.375
r144 1 73 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.37 $X2=1.16 $Y2=0.45
.ends


* File: sky130_fd_sc_ms__o32ai_4.spice
* Created: Wed Sep  2 12:26:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o32ai_4.pex.spice"
.subckt sky130_fd_sc_ms__o32ai_4  VNB VPB B2 B1 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1022 N_A_27_74#_M1022_d N_B2_M1022_g N_Y_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75010 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_74#_M1030_d N_B2_M1030_g N_Y_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75009.6 A=0.111 P=1.78 MULT=1
MM1031 N_A_27_74#_M1030_d N_B2_M1031_g N_Y_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.10915 PD=1.09 PS=1.035 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75009.1 A=0.111 P=1.78 MULT=1
MM1032 N_A_27_74#_M1032_d N_B2_M1032_g N_Y_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12395 AS=0.10915 PD=1.075 PS=1.035 NRD=8.916 NRS=2.424 M=1 R=4.93333
+ SA=75001.6 SB=75008.6 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_74#_M1032_d N_B1_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12395 AS=0.1295 PD=1.075 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75008.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1004_d N_B1_M1004_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75007.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1004_d N_B1_M1011_g N_Y_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.1
+ SB=75007.1 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_B1_M1014_g N_Y_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75006.6 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_74#_M1014_d N_A3_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1773 PD=1.09 PS=1.28 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75004.1
+ SB=75006.1 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1033_d N_A3_M1033_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12765 AS=0.1773 PD=1.085 PS=1.28 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75004.7 SB=75005.6 A=0.111 P=1.78 MULT=1
MM1036 N_A_27_74#_M1033_d N_A3_M1036_g N_VGND_M1036_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12765 AS=0.10545 PD=1.085 PS=1.025 NRD=10.536 NRS=0.804 M=1 R=4.93333
+ SA=75005.2 SB=75005.1 A=0.111 P=1.78 MULT=1
MM1038 N_A_27_74#_M1038_d N_A3_M1038_g N_VGND_M1036_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2626 AS=0.10545 PD=1.455 PS=1.025 NRD=33.24 NRS=0 M=1 R=4.93333
+ SA=75005.6 SB=75004.6 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_27_74#_M1038_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2626 PD=1.16 PS=1.455 NRD=11.34 NRS=34.044 M=1 R=4.93333
+ SA=75006.4 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1005_d N_A2_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A2_M1017_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1034 N_VGND_M1017_d N_A2_M1034_g N_A_27_74#_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1295 PD=1.16 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75008
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_27_74#_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75008.5
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1002_d N_A1_M1018_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75009
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A1_M1027_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75009.4
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1039 N_VGND_M1027_d N_A1_M1039_g N_A_27_74#_M1039_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2627 PD=1.09 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75009.9
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1015_d N_B2_M1015_g N_A_27_368#_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1016 N_Y_M1015_d N_B2_M1016_g N_A_27_368#_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1019 N_Y_M1019_d N_B2_M1019_g N_A_27_368#_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1020 N_Y_M1019_d N_B2_M1020_g N_A_27_368#_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1012 N_A_27_368#_M1020_s N_B1_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1023 N_A_27_368#_M1023_d N_B1_M1023_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1025 N_A_27_368#_M1023_d N_B1_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1028 N_A_27_368#_M1028_d N_B1_M1028_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1568 PD=2.8 PS=1.4 NRD=0 NRS=0.8668 M=1 R=6.22222 SA=90003.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_A3_M1006_g N_A_861_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.6 A=0.2016 P=2.6 MULT=1
MM1013 N_Y_M1006_d N_A3_M1013_g N_A_861_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1029 N_Y_M1029_d N_A3_M1029_g N_A_861_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1037 N_Y_M1029_d N_A3_M1037_g N_A_861_368#_M1037_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.5
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1003 N_A_1333_368#_M1003_d N_A2_M1003_g N_A_861_368#_M1037_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.1 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1007 N_A_1333_368#_M1003_d N_A2_M1007_g N_A_861_368#_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.5 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1009 N_A_1333_368#_M1009_d N_A2_M1009_g N_A_861_368#_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90003 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1010 N_A_1333_368#_M1009_d N_A2_M1010_g N_A_861_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.3696 PD=1.44 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90003.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1021 N_A_1333_368#_M1021_d N_A1_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1024 N_A_1333_368#_M1021_d N_A1_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.6 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1026 N_A_1333_368#_M1026_d N_A1_M1026_g N_VPWR_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1035 N_A_1333_368#_M1026_d N_A1_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=21.2412 P=26.56
*
.include "sky130_fd_sc_ms__o32ai_4.pxi.spice"
*
.ends
*
*

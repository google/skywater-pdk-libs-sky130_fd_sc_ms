* File: sky130_fd_sc_ms__edfxtp_1.spice
* Created: Wed Sep  2 12:08:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__edfxtp_1.pex.spice"
.subckt sky130_fd_sc_ms__edfxtp_1  VNB VPB D DE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1009 A_131_74# N_D_M1009_g N_A_27_508#_M1009_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_DE_M1006_g A_131_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1176
+ AS=0.0504 PD=1.4 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_DE_M1010_g N_A_159_446#_M1010_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1021 A_491_87# N_A_159_446#_M1021_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_27_508#_M1022_d N_A_533_61#_M1022_g A_491_87# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_763_74#_M1011_d N_CLK_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.2109 PD=2.03 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_A_958_74#_M1033_d N_A_763_74#_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2072 PD=2.05 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_1156_90#_M1024_d N_A_763_74#_M1024_g N_A_27_508#_M1024_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.17115 AS=0.1197 PD=1.235 PS=1.41 NRD=134.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1028 A_1349_90# N_A_958_74#_M1028_g N_A_1156_90#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.063 AS=0.17115 PD=0.72 PS=1.235 NRD=27.132 NRS=18.564 M=1 R=2.8
+ SA=75001.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1409_64#_M1001_g A_1349_90# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109992 AS=0.063 PD=0.92717 PS=0.72 NRD=0 NRS=27.132 M=1 R=2.8 SA=75001.6
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_1409_64#_M1004_d N_A_1156_90#_M1004_g N_VGND_M1001_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.167608 PD=1.85 PS=1.41283 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 A_1797_74# N_A_1409_64#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2109 PD=1.08 PS=2.05 NRD=18.648 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1029 N_A_1895_74#_M1029_d N_A_958_74#_M1029_g A_1797_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.154634 AS=0.1258 PD=1.40345 PS=1.08 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75000.7 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1007 A_1997_74# N_A_763_74#_M1007_g N_A_1895_74#_M1029_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0877655 PD=0.66 PS=0.796552 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_533_61#_M1002_g A_1997_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20055 AS=0.0504 PD=1.375 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_533_61#_M1003_d N_A_1895_74#_M1003_g N_VGND_M1002_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.20055 PD=1.41 PS=1.375 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_1895_74#_M1019_g N_Q_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 A_117_508# N_D_M1008_g N_A_27_508#_M1008_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0441 AS=0.1134 PD=0.63 PS=1.38 NRD=23.443 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_A_159_446#_M1015_g A_117_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333 SA=90000.6
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1032 N_VPWR_M1032_d N_DE_M1032_g N_A_159_446#_M1032_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.3766 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1016 A_557_436# N_DE_M1016_g N_VPWR_M1032_d VPB PSHORT L=0.18 W=0.42 AD=0.0441
+ AS=0.105 PD=0.63 PS=0.903396 NRD=23.443 NRS=0 M=1 R=2.33333 SA=90000.9
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1027 N_A_27_508#_M1027_d N_A_533_61#_M1027_g A_557_436# VPB PSHORT L=0.18
+ W=0.42 AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333
+ SA=90001.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1025 N_A_763_74#_M1025_d N_CLK_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2968 PD=2.76 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1005 N_A_958_74#_M1005_d N_A_763_74#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1013 N_A_1156_90#_M1013_d N_A_958_74#_M1013_g N_A_27_508#_M1013_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1113 PD=0.69 PS=1.37 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1017 A_1385_508# N_A_763_74#_M1017_g N_A_1156_90#_M1013_d VPB PSHORT L=0.18
+ W=0.42 AD=0.06825 AS=0.0567 PD=0.745 PS=0.69 NRD=50.4123 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1409_64#_M1020_g A_1385_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0916417 AS=0.06825 PD=0.866667 PS=0.745 NRD=2.3443 NRS=50.4123 M=1
+ R=2.33333 SA=90001.1 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1023 N_A_1409_64#_M1023_d N_A_1156_90#_M1023_g N_VPWR_M1020_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.183283 PD=2.24 PS=1.73333 NRD=0 NRS=19.9167 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1018 A_1797_392# N_A_1409_64#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.3775 AS=0.28 PD=1.755 PS=2.56 NRD=63.5128 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1030 N_A_1895_74#_M1030_d N_A_763_74#_M1030_g A_1797_392# VPB PSHORT L=0.18
+ W=1 AD=0.219366 AS=0.3775 PD=1.90845 PS=1.755 NRD=0 NRS=63.5128 M=1 R=5.55556
+ SA=90001.1 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1026 A_2091_502# N_A_958_74#_M1026_g N_A_1895_74#_M1030_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0921338 PD=0.66 PS=0.801549 NRD=30.4759 NRS=38.6908 M=1
+ R=2.33333 SA=90001.7 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_533_61#_M1000_g A_2091_502# VPB PSHORT L=0.18 W=0.42
+ AD=0.109992 AS=0.0504 PD=0.92717 PS=0.66 NRD=58.6272 NRS=30.4759 M=1 R=2.33333
+ SA=90002.1 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1014 N_A_533_61#_M1014_d N_A_1895_74#_M1014_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1664 AS=0.167608 PD=1.8 PS=1.41283 NRD=0 NRS=38.4741 M=1 R=3.55556
+ SA=90001.9 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1031 N_VPWR_M1031_d N_A_1895_74#_M1031_g N_Q_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.2912 PD=2.78 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=24.8976 P=30.56
c_143 VNB 0 4.56061e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__edfxtp_1.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ms__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__nand3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 4.195000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.430000 1.795000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.232000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.260000 1.950000 3.695000 2.120000 ;
        RECT 1.260000 2.120000 1.635000 2.980000 ;
        RECT 2.335000 2.120000 2.585000 2.980000 ;
        RECT 2.470000 1.010000 2.800000 1.180000 ;
        RECT 2.525000 1.180000 2.800000 1.950000 ;
        RECT 3.365000 2.120000 3.695000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 4.320000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 4.510000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.100000  0.450000 0.350000 1.090000 ;
      RECT 0.100000  1.090000 2.195000 1.260000 ;
      RECT 0.305000  1.950000 0.890000 2.120000 ;
      RECT 0.305000  2.120000 0.635000 2.980000 ;
      RECT 0.530000  0.085000 0.820000 0.910000 ;
      RECT 0.720000  1.260000 0.890000 1.950000 ;
      RECT 0.830000  2.290000 1.075000 3.245000 ;
      RECT 1.005000  0.330000 1.255000 0.750000 ;
      RECT 1.005000  0.750000 3.790000 0.840000 ;
      RECT 1.005000  0.840000 2.105000 0.920000 ;
      RECT 1.435000  0.085000 1.765000 0.580000 ;
      RECT 1.805000  2.290000 2.135000 3.245000 ;
      RECT 1.935000  0.670000 3.790000 0.750000 ;
      RECT 1.975000  0.330000 4.220000 0.500000 ;
      RECT 2.025000  1.260000 2.195000 1.350000 ;
      RECT 2.025000  1.350000 2.355000 1.680000 ;
      RECT 2.790000  2.290000 3.120000 3.245000 ;
      RECT 2.970000  0.840000 3.790000 1.180000 ;
      RECT 3.875000  1.950000 4.205000 3.245000 ;
      RECT 3.960000  0.500000 4.220000 1.180000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__nand3b_2
END LIBRARY

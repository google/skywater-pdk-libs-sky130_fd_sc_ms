* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_300_387# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 a_300_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_27_125# B1 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_114_125# A2 a_766_387# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_300_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 X a_114_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 X a_114_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_114_125# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 a_27_125# B2 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VPWR A1 a_766_387# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X10 VGND A2 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VGND a_114_125# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_114_125# B2 a_300_387# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 VPWR C1 a_114_125# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 VPWR B1 a_300_387# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 a_300_125# B1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_300_125# B2 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 VPWR a_114_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 X a_114_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 a_27_125# C1 a_114_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 X a_114_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VGND A1 a_300_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 VGND a_114_125# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_766_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X24 a_114_125# C1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X25 VPWR a_114_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 a_300_387# B2 a_114_125# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X27 a_766_387# A2 a_114_125# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__nand4_4.pxi.spice
* Created: Fri Aug 28 17:44:57 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4_4%D N_D_M1006_g N_D_M1008_g N_D_c_109_n N_D_M1014_g
+ N_D_M1005_g N_D_M1019_g N_D_M1007_g N_D_c_112_n N_D_c_113_n N_D_c_114_n D D D
+ D D N_D_c_116_n PM_SKY130_FD_SC_MS__NAND4_4%D
x_PM_SKY130_FD_SC_MS__NAND4_4%C N_C_M1001_g N_C_M1009_g N_C_M1010_g N_C_M1018_g
+ N_C_M1011_g N_C_M1020_g C C C C N_C_c_186_n PM_SKY130_FD_SC_MS__NAND4_4%C
x_PM_SKY130_FD_SC_MS__NAND4_4%B N_B_M1000_g N_B_M1003_g N_B_M1017_g N_B_M1004_g
+ N_B_M1016_g N_B_M1021_g B B B B N_B_c_244_n PM_SKY130_FD_SC_MS__NAND4_4%B
x_PM_SKY130_FD_SC_MS__NAND4_4%A N_A_M1002_g N_A_M1012_g N_A_M1013_g N_A_M1015_g
+ N_A_M1022_g N_A_M1023_g N_A_c_308_n N_A_c_309_n A A A N_A_c_310_n
+ PM_SKY130_FD_SC_MS__NAND4_4%A
x_PM_SKY130_FD_SC_MS__NAND4_4%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_M1018_s
+ N_VPWR_M1017_d N_VPWR_M1022_d N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n
+ N_VPWR_c_375_n N_VPWR_c_376_n VPWR N_VPWR_c_377_n N_VPWR_c_378_n
+ N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n
+ N_VPWR_c_371_n PM_SKY130_FD_SC_MS__NAND4_4%VPWR
x_PM_SKY130_FD_SC_MS__NAND4_4%Y N_Y_M1002_d N_Y_M1015_d N_Y_M1005_s N_Y_M1009_d
+ N_Y_M1000_s N_Y_M1013_s N_Y_c_448_n N_Y_c_442_n N_Y_c_453_n N_Y_c_443_n
+ N_Y_c_459_n N_Y_c_444_n N_Y_c_468_n N_Y_c_437_n N_Y_c_445_n N_Y_c_438_n
+ N_Y_c_446_n N_Y_c_462_n N_Y_c_472_n N_Y_c_485_n N_Y_c_439_n N_Y_c_440_n Y Y
+ PM_SKY130_FD_SC_MS__NAND4_4%Y
x_PM_SKY130_FD_SC_MS__NAND4_4%A_27_74# N_A_27_74#_M1006_s N_A_27_74#_M1008_s
+ N_A_27_74#_M1019_s N_A_27_74#_M1010_s N_A_27_74#_M1020_s N_A_27_74#_c_533_n
+ N_A_27_74#_c_534_n N_A_27_74#_c_535_n N_A_27_74#_c_536_n N_A_27_74#_c_537_n
+ N_A_27_74#_c_538_n N_A_27_74#_c_557_n N_A_27_74#_c_539_n N_A_27_74#_c_540_n
+ PM_SKY130_FD_SC_MS__NAND4_4%A_27_74#
x_PM_SKY130_FD_SC_MS__NAND4_4%VGND N_VGND_M1006_d N_VGND_M1014_d N_VGND_c_595_n
+ N_VGND_c_596_n N_VGND_c_597_n VGND N_VGND_c_598_n N_VGND_c_599_n
+ N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n PM_SKY130_FD_SC_MS__NAND4_4%VGND
x_PM_SKY130_FD_SC_MS__NAND4_4%A_554_74# N_A_554_74#_M1001_d N_A_554_74#_M1011_d
+ N_A_554_74#_M1003_s N_A_554_74#_M1016_s N_A_554_74#_c_663_n
+ N_A_554_74#_c_664_n N_A_554_74#_c_665_n N_A_554_74#_c_666_n
+ N_A_554_74#_c_667_n PM_SKY130_FD_SC_MS__NAND4_4%A_554_74#
x_PM_SKY130_FD_SC_MS__NAND4_4%A_923_74# N_A_923_74#_M1003_d N_A_923_74#_M1004_d
+ N_A_923_74#_M1021_d N_A_923_74#_M1012_s N_A_923_74#_M1023_s
+ N_A_923_74#_c_703_n N_A_923_74#_c_704_n N_A_923_74#_c_705_n
+ N_A_923_74#_c_706_n N_A_923_74#_c_707_n N_A_923_74#_c_708_n
+ N_A_923_74#_c_709_n N_A_923_74#_c_710_n N_A_923_74#_c_711_n
+ PM_SKY130_FD_SC_MS__NAND4_4%A_923_74#
cc_1 VNB N_D_M1006_g 0.0336211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_D_M1008_g 0.024496f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_D_c_109_n 0.0155552f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.515
cc_4 VNB N_D_M1014_g 0.0272963f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_5 VNB N_D_M1019_g 0.0277516f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_6 VNB N_D_c_112_n 0.0137535f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.515
cc_7 VNB N_D_c_113_n 0.0155576f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_8 VNB N_D_c_114_n 0.004935f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_9 VNB D 0.0166475f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_10 VNB N_D_c_116_n 0.0480683f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.515
cc_11 VNB N_C_M1001_g 0.0250243f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_12 VNB N_C_M1010_g 0.0234232f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.35
cc_13 VNB N_C_M1011_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.35
cc_14 VNB N_C_M1020_g 0.0337355f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.68
cc_15 VNB C 0.00704574f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_16 VNB N_C_c_186_n 0.0644659f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.515
cc_17 VNB N_B_M1003_g 0.0336884f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_18 VNB N_B_M1004_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.68
cc_19 VNB N_B_M1016_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.35
cc_20 VNB N_B_M1021_g 0.0241156f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.68
cc_21 VNB B 0.00267486f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_22 VNB N_B_c_244_n 0.0920128f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.515
cc_23 VNB N_A_M1002_g 0.0241156f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_24 VNB N_A_M1012_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_25 VNB N_A_M1015_g 0.0255586f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.68
cc_26 VNB N_A_M1023_g 0.0301963f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.68
cc_27 VNB N_A_c_308_n 0.0199665f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_28 VNB N_A_c_309_n 0.0136818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_c_310_n 0.0445768f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_30 VNB N_VPWR_c_371_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_437_n 0.00204539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_438_n 0.0145179f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_33 VNB N_Y_c_439_n 0.00408444f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.565
cc_34 VNB N_Y_c_440_n 0.00133991f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_35 VNB Y 0.0265321f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_36 VNB N_A_27_74#_c_533_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_534_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_38 VNB N_A_27_74#_c_535_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_39 VNB N_A_27_74#_c_536_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_40 VNB N_A_27_74#_c_537_n 0.0136988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_538_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_42 VNB N_A_27_74#_c_539_n 0.0136639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_540_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_595_n 0.00586453f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.515
cc_45 VNB N_VGND_c_596_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.35
cc_46 VNB N_VGND_c_597_n 0.00916033f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.68
cc_47 VNB N_VGND_c_598_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.35
cc_48 VNB N_VGND_c_599_n 0.168013f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_49 VNB N_VGND_c_600_n 0.467293f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_50 VNB N_VGND_c_601_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_51 VNB N_VGND_c_602_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_554_74#_c_663_n 0.00641753f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_53 VNB N_A_554_74#_c_664_n 0.0062129f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_54 VNB N_A_554_74#_c_665_n 0.00108276f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.68
cc_55 VNB N_A_554_74#_c_666_n 0.0265392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_554_74#_c_667_n 0.00159267f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.515
cc_57 VNB N_A_923_74#_c_703_n 0.00374122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_923_74#_c_704_n 0.00643668f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_59 VNB N_A_923_74#_c_705_n 0.002345f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_60 VNB N_A_923_74#_c_706_n 0.00237781f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_61 VNB N_A_923_74#_c_707_n 0.002345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_923_74#_c_708_n 0.00237781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_923_74#_c_709_n 0.002345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_923_74#_c_710_n 0.00237781f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.515
cc_65 VNB N_A_923_74#_c_711_n 0.0171072f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.515
cc_66 VPB N_D_c_109_n 0.0106787f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.515
cc_67 VPB N_D_M1005_g 0.0252124f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=2.4
cc_68 VPB N_D_M1007_g 0.0211634f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.4
cc_69 VPB N_D_c_112_n 0.00517001f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.515
cc_70 VPB N_D_c_113_n 0.0106787f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_71 VPB N_D_c_114_n 0.00459923f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_72 VPB D 0.0233118f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_73 VPB N_D_c_116_n 0.013497f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=1.515
cc_74 VPB N_C_M1009_g 0.023379f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_75 VPB N_C_M1018_g 0.0287153f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=1.68
cc_76 VPB C 0.0139215f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_77 VPB N_C_c_186_n 0.0293676f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.515
cc_78 VPB N_B_M1000_g 0.0287153f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_79 VPB N_B_M1017_g 0.0287439f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=1.35
cc_80 VPB B 0.0154502f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_81 VPB N_B_c_244_n 0.0425974f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.515
cc_82 VPB N_A_M1013_g 0.0322708f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=1.35
cc_83 VPB N_A_M1022_g 0.0299648f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.35
cc_84 VPB N_A_c_308_n 0.0099814f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.4
cc_85 VPB N_A_c_309_n 8.82697e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB A 0.0120739f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_87 VPB N_A_c_310_n 0.0236005f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_88 VPB N_VPWR_c_372_n 0.00341267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_373_n 0.0251016f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=0.74
cc_90 VPB N_VPWR_c_374_n 0.0090297f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.4
cc_91 VPB N_VPWR_c_375_n 0.0121562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_376_n 0.0355096f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_93 VPB N_VPWR_c_377_n 0.0185368f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_94 VPB N_VPWR_c_378_n 0.10355f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_95 VPB N_VPWR_c_379_n 0.027658f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.515
cc_96 VPB N_VPWR_c_380_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_381_n 0.016897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_382_n 0.0251007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_383_n 0.0494568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_371_n 0.0711077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_Y_c_442_n 0.00275675f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=0.74
cc_102 VPB N_Y_c_443_n 0.00587533f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.515
cc_103 VPB N_Y_c_444_n 0.00587443f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_104 VPB N_Y_c_445_n 0.00663712f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.515
cc_105 VPB N_Y_c_446_n 0.00714919f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.515
cc_106 VPB Y 0.0128922f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_107 N_D_M1019_g N_C_M1001_g 0.0255149f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_108 N_D_M1007_g N_C_M1009_g 0.0249033f $X=2.26 $Y=2.4 $X2=0 $Y2=0
cc_109 D C 0.0285068f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_110 N_D_c_116_n C 0.00366877f $X=2.26 $Y=1.515 $X2=0 $Y2=0
cc_111 D N_C_c_186_n 4.14707e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_112 N_D_c_116_n N_C_c_186_n 0.0249033f $X=2.26 $Y=1.515 $X2=0 $Y2=0
cc_113 N_D_M1005_g N_VPWR_c_372_n 5.17373e-19 $X=1.76 $Y=2.4 $X2=0 $Y2=0
cc_114 N_D_M1007_g N_VPWR_c_372_n 0.0125259f $X=2.26 $Y=2.4 $X2=0 $Y2=0
cc_115 N_D_M1005_g N_VPWR_c_377_n 0.005209f $X=1.76 $Y=2.4 $X2=0 $Y2=0
cc_116 N_D_M1007_g N_VPWR_c_377_n 0.00460063f $X=2.26 $Y=2.4 $X2=0 $Y2=0
cc_117 N_D_M1005_g N_VPWR_c_378_n 0.00419671f $X=1.76 $Y=2.4 $X2=0 $Y2=0
cc_118 N_D_c_112_n N_VPWR_c_378_n 0.00741187f $X=0.57 $Y=1.515 $X2=0 $Y2=0
cc_119 D N_VPWR_c_378_n 0.133163f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_120 N_D_M1005_g N_VPWR_c_371_n 0.00987193f $X=1.76 $Y=2.4 $X2=0 $Y2=0
cc_121 N_D_M1007_g N_VPWR_c_371_n 0.00909043f $X=2.26 $Y=2.4 $X2=0 $Y2=0
cc_122 N_D_M1005_g N_Y_c_448_n 0.00241985f $X=1.76 $Y=2.4 $X2=0 $Y2=0
cc_123 D N_Y_c_448_n 0.0246996f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_124 N_D_c_116_n N_Y_c_448_n 8.59451e-19 $X=2.26 $Y=1.515 $X2=0 $Y2=0
cc_125 N_D_M1005_g N_Y_c_442_n 0.0106812f $X=1.76 $Y=2.4 $X2=0 $Y2=0
cc_126 N_D_M1007_g N_Y_c_442_n 2.25304e-19 $X=2.26 $Y=2.4 $X2=0 $Y2=0
cc_127 N_D_M1007_g N_Y_c_453_n 0.0163757f $X=2.26 $Y=2.4 $X2=0 $Y2=0
cc_128 D N_Y_c_453_n 0.00849394f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_129 N_D_M1006_g N_A_27_74#_c_533_n 0.0102216f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_D_M1008_g N_A_27_74#_c_533_n 6.38603e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_131 N_D_M1006_g N_A_27_74#_c_534_n 0.0115433f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_D_M1008_g N_A_27_74#_c_534_n 0.0151263f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_133 N_D_c_113_n N_A_27_74#_c_534_n 0.00381149f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_134 D N_A_27_74#_c_534_n 0.0501792f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_D_M1006_g N_A_27_74#_c_535_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_136 D N_A_27_74#_c_535_n 0.0286342f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_137 N_D_M1008_g N_A_27_74#_c_536_n 0.00350341f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_138 N_D_M1014_g N_A_27_74#_c_536_n 0.010082f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_139 N_D_M1019_g N_A_27_74#_c_536_n 7.91979e-19 $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_140 N_D_M1014_g N_A_27_74#_c_537_n 0.0123334f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_141 N_D_M1019_g N_A_27_74#_c_537_n 0.013916f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_142 D N_A_27_74#_c_537_n 0.062829f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_D_c_116_n N_A_27_74#_c_537_n 0.0131245f $X=2.26 $Y=1.515 $X2=0 $Y2=0
cc_144 N_D_M1019_g N_A_27_74#_c_538_n 0.00502264f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_145 N_D_M1014_g N_A_27_74#_c_557_n 7.59304e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_146 N_D_M1019_g N_A_27_74#_c_557_n 0.00666311f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_147 N_D_c_109_n N_A_27_74#_c_540_n 0.00396026f $X=1.42 $Y=1.515 $X2=0 $Y2=0
cc_148 N_D_M1014_g N_A_27_74#_c_540_n 0.00173883f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_149 D N_A_27_74#_c_540_n 0.0281948f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_D_M1006_g N_VGND_c_595_n 0.00571035f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_151 N_D_M1008_g N_VGND_c_595_n 0.0109084f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_152 N_D_M1014_g N_VGND_c_595_n 4.99121e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_153 N_D_M1008_g N_VGND_c_596_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_154 N_D_M1014_g N_VGND_c_596_n 0.00434272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_155 N_D_M1014_g N_VGND_c_597_n 0.00572004f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_156 N_D_M1019_g N_VGND_c_597_n 0.00777206f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_157 N_D_M1006_g N_VGND_c_598_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_158 N_D_M1019_g N_VGND_c_599_n 0.00433139f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_159 N_D_M1006_g N_VGND_c_600_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_160 N_D_M1008_g N_VGND_c_600_n 0.00758198f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_161 N_D_M1014_g N_VGND_c_600_n 0.00822835f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_162 N_D_M1019_g N_VGND_c_600_n 0.0082043f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_163 C B 0.0305568f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_164 N_C_c_186_n B 0.00116481f $X=3.985 $Y=1.515 $X2=0 $Y2=0
cc_165 C N_B_c_244_n 0.00216742f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_166 N_C_c_186_n N_B_c_244_n 0.00895304f $X=3.985 $Y=1.515 $X2=0 $Y2=0
cc_167 N_C_M1009_g N_VPWR_c_372_n 0.0153239f $X=2.71 $Y=2.4 $X2=0 $Y2=0
cc_168 N_C_M1009_g N_VPWR_c_373_n 0.00460063f $X=2.71 $Y=2.4 $X2=0 $Y2=0
cc_169 N_C_M1018_g N_VPWR_c_373_n 0.00460063f $X=3.54 $Y=2.4 $X2=0 $Y2=0
cc_170 N_C_M1018_g N_VPWR_c_374_n 0.0176127f $X=3.54 $Y=2.4 $X2=0 $Y2=0
cc_171 N_C_M1009_g N_VPWR_c_371_n 0.00911317f $X=2.71 $Y=2.4 $X2=0 $Y2=0
cc_172 N_C_M1018_g N_VPWR_c_371_n 0.00911317f $X=3.54 $Y=2.4 $X2=0 $Y2=0
cc_173 N_C_M1009_g N_Y_c_453_n 0.0142175f $X=2.71 $Y=2.4 $X2=0 $Y2=0
cc_174 C N_Y_c_453_n 0.019463f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_175 N_C_M1009_g N_Y_c_443_n 3.56899e-19 $X=2.71 $Y=2.4 $X2=0 $Y2=0
cc_176 N_C_M1018_g N_Y_c_443_n 3.56899e-19 $X=3.54 $Y=2.4 $X2=0 $Y2=0
cc_177 N_C_M1018_g N_Y_c_459_n 0.0163793f $X=3.54 $Y=2.4 $X2=0 $Y2=0
cc_178 C N_Y_c_459_n 0.0568989f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_179 N_C_c_186_n N_Y_c_459_n 0.00221855f $X=3.985 $Y=1.515 $X2=0 $Y2=0
cc_180 C N_Y_c_462_n 0.0506009f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_181 N_C_c_186_n N_Y_c_462_n 0.00287383f $X=3.985 $Y=1.515 $X2=0 $Y2=0
cc_182 N_C_M1001_g N_A_27_74#_c_537_n 0.00237285f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_183 C N_A_27_74#_c_537_n 0.00450841f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_184 N_C_M1001_g N_A_27_74#_c_539_n 0.0186789f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_185 N_C_M1010_g N_A_27_74#_c_539_n 0.0123211f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_186 N_C_M1011_g N_A_27_74#_c_539_n 0.0123211f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_187 N_C_M1020_g N_A_27_74#_c_539_n 0.0126246f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_188 C N_A_27_74#_c_539_n 0.00379054f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_189 N_C_M1001_g N_VGND_c_599_n 0.00291649f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_190 N_C_M1010_g N_VGND_c_599_n 0.00291649f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_191 N_C_M1011_g N_VGND_c_599_n 0.00291649f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_192 N_C_M1020_g N_VGND_c_599_n 0.00291649f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_193 N_C_M1001_g N_VGND_c_600_n 0.00359833f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_194 N_C_M1010_g N_VGND_c_600_n 0.00359121f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_195 N_C_M1011_g N_VGND_c_600_n 0.00359121f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_196 N_C_M1020_g N_VGND_c_600_n 0.0036412f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_197 N_C_M1001_g N_A_554_74#_c_663_n 0.00380276f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_198 N_C_M1010_g N_A_554_74#_c_663_n 0.0119209f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_199 N_C_M1011_g N_A_554_74#_c_663_n 0.0119209f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_200 C N_A_554_74#_c_663_n 0.0936883f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_201 N_C_c_186_n N_A_554_74#_c_663_n 0.00681933f $X=3.985 $Y=1.515 $X2=0 $Y2=0
cc_202 N_C_M1020_g N_A_554_74#_c_665_n 0.00288027f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_203 N_C_M1020_g N_A_554_74#_c_666_n 0.0127268f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_204 N_C_M1020_g N_A_923_74#_c_704_n 6.08634e-19 $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_M1021_g N_A_M1002_g 0.0255996f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_206 B A 0.0140912f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_207 N_B_c_244_n A 0.00131406f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_208 B N_A_c_310_n 0.00116053f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_209 N_B_c_244_n N_A_c_310_n 0.0255996f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_210 N_B_M1000_g N_VPWR_c_374_n 0.0176127f $X=4.56 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B_M1000_g N_VPWR_c_382_n 0.00460063f $X=4.56 $Y=2.4 $X2=0 $Y2=0
cc_212 N_B_M1017_g N_VPWR_c_382_n 0.00460063f $X=5.39 $Y=2.4 $X2=0 $Y2=0
cc_213 N_B_M1017_g N_VPWR_c_383_n 0.0176762f $X=5.39 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B_M1000_g N_VPWR_c_371_n 0.00911317f $X=4.56 $Y=2.4 $X2=0 $Y2=0
cc_215 N_B_M1017_g N_VPWR_c_371_n 0.0090668f $X=5.39 $Y=2.4 $X2=0 $Y2=0
cc_216 N_B_M1000_g N_Y_c_459_n 0.0163793f $X=4.56 $Y=2.4 $X2=0 $Y2=0
cc_217 B N_Y_c_459_n 0.0150495f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_218 N_B_M1000_g N_Y_c_444_n 3.56899e-19 $X=4.56 $Y=2.4 $X2=0 $Y2=0
cc_219 N_B_M1017_g N_Y_c_444_n 3.56489e-19 $X=5.39 $Y=2.4 $X2=0 $Y2=0
cc_220 N_B_M1017_g N_Y_c_468_n 0.0163499f $X=5.39 $Y=2.4 $X2=0 $Y2=0
cc_221 B N_Y_c_468_n 0.0660586f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B_c_244_n N_Y_c_468_n 0.0102833f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_223 N_B_M1021_g N_Y_c_437_n 7.32989e-19 $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_224 B N_Y_c_472_n 0.0506009f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B_c_244_n N_Y_c_472_n 0.0028802f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_226 N_B_M1003_g N_A_27_74#_c_539_n 7.21241e-19 $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B_M1003_g N_VGND_c_599_n 0.00292759f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B_M1004_g N_VGND_c_599_n 0.00291649f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B_M1016_g N_VGND_c_599_n 0.00291649f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B_M1021_g N_VGND_c_599_n 0.00291649f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B_M1003_g N_VGND_c_600_n 0.00363156f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B_M1004_g N_VGND_c_600_n 0.00359121f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B_M1016_g N_VGND_c_600_n 0.00359121f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B_M1021_g N_VGND_c_600_n 0.00359219f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B_M1004_g N_A_554_74#_c_664_n 0.0120015f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B_M1016_g N_A_554_74#_c_664_n 0.0131801f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B_M1021_g N_A_554_74#_c_664_n 0.00620273f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_238 B N_A_554_74#_c_664_n 0.0136738f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B_c_244_n N_A_554_74#_c_664_n 0.00440417f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_240 N_B_M1003_g N_A_554_74#_c_666_n 0.0149988f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_241 B N_A_554_74#_c_666_n 0.0967792f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B_c_244_n N_A_554_74#_c_666_n 0.0104341f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_243 N_B_c_244_n N_A_554_74#_c_667_n 0.00232225f $X=6.265 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B_M1003_g N_A_923_74#_c_704_n 0.00509819f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B_M1004_g N_A_923_74#_c_704_n 6.42481e-19 $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B_M1003_g N_A_923_74#_c_705_n 0.00833016f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B_M1004_g N_A_923_74#_c_705_n 0.00775417f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B_M1003_g N_A_923_74#_c_706_n 5.57235e-19 $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B_M1004_g N_A_923_74#_c_706_n 0.00449305f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B_M1016_g N_A_923_74#_c_706_n 0.00448992f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B_M1021_g N_A_923_74#_c_706_n 5.57001e-19 $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B_M1016_g N_A_923_74#_c_707_n 0.00674334f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B_M1021_g N_A_923_74#_c_707_n 0.00792254f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B_M1016_g N_A_923_74#_c_708_n 5.57001e-19 $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B_M1021_g N_A_923_74#_c_708_n 0.00530316f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_M1022_g N_VPWR_c_376_n 0.0168357f $X=8.13 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A_M1013_g N_VPWR_c_379_n 0.00460063f $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A_M1022_g N_VPWR_c_379_n 0.00460063f $X=8.13 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A_M1013_g N_VPWR_c_383_n 0.0178544f $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_M1013_g N_VPWR_c_371_n 0.0090905f $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A_M1022_g N_VPWR_c_371_n 0.00913687f $X=8.13 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_M1013_g N_Y_c_468_n 0.0163499f $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_263 A N_Y_c_468_n 0.0421985f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A_c_310_n N_Y_c_468_n 0.00621082f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_265 N_A_M1002_g N_Y_c_437_n 0.00550051f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_266 A N_Y_c_437_n 0.0171684f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_267 N_A_c_310_n N_Y_c_437_n 0.00221206f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A_M1013_g N_Y_c_445_n 6.96309e-19 $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A_M1022_g N_Y_c_445_n 6.96717e-19 $X=8.13 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A_M1023_g N_Y_c_438_n 0.0220597f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_M1022_g N_Y_c_446_n 0.0198033f $X=8.13 $Y=2.4 $X2=0 $Y2=0
cc_272 A N_Y_c_446_n 0.00454949f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_273 A N_Y_c_485_n 0.0585703f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_274 N_A_c_310_n N_Y_c_485_n 0.00348667f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_275 N_A_M1012_g N_Y_c_439_n 0.0131801f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_M1015_g N_Y_c_439_n 0.0159744f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A_c_308_n N_Y_c_439_n 0.00584045f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_278 A N_Y_c_439_n 0.0691561f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A_c_310_n N_Y_c_439_n 0.00252813f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_280 N_A_M1015_g N_Y_c_440_n 0.0019074f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_M1023_g N_Y_c_440_n 0.0019074f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_M1023_g Y 0.0279739f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_283 A Y 0.0308719f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_284 N_A_M1002_g N_VGND_c_599_n 0.00291649f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_M1012_g N_VGND_c_599_n 0.00291649f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_M1015_g N_VGND_c_599_n 0.00291649f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_M1023_g N_VGND_c_599_n 0.00292759f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_M1002_g N_VGND_c_600_n 0.00359219f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A_M1012_g N_VGND_c_600_n 0.00359121f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_M1015_g N_VGND_c_600_n 0.00360505f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A_M1023_g N_VGND_c_600_n 0.00363199f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A_M1002_g N_A_554_74#_c_664_n 7.32989e-19 $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A_M1015_g N_A_923_74#_c_703_n 0.00855567f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A_M1023_g N_A_923_74#_c_703_n 0.00913165f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A_M1002_g N_A_923_74#_c_708_n 0.00530316f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_M1012_g N_A_923_74#_c_708_n 5.57001e-19 $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_M1002_g N_A_923_74#_c_709_n 0.00792254f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_M1012_g N_A_923_74#_c_709_n 0.00674334f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_M1002_g N_A_923_74#_c_710_n 5.57001e-19 $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_M1012_g N_A_923_74#_c_710_n 0.00448992f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_M1015_g N_A_923_74#_c_710_n 0.00510671f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_M1023_g N_A_923_74#_c_710_n 8.54686e-19 $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_M1015_g N_A_923_74#_c_711_n 9.39838e-19 $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_M1023_g N_A_923_74#_c_711_n 0.00577613f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_305 N_VPWR_c_372_n N_Y_c_442_n 0.0266809f $X=2.485 $Y=2.455 $X2=0 $Y2=0
cc_306 N_VPWR_c_377_n N_Y_c_442_n 0.014549f $X=2.32 $Y=3.33 $X2=0 $Y2=0
cc_307 N_VPWR_c_378_n N_Y_c_442_n 0.0332705f $X=1.65 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_371_n N_Y_c_442_n 0.0119743f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_M1007_d N_Y_c_453_n 0.0065656f $X=2.35 $Y=1.84 $X2=0 $Y2=0
cc_310 N_VPWR_c_372_n N_Y_c_453_n 0.0170259f $X=2.485 $Y=2.455 $X2=0 $Y2=0
cc_311 N_VPWR_c_372_n N_Y_c_443_n 0.0267578f $X=2.485 $Y=2.455 $X2=0 $Y2=0
cc_312 N_VPWR_c_373_n N_Y_c_443_n 0.0271295f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_c_374_n N_Y_c_443_n 0.0297956f $X=4.335 $Y=2.415 $X2=0 $Y2=0
cc_314 N_VPWR_c_371_n N_Y_c_443_n 0.0224555f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_M1018_s N_Y_c_459_n 0.025179f $X=3.63 $Y=1.84 $X2=0 $Y2=0
cc_316 N_VPWR_c_374_n N_Y_c_459_n 0.0634002f $X=4.335 $Y=2.415 $X2=0 $Y2=0
cc_317 N_VPWR_c_374_n N_Y_c_444_n 0.0297956f $X=4.335 $Y=2.415 $X2=0 $Y2=0
cc_318 N_VPWR_c_382_n N_Y_c_444_n 0.0271295f $X=5.45 $Y=2.852 $X2=0 $Y2=0
cc_319 N_VPWR_c_383_n N_Y_c_444_n 0.0298945f $X=7.14 $Y=2.852 $X2=0 $Y2=0
cc_320 N_VPWR_c_371_n N_Y_c_444_n 0.0224555f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_321 N_VPWR_M1017_d N_Y_c_468_n 0.0505215f $X=5.48 $Y=1.84 $X2=0 $Y2=0
cc_322 N_VPWR_c_383_n N_Y_c_468_n 0.127264f $X=7.14 $Y=2.852 $X2=0 $Y2=0
cc_323 N_VPWR_c_376_n N_Y_c_445_n 0.0255792f $X=8.355 $Y=2.415 $X2=0 $Y2=0
cc_324 N_VPWR_c_379_n N_Y_c_445_n 0.0306992f $X=8.19 $Y=3.33 $X2=0 $Y2=0
cc_325 N_VPWR_c_383_n N_Y_c_445_n 0.0285676f $X=7.14 $Y=2.852 $X2=0 $Y2=0
cc_326 N_VPWR_c_371_n N_Y_c_445_n 0.0254101f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_M1022_d N_Y_c_446_n 0.00365063f $X=8.22 $Y=1.84 $X2=0 $Y2=0
cc_328 N_VPWR_c_376_n N_Y_c_446_n 0.0234797f $X=8.355 $Y=2.415 $X2=0 $Y2=0
cc_329 N_VPWR_M1022_d Y 0.00184872f $X=8.22 $Y=1.84 $X2=0 $Y2=0
cc_330 N_Y_c_437_n N_A_554_74#_c_664_n 0.00828756f $X=7.005 $Y=1.005 $X2=0 $Y2=0
cc_331 N_Y_c_439_n N_A_923_74#_M1012_s 0.00179007f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_332 N_Y_c_438_n N_A_923_74#_M1023_s 0.0030137f $X=8.285 $Y=1.005 $X2=0 $Y2=0
cc_333 N_Y_M1015_d N_A_923_74#_c_703_n 0.00526523f $X=7.63 $Y=0.37 $X2=0 $Y2=0
cc_334 N_Y_c_438_n N_A_923_74#_c_703_n 0.00768836f $X=8.285 $Y=1.005 $X2=0 $Y2=0
cc_335 N_Y_c_439_n N_A_923_74#_c_703_n 0.00766981f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_336 N_Y_c_440_n N_A_923_74#_c_703_n 0.0091307f $X=7.945 $Y=0.965 $X2=0 $Y2=0
cc_337 N_Y_M1002_d N_A_923_74#_c_709_n 0.00221561f $X=6.77 $Y=0.37 $X2=0 $Y2=0
cc_338 N_Y_c_437_n N_A_923_74#_c_709_n 0.00894405f $X=7.005 $Y=1.005 $X2=0 $Y2=0
cc_339 N_Y_c_439_n N_A_923_74#_c_709_n 0.0028488f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_340 N_Y_c_439_n N_A_923_74#_c_710_n 0.0167547f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_341 N_Y_c_438_n N_A_923_74#_c_711_n 0.0222972f $X=8.285 $Y=1.005 $X2=0 $Y2=0
cc_342 N_A_27_74#_c_534_n N_VGND_M1006_d 0.00250873f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_343 N_A_27_74#_c_537_n N_VGND_M1014_d 0.00895142f $X=2.245 $Y=1.095 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_533_n N_VGND_c_595_n 0.0191765f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_345 N_A_27_74#_c_534_n N_VGND_c_595_n 0.0209867f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_536_n N_VGND_c_595_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_347 N_A_27_74#_c_536_n N_VGND_c_596_n 0.0145639f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_348 N_A_27_74#_c_536_n N_VGND_c_597_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_349 N_A_27_74#_c_537_n N_VGND_c_597_n 0.0257907f $X=2.245 $Y=1.095 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_538_n N_VGND_c_597_n 0.0175755f $X=2.41 $Y=0.68 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_557_n N_VGND_c_597_n 0.00801271f $X=2.41 $Y=0.965 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_533_n N_VGND_c_598_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_353 N_A_27_74#_c_538_n N_VGND_c_599_n 0.0146502f $X=2.41 $Y=0.68 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_539_n N_VGND_c_599_n 0.0738988f $X=4.2 $Y=0.515 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_533_n N_VGND_c_600_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_536_n N_VGND_c_600_n 0.0119984f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_538_n N_VGND_c_600_n 0.0120674f $X=2.41 $Y=0.68 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_539_n N_VGND_c_600_n 0.0616452f $X=4.2 $Y=0.515 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_539_n N_A_554_74#_M1001_d 0.00172862f $X=4.2 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_360 N_A_27_74#_c_539_n N_A_554_74#_M1011_d 0.00172862f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_M1010_s N_A_554_74#_c_663_n 0.00177318f $X=3.2 $Y=0.37 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_537_n N_A_554_74#_c_663_n 0.00587942f $X=2.245 $Y=1.095
+ $X2=0 $Y2=0
cc_363 N_A_27_74#_c_539_n N_A_554_74#_c_663_n 0.0636023f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_M1020_s N_A_554_74#_c_666_n 0.00311853f $X=4.06 $Y=0.37 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_c_539_n N_A_554_74#_c_666_n 0.0254477f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_539_n N_A_923_74#_c_704_n 0.0234648f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_VGND_c_599_n N_A_923_74#_c_704_n 0.0139208f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_600_n N_A_923_74#_c_704_n 0.0117508f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_599_n N_A_923_74#_c_705_n 0.131762f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_600_n N_A_923_74#_c_705_n 0.111189f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_599_n N_A_923_74#_c_711_n 0.0139208f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_600_n N_A_923_74#_c_711_n 0.0117508f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_373 N_A_554_74#_c_666_n N_A_923_74#_M1003_d 0.00296342f $X=5.095 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_374 N_A_554_74#_c_664_n N_A_923_74#_M1004_d 0.00179007f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
cc_375 N_A_554_74#_c_666_n N_A_923_74#_c_704_n 0.0214875f $X=5.095 $Y=0.965
+ $X2=0 $Y2=0
cc_376 N_A_554_74#_M1003_s N_A_923_74#_c_705_n 0.00221951f $X=5.05 $Y=0.37 $X2=0
+ $Y2=0
cc_377 N_A_554_74#_c_664_n N_A_923_74#_c_705_n 0.00474257f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
cc_378 N_A_554_74#_c_666_n N_A_923_74#_c_705_n 0.00476112f $X=5.095 $Y=0.965
+ $X2=0 $Y2=0
cc_379 N_A_554_74#_c_667_n N_A_923_74#_c_705_n 0.00797735f $X=5.285 $Y=0.965
+ $X2=0 $Y2=0
cc_380 N_A_554_74#_c_664_n N_A_923_74#_c_706_n 0.0167547f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
cc_381 N_A_554_74#_M1016_s N_A_923_74#_c_707_n 0.00221561f $X=5.91 $Y=0.37 $X2=0
+ $Y2=0
cc_382 N_A_554_74#_c_664_n N_A_923_74#_c_707_n 0.0117928f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0

* File: sky130_fd_sc_ms__ebufn_1.pxi.spice
* Created: Fri Aug 28 17:31:45 2020
* 
x_PM_SKY130_FD_SC_MS__EBUFN_1%TE_B N_TE_B_M1000_g N_TE_B_M1007_g N_TE_B_c_72_n
+ N_TE_B_c_73_n N_TE_B_c_79_n N_TE_B_M1001_g N_TE_B_c_80_n N_TE_B_c_81_n
+ N_TE_B_c_82_n N_TE_B_c_106_p N_TE_B_c_83_n N_TE_B_c_84_n TE_B N_TE_B_c_75_n
+ PM_SKY130_FD_SC_MS__EBUFN_1%TE_B
x_PM_SKY130_FD_SC_MS__EBUFN_1%A N_A_M1002_g N_A_M1003_g N_A_c_164_n A A
+ N_A_c_166_n PM_SKY130_FD_SC_MS__EBUFN_1%A
x_PM_SKY130_FD_SC_MS__EBUFN_1%A_27_404# N_A_27_404#_M1007_s N_A_27_404#_M1000_s
+ N_A_27_404#_c_201_n N_A_27_404#_c_202_n N_A_27_404#_M1005_g
+ N_A_27_404#_c_203_n N_A_27_404#_c_204_n N_A_27_404#_c_209_n
+ N_A_27_404#_c_205_n N_A_27_404#_c_206_n N_A_27_404#_c_207_n
+ N_A_27_404#_c_208_n PM_SKY130_FD_SC_MS__EBUFN_1%A_27_404#
x_PM_SKY130_FD_SC_MS__EBUFN_1%A_229_74# N_A_229_74#_M1002_d N_A_229_74#_M1003_d
+ N_A_229_74#_M1006_g N_A_229_74#_M1004_g N_A_229_74#_c_264_n
+ N_A_229_74#_c_272_n N_A_229_74#_c_265_n N_A_229_74#_c_266_n
+ N_A_229_74#_c_273_n N_A_229_74#_c_267_n N_A_229_74#_c_268_n
+ N_A_229_74#_c_269_n N_A_229_74#_c_274_n N_A_229_74#_c_275_n
+ N_A_229_74#_c_276_n N_A_229_74#_c_270_n PM_SKY130_FD_SC_MS__EBUFN_1%A_229_74#
x_PM_SKY130_FD_SC_MS__EBUFN_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_s N_VPWR_c_358_n
+ N_VPWR_c_359_n VPWR N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_357_n
+ N_VPWR_c_363_n N_VPWR_c_364_n PM_SKY130_FD_SC_MS__EBUFN_1%VPWR
x_PM_SKY130_FD_SC_MS__EBUFN_1%Z N_Z_M1006_d N_Z_M1004_d N_Z_c_406_n N_Z_c_407_n
+ N_Z_c_404_n Z Z N_Z_c_405_n PM_SKY130_FD_SC_MS__EBUFN_1%Z
x_PM_SKY130_FD_SC_MS__EBUFN_1%VGND N_VGND_M1007_d N_VGND_M1005_s N_VGND_c_431_n
+ N_VGND_c_432_n VGND N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ N_VGND_c_436_n N_VGND_c_437_n PM_SKY130_FD_SC_MS__EBUFN_1%VGND
cc_1 VNB N_TE_B_M1007_g 0.0507161f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.645
cc_2 VNB N_TE_B_c_72_n 0.0118248f $X=-0.19 $Y=-0.245 $X2=2.665 $Y2=1.69
cc_3 VNB N_TE_B_c_73_n 0.0043072f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.69
cc_4 VNB TE_B 0.00341842f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_TE_B_c_75_n 0.0168752f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_6 VNB N_A_M1002_g 0.0580975f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.44
cc_7 VNB N_A_c_164_n 0.00848377f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=2.34
cc_8 VNB A 0.00358455f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.69
cc_9 VNB N_A_c_166_n 0.0229517f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.505
cc_10 VNB N_A_27_404#_c_201_n 0.0395168f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.645
cc_11 VNB N_A_27_404#_c_202_n 0.0172236f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=1.765
cc_12 VNB N_A_27_404#_c_203_n 0.0365396f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_13 VNB N_A_27_404#_c_204_n 0.0118865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_404#_c_205_n 0.0162952f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.505
cc_15 VNB N_A_27_404#_c_206_n 9.95647e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_A_27_404#_c_207_n 0.0271006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_404#_c_208_n 0.0424548f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_18 VNB N_A_229_74#_M1006_g 0.0284822f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=1.765
cc_19 VNB N_A_229_74#_M1004_g 5.55278e-19 $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=1.765
cc_20 VNB N_A_229_74#_c_264_n 0.0139199f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.34
cc_21 VNB N_A_229_74#_c_265_n 0.029099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_229_74#_c_266_n 0.00347683f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.465
cc_23 VNB N_A_229_74#_c_267_n 0.00135177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_229_74#_c_268_n 0.00449629f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_25 VNB N_A_229_74#_c_269_n 0.0363898f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.5
cc_26 VNB N_A_229_74#_c_270_n 0.0147135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_357_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_28 VNB N_Z_c_404_n 0.0252276f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_29 VNB N_Z_c_405_n 0.0503455f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.505
cc_30 VNB N_VGND_c_431_n 0.00944084f $X=-0.19 $Y=-0.245 $X2=2.665 $Y2=1.69
cc_31 VNB N_VGND_c_432_n 0.0203845f $X=-0.19 $Y=-0.245 $X2=2.755 $Y2=2.4
cc_32 VNB N_VGND_c_433_n 0.042784f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.42
cc_33 VNB N_VGND_c_434_n 0.033384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_435_n 0.24203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_436_n 0.0270337f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.665
cc_36 VNB N_VGND_c_437_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_37 VPB N_TE_B_M1000_g 0.030166f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.44
cc_38 VPB N_TE_B_c_72_n 0.0167129f $X=-0.19 $Y=1.66 $X2=2.665 $Y2=1.69
cc_39 VPB N_TE_B_c_73_n 0.00373927f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.69
cc_40 VPB N_TE_B_c_79_n 0.0175945f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_41 VPB N_TE_B_c_80_n 0.0393321f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.34
cc_42 VPB N_TE_B_c_81_n 0.00339826f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.42
cc_43 VPB N_TE_B_c_82_n 0.00956627f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.505
cc_44 VPB N_TE_B_c_83_n 0.00739652f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_45 VPB N_TE_B_c_84_n 0.0719223f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_46 VPB TE_B 0.00363527f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_47 VPB N_TE_B_c_75_n 0.0167615f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.665
cc_48 VPB N_A_M1003_g 0.0313773f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.645
cc_49 VPB N_A_c_164_n 0.00846445f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=2.34
cc_50 VPB A 0.00240167f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.69
cc_51 VPB N_A_c_166_n 0.022161f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_52 VPB N_A_27_404#_c_209_n 0.0406343f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.465
cc_53 VPB N_A_27_404#_c_205_n 0.0158855f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_54 VPB N_A_229_74#_M1004_g 0.0289004f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=1.765
cc_55 VPB N_A_229_74#_c_272_n 0.00334574f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.42
cc_56 VPB N_A_229_74#_c_273_n 0.00833716f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.505
cc_57 VPB N_A_229_74#_c_274_n 0.0039456f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_58 VPB N_A_229_74#_c_275_n 0.00831023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_229_74#_c_276_n 0.00604866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_229_74#_c_270_n 0.00163048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_358_n 0.016053f $X=-0.19 $Y=1.66 $X2=2.665 $Y2=1.69
cc_62 VPB N_VPWR_c_359_n 0.0151141f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_63 VPB N_VPWR_c_360_n 0.0380943f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.505
cc_64 VPB N_VPWR_c_361_n 0.0343749f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.665
cc_65 VPB N_VPWR_c_357_n 0.0861643f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.665
cc_66 VPB N_VPWR_c_363_n 0.02685f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.83
cc_67 VPB N_VPWR_c_364_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_Z_c_406_n 0.0466392f $X=-0.19 $Y=1.66 $X2=2.12 $Y2=1.765
cc_69 VPB N_Z_c_407_n 0.0201226f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_70 VPB N_Z_c_404_n 0.007785f $X=-0.19 $Y=1.66 $X2=2.755 $Y2=2.4
cc_71 N_TE_B_M1007_g N_A_M1002_g 0.0347876f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_72 N_TE_B_M1000_g N_A_M1003_g 0.0238284f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_73 N_TE_B_c_81_n N_A_M1003_g 0.00955527f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_74 N_TE_B_c_82_n N_A_M1003_g 0.0174187f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_75 N_TE_B_c_83_n N_A_M1003_g 0.00230471f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_76 N_TE_B_c_84_n N_A_M1003_g 0.0109557f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_77 TE_B N_A_c_164_n 0.00231785f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_78 N_TE_B_c_75_n N_A_c_164_n 0.018318f $X=0.59 $Y=1.665 $X2=0 $Y2=0
cc_79 N_TE_B_c_73_n A 0.00172831f $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_80 N_TE_B_c_82_n A 0.00423629f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_81 TE_B A 0.0279811f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_82 N_TE_B_c_75_n A 3.47969e-19 $X=0.59 $Y=1.665 $X2=0 $Y2=0
cc_83 N_TE_B_c_73_n N_A_c_166_n 0.00676649f $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_84 N_TE_B_c_72_n N_A_27_404#_c_201_n 0.0258375f $X=2.665 $Y=1.69 $X2=0 $Y2=0
cc_85 N_TE_B_M1007_g N_A_27_404#_c_203_n 0.0112033f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_86 TE_B N_A_27_404#_c_204_n 0.00843991f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_87 N_TE_B_c_75_n N_A_27_404#_c_204_n 0.0011791f $X=0.59 $Y=1.665 $X2=0 $Y2=0
cc_88 N_TE_B_M1000_g N_A_27_404#_c_209_n 0.0176045f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_89 N_TE_B_c_81_n N_A_27_404#_c_209_n 0.0255665f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_90 N_TE_B_c_106_p N_A_27_404#_c_209_n 0.0115775f $X=0.835 $Y=2.505 $X2=0
+ $Y2=0
cc_91 TE_B N_A_27_404#_c_209_n 0.00144434f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_92 N_TE_B_M1007_g N_A_27_404#_c_205_n 0.00389989f $X=0.62 $Y=0.645 $X2=0
+ $Y2=0
cc_93 N_TE_B_c_81_n N_A_27_404#_c_205_n 0.00487261f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_94 TE_B N_A_27_404#_c_205_n 0.0252195f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_95 N_TE_B_c_75_n N_A_27_404#_c_205_n 0.010238f $X=0.59 $Y=1.665 $X2=0 $Y2=0
cc_96 N_TE_B_c_73_n N_A_27_404#_c_206_n 5.97257e-19 $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_97 N_TE_B_M1007_g N_A_27_404#_c_207_n 0.0169119f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_98 TE_B N_A_27_404#_c_207_n 0.0224553f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_99 N_TE_B_c_75_n N_A_27_404#_c_207_n 5.1855e-19 $X=0.59 $Y=1.665 $X2=0 $Y2=0
cc_100 N_TE_B_c_73_n N_A_27_404#_c_208_n 0.0258375f $X=2.195 $Y=1.69 $X2=0 $Y2=0
cc_101 N_TE_B_c_82_n N_A_229_74#_M1003_d 0.00782008f $X=1.865 $Y=2.505 $X2=0
+ $Y2=0
cc_102 N_TE_B_c_79_n N_A_229_74#_M1004_g 0.0378105f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_81_n N_A_229_74#_c_272_n 0.0110923f $X=0.75 $Y=2.42 $X2=0 $Y2=0
cc_104 N_TE_B_c_82_n N_A_229_74#_c_272_n 0.0341849f $X=1.865 $Y=2.505 $X2=0
+ $Y2=0
cc_105 N_TE_B_c_80_n N_A_229_74#_c_273_n 0.00126228f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_106 N_TE_B_c_82_n N_A_229_74#_c_273_n 0.00972763f $X=1.865 $Y=2.505 $X2=0
+ $Y2=0
cc_107 N_TE_B_c_83_n N_A_229_74#_c_273_n 0.0079822f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_108 N_TE_B_c_84_n N_A_229_74#_c_273_n 6.96394e-19 $X=2.03 $Y=2.505 $X2=0
+ $Y2=0
cc_109 N_TE_B_c_72_n N_A_229_74#_c_269_n 0.0378105f $X=2.665 $Y=1.69 $X2=0 $Y2=0
cc_110 N_TE_B_c_80_n N_A_229_74#_c_274_n 0.00163127f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_111 N_TE_B_c_73_n N_A_229_74#_c_275_n 0.00203925f $X=2.195 $Y=1.69 $X2=0
+ $Y2=0
cc_112 N_TE_B_c_79_n N_A_229_74#_c_275_n 6.12337e-19 $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_TE_B_c_80_n N_A_229_74#_c_275_n 0.014524f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_114 N_TE_B_c_83_n N_A_229_74#_c_275_n 0.0141324f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_115 N_TE_B_c_84_n N_A_229_74#_c_275_n 5.95224e-19 $X=2.03 $Y=2.505 $X2=0
+ $Y2=0
cc_116 N_TE_B_c_72_n N_A_229_74#_c_276_n 0.00771499f $X=2.665 $Y=1.69 $X2=0
+ $Y2=0
cc_117 N_TE_B_c_73_n N_A_229_74#_c_276_n 0.00114693f $X=2.195 $Y=1.69 $X2=0
+ $Y2=0
cc_118 N_TE_B_c_80_n N_A_229_74#_c_276_n 0.00437206f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_119 N_TE_B_c_83_n N_A_229_74#_c_276_n 0.00203003f $X=2.03 $Y=2.505 $X2=0
+ $Y2=0
cc_120 N_TE_B_c_72_n N_A_229_74#_c_270_n 0.0144694f $X=2.665 $Y=1.69 $X2=0 $Y2=0
cc_121 N_TE_B_c_79_n N_A_229_74#_c_270_n 0.012865f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_122 N_TE_B_c_81_n N_VPWR_M1000_d 0.011927f $X=0.75 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_123 N_TE_B_c_82_n N_VPWR_M1000_d 0.00706944f $X=1.865 $Y=2.505 $X2=-0.19
+ $Y2=-0.245
cc_124 N_TE_B_c_106_p N_VPWR_M1000_d 0.00501257f $X=0.835 $Y=2.505 $X2=-0.19
+ $Y2=-0.245
cc_125 N_TE_B_M1000_g N_VPWR_c_358_n 0.00407444f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_126 N_TE_B_c_82_n N_VPWR_c_358_n 0.0111946f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_127 N_TE_B_c_106_p N_VPWR_c_358_n 0.0146637f $X=0.835 $Y=2.505 $X2=0 $Y2=0
cc_128 N_TE_B_c_72_n N_VPWR_c_359_n 0.0012721f $X=2.665 $Y=1.69 $X2=0 $Y2=0
cc_129 N_TE_B_c_79_n N_VPWR_c_359_n 0.0225918f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_130 N_TE_B_c_80_n N_VPWR_c_359_n 0.00440568f $X=2.03 $Y=2.34 $X2=0 $Y2=0
cc_131 N_TE_B_c_83_n N_VPWR_c_359_n 0.0537867f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_132 N_TE_B_c_84_n N_VPWR_c_359_n 0.00470851f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_133 N_TE_B_c_82_n N_VPWR_c_360_n 0.011737f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_134 N_TE_B_c_83_n N_VPWR_c_360_n 0.015584f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_135 N_TE_B_c_84_n N_VPWR_c_360_n 0.00192529f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_136 N_TE_B_c_79_n N_VPWR_c_361_n 0.00460063f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_137 N_TE_B_M1000_g N_VPWR_c_357_n 0.00617325f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_138 N_TE_B_c_79_n N_VPWR_c_357_n 0.00908371f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_139 N_TE_B_c_82_n N_VPWR_c_357_n 0.0236758f $X=1.865 $Y=2.505 $X2=0 $Y2=0
cc_140 N_TE_B_c_106_p N_VPWR_c_357_n 7.17789e-19 $X=0.835 $Y=2.505 $X2=0 $Y2=0
cc_141 N_TE_B_c_83_n N_VPWR_c_357_n 0.0120766f $X=2.03 $Y=2.505 $X2=0 $Y2=0
cc_142 N_TE_B_M1000_g N_VPWR_c_363_n 0.00582418f $X=0.505 $Y=2.44 $X2=0 $Y2=0
cc_143 N_TE_B_c_79_n N_Z_c_407_n 0.00348457f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_144 N_TE_B_M1007_g N_VGND_c_431_n 0.00408774f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_145 N_TE_B_M1007_g N_VGND_c_435_n 0.00911508f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_146 N_TE_B_M1007_g N_VGND_c_436_n 0.00461464f $X=0.62 $Y=0.645 $X2=0 $Y2=0
cc_147 N_A_M1003_g N_A_27_404#_c_209_n 8.92556e-19 $X=1.125 $Y=2.44 $X2=0 $Y2=0
cc_148 N_A_M1002_g N_A_27_404#_c_207_n 0.0175221f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_149 N_A_c_164_n N_A_27_404#_c_207_n 0.0120594f $X=1.105 $Y=1.665 $X2=0 $Y2=0
cc_150 A N_A_27_404#_c_207_n 0.0568065f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A_M1003_g N_A_229_74#_c_272_n 0.00515596f $X=1.125 $Y=2.44 $X2=0 $Y2=0
cc_152 A N_A_229_74#_c_272_n 0.0472651f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A_c_166_n N_A_229_74#_c_272_n 0.0103846f $X=1.51 $Y=1.665 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_A_229_74#_c_266_n 0.00357394f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_155 A N_A_229_74#_c_275_n 0.0100487f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A_c_166_n N_A_229_74#_c_275_n 2.98913e-19 $X=1.51 $Y=1.665 $X2=0 $Y2=0
cc_157 A N_A_229_74#_c_270_n 0.00704617f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_VPWR_c_358_n 0.00443659f $X=1.125 $Y=2.44 $X2=0 $Y2=0
cc_159 N_A_M1003_g N_VPWR_c_360_n 0.00477315f $X=1.125 $Y=2.44 $X2=0 $Y2=0
cc_160 N_A_M1003_g N_VPWR_c_357_n 0.00617325f $X=1.125 $Y=2.44 $X2=0 $Y2=0
cc_161 N_A_M1002_g N_VGND_c_431_n 0.00405933f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_162 N_A_M1002_g N_VGND_c_433_n 0.00461464f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_163 N_A_M1002_g N_VGND_c_435_n 0.00912604f $X=1.07 $Y=0.645 $X2=0 $Y2=0
cc_164 N_A_27_404#_c_202_n N_A_229_74#_M1006_g 0.0303584f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_165 N_A_27_404#_c_201_n N_A_229_74#_c_265_n 0.00892394f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_166 N_A_27_404#_c_207_n N_A_229_74#_c_265_n 0.0553447f $X=1.87 $Y=1.245 $X2=0
+ $Y2=0
cc_167 N_A_27_404#_c_208_n N_A_229_74#_c_265_n 0.00808505f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_168 N_A_27_404#_c_203_n N_A_229_74#_c_266_n 0.00210758f $X=0.405 $Y=0.645
+ $X2=0 $Y2=0
cc_169 N_A_27_404#_c_207_n N_A_229_74#_c_266_n 0.0243942f $X=1.87 $Y=1.245 $X2=0
+ $Y2=0
cc_170 N_A_27_404#_c_206_n N_A_229_74#_c_273_n 0.00244148f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_171 N_A_27_404#_c_208_n N_A_229_74#_c_273_n 0.0015619f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_172 N_A_27_404#_c_201_n N_A_229_74#_c_267_n 0.0117554f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_173 N_A_27_404#_c_202_n N_A_229_74#_c_267_n 0.00393509f $X=2.77 $Y=1.185
+ $X2=0 $Y2=0
cc_174 N_A_27_404#_c_206_n N_A_229_74#_c_267_n 0.00939079f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_175 N_A_27_404#_c_208_n N_A_229_74#_c_267_n 0.00179597f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_176 N_A_27_404#_c_201_n N_A_229_74#_c_269_n 0.0303584f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_177 N_A_27_404#_c_206_n N_A_229_74#_c_275_n 0.00701624f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_178 N_A_27_404#_c_208_n N_A_229_74#_c_275_n 0.00200399f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_179 N_A_27_404#_c_206_n N_A_229_74#_c_276_n 0.00236052f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_180 N_A_27_404#_c_208_n N_A_229_74#_c_276_n 0.00164906f $X=2.2 $Y=1.24 $X2=0
+ $Y2=0
cc_181 N_A_27_404#_c_201_n N_A_229_74#_c_270_n 0.0207665f $X=2.695 $Y=1.295
+ $X2=0 $Y2=0
cc_182 N_A_27_404#_c_206_n N_A_229_74#_c_270_n 0.00102519f $X=2.035 $Y=1.24
+ $X2=0 $Y2=0
cc_183 N_A_27_404#_c_209_n N_VPWR_c_358_n 0.00462123f $X=0.28 $Y=2.165 $X2=0
+ $Y2=0
cc_184 N_A_27_404#_c_209_n N_VPWR_c_357_n 0.0123694f $X=0.28 $Y=2.165 $X2=0
+ $Y2=0
cc_185 N_A_27_404#_c_209_n N_VPWR_c_363_n 0.0112883f $X=0.28 $Y=2.165 $X2=0
+ $Y2=0
cc_186 N_A_27_404#_c_202_n N_Z_c_405_n 0.00258266f $X=2.77 $Y=1.185 $X2=0 $Y2=0
cc_187 N_A_27_404#_c_207_n N_VGND_c_431_n 0.0126908f $X=1.87 $Y=1.245 $X2=0
+ $Y2=0
cc_188 N_A_27_404#_c_201_n N_VGND_c_432_n 8.1259e-19 $X=2.695 $Y=1.295 $X2=0
+ $Y2=0
cc_189 N_A_27_404#_c_202_n N_VGND_c_432_n 0.0110763f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_190 N_A_27_404#_c_202_n N_VGND_c_434_n 0.00383152f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_191 N_A_27_404#_c_202_n N_VGND_c_435_n 0.0075725f $X=2.77 $Y=1.185 $X2=0
+ $Y2=0
cc_192 N_A_27_404#_c_203_n N_VGND_c_435_n 0.0152899f $X=0.405 $Y=0.645 $X2=0
+ $Y2=0
cc_193 N_A_27_404#_c_203_n N_VGND_c_436_n 0.0129976f $X=0.405 $Y=0.645 $X2=0
+ $Y2=0
cc_194 N_A_229_74#_c_276_n N_VPWR_M1001_s 7.86634e-19 $X=2.46 $Y=1.6 $X2=0 $Y2=0
cc_195 N_A_229_74#_c_270_n N_VPWR_M1001_s 0.00163196f $X=3.065 $Y=1.6 $X2=0
+ $Y2=0
cc_196 N_A_229_74#_M1004_g N_VPWR_c_359_n 0.00318011f $X=3.175 $Y=2.4 $X2=0
+ $Y2=0
cc_197 N_A_229_74#_c_274_n N_VPWR_c_359_n 0.00258243f $X=1.695 $Y=2.125 $X2=0
+ $Y2=0
cc_198 N_A_229_74#_c_275_n N_VPWR_c_359_n 0.00723556f $X=2.05 $Y=1.795 $X2=0
+ $Y2=0
cc_199 N_A_229_74#_c_276_n N_VPWR_c_359_n 0.0231278f $X=2.46 $Y=1.6 $X2=0 $Y2=0
cc_200 N_A_229_74#_M1004_g N_VPWR_c_361_n 0.005209f $X=3.175 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_229_74#_M1004_g N_VPWR_c_357_n 0.00987364f $X=3.175 $Y=2.4 $X2=0
+ $Y2=0
cc_202 N_A_229_74#_c_270_n A_569_368# 0.0055509f $X=3.065 $Y=1.6 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_229_74#_M1004_g N_Z_c_406_n 0.0184881f $X=3.175 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_229_74#_M1004_g N_Z_c_407_n 0.00539711f $X=3.175 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_229_74#_c_268_n N_Z_c_407_n 0.0149649f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_206 N_A_229_74#_c_269_n N_Z_c_407_n 0.00349435f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_207 N_A_229_74#_c_270_n N_Z_c_407_n 0.00327027f $X=3.065 $Y=1.6 $X2=0 $Y2=0
cc_208 N_A_229_74#_M1006_g N_Z_c_404_n 0.00394404f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_229_74#_M1004_g N_Z_c_404_n 0.00231906f $X=3.175 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_229_74#_c_268_n N_Z_c_404_n 0.0262124f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_211 N_A_229_74#_c_269_n N_Z_c_404_n 0.00231223f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_212 N_A_229_74#_c_270_n N_Z_c_404_n 0.00459991f $X=3.065 $Y=1.6 $X2=0 $Y2=0
cc_213 N_A_229_74#_M1006_g N_Z_c_405_n 0.0164306f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_229_74#_c_267_n N_Z_c_405_n 0.00263651f $X=2.56 $Y=1.32 $X2=0 $Y2=0
cc_215 N_A_229_74#_c_268_n N_Z_c_405_n 0.0157141f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_216 N_A_229_74#_c_269_n N_Z_c_405_n 0.0042671f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_217 N_A_229_74#_c_265_n N_VGND_M1005_s 0.00506875f $X=2.46 $Y=0.895 $X2=0
+ $Y2=0
cc_218 N_A_229_74#_c_267_n N_VGND_M1005_s 0.00433646f $X=2.56 $Y=1.32 $X2=0
+ $Y2=0
cc_219 N_A_229_74#_M1006_g N_VGND_c_432_n 0.00138195f $X=3.16 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_229_74#_c_265_n N_VGND_c_432_n 0.0207988f $X=2.46 $Y=0.895 $X2=0
+ $Y2=0
cc_221 N_A_229_74#_c_264_n N_VGND_c_433_n 0.00811823f $X=1.285 $Y=0.645 $X2=0
+ $Y2=0
cc_222 N_A_229_74#_M1006_g N_VGND_c_434_n 0.00434272f $X=3.16 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_229_74#_M1006_g N_VGND_c_435_n 0.00825123f $X=3.16 $Y=0.74 $X2=0
+ $Y2=0
cc_224 N_A_229_74#_c_264_n N_VGND_c_435_n 0.0100099f $X=1.285 $Y=0.645 $X2=0
+ $Y2=0
cc_225 N_A_229_74#_c_265_n N_VGND_c_435_n 0.0343415f $X=2.46 $Y=0.895 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_361_n N_Z_c_406_n 0.0230269f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_227 N_VPWR_c_357_n N_Z_c_406_n 0.0189916f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_228 N_VPWR_c_359_n N_Z_c_407_n 0.0280012f $X=2.53 $Y=2.135 $X2=0 $Y2=0
cc_229 N_Z_c_405_n N_VGND_c_432_n 0.00955365f $X=3.375 $Y=0.515 $X2=0 $Y2=0
cc_230 N_Z_c_405_n N_VGND_c_434_n 0.0241574f $X=3.375 $Y=0.515 $X2=0 $Y2=0
cc_231 N_Z_c_405_n N_VGND_c_435_n 0.019939f $X=3.375 $Y=0.515 $X2=0 $Y2=0

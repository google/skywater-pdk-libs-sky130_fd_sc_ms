* File: sky130_fd_sc_ms__a32o_4.pex.spice
* Created: Fri Aug 28 17:08:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A32O_4%A_83_283# 1 2 3 4 15 17 19 20 22 25 29 33 37
+ 41 43 52 53 54 57 60 63 64 66 71 73 85
c176 73 0 1.2831e-19 $X=5.965 $Y=1.1
c177 71 0 7.5232e-20 $X=4.19 $Y=2.115
c178 64 0 7.32746e-20 $X=4.055 $Y=1.195
c179 63 0 1.79774e-20 $X=5.8 $Y=1.195
r180 79 80 2.02521 $w=3.57e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.472
+ $X2=0.955 $Y2=1.472
r181 78 79 58.7311 $w=3.57e-07 $l=4.35e-07 $layer=POLY_cond $X=0.505 $Y=1.472
+ $X2=0.94 $Y2=1.472
r182 77 78 1.35014 $w=3.57e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.472
+ $X2=0.505 $Y2=1.472
r183 73 75 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.965 $Y=1.1
+ $X2=5.965 $Y2=1.195
r184 68 69 26.5367 $w=1.77e-07 $l=3.85e-07 $layer=LI1_cond $X=3.585 $Y=1.187
+ $X2=3.97 $Y2=1.187
r185 64 69 5.85876 $w=1.77e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.055 $Y=1.195
+ $X2=3.97 $Y2=1.187
r186 63 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=1.195
+ $X2=5.965 $Y2=1.195
r187 63 64 113.845 $w=1.68e-07 $l=1.745e-06 $layer=LI1_cond $X=5.8 $Y=1.195
+ $X2=4.055 $Y2=1.195
r188 60 71 3.70735 $w=2.5e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.97 $Y=1.95
+ $X2=4.12 $Y2=2.035
r189 59 69 0.961343 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=3.97 $Y=1.28
+ $X2=3.97 $Y2=1.187
r190 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.97 $Y=1.28
+ $X2=3.97 $Y2=1.95
r191 58 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=2.035
+ $X2=3.19 $Y2=2.035
r192 57 71 2.76166 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.885 $Y=2.035
+ $X2=4.12 $Y2=2.035
r193 57 58 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.885 $Y=2.035
+ $X2=3.355 $Y2=2.035
r194 53 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=3.19 $Y2=2.035
r195 53 54 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=2.185 $Y2=2.035
r196 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.1 $Y=1.95
+ $X2=2.185 $Y2=2.035
r197 51 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.1 $Y=1.68 $X2=2.1
+ $Y2=1.95
r198 50 85 10.126 $w=3.57e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.472
+ $X2=1.905 $Y2=1.472
r199 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.515 $X2=1.83 $Y2=1.515
r200 46 82 41.1793 $w=3.57e-07 $l=3.05e-07 $layer=POLY_cond $X=1.15 $Y=1.472
+ $X2=1.455 $Y2=1.472
r201 46 80 26.3277 $w=3.57e-07 $l=1.95e-07 $layer=POLY_cond $X=1.15 $Y=1.472
+ $X2=0.955 $Y2=1.472
r202 45 49 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.15 $Y=1.515
+ $X2=1.83 $Y2=1.515
r203 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.515 $X2=1.15 $Y2=1.515
r204 43 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=1.515
+ $X2=2.1 $Y2=1.68
r205 43 49 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.015 $Y=1.515
+ $X2=1.83 $Y2=1.515
r206 39 85 6.07563 $w=3.57e-07 $l=4.5e-08 $layer=POLY_cond $X=1.95 $Y=1.472
+ $X2=1.905 $Y2=1.472
r207 39 41 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.95 $Y=1.35
+ $X2=1.95 $Y2=0.82
r208 35 85 18.7718 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=1.472
r209 35 37 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=2.4
r210 31 50 41.8543 $w=3.57e-07 $l=3.1e-07 $layer=POLY_cond $X=1.52 $Y=1.472
+ $X2=1.83 $Y2=1.472
r211 31 82 8.77591 $w=3.57e-07 $l=6.5e-08 $layer=POLY_cond $X=1.52 $Y=1.472
+ $X2=1.455 $Y2=1.472
r212 31 33 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.52 $Y=1.35
+ $X2=1.52 $Y2=0.82
r213 27 82 18.7718 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.472
r214 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r215 23 80 18.7718 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.472
r216 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r217 20 79 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=1.265
+ $X2=0.94 $Y2=1.472
r218 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.94 $Y=1.265
+ $X2=0.94 $Y2=0.82
r219 17 77 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.265
+ $X2=0.495 $Y2=1.472
r220 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.265
+ $X2=0.495 $Y2=0.82
r221 13 78 18.7718 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.472
r222 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
r223 4 71 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=4.005
+ $Y=1.96 $X2=4.19 $Y2=2.115
r224 3 66 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=3.005
+ $Y=1.96 $X2=3.19 $Y2=2.115
r225 2 73 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.825
+ $Y=0.61 $X2=5.965 $Y2=1.1
r226 1 68 182 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.55 $X2=3.585 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%B2 3 7 9 11 12 14 15 18 20 23 27 31 32 33 39
+ 46 51 53
c107 51 0 6.39601e-20 $X=4.415 $Y=0.42
c108 33 0 1.33336e-19 $X=4.25 $Y=0.34
c109 20 0 1.0936e-19 $X=4.81 $Y=1.08
c110 12 0 7.57553e-20 $X=4.415 $Y=1.855
c111 9 0 7.32746e-20 $X=4.23 $Y=0.585
r112 45 46 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.86 $Y=1.615
+ $X2=2.915 $Y2=1.615
r113 42 45 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.67 $Y=1.615
+ $X2=2.86 $Y2=1.615
r114 39 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=1.615
+ $X2=2.67 $Y2=1.45
r115 39 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.615 $X2=2.67 $Y2=1.615
r116 37 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=0.42
+ $X2=4.415 $Y2=0.42
r117 37 48 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.25 $Y=0.42 $X2=4.23
+ $Y2=0.42
r118 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=0.42 $X2=4.25 $Y2=0.42
r119 33 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.25 $Y=0.34 $X2=4.25
+ $Y2=0.42
r120 31 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=4.25 $Y2=0.34
r121 31 32 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=2.74 $Y2=0.34
r122 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.74 $Y2=0.34
r123 29 53 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.655 $Y2=1.45
r124 25 27 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=4.705 $Y=1.155
+ $X2=4.81 $Y2=1.155
r125 20 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.81 $Y=1.08
+ $X2=4.81 $Y2=1.155
r126 19 20 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.81 $Y=0.585
+ $X2=4.81 $Y2=1.08
r127 18 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=1.705
+ $X2=4.705 $Y2=1.78
r128 17 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.705 $Y=1.23
+ $X2=4.705 $Y2=1.155
r129 17 18 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.705 $Y=1.23
+ $X2=4.705 $Y2=1.705
r130 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.735 $Y=0.51
+ $X2=4.81 $Y2=0.585
r131 15 51 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.735 $Y=0.51
+ $X2=4.415 $Y2=0.51
r132 12 23 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.415 $Y=1.78
+ $X2=4.705 $Y2=1.78
r133 12 14 162.006 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=4.415 $Y=1.855
+ $X2=4.415 $Y2=2.46
r134 9 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=0.585
+ $X2=4.23 $Y2=0.42
r135 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.23 $Y=0.585
+ $X2=4.23 $Y2=1.015
r136 5 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.78
+ $X2=2.915 $Y2=1.615
r137 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.915 $Y=1.78
+ $X2=2.915 $Y2=2.46
r138 1 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.86 $Y=1.45
+ $X2=2.86 $Y2=1.615
r139 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.86 $Y=1.45 $X2=2.86
+ $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%B1 3 5 7 8 10 11 13 14 15 23
c56 23 0 8.37829e-20 $X=3.8 $Y=1.652
c57 8 0 1.33336e-19 $X=3.8 $Y=1.45
r58 21 23 45.6942 $w=3.27e-07 $l=3.1e-07 $layer=POLY_cond $X=3.49 $Y=1.652
+ $X2=3.8 $Y2=1.652
r59 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.615 $X2=3.49 $Y2=1.615
r60 19 21 11.055 $w=3.27e-07 $l=7.5e-08 $layer=POLY_cond $X=3.415 $Y=1.652
+ $X2=3.49 $Y2=1.652
r61 15 22 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.6 $Y=1.615
+ $X2=3.49 $Y2=1.615
r62 14 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.615
+ $X2=3.49 $Y2=1.615
r63 11 23 16.9511 $w=3.27e-07 $l=2.54075e-07 $layer=POLY_cond $X=3.915 $Y=1.855
+ $X2=3.8 $Y2=1.652
r64 11 13 162.006 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=3.915 $Y=1.855
+ $X2=3.915 $Y2=2.46
r65 8 23 21.0057 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=3.8 $Y=1.45 $X2=3.8
+ $Y2=1.652
r66 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.8 $Y=1.45 $X2=3.8
+ $Y2=1.015
r67 5 19 16.7191 $w=1.8e-07 $l=2.03e-07 $layer=POLY_cond $X=3.415 $Y=1.855
+ $X2=3.415 $Y2=1.652
r68 5 7 162.006 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=3.415 $Y=1.855
+ $X2=3.415 $Y2=2.46
r69 1 19 18.4251 $w=3.27e-07 $l=2.5701e-07 $layer=POLY_cond $X=3.29 $Y=1.45
+ $X2=3.415 $Y2=1.652
r70 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.29 $Y=1.45 $X2=3.29
+ $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A2 3 7 11 15 17 18 19 20 22 23 30 31 33 38
c108 30 0 6.33061e-20 $X=6.66 $Y=1.605
c109 23 0 8.37829e-20 $X=5.18 $Y=1.63
c110 20 0 7.57553e-20 $X=5.35 $Y=2.035
c111 15 0 3.15576e-20 $X=6.705 $Y=2.46
c112 11 0 3.2498e-19 $X=6.69 $Y=0.93
c113 7 0 1.13206e-20 $X=5.32 $Y=0.93
c114 3 0 7.5232e-20 $X=5.11 $Y=2.46
r115 31 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.605
+ $X2=6.66 $Y2=1.77
r116 31 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.605
+ $X2=6.66 $Y2=1.44
r117 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.605 $X2=6.66 $Y2=1.605
r118 27 30 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.51 $Y=1.605
+ $X2=6.66 $Y2=1.605
r119 26 38 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.185 $Y=1.635
+ $X2=5.32 $Y2=1.635
r120 26 35 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.185 $Y=1.635
+ $X2=5.11 $Y2=1.635
r121 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.185
+ $Y=1.635 $X2=5.185 $Y2=1.635
r122 23 33 5.3375 $w=3.2e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=1.63 $X2=5.04
+ $Y2=1.63
r123 23 25 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=1.63
+ $X2=5.265 $Y2=1.63
r124 21 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.51 $Y=1.77
+ $X2=6.51 $Y2=1.605
r125 21 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.51 $Y=1.77
+ $X2=6.51 $Y2=1.95
r126 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=6.51 $Y2=1.95
r127 19 20 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=5.35 $Y2=2.035
r128 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.265 $Y=1.95
+ $X2=5.35 $Y2=2.035
r129 17 25 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.265 $Y=1.79
+ $X2=5.265 $Y2=1.63
r130 17 18 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.265 $Y=1.79
+ $X2=5.265 $Y2=1.95
r131 15 42 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.705 $Y=2.46
+ $X2=6.705 $Y2=1.77
r132 11 41 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.69 $Y=0.93
+ $X2=6.69 $Y2=1.44
r133 5 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.47
+ $X2=5.32 $Y2=1.635
r134 5 7 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.32 $Y=1.47 $X2=5.32
+ $Y2=0.93
r135 1 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.11 $Y=1.8
+ $X2=5.11 $Y2=1.635
r136 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.11 $Y=1.8 $X2=5.11
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A1 3 7 11 15 17 26
c53 15 0 1.10938e-19 $X=6.195 $Y=2.46
c54 11 0 1.83396e-19 $X=6.18 $Y=0.93
c55 7 0 2.77406e-20 $X=5.75 $Y=0.93
r56 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.18 $Y=1.615
+ $X2=6.195 $Y2=1.615
r57 23 25 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=5.8 $Y=1.615
+ $X2=6.18 $Y2=1.615
r58 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.8
+ $Y=1.615 $X2=5.8 $Y2=1.615
r59 21 23 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=5.75 $Y=1.615 $X2=5.8
+ $Y2=1.615
r60 19 21 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.725 $Y=1.615
+ $X2=5.75 $Y2=1.615
r61 17 24 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6 $Y=1.615 $X2=5.8
+ $Y2=1.615
r62 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.78
+ $X2=6.195 $Y2=1.615
r63 13 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.195 $Y=1.78
+ $X2=6.195 $Y2=2.46
r64 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.45
+ $X2=6.18 $Y2=1.615
r65 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.18 $Y=1.45 $X2=6.18
+ $Y2=0.93
r66 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.75 $Y=1.45
+ $X2=5.75 $Y2=1.615
r67 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.75 $Y=1.45 $X2=5.75
+ $Y2=0.93
r68 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=1.78
+ $X2=5.725 $Y2=1.615
r69 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.725 $Y=1.78
+ $X2=5.725 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A3 3 7 11 15 17 18 28
c50 18 0 3.15576e-20 $X=7.92 $Y=1.665
c51 3 0 6.33061e-20 $X=7.14 $Y=0.93
r52 27 28 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=7.655 $Y=1.615
+ $X2=7.665 $Y2=1.615
r53 25 27 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.65 $Y=1.615
+ $X2=7.655 $Y2=1.615
r54 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.65
+ $Y=1.615 $X2=7.65 $Y2=1.615
r55 23 25 86.5563 $w=3.3e-07 $l=4.95e-07 $layer=POLY_cond $X=7.155 $Y=1.615
+ $X2=7.65 $Y2=1.615
r56 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.14 $Y=1.615
+ $X2=7.155 $Y2=1.615
r57 18 26 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.92 $Y=1.615
+ $X2=7.65 $Y2=1.615
r58 17 26 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.65 $Y2=1.615
r59 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.45
+ $X2=7.665 $Y2=1.615
r60 13 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.665 $Y=1.45
+ $X2=7.665 $Y2=0.93
r61 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.78
+ $X2=7.655 $Y2=1.615
r62 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.655 $Y=1.78
+ $X2=7.655 $Y2=2.46
r63 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.78
+ $X2=7.155 $Y2=1.615
r64 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.155 $Y=1.78
+ $X2=7.155 $Y2=2.46
r65 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.14 $Y=1.45
+ $X2=7.14 $Y2=1.615
r66 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.14 $Y=1.45 $X2=7.14
+ $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 43 45 47
+ 52 57 65 70 77 78 84 87 90 93 96
r111 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r116 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r117 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r119 75 96 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.405 $Y2=3.33
r120 75 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 74 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 74 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 71 93 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.465 $Y2=3.33
r125 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.645 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 70 96 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.405 $Y2=3.33
r127 70 73 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r128 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r129 69 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r130 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r131 66 90 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.615 $Y=3.33
+ $X2=5.412 $Y2=3.33
r132 66 68 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.615 $Y=3.33
+ $X2=6 $Y2=3.33
r133 65 93 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.285 $Y=3.33
+ $X2=6.465 $Y2=3.33
r134 65 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.285 $Y=3.33
+ $X2=6 $Y2=3.33
r135 64 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r136 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r137 61 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 60 63 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r139 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 58 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.13 $Y2=3.33
r141 58 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r142 57 90 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.412 $Y2=3.33
r143 57 63 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 56 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 56 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r147 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r148 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r149 52 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.13 $Y2=3.33
r150 52 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 51 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 51 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 48 81 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r155 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r156 47 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r157 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r158 45 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r159 45 61 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r160 41 96 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=3.33
r161 41 43 32.5154 $w=2.78e-07 $l=7.9e-07 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=2.455
r162 37 93 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.465 $Y=3.245
+ $X2=6.465 $Y2=3.33
r163 37 39 14.4055 $w=3.58e-07 $l=4.5e-07 $layer=LI1_cond $X=6.465 $Y=3.245
+ $X2=6.465 $Y2=2.795
r164 33 90 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.412 $Y=3.245
+ $X2=5.412 $Y2=3.33
r165 33 35 13.9431 $w=4.03e-07 $l=4.9e-07 $layer=LI1_cond $X=5.412 $Y=3.245
+ $X2=5.412 $Y2=2.755
r166 29 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=3.33
r167 29 31 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=2.405
r168 25 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r169 25 27 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.295
r170 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r171 19 81 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r172 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r173 6 43 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=7.245
+ $Y=1.96 $X2=7.38 $Y2=2.455
r174 5 39 600 $w=1.7e-07 $l=9.20611e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.96 $X2=6.465 $Y2=2.795
r175 4 35 600 $w=1.7e-07 $l=8.84915e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.96 $X2=5.39 $Y2=2.755
r176 3 31 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.84 $X2=2.13 $Y2=2.405
r177 2 27 300 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.295
r178 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r179 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%X 1 2 3 4 13 14 15 16 18 21 25 27 29 31 33 37
+ 42 44 47
c69 47 0 1.55137e-19 $X=0.24 $Y=1.295
c70 13 0 1.58808e-19 $X=0.615 $Y=1.055
r71 40 47 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.24 $Y2=1.295
r72 39 47 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r73 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.735 $Y=0.93
+ $X2=1.735 $Y2=0.595
r74 31 46 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=2.02
+ $X2=1.655 $Y2=1.935
r75 31 33 33.5443 $w=2.78e-07 $l=8.15e-07 $layer=LI1_cond $X=1.655 $Y=2.02
+ $X2=1.655 $Y2=2.835
r76 30 44 4.36636 $w=2.5e-07 $l=1.03e-07 $layer=LI1_cond $X=0.82 $Y=1.055
+ $X2=0.717 $Y2=1.055
r77 29 35 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=1.57 $Y=1.055
+ $X2=1.735 $Y2=0.93
r78 29 30 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=1.57 $Y=1.055
+ $X2=0.82 $Y2=1.055
r79 28 42 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=1.935
+ $X2=0.69 $Y2=1.935
r80 27 46 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.515 $Y=1.935
+ $X2=1.655 $Y2=1.935
r81 27 28 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.515 $Y=1.935
+ $X2=0.815 $Y2=1.935
r82 23 44 2.066 $w=2.05e-07 $l=1.25e-07 $layer=LI1_cond $X=0.717 $Y=0.93
+ $X2=0.717 $Y2=1.055
r83 23 25 19.2062 $w=2.03e-07 $l=3.55e-07 $layer=LI1_cond $X=0.717 $Y=0.93
+ $X2=0.717 $Y2=0.575
r84 19 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.02 $X2=0.69
+ $Y2=1.935
r85 19 21 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=0.69 $Y=2.02
+ $X2=0.69 $Y2=2.815
r86 18 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.85 $X2=0.69
+ $Y2=1.935
r87 17 18 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=0.69 $Y=1.65 $X2=0.69
+ $Y2=1.85
r88 16 40 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.565
+ $X2=0.24 $Y2=1.48
r89 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.69 $Y2=1.65
r90 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.355 $Y2=1.565
r91 14 39 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=0.355 $Y=1.055
+ $X2=0.24 $Y2=1.18
r92 13 44 4.36636 $w=2.5e-07 $l=1.02e-07 $layer=LI1_cond $X=0.615 $Y=1.055
+ $X2=0.717 $Y2=1.055
r93 13 14 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.055
+ $X2=0.355 $Y2=1.055
r94 4 46 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.015
r95 4 33 400 $w=1.7e-07 $l=1.06035e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.835
r96 3 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r97 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r98 2 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.595
+ $Y=0.45 $X2=1.735 $Y2=0.595
r99 1 44 182 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.45 $X2=0.715 $Y2=1.065
r100 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.45 $X2=0.715 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A_509_392# 1 2 3 4 5 6 21 23 24 27 29 33 37
+ 39 40 43 45 47 49 51 53 59 62
c107 39 0 1.10938e-19 $X=6.93 $Y=2.12
r108 55 57 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=4.76 $Y=2.375
+ $X2=4.76 $Y2=2.435
r109 53 55 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.76 $Y=2.085
+ $X2=4.76 $Y2=2.375
r110 47 64 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=2.12 $X2=7.88
+ $Y2=2.035
r111 47 49 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.88 $Y=2.12
+ $X2=7.88 $Y2=2.815
r112 46 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=2.035
+ $X2=6.93 $Y2=2.035
r113 45 64 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=2.035
+ $X2=7.88 $Y2=2.035
r114 45 46 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.715 $Y=2.035
+ $X2=7.095 $Y2=2.035
r115 41 62 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.955 $Y=2.46
+ $X2=6.93 $Y2=2.375
r116 41 43 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=6.955 $Y=2.46
+ $X2=6.955 $Y2=2.465
r117 40 62 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=2.29
+ $X2=6.93 $Y2=2.375
r118 39 61 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=2.12 $X2=6.93
+ $Y2=2.035
r119 39 40 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.93 $Y=2.12
+ $X2=6.93 $Y2=2.29
r120 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=2.375
+ $X2=5.95 $Y2=2.375
r121 37 62 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=2.375
+ $X2=6.93 $Y2=2.375
r122 37 38 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.765 $Y=2.375
+ $X2=6.115 $Y2=2.375
r123 34 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=2.375
+ $X2=4.76 $Y2=2.375
r124 33 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=2.375
+ $X2=5.95 $Y2=2.375
r125 33 34 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.785 $Y=2.375
+ $X2=4.925 $Y2=2.375
r126 31 57 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.76 $Y=2.46
+ $X2=4.76 $Y2=2.435
r127 31 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.76 $Y=2.46
+ $X2=4.76 $Y2=2.905
r128 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.99
+ $X2=3.69 $Y2=2.99
r129 29 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.595 $Y=2.99
+ $X2=4.76 $Y2=2.905
r130 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.595 $Y=2.99
+ $X2=3.855 $Y2=2.99
r131 25 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.905
+ $X2=3.69 $Y2=2.99
r132 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.69 $Y=2.905
+ $X2=3.69 $Y2=2.405
r133 23 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=3.69 $Y2=2.99
r134 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=2.855 $Y2=2.99
r135 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.69 $Y=2.905
+ $X2=2.855 $Y2=2.99
r136 19 21 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.69 $Y=2.905
+ $X2=2.69 $Y2=2.405
r137 6 64 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.96 $X2=7.88 $Y2=2.115
r138 6 49 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.96 $X2=7.88 $Y2=2.815
r139 5 61 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.96 $X2=6.93 $Y2=2.085
r140 5 43 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=6.795
+ $Y=1.96 $X2=6.93 $Y2=2.465
r141 4 59 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=5.815
+ $Y=1.96 $X2=5.95 $Y2=2.375
r142 3 57 300 $w=1.7e-07 $l=5.88855e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=1.96 $X2=4.76 $Y2=2.435
r143 3 53 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.96 $X2=4.76 $Y2=2.085
r144 2 27 300 $w=1.7e-07 $l=5.29481e-07 $layer=licon1_PDIFF $count=2 $X=3.505
+ $Y=1.96 $X2=3.69 $Y2=2.405
r145 1 21 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.96 $X2=2.69 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%VGND 1 2 3 4 5 16 18 22 26 29 32 40 41 42 44
+ 49 61 70 71 77 80 83
c89 71 0 6.39601e-20 $X=7.92 $Y=0
c90 40 0 1.36109e-20 $X=4.585 $Y=0
c91 32 0 1.9667e-19 $X=7.365 $Y=0.755
c92 1 0 3.13945e-19 $X=0.135 $Y=0.45
r93 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r94 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r95 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r96 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 71 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r98 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r99 68 83 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=7.545 $Y=0 $X2=7.367
+ $Y2=0
r100 68 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.92 $Y2=0
r101 67 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r102 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r103 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r104 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r105 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r106 61 83 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.19 $Y=0 $X2=7.367
+ $Y2=0
r107 61 66 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.19 $Y=0 $X2=6.96
+ $Y2=0
r108 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r109 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r110 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r111 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r112 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r113 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r114 54 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r115 53 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r116 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r117 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r118 50 77 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.195
+ $Y2=0
r119 50 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.68
+ $Y2=0
r120 49 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.235
+ $Y2=0
r121 49 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.68
+ $Y2=0
r122 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r123 48 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r124 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r125 45 74 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r126 45 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r127 44 77 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.195
+ $Y2=0
r128 44 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r129 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r130 42 57 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r131 40 59 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.56
+ $Y2=0
r132 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.67
+ $Y2=0
r133 39 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=5.04 $Y2=0
r134 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.67
+ $Y2=0
r135 30 83 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.367 $Y=0.085
+ $X2=7.367 $Y2=0
r136 30 32 21.7503 $w=3.53e-07 $l=6.7e-07 $layer=LI1_cond $X=7.367 $Y=0.085
+ $X2=7.367 $Y2=0.755
r137 29 35 9.29238 $w=1.83e-07 $l=1.55e-07 $layer=LI1_cond $X=4.67 $Y=0.847
+ $X2=4.515 $Y2=0.847
r138 28 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0
r139 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0.755
r140 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r141 24 26 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.675
r142 20 77 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r143 20 22 14.3353 $w=4.08e-07 $l=5.1e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.595
r144 16 74 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r145 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.595
r146 5 32 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=7.215
+ $Y=0.61 $X2=7.365 $Y2=0.755
r147 4 35 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.695 $X2=4.515 $Y2=0.845
r148 3 26 91 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.45 $X2=2.235 $Y2=0.675
r149 2 22 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.45 $X2=1.195 $Y2=0.595
r150 1 18 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.45 $X2=0.28 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A_587_110# 1 2 9 12
c23 9 0 1.22971e-19 $X=4.015 $Y=0.84
r24 12 14 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.075 $Y=0.705
+ $X2=3.075 $Y2=0.84
r25 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0.84
+ $X2=3.075 $Y2=0.84
r26 7 9 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.24 $Y=0.84
+ $X2=4.015 $Y2=0.84
r27 2 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.695 $X2=4.015 $Y2=0.84
r28 1 12 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=2.935
+ $Y=0.55 $X2=3.075 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A_992_122# 1 2 3 12 14 15 19 20 21 24
r48 22 24 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=7.88 $Y=1.1
+ $X2=7.88 $Y2=0.755
r49 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=1.185
+ $X2=7.88 $Y2=1.1
r50 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.715 $Y=1.185
+ $X2=6.99 $Y2=1.185
r51 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.865 $Y=1.1
+ $X2=6.99 $Y2=1.185
r52 17 19 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=6.865 $Y=1.1
+ $X2=6.865 $Y2=0.755
r53 16 19 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=6.865 $Y=0.425
+ $X2=6.865 $Y2=0.755
r54 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.74 $Y=0.34
+ $X2=6.865 $Y2=0.425
r55 14 15 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=6.74 $Y=0.34
+ $X2=5.19 $Y2=0.34
r56 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.065 $Y=0.425
+ $X2=5.19 $Y2=0.34
r57 10 12 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.065 $Y=0.425
+ $X2=5.065 $Y2=0.765
r58 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.61 $X2=7.88 $Y2=0.755
r59 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.61 $X2=6.905 $Y2=0.755
r60 1 12 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=4.96
+ $Y=0.61 $X2=5.105 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_4%A_1079_122# 1 2 7 13 16
c21 16 0 1.65419e-19 $X=6.395 $Y=0.76
c22 13 0 2.77406e-20 $X=5.535 $Y=0.765
c23 7 0 1.13206e-20 $X=6.31 $Y=0.68
r24 8 13 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.62 $Y=0.68
+ $X2=5.495 $Y2=0.68
r25 7 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.31 $Y=0.68
+ $X2=6.435 $Y2=0.68
r26 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.31 $Y=0.68 $X2=5.62
+ $Y2=0.68
r27 2 16 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=6.255
+ $Y=0.61 $X2=6.395 $Y2=0.76
r28 1 13 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.61 $X2=5.535 $Y2=0.765
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o32ai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o32ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.071000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.610000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 3.095000 1.180000 ;
        RECT 0.565000 1.950000 3.255000 2.120000 ;
        RECT 0.565000 2.120000 0.895000 2.735000 ;
        RECT 1.545000 0.610000 1.875000 1.010000 ;
        RECT 2.925000 1.180000 3.095000 1.820000 ;
        RECT 2.925000 1.820000 3.255000 1.950000 ;
        RECT 2.925000 2.120000 3.255000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.240000 0.085000 ;
        RECT 2.555000  0.085000 3.125000 0.500000 ;
        RECT 3.805000  0.085000 4.135000 0.800000 ;
        RECT 4.805000  0.085000 5.625000 0.805000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.240000 3.415000 ;
        RECT 1.465000 2.630000 1.715000 3.245000 ;
        RECT 4.835000 2.290000 5.165000 3.245000 ;
        RECT 5.870000 1.950000 6.120000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.255000 2.375000 0.425000 ;
      RECT 0.115000 0.425000 0.365000 1.130000 ;
      RECT 0.115000 1.950000 0.365000 2.905000 ;
      RECT 0.115000 2.905000 1.265000 3.075000 ;
      RECT 1.045000 0.425000 1.375000 0.825000 ;
      RECT 1.095000 2.290000 2.245000 2.460000 ;
      RECT 1.095000 2.460000 1.265000 2.905000 ;
      RECT 1.915000 2.460000 2.245000 2.980000 ;
      RECT 2.045000 0.425000 2.375000 0.670000 ;
      RECT 2.045000 0.670000 3.635000 0.840000 ;
      RECT 2.475000 2.290000 2.725000 2.905000 ;
      RECT 2.475000 2.905000 4.605000 3.075000 ;
      RECT 3.305000 0.350000 3.635000 0.670000 ;
      RECT 3.305000 0.840000 3.635000 1.010000 ;
      RECT 3.305000 1.010000 6.125000 1.180000 ;
      RECT 3.455000 1.950000 3.625000 2.905000 ;
      RECT 3.825000 1.950000 5.670000 2.120000 ;
      RECT 3.825000 2.120000 4.075000 2.735000 ;
      RECT 4.275000 2.290000 4.605000 2.905000 ;
      RECT 4.305000 0.350000 4.635000 1.010000 ;
      RECT 5.335000 2.120000 5.670000 2.980000 ;
      RECT 5.795000 0.350000 6.125000 1.010000 ;
  END
END sky130_fd_sc_ms__o32ai_2

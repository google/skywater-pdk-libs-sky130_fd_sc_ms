* File: sky130_fd_sc_ms__or3_1.pex.spice
* Created: Wed Sep  2 12:28:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR3_1%C 1 3 6 8 12
c27 12 0 1.21053e-19 $X=0.405 $Y=1.515
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.515 $X2=0.405 $Y2=1.515
r29 8 12 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.405 $Y2=1.565
r30 4 11 38.5662 $w=2.97e-07 $l=2.00237e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.417 $Y2=1.515
r31 4 6 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.495 $Y=1.35 $X2=0.495
+ $Y2=0.645
r32 1 11 48.8089 $w=2.97e-07 $l=2.95745e-07 $layer=POLY_cond $X=0.505 $Y=1.77
+ $X2=0.417 $Y2=1.515
r33 1 3 152.633 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=0.505 $Y=1.77
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_1%B 3 7 9 12
c33 3 0 1.94824e-19 $X=0.925 $Y=2.34
r34 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.515 $X2=1
+ $Y2=1.68
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.515 $X2=1
+ $Y2=1.35
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.515
+ $X2=1 $Y2=1.515
r37 9 13 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1
+ $Y2=1.565
r38 7 14 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.995 $Y=0.645
+ $X2=0.995 $Y2=1.35
r39 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=2.34
+ $X2=0.925 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_1%A 3 7 9 15 16
c36 15 0 7.37712e-20 $X=1.65 $Y=1.515
c37 7 0 7.84672e-20 $X=1.81 $Y=0.645
r38 14 16 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.65 $Y=1.515
+ $X2=1.81 $Y2=1.515
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r40 11 14 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.495 $Y=1.515
+ $X2=1.65 $Y2=1.515
r41 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r42 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.81 $Y2=1.515
r43 5 7 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.81 $Y=1.35 $X2=1.81
+ $Y2=0.645
r44 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.68
+ $X2=1.495 $Y2=1.515
r45 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.495 $Y=1.68
+ $X2=1.495 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_1%A_27_74# 1 2 3 12 16 20 25 26 28 30 31 33 36
+ 37 41
r87 41 44 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.465
+ $X2=2.295 $Y2=1.63
r88 41 43 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.465
+ $X2=2.295 $Y2=1.3
r89 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.465 $X2=2.29 $Y2=1.465
r90 35 37 10.9648 $w=7.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.595 $Y=0.817
+ $X2=1.76 $Y2=0.817
r91 35 36 17.3164 $w=7.23e-07 $l=5.5e-07 $layer=LI1_cond $X=1.595 $Y=0.817
+ $X2=1.045 $Y2=0.817
r92 30 40 9.1003 $w=2.73e-07 $l=2.07918e-07 $layer=LI1_cond $X=2.175 $Y=1.63
+ $X2=2.272 $Y2=1.465
r93 30 31 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.175 $Y=1.63
+ $X2=2.175 $Y2=1.95
r94 28 40 16.5348 $w=2.73e-07 $l=4.51929e-07 $layer=LI1_cond $X=2.09 $Y=1.095
+ $X2=2.272 $Y2=1.465
r95 28 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.09 $Y=1.095
+ $X2=1.76 $Y2=1.095
r96 27 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r97 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.09 $Y=2.035
+ $X2=2.175 $Y2=1.95
r98 26 27 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=2.09 $Y=2.035
+ $X2=0.445 $Y2=2.035
r99 25 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.365 $Y=1.095
+ $X2=1.045 $Y2=1.095
r100 18 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r101 18 20 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.645
r102 16 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.38 $Y=0.74
+ $X2=2.38 $Y2=1.3
r103 12 44 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.375 $Y=2.4
+ $X2=2.375 $Y2=1.63
r104 3 33 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r105 2 35 91 $w=1.7e-07 $l=6.37868e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.595 $Y2=0.62
r106 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_1%VPWR 1 6 8 10 20 21 24
r27 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 18 24 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=1.935 $Y2=3.33
r31 18 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 13 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 10 24 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.935 $Y2=3.33
r37 10 16 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r38 8 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 4 24 3.03114 $w=7.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=3.245
+ $X2=1.935 $Y2=3.33
r41 4 6 13.6919 $w=7.58e-07 $l=8.7e-07 $layer=LI1_cond $X=1.935 $Y=3.245
+ $X2=1.935 $Y2=2.375
r42 1 6 150 $w=1.7e-07 $l=7.88353e-07 $layer=licon1_PDIFF $count=4 $X=1.585
+ $Y=1.84 $X2=2.15 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_1%X 1 2 7 9 15 16 17 28
c24 17 0 7.84672e-20 $X=2.555 $Y=0.84
r25 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=2.612 $Y=0.948
+ $X2=2.612 $Y2=0.925
r26 17 30 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=2.612 $Y=0.979
+ $X2=2.612 $Y2=1.13
r27 17 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=2.612 $Y=0.979
+ $X2=2.612 $Y2=0.948
r28 17 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=2.612 $Y=0.894
+ $X2=2.612 $Y2=0.925
r29 16 17 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=2.612 $Y=0.515
+ $X2=2.612 $Y2=0.894
r30 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.71 $Y=1.82 $X2=2.71
+ $Y2=1.13
r31 9 11 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.655 $Y=1.985
+ $X2=2.655 $Y2=2.815
r32 7 15 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.655 $Y=1.96
+ $X2=2.655 $Y2=1.82
r33 7 9 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.655 $Y=1.96
+ $X2=2.655 $Y2=1.985
r34 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=2.815
r35 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=1.985
r36 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.455
+ $Y=0.37 $X2=2.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.095
+ $Y2=0
r39 27 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.64
+ $Y2=0
r40 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r42 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r43 23 25 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.68
+ $Y2=0
r44 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.095
+ $Y2=0
r45 22 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.68
+ $Y2=0
r46 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r49 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r50 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r51 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r52 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r53 11 13 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.645
r54 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r55 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.645
r56 2 13 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.37 $X2=2.095 $Y2=0.645
r57 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.645
.ends


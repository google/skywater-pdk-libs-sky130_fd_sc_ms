* File: sky130_fd_sc_ms__buf_1.pxi.spice
* Created: Wed Sep  2 11:59:21 2020
* 
x_PM_SKY130_FD_SC_MS__BUF_1%A N_A_M1002_g N_A_M1001_g N_A_c_39_n N_A_c_40_n A A
+ PM_SKY130_FD_SC_MS__BUF_1%A
x_PM_SKY130_FD_SC_MS__BUF_1%A_27_164# N_A_27_164#_M1002_s N_A_27_164#_M1001_s
+ N_A_27_164#_M1000_g N_A_27_164#_M1003_g N_A_27_164#_c_83_n N_A_27_164#_c_77_n
+ N_A_27_164#_c_84_n N_A_27_164#_c_85_n N_A_27_164#_c_78_n N_A_27_164#_c_79_n
+ N_A_27_164#_c_80_n N_A_27_164#_c_81_n PM_SKY130_FD_SC_MS__BUF_1%A_27_164#
x_PM_SKY130_FD_SC_MS__BUF_1%VPWR N_VPWR_M1001_d N_VPWR_c_138_n VPWR
+ N_VPWR_c_139_n N_VPWR_c_140_n N_VPWR_c_137_n N_VPWR_c_142_n
+ PM_SKY130_FD_SC_MS__BUF_1%VPWR
x_PM_SKY130_FD_SC_MS__BUF_1%X N_X_M1003_d N_X_M1000_d N_X_c_159_n N_X_c_160_n X
+ X X X N_X_c_161_n PM_SKY130_FD_SC_MS__BUF_1%X
x_PM_SKY130_FD_SC_MS__BUF_1%VGND N_VGND_M1002_d N_VGND_c_184_n VGND
+ N_VGND_c_185_n N_VGND_c_186_n N_VGND_c_187_n N_VGND_c_188_n
+ PM_SKY130_FD_SC_MS__BUF_1%VGND
cc_1 VNB N_A_M1002_g 0.0400717f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.835
cc_2 VNB N_A_c_39_n 0.0305395f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.615
cc_3 VNB N_A_c_40_n 0.00733759f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.45
cc_4 VNB A 0.00958066f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_A_27_164#_M1000_g 0.00187089f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.615
cc_6 VNB N_A_27_164#_M1003_g 0.0286459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_164#_c_77_n 0.00640208f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_8 VNB N_A_27_164#_c_78_n 0.00728026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_164#_c_79_n 4.08398e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_164#_c_80_n 0.0351504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_164#_c_81_n 0.0336658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_137_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_X_c_159_n 0.0265168f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.615
cc_14 VNB N_X_c_160_n 0.0135379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_X_c_161_n 0.0246538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_184_n 0.0169218f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.54
cc_17 VNB N_VGND_c_185_n 0.0331697f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.45
cc_18 VNB N_VGND_c_186_n 0.0189562f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.615
cc_19 VNB N_VGND_c_187_n 0.146496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_188_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VPB N_A_M1001_g 0.0273665f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=2.54
cc_22 VPB N_A_c_39_n 0.0290939f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.615
cc_23 VPB N_A_c_40_n 0.0213385f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.45
cc_24 VPB A 0.00913245f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_25 VPB N_A_27_164#_M1000_g 0.0301494f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.615
cc_26 VPB N_A_27_164#_c_83_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.615
cc_27 VPB N_A_27_164#_c_84_n 0.00345358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_A_27_164#_c_85_n 0.00948019f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_29 VPB N_A_27_164#_c_79_n 0.00294881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_138_n 0.00969617f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=2.54
cc_31 VPB N_VPWR_c_139_n 0.0304483f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.45
cc_32 VPB N_VPWR_c_140_n 0.0190763f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.615
cc_33 VPB N_VPWR_c_137_n 0.0656471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_142_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB X 0.0136968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB X 0.0415472f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_X_c_161_n 0.00750262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 N_A_c_40_n N_A_27_164#_M1000_g 0.0195122f $X=0.77 $Y=1.45 $X2=0 $Y2=0
cc_39 N_A_M1002_g N_A_27_164#_M1003_g 0.0174961f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_40 N_A_M1001_g N_A_27_164#_c_83_n 0.0153149f $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_41 N_A_M1002_g N_A_27_164#_c_77_n 0.0116849f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_42 N_A_c_40_n N_A_27_164#_c_77_n 5.73673e-19 $X=0.77 $Y=1.45 $X2=0 $Y2=0
cc_43 N_A_M1001_g N_A_27_164#_c_84_n 0.0108741f $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_44 N_A_c_40_n N_A_27_164#_c_84_n 0.00259237f $X=0.77 $Y=1.45 $X2=0 $Y2=0
cc_45 A N_A_27_164#_c_84_n 0.00782149f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_46 N_A_M1001_g N_A_27_164#_c_85_n 0.00362915f $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_47 N_A_c_39_n N_A_27_164#_c_85_n 0.00696845f $X=0.77 $Y=1.615 $X2=0 $Y2=0
cc_48 N_A_c_40_n N_A_27_164#_c_85_n 6.64394e-19 $X=0.77 $Y=1.45 $X2=0 $Y2=0
cc_49 A N_A_27_164#_c_85_n 0.027657f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A_M1002_g N_A_27_164#_c_78_n 0.00504032f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_51 A N_A_27_164#_c_78_n 0.0124978f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_52 N_A_c_40_n N_A_27_164#_c_79_n 0.0048699f $X=0.77 $Y=1.45 $X2=0 $Y2=0
cc_53 A N_A_27_164#_c_79_n 0.00976617f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A_M1002_g N_A_27_164#_c_80_n 0.0105457f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_55 N_A_c_39_n N_A_27_164#_c_80_n 0.0121759f $X=0.77 $Y=1.615 $X2=0 $Y2=0
cc_56 A N_A_27_164#_c_80_n 0.0631563f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_A_27_164#_c_81_n 0.0175909f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_58 A N_A_27_164#_c_81_n 2.10849e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_138_n 0.00343717f $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_60 N_A_M1001_g N_VPWR_c_139_n 0.005209f $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_VPWR_c_137_n 0.00987709f $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_X_c_159_n 8.70516e-19 $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_63 N_A_M1001_g X 6.56662e-19 $X=0.86 $Y=2.54 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_VGND_c_184_n 0.0060489f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_65 N_A_M1002_g N_VGND_c_185_n 0.00451272f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_66 N_A_M1002_g N_VGND_c_187_n 0.00487769f $X=0.845 $Y=0.835 $X2=0 $Y2=0
cc_67 N_A_27_164#_c_84_n N_VPWR_M1001_d 0.00452164f $X=1.13 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_68 N_A_27_164#_c_79_n N_VPWR_M1001_d 0.00207688f $X=1.215 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_27_164#_M1000_g N_VPWR_c_138_n 0.00343717f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A_27_164#_c_83_n N_VPWR_c_138_n 0.0266809f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_71 N_A_27_164#_c_84_n N_VPWR_c_138_n 0.023362f $X=1.13 $Y=2.035 $X2=0 $Y2=0
cc_72 N_A_27_164#_c_81_n N_VPWR_c_138_n 3.74259e-19 $X=1.325 $Y=1.465 $X2=0
+ $Y2=0
cc_73 N_A_27_164#_c_83_n N_VPWR_c_139_n 0.014549f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_74 N_A_27_164#_M1000_g N_VPWR_c_140_n 0.005209f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_75 N_A_27_164#_M1000_g N_VPWR_c_137_n 0.00986335f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A_27_164#_c_83_n N_VPWR_c_137_n 0.0119743f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_77 N_A_27_164#_M1003_g N_X_c_159_n 0.00823464f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A_27_164#_M1003_g N_X_c_160_n 0.00455868f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_79 N_A_27_164#_c_78_n N_X_c_160_n 0.00278159f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_80 N_A_27_164#_M1000_g X 0.00323703f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A_27_164#_c_78_n X 0.00139316f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_82 N_A_27_164#_c_79_n X 0.00565814f $X=1.215 $Y=1.95 $X2=0 $Y2=0
cc_83 N_A_27_164#_M1000_g X 0.0144831f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_27_164#_c_83_n X 0.0040668f $X=0.635 $Y=2.265 $X2=0 $Y2=0
cc_85 N_A_27_164#_M1003_g N_X_c_161_n 0.0131732f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_27_164#_c_78_n N_X_c_161_n 0.0309827f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_87 N_A_27_164#_c_79_n N_X_c_161_n 0.00622921f $X=1.215 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_27_164#_c_78_n N_VGND_M1002_d 0.00188126f $X=1.215 $Y=1.63 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_27_164#_M1003_g N_VGND_c_184_n 0.00941074f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_90 N_A_27_164#_c_77_n N_VGND_c_184_n 0.0126515f $X=1.13 $Y=1.195 $X2=0 $Y2=0
cc_91 N_A_27_164#_c_78_n N_VGND_c_184_n 0.0150119f $X=1.215 $Y=1.63 $X2=0 $Y2=0
cc_92 N_A_27_164#_c_81_n N_VGND_c_184_n 6.97737e-19 $X=1.325 $Y=1.465 $X2=0
+ $Y2=0
cc_93 N_A_27_164#_M1003_g N_VGND_c_186_n 0.00434272f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_94 N_A_27_164#_M1003_g N_VGND_c_187_n 0.00828717f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_95 N_A_27_164#_c_80_n N_VGND_c_187_n 0.0266705f $X=0.795 $Y=1.04 $X2=0 $Y2=0
cc_96 N_VPWR_c_138_n X 0.027028f $X=1.135 $Y=2.455 $X2=0 $Y2=0
cc_97 N_VPWR_c_140_n X 0.0158876f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_98 N_VPWR_c_137_n X 0.0130823f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_99 N_X_c_159_n N_VGND_c_184_n 0.0231775f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_100 N_X_c_159_n N_VGND_c_186_n 0.0156794f $X=1.64 $Y=0.515 $X2=0 $Y2=0
cc_101 N_X_c_159_n N_VGND_c_187_n 0.0129217f $X=1.64 $Y=0.515 $X2=0 $Y2=0

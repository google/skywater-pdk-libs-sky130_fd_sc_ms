# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__nor4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295000 1.350000 4.195000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.470000 0.865000 1.800000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.290300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.250000 0.330000 1.580000 0.790000 ;
        RECT 1.250000 0.790000 2.770000 0.960000 ;
        RECT 1.655000 1.820000 1.825000 1.950000 ;
        RECT 1.655000 1.950000 3.095000 2.120000 ;
        RECT 1.655000 2.120000 1.825000 2.735000 ;
        RECT 2.440000 0.350000 2.770000 0.790000 ;
        RECT 2.440000 0.960000 2.770000 1.010000 ;
        RECT 2.440000 1.010000 5.145000 1.180000 ;
        RECT 2.925000 1.180000 3.095000 1.950000 ;
        RECT 3.440000 0.350000 3.770000 1.010000 ;
        RECT 4.815000 0.350000 5.145000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.580000 1.130000 ;
      RECT 0.115000  1.130000 1.775000 1.300000 ;
      RECT 0.115000  1.300000 0.365000 2.980000 ;
      RECT 0.565000  1.970000 0.895000 3.245000 ;
      RECT 0.750000  0.085000 1.080000 0.960000 ;
      RECT 1.105000  1.300000 1.775000 1.550000 ;
      RECT 1.125000  1.820000 1.455000 2.905000 ;
      RECT 1.125000  2.905000 2.275000 3.075000 ;
      RECT 1.750000  0.085000 2.270000 0.600000 ;
      RECT 2.025000  2.290000 3.255000 2.460000 ;
      RECT 2.025000  2.460000 2.275000 2.905000 ;
      RECT 2.475000  2.630000 2.805000 2.905000 ;
      RECT 2.475000  2.905000 4.265000 3.075000 ;
      RECT 2.940000  0.085000 3.270000 0.840000 ;
      RECT 3.005000  2.460000 3.255000 2.735000 ;
      RECT 3.485000  1.950000 5.625000 2.120000 ;
      RECT 3.485000  2.120000 3.735000 2.735000 ;
      RECT 3.935000  2.290000 4.265000 2.905000 ;
      RECT 3.940000  0.085000 4.645000 0.790000 ;
      RECT 4.465000  2.120000 4.635000 2.980000 ;
      RECT 4.835000  2.290000 5.165000 3.245000 ;
      RECT 5.315000  0.085000 5.645000 1.130000 ;
      RECT 5.375000  2.120000 5.625000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__nor4b_2
END LIBRARY

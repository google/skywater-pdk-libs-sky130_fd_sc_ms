* File: sky130_fd_sc_ms__a31oi_4.pxi.spice
* Created: Wed Sep  2 11:55:34 2020
* 
x_PM_SKY130_FD_SC_MS__A31OI_4%A3 N_A3_M1008_g N_A3_M1015_g N_A3_M1021_g
+ N_A3_M1009_g N_A3_M1028_g N_A3_M1011_g N_A3_M1013_g N_A3_M1029_g A3 A3 A3
+ N_A3_c_127_n N_A3_c_128_n PM_SKY130_FD_SC_MS__A31OI_4%A3
x_PM_SKY130_FD_SC_MS__A31OI_4%A2 N_A2_M1014_g N_A2_M1003_g N_A2_M1012_g
+ N_A2_M1016_g N_A2_M1022_g N_A2_M1019_g N_A2_M1026_g N_A2_M1020_g A2 A2 A2 A2
+ N_A2_c_207_n PM_SKY130_FD_SC_MS__A31OI_4%A2
x_PM_SKY130_FD_SC_MS__A31OI_4%A1 N_A1_c_299_n N_A1_M1002_g N_A1_c_290_n
+ N_A1_c_291_n N_A1_M1000_g N_A1_c_302_n N_A1_M1006_g N_A1_c_293_n N_A1_M1005_g
+ N_A1_M1017_g N_A1_M1024_g N_A1_M1018_g N_A1_M1025_g N_A1_c_297_n A1 A1 A1
+ N_A1_c_298_n PM_SKY130_FD_SC_MS__A31OI_4%A1
x_PM_SKY130_FD_SC_MS__A31OI_4%B1 N_B1_M1001_g N_B1_M1023_g N_B1_M1004_g
+ N_B1_M1007_g N_B1_M1010_g N_B1_M1027_g B1 B1 B1 B1 B1 N_B1_c_404_n
+ PM_SKY130_FD_SC_MS__A31OI_4%B1
x_PM_SKY130_FD_SC_MS__A31OI_4%A_27_368# N_A_27_368#_M1008_s N_A_27_368#_M1009_s
+ N_A_27_368#_M1013_s N_A_27_368#_M1016_d N_A_27_368#_M1020_d
+ N_A_27_368#_M1006_d N_A_27_368#_M1018_d N_A_27_368#_M1004_s
+ N_A_27_368#_M1010_s N_A_27_368#_c_464_n N_A_27_368#_c_465_n
+ N_A_27_368#_c_476_n N_A_27_368#_c_549_p N_A_27_368#_c_480_n
+ N_A_27_368#_c_466_n N_A_27_368#_c_547_p N_A_27_368#_c_490_n
+ N_A_27_368#_c_467_n N_A_27_368#_c_498_n N_A_27_368#_c_502_n
+ N_A_27_368#_c_508_n N_A_27_368#_c_510_n N_A_27_368#_c_512_n
+ N_A_27_368#_c_513_n N_A_27_368#_c_468_n N_A_27_368#_c_469_n
+ N_A_27_368#_c_576_p N_A_27_368#_c_470_n N_A_27_368#_c_471_n
+ N_A_27_368#_c_486_n N_A_27_368#_c_503_n N_A_27_368#_c_472_n
+ N_A_27_368#_c_518_n N_A_27_368#_c_521_n N_A_27_368#_c_473_n
+ PM_SKY130_FD_SC_MS__A31OI_4%A_27_368#
x_PM_SKY130_FD_SC_MS__A31OI_4%VPWR N_VPWR_M1008_d N_VPWR_M1011_d N_VPWR_M1014_s
+ N_VPWR_M1019_s N_VPWR_M1002_s N_VPWR_M1017_s N_VPWR_c_584_n N_VPWR_c_585_n
+ N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n
+ N_VPWR_c_591_n VPWR N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n
+ N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_583_n N_VPWR_c_599_n
+ N_VPWR_c_600_n N_VPWR_c_601_n N_VPWR_c_602_n N_VPWR_c_603_n
+ PM_SKY130_FD_SC_MS__A31OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A31OI_4%Y N_Y_M1000_d N_Y_M1005_d N_Y_M1025_d N_Y_M1027_d
+ N_Y_M1001_d N_Y_M1007_d N_Y_c_694_n N_Y_c_712_n N_Y_c_718_n N_Y_c_720_n
+ N_Y_c_695_n N_Y_c_696_n N_Y_c_697_n N_Y_c_749_n N_Y_c_698_n N_Y_c_699_n
+ N_Y_c_700_n N_Y_c_701_n N_Y_c_733_n N_Y_c_762_n Y Y
+ PM_SKY130_FD_SC_MS__A31OI_4%Y
x_PM_SKY130_FD_SC_MS__A31OI_4%A_30_74# N_A_30_74#_M1015_d N_A_30_74#_M1021_d
+ N_A_30_74#_M1029_d N_A_30_74#_M1012_s N_A_30_74#_M1026_s N_A_30_74#_c_808_n
+ N_A_30_74#_c_809_n N_A_30_74#_c_810_n N_A_30_74#_c_811_n N_A_30_74#_c_812_n
+ N_A_30_74#_c_813_n N_A_30_74#_c_814_n N_A_30_74#_c_842_n N_A_30_74#_c_815_n
+ N_A_30_74#_c_816_n N_A_30_74#_c_817_n N_A_30_74#_c_818_n N_A_30_74#_c_819_n
+ PM_SKY130_FD_SC_MS__A31OI_4%A_30_74#
x_PM_SKY130_FD_SC_MS__A31OI_4%VGND N_VGND_M1015_s N_VGND_M1028_s N_VGND_M1023_s
+ N_VGND_c_885_n N_VGND_c_886_n VGND N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n
+ N_VGND_c_894_n PM_SKY130_FD_SC_MS__A31OI_4%VGND
x_PM_SKY130_FD_SC_MS__A31OI_4%A_475_74# N_A_475_74#_M1003_d N_A_475_74#_M1022_d
+ N_A_475_74#_M1000_s N_A_475_74#_M1024_s N_A_475_74#_c_974_n
+ N_A_475_74#_c_967_n N_A_475_74#_c_968_n N_A_475_74#_c_1011_n
+ N_A_475_74#_c_969_n N_A_475_74#_c_980_n N_A_475_74#_c_970_n
+ N_A_475_74#_c_985_n N_A_475_74#_c_971_n N_A_475_74#_c_972_n
+ PM_SKY130_FD_SC_MS__A31OI_4%A_475_74#
cc_1 VNB N_A3_M1015_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_2 VNB N_A3_M1021_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_3 VNB N_A3_M1028_g 0.0234867f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_4 VNB N_A3_M1029_g 0.0244051f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_5 VNB N_A3_c_127_n 0.0166903f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.515
cc_6 VNB N_A3_c_128_n 0.0749748f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.515
cc_7 VNB N_A2_M1003_g 0.0233537f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_8 VNB N_A2_M1012_g 0.0223644f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_9 VNB N_A2_M1022_g 0.0240746f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_10 VNB N_A2_M1026_g 0.0295412f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_11 VNB A2 0.00842528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_207_n 0.0797328f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.515
cc_13 VNB N_A1_c_290_n 0.0108178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_291_n 0.0106752f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.35
cc_15 VNB N_A1_M1000_g 0.0285005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_293_n 0.0288001f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_17 VNB N_A1_M1005_g 0.0246283f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.35
cc_18 VNB N_A1_M1024_g 0.0215982f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.68
cc_19 VNB N_A1_M1025_g 0.0224969f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_A1_c_297_n 0.0149141f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_21 VNB N_A1_c_298_n 0.0512459f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.515
cc_22 VNB N_B1_M1023_g 0.031167f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_23 VNB N_B1_M1027_g 0.0393239f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_24 VNB B1 0.0185476f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_25 VNB N_B1_c_404_n 0.091258f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.515
cc_26 VNB N_VPWR_c_583_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_694_n 0.00688419f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_28 VNB N_Y_c_695_n 0.00592048f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_29 VNB N_Y_c_696_n 0.00280366f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_30 VNB N_Y_c_697_n 0.0193773f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_Y_c_698_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.515
cc_32 VNB N_Y_c_699_n 0.00599341f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.515
cc_33 VNB N_Y_c_700_n 0.00228316f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.515
cc_34 VNB N_Y_c_701_n 0.002409f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=1.515
cc_35 VNB Y 0.00520045f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_36 VNB N_A_30_74#_c_808_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_37 VNB N_A_30_74#_c_809_n 0.00318294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_30_74#_c_810_n 0.00966224f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.68
cc_39 VNB N_A_30_74#_c_811_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_30_74#_c_812_n 0.00442934f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_41 VNB N_A_30_74#_c_813_n 0.00215292f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_42 VNB N_A_30_74#_c_814_n 0.00423139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_30_74#_c_815_n 0.00785609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_30_74#_c_816_n 0.0052509f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.515
cc_45 VNB N_A_30_74#_c_817_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.515
cc_46 VNB N_A_30_74#_c_818_n 0.00380807f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.515
cc_47 VNB N_A_30_74#_c_819_n 0.00219532f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.515
cc_48 VNB N_VGND_c_885_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_886_n 0.00555557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_887_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_888_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.68
cc_52 VNB N_VGND_c_889_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_890_n 0.457781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_891_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_55 VNB N_VGND_c_892_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.515
cc_56 VNB N_VGND_c_893_n 0.124154f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.515
cc_57 VNB N_VGND_c_894_n 0.0365846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_475_74#_c_967_n 0.00237099f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.35
cc_59 VNB N_A_475_74#_c_968_n 0.00202581f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_60 VNB N_A_475_74#_c_969_n 0.0191972f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_61 VNB N_A_475_74#_c_970_n 0.0053724f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_62 VNB N_A_475_74#_c_971_n 0.0026368f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_63 VNB N_A_475_74#_c_972_n 0.00327156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_A3_M1008_g 0.026777f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_65 VPB N_A3_M1009_g 0.0198975f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_66 VPB N_A3_M1011_g 0.0198963f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_67 VPB N_A3_M1013_g 0.0209948f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_68 VPB N_A3_c_127_n 0.0163699f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.515
cc_69 VPB N_A3_c_128_n 0.0119282f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.515
cc_70 VPB N_A2_M1014_g 0.0213574f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_71 VPB N_A2_M1016_g 0.0208299f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_72 VPB N_A2_M1019_g 0.021006f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_73 VPB N_A2_M1020_g 0.0213737f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_74 VPB A2 0.0122026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A2_c_207_n 0.0152437f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.515
cc_76 VPB N_A1_c_299_n 0.0178012f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.68
cc_77 VPB N_A1_c_290_n 0.00755414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A1_c_291_n 0.00356618f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.35
cc_79 VPB N_A1_c_302_n 0.022202f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.74
cc_80 VPB N_A1_c_293_n 0.0139719f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_81 VPB N_A1_M1017_g 0.0290858f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.68
cc_82 VPB N_A1_M1018_g 0.0220532f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.35
cc_83 VPB N_A1_c_297_n 0.00412943f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_84 VPB A1 0.0107483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A1_c_298_n 0.0126574f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.515
cc_86 VPB N_B1_M1001_g 0.0203537f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_87 VPB N_B1_M1004_g 0.0198792f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.74
cc_88 VPB N_B1_M1007_g 0.0196385f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_89 VPB N_B1_M1010_g 0.0252952f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=0.74
cc_90 VPB B1 0.0194751f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.35
cc_91 VPB N_B1_c_404_n 0.0124281f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.515
cc_92 VPB N_A_27_368#_c_464_n 0.0075506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_368#_c_465_n 0.0346591f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_94 VPB N_A_27_368#_c_466_n 0.00455826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_368#_c_467_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.515
cc_96 VPB N_A_27_368#_c_468_n 0.00241371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_368#_c_469_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=1.565
cc_98 VPB N_A_27_368#_c_470_n 0.0117045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_368#_c_471_n 0.0358214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_368#_c_472_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_368#_c_473_n 0.00145593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_584_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.68
cc_103 VPB N_VPWR_c_585_n 0.00261791f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.68
cc_104 VPB N_VPWR_c_586_n 0.00498646f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.35
cc_105 VPB N_VPWR_c_587_n 0.00510895f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_106 VPB N_VPWR_c_588_n 0.00565985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_589_n 0.0093624f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.515
cc_108 VPB N_VPWR_c_590_n 0.0160795f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.515
cc_109 VPB N_VPWR_c_591_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.515
cc_110 VPB N_VPWR_c_592_n 0.017793f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.515
cc_111 VPB N_VPWR_c_593_n 0.0161283f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.515
cc_112 VPB N_VPWR_c_594_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_595_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_596_n 0.0306486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_597_n 0.0594276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_583_n 0.0828425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_599_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_600_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_601_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_602_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_603_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB Y 6.81854e-19 $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_123 N_A3_M1013_g N_A2_M1014_g 0.0123893f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A3_M1029_g N_A2_M1003_g 0.0145382f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A3_c_127_n A2 0.0122223f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A3_c_128_n A2 0.00116522f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A3_c_127_n N_A2_c_207_n 0.00114368f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A3_c_128_n N_A2_c_207_n 0.0269275f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A3_c_127_n N_A_27_368#_c_464_n 0.0222244f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A3_M1008_g N_A_27_368#_c_465_n 6.86474e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A3_M1008_g N_A_27_368#_c_476_n 0.0142562f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A3_M1009_g N_A_27_368#_c_476_n 0.0142562f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A3_c_127_n N_A_27_368#_c_476_n 0.045298f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A3_c_128_n N_A_27_368#_c_476_n 4.90767e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A3_M1011_g N_A_27_368#_c_480_n 0.0142562f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A3_M1013_g N_A_27_368#_c_480_n 0.0165948f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A3_c_127_n N_A_27_368#_c_480_n 0.0304652f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A3_c_128_n N_A_27_368#_c_480_n 4.90767e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A3_M1011_g N_A_27_368#_c_466_n 6.1989e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A3_M1013_g N_A_27_368#_c_466_n 0.00541281f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A3_c_127_n N_A_27_368#_c_486_n 0.0170101f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A3_c_128_n N_A_27_368#_c_486_n 5.53363e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A3_M1008_g N_VPWR_c_584_n 0.0161703f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A3_M1009_g N_VPWR_c_584_n 0.0134815f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A3_M1011_g N_VPWR_c_584_n 5.76765e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A3_M1009_g N_VPWR_c_585_n 5.76765e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A3_M1011_g N_VPWR_c_585_n 0.0134815f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A3_M1013_g N_VPWR_c_585_n 0.0133619f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A3_M1013_g N_VPWR_c_586_n 5.60684e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A3_M1013_g N_VPWR_c_590_n 0.00460063f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A3_M1008_g N_VPWR_c_592_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A3_M1009_g N_VPWR_c_593_n 0.00460063f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A3_M1011_g N_VPWR_c_593_n 0.00460063f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A3_M1008_g N_VPWR_c_583_n 0.00912296f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A3_M1009_g N_VPWR_c_583_n 0.00908554f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A3_M1011_g N_VPWR_c_583_n 0.00908554f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A3_M1013_g N_VPWR_c_583_n 0.00908665f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A3_M1015_g N_A_30_74#_c_808_n 0.00159319f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A3_M1015_g N_A_30_74#_c_809_n 0.0136535f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A3_M1021_g N_A_30_74#_c_809_n 0.0130918f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A3_c_127_n N_A_30_74#_c_809_n 0.051883f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A3_c_128_n N_A_30_74#_c_809_n 0.00280866f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A3_c_127_n N_A_30_74#_c_810_n 0.0225421f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A3_M1021_g N_A_30_74#_c_811_n 3.92313e-19 $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A3_M1028_g N_A_30_74#_c_811_n 3.92313e-19 $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A3_M1028_g N_A_30_74#_c_812_n 0.0134851f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A3_M1029_g N_A_30_74#_c_812_n 0.0151535f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A3_c_127_n N_A_30_74#_c_812_n 0.0381409f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A3_c_128_n N_A_30_74#_c_812_n 0.00412669f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A3_M1028_g N_A_30_74#_c_813_n 9.2425e-19 $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A3_M1029_g N_A_30_74#_c_813_n 0.00986519f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A3_c_127_n N_A_30_74#_c_817_n 0.0146029f $X=1.62 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A3_c_128_n N_A_30_74#_c_817_n 0.00244789f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A3_M1029_g N_A_30_74#_c_818_n 0.00194714f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A3_M1015_g N_VGND_c_885_n 0.0137191f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A3_M1021_g N_VGND_c_885_n 0.0106755f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A3_M1028_g N_VGND_c_885_n 4.71636e-19 $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A3_M1021_g N_VGND_c_886_n 4.71636e-19 $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A3_M1028_g N_VGND_c_886_n 0.0106899f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A3_M1029_g N_VGND_c_886_n 0.00430002f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A3_M1015_g N_VGND_c_887_n 0.00383152f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A3_M1021_g N_VGND_c_888_n 0.00383152f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A3_M1028_g N_VGND_c_888_n 0.00383152f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A3_M1015_g N_VGND_c_890_n 0.00761248f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A3_M1021_g N_VGND_c_890_n 0.0075754f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A3_M1028_g N_VGND_c_890_n 0.0075754f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A3_M1029_g N_VGND_c_890_n 0.0082051f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A3_M1029_g N_VGND_c_893_n 0.00433834f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A3_M1029_g N_A_475_74#_c_968_n 2.72169e-19 $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A2_M1020_g N_A1_c_299_n 0.00701809f $X=3.755 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_191 A2 N_A1_c_299_n 7.6843e-19 $X=3.995 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_192 A2 N_A1_c_291_n 0.00568469f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_c_207_n N_A1_c_291_n 0.00701809f $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_194 A2 N_A1_c_297_n 0.0012834f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A2_M1014_g N_A_27_368#_c_466_n 0.00555244f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A2_M1016_g N_A_27_368#_c_466_n 6.08944e-19 $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A2_M1014_g N_A_27_368#_c_490_n 0.0179409f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A2_M1016_g N_A_27_368#_c_490_n 0.0141879f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_199 A2 N_A_27_368#_c_490_n 0.0317045f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A2_c_207_n N_A_27_368#_c_490_n 7.78314e-19 $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_201 N_A2_M1014_g N_A_27_368#_c_467_n 4.56122e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A2_M1016_g N_A_27_368#_c_467_n 0.0116548f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A2_M1019_g N_A_27_368#_c_467_n 0.0113654f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A2_M1020_g N_A_27_368#_c_467_n 3.83869e-19 $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A2_M1019_g N_A_27_368#_c_498_n 0.0132272f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A2_M1020_g N_A_27_368#_c_498_n 0.0145524f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_207 A2 N_A_27_368#_c_498_n 0.046225f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A2_c_207_n N_A_27_368#_c_498_n 7.63416e-19 $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_209 A2 N_A_27_368#_c_502_n 0.0246997f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A2_M1016_g N_A_27_368#_c_503_n 9.66537e-19 $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A2_M1019_g N_A_27_368#_c_503_n 0.00151375f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_212 A2 N_A_27_368#_c_503_n 0.0235495f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A2_c_207_n N_A_27_368#_c_503_n 5.49827e-19 $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_214 N_A2_M1014_g N_VPWR_c_585_n 5.68836e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A2_M1014_g N_VPWR_c_586_n 0.0126294f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A2_M1016_g N_VPWR_c_586_n 0.00216202f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A2_M1019_g N_VPWR_c_587_n 0.00232104f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A2_M1020_g N_VPWR_c_587_n 0.0133144f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A2_M1014_g N_VPWR_c_590_n 0.00460063f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A2_M1016_g N_VPWR_c_594_n 0.005209f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A2_M1019_g N_VPWR_c_594_n 0.005209f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A2_M1020_g N_VPWR_c_595_n 0.00460063f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A2_M1014_g N_VPWR_c_583_n 0.00908665f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A2_M1016_g N_VPWR_c_583_n 0.00982082f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A2_M1019_g N_VPWR_c_583_n 0.00982082f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A2_M1020_g N_VPWR_c_583_n 0.00909121f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A2_M1026_g N_Y_c_699_n 0.00128862f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A2_M1026_g Y 0.00378125f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_229 A2 Y 0.0268823f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_230 N_A2_c_207_n Y 9.72953e-19 $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_231 N_A2_M1003_g N_A_30_74#_c_813_n 7.13357e-19 $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A2_M1003_g N_A_30_74#_c_814_n 0.0173943f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A2_M1012_g N_A_30_74#_c_814_n 0.0125402f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_234 A2 N_A_30_74#_c_814_n 0.0308532f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A2_c_207_n N_A_30_74#_c_814_n 0.00280982f $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_236 N_A2_M1022_g N_A_30_74#_c_842_n 0.0068333f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A2_M1026_g N_A_30_74#_c_842_n 5.80602e-19 $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A2_M1022_g N_A_30_74#_c_815_n 0.00972446f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A2_M1026_g N_A_30_74#_c_815_n 0.0139049f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_240 A2 N_A_30_74#_c_815_n 0.0795886f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A2_c_207_n N_A_30_74#_c_815_n 0.00593584f $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_242 N_A2_M1022_g N_A_30_74#_c_816_n 5.80141e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A2_M1026_g N_A_30_74#_c_816_n 0.0073896f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1022_g N_A_30_74#_c_819_n 0.00277633f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_245 A2 N_A_30_74#_c_819_n 0.024925f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_207_n N_A_30_74#_c_819_n 0.002631f $X=3.74 $Y=1.517 $X2=0 $Y2=0
cc_247 N_A2_M1003_g N_VGND_c_890_n 0.00816865f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1012_g N_VGND_c_890_n 0.00353528f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1022_g N_VGND_c_890_n 0.00354662f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_M1026_g N_VGND_c_890_n 0.00359661f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1003_g N_VGND_c_893_n 0.00430908f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1012_g N_VGND_c_893_n 0.00278271f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1022_g N_VGND_c_893_n 0.00278271f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1026_g N_VGND_c_893_n 0.00278271f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A2_M1003_g N_A_475_74#_c_974_n 0.00517057f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_M1012_g N_A_475_74#_c_967_n 0.0112351f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A2_M1022_g N_A_475_74#_c_967_n 0.0115476f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A2_M1003_g N_A_475_74#_c_968_n 0.00460758f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1026_g N_A_475_74#_c_969_n 0.0135881f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A1_M1018_g N_B1_M1001_g 0.0194599f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A1_M1025_g N_B1_M1023_g 0.0244181f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A1_M1018_g B1 0.00252869f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_263 A1 B1 0.0269702f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A1_c_298_n B1 0.0141744f $X=6.285 $Y=1.5 $X2=0 $Y2=0
cc_265 N_A1_c_298_n N_B1_c_404_n 0.0273272f $X=6.285 $Y=1.5 $X2=0 $Y2=0
cc_266 N_A1_c_299_n N_A_27_368#_c_502_n 0.00265729f $X=4.255 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A1_c_299_n N_A_27_368#_c_508_n 0.00350217f $X=4.255 $Y=1.765 $X2=0
+ $Y2=0
cc_268 N_A1_c_302_n N_A_27_368#_c_508_n 7.90167e-19 $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_269 N_A1_M1017_g N_A_27_368#_c_510_n 0.0132511f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A1_M1018_g N_A_27_368#_c_510_n 0.0132511f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A1_M1018_g N_A_27_368#_c_512_n 8.84614e-19 $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A1_M1017_g N_A_27_368#_c_513_n 4.40686e-19 $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A1_M1018_g N_A_27_368#_c_513_n 0.00745636f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_274 N_A1_M1018_g N_A_27_368#_c_469_n 0.00350772f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A1_c_299_n N_A_27_368#_c_472_n 0.00844309f $X=4.255 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A1_c_302_n N_A_27_368#_c_472_n 4.7829e-19 $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A1_c_299_n N_A_27_368#_c_518_n 0.0173474f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A1_c_290_n N_A_27_368#_c_518_n 6.82751e-19 $X=4.665 $Y=1.69 $X2=0 $Y2=0
cc_279 N_A1_c_302_n N_A_27_368#_c_518_n 0.0143011f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A1_M1017_g N_A_27_368#_c_521_n 0.00825833f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A1_M1018_g N_A_27_368#_c_521_n 4.43595e-19 $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_282 N_A1_c_299_n N_VPWR_c_587_n 5.12947e-19 $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A1_c_299_n N_VPWR_c_588_n 0.00194999f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A1_c_302_n N_VPWR_c_588_n 0.0128966f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A1_M1017_g N_VPWR_c_589_n 0.00382308f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A1_M1018_g N_VPWR_c_589_n 0.00150551f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A1_c_299_n N_VPWR_c_595_n 0.005209f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A1_c_302_n N_VPWR_c_596_n 0.00460063f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A1_M1017_g N_VPWR_c_596_n 0.00521123f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A1_M1018_g N_VPWR_c_597_n 0.00517089f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A1_c_299_n N_VPWR_c_583_n 0.00982648f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A1_c_302_n N_VPWR_c_583_n 0.00913687f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A1_M1017_g N_VPWR_c_583_n 0.00985277f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A1_M1018_g N_VPWR_c_583_n 0.00978126f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_295 N_A1_M1000_g N_Y_c_694_n 0.0154768f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A1_c_293_n N_Y_c_694_n 0.00971014f $X=5.385 $Y=1.5 $X2=0 $Y2=0
cc_297 N_A1_M1005_g N_Y_c_694_n 0.0115559f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_298 A1 N_Y_c_694_n 0.0451166f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_299 N_A1_c_302_n N_Y_c_712_n 0.0154227f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_300 N_A1_c_293_n N_Y_c_712_n 0.00335607f $X=5.385 $Y=1.5 $X2=0 $Y2=0
cc_301 N_A1_M1017_g N_Y_c_712_n 0.0143417f $X=5.735 $Y=2.4 $X2=0 $Y2=0
cc_302 N_A1_M1018_g N_Y_c_712_n 0.0174995f $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_303 A1 N_Y_c_712_n 0.0894406f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_304 N_A1_c_298_n N_Y_c_712_n 0.00127178f $X=6.285 $Y=1.5 $X2=0 $Y2=0
cc_305 N_A1_c_299_n N_Y_c_718_n 0.00161168f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_306 N_A1_c_302_n N_Y_c_718_n 0.00242711f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_307 N_A1_M1000_g N_Y_c_720_n 7.50704e-19 $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A1_M1005_g N_Y_c_720_n 0.00672007f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A1_M1024_g N_Y_c_695_n 0.0125269f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A1_M1025_g N_Y_c_695_n 0.0161994f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_311 A1 N_Y_c_695_n 0.0204973f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_312 N_A1_c_298_n N_Y_c_695_n 0.00428771f $X=6.285 $Y=1.5 $X2=0 $Y2=0
cc_313 N_A1_M1025_g N_Y_c_696_n 0.00350307f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A1_c_290_n N_Y_c_699_n 0.00300811f $X=4.665 $Y=1.69 $X2=0 $Y2=0
cc_315 N_A1_M1000_g N_Y_c_699_n 0.00646341f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A1_M1005_g N_Y_c_699_n 7.12864e-19 $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A1_M1005_g N_Y_c_700_n 0.00382108f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_318 A1 N_Y_c_700_n 0.0278934f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A1_c_298_n N_Y_c_700_n 0.00477338f $X=6.285 $Y=1.5 $X2=0 $Y2=0
cc_320 N_A1_M1018_g N_Y_c_733_n 6.69372e-19 $X=6.285 $Y=2.4 $X2=0 $Y2=0
cc_321 N_A1_c_299_n Y 0.00434248f $X=4.255 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A1_c_290_n Y 0.0135794f $X=4.665 $Y=1.69 $X2=0 $Y2=0
cc_323 N_A1_M1000_g Y 0.00562378f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A1_c_302_n Y 0.00918269f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A1_M1005_g Y 5.82457e-19 $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A1_c_297_n Y 0.0143137f $X=4.755 $Y=1.542 $X2=0 $Y2=0
cc_327 A1 Y 0.0262176f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_328 N_A1_M1000_g N_A_30_74#_c_815_n 5.33994e-19 $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_M1000_g N_A_30_74#_c_816_n 0.0043775f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1000_g N_VGND_c_890_n 0.00360662f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1005_g N_VGND_c_890_n 0.00356321f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1024_g N_VGND_c_890_n 0.00354085f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1025_g N_VGND_c_890_n 0.0081738f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1000_g N_VGND_c_893_n 0.00278271f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A1_M1005_g N_VGND_c_893_n 0.00278271f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A1_M1024_g N_VGND_c_893_n 0.00278247f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1025_g N_VGND_c_893_n 0.00430908f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1000_g N_A_475_74#_c_969_n 0.0141742f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1000_g N_A_475_74#_c_980_n 0.00991621f $X=4.74 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1005_g N_A_475_74#_c_980_n 0.00687235f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A1_M1005_g N_A_475_74#_c_970_n 0.0123233f $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A1_M1024_g N_A_475_74#_c_970_n 0.0108687f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A1_M1025_g N_A_475_74#_c_970_n 0.00483594f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A1_M1005_g N_A_475_74#_c_985_n 7.30686e-19 $X=5.46 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A1_M1024_g N_A_475_74#_c_985_n 0.00674664f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A1_M1025_g N_A_475_74#_c_985_n 0.00520362f $X=6.39 $Y=0.74 $X2=0 $Y2=0
cc_347 N_B1_M1001_g N_A_27_368#_c_468_n 0.0134336f $X=6.765 $Y=2.4 $X2=0 $Y2=0
cc_348 N_B1_M1004_g N_A_27_368#_c_468_n 0.0141454f $X=7.235 $Y=2.4 $X2=0 $Y2=0
cc_349 N_B1_M1001_g N_A_27_368#_c_469_n 0.00140005f $X=6.765 $Y=2.4 $X2=0 $Y2=0
cc_350 N_B1_M1007_g N_A_27_368#_c_470_n 0.0140221f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_351 N_B1_M1010_g N_A_27_368#_c_470_n 0.0149887f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_352 B1 N_A_27_368#_c_471_n 0.0217457f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_353 N_B1_M1001_g N_VPWR_c_597_n 0.00333926f $X=6.765 $Y=2.4 $X2=0 $Y2=0
cc_354 N_B1_M1004_g N_VPWR_c_597_n 0.00333926f $X=7.235 $Y=2.4 $X2=0 $Y2=0
cc_355 N_B1_M1007_g N_VPWR_c_597_n 0.00333926f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_356 N_B1_M1010_g N_VPWR_c_597_n 0.00333926f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_357 N_B1_M1001_g N_VPWR_c_583_n 0.00423277f $X=6.765 $Y=2.4 $X2=0 $Y2=0
cc_358 N_B1_M1004_g N_VPWR_c_583_n 0.00422888f $X=7.235 $Y=2.4 $X2=0 $Y2=0
cc_359 N_B1_M1007_g N_VPWR_c_583_n 0.00422687f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_360 N_B1_M1010_g N_VPWR_c_583_n 0.00426429f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_361 N_B1_M1001_g N_Y_c_712_n 0.0145431f $X=6.765 $Y=2.4 $X2=0 $Y2=0
cc_362 B1 N_Y_c_712_n 0.0328548f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_363 B1 N_Y_c_695_n 0.010903f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_364 N_B1_M1023_g N_Y_c_696_n 0.0137567f $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_365 N_B1_M1023_g N_Y_c_697_n 0.0131906f $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_366 N_B1_M1027_g N_Y_c_697_n 0.0153378f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_367 B1 N_Y_c_697_n 0.131572f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_368 N_B1_c_404_n N_Y_c_697_n 0.0237f $X=8.135 $Y=1.515 $X2=0 $Y2=0
cc_369 N_B1_M1004_g N_Y_c_749_n 0.012931f $X=7.235 $Y=2.4 $X2=0 $Y2=0
cc_370 N_B1_M1007_g N_Y_c_749_n 0.012931f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_371 B1 N_Y_c_749_n 0.0391869f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_372 N_B1_c_404_n N_Y_c_749_n 4.90767e-19 $X=8.135 $Y=1.515 $X2=0 $Y2=0
cc_373 N_B1_M1027_g N_Y_c_698_n 0.0144033f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_374 N_B1_M1023_g N_Y_c_701_n 0.00171391f $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_375 B1 N_Y_c_701_n 0.0289371f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_376 N_B1_c_404_n N_Y_c_701_n 0.00381358f $X=8.135 $Y=1.515 $X2=0 $Y2=0
cc_377 N_B1_M1001_g N_Y_c_733_n 0.0106423f $X=6.765 $Y=2.4 $X2=0 $Y2=0
cc_378 N_B1_M1004_g N_Y_c_733_n 0.0119137f $X=7.235 $Y=2.4 $X2=0 $Y2=0
cc_379 N_B1_M1007_g N_Y_c_733_n 5.73047e-19 $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_380 B1 N_Y_c_733_n 0.0236897f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_381 N_B1_c_404_n N_Y_c_733_n 6.70282e-19 $X=8.135 $Y=1.515 $X2=0 $Y2=0
cc_382 N_B1_M1004_g N_Y_c_762_n 5.53268e-19 $X=7.235 $Y=2.4 $X2=0 $Y2=0
cc_383 N_B1_M1007_g N_Y_c_762_n 0.0114812f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_384 N_B1_M1010_g N_Y_c_762_n 0.0122203f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_385 B1 N_Y_c_762_n 0.0235495f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_386 N_B1_c_404_n N_Y_c_762_n 5.54777e-19 $X=8.135 $Y=1.515 $X2=0 $Y2=0
cc_387 N_B1_M1027_g N_VGND_c_889_n 0.00434272f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_388 N_B1_M1023_g N_VGND_c_890_n 0.00825748f $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_389 N_B1_M1027_g N_VGND_c_890_n 0.00828694f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_390 N_B1_M1023_g N_VGND_c_893_n 0.00434272f $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_391 N_B1_M1023_g N_VGND_c_894_n 0.00628433f $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_392 N_B1_M1027_g N_VGND_c_894_n 0.00772874f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_393 N_B1_M1023_g N_A_475_74#_c_970_n 3.238e-19 $X=6.89 $Y=0.74 $X2=0 $Y2=0
cc_394 N_A_27_368#_c_476_n N_VPWR_M1008_d 0.00314376f $X=1.065 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_395 N_A_27_368#_c_480_n N_VPWR_M1011_d 0.00314376f $X=1.915 $Y=2.035 $X2=0
+ $Y2=0
cc_396 N_A_27_368#_c_490_n N_VPWR_M1014_s 0.004128f $X=2.865 $Y=2.05 $X2=0 $Y2=0
cc_397 N_A_27_368#_c_498_n N_VPWR_M1019_s 0.00410979f $X=3.865 $Y=2.035 $X2=0
+ $Y2=0
cc_398 N_A_27_368#_c_518_n N_VPWR_M1002_s 0.00518551f $X=4.865 $Y=2.61 $X2=0
+ $Y2=0
cc_399 N_A_27_368#_c_510_n N_VPWR_M1017_s 0.00537357f $X=6.345 $Y=2.375 $X2=0
+ $Y2=0
cc_400 N_A_27_368#_c_465_n N_VPWR_c_584_n 0.0266615f $X=0.28 $Y=2.435 $X2=0
+ $Y2=0
cc_401 N_A_27_368#_c_476_n N_VPWR_c_584_n 0.0170259f $X=1.065 $Y=2.035 $X2=0
+ $Y2=0
cc_402 N_A_27_368#_c_480_n N_VPWR_c_585_n 0.0170259f $X=1.915 $Y=2.035 $X2=0
+ $Y2=0
cc_403 N_A_27_368#_c_490_n N_VPWR_c_586_n 0.0191372f $X=2.865 $Y=2.05 $X2=0
+ $Y2=0
cc_404 N_A_27_368#_c_467_n N_VPWR_c_586_n 0.0255552f $X=3.03 $Y=2.815 $X2=0
+ $Y2=0
cc_405 N_A_27_368#_c_467_n N_VPWR_c_587_n 0.0266809f $X=3.03 $Y=2.815 $X2=0
+ $Y2=0
cc_406 N_A_27_368#_c_498_n N_VPWR_c_587_n 0.0189268f $X=3.865 $Y=2.035 $X2=0
+ $Y2=0
cc_407 N_A_27_368#_c_472_n N_VPWR_c_587_n 0.0203021f $X=4.03 $Y=2.44 $X2=0 $Y2=0
cc_408 N_A_27_368#_c_472_n N_VPWR_c_588_n 0.0139233f $X=4.03 $Y=2.44 $X2=0 $Y2=0
cc_409 N_A_27_368#_c_518_n N_VPWR_c_588_n 0.0189268f $X=4.865 $Y=2.61 $X2=0
+ $Y2=0
cc_410 N_A_27_368#_c_510_n N_VPWR_c_589_n 0.0208278f $X=6.345 $Y=2.375 $X2=0
+ $Y2=0
cc_411 N_A_27_368#_c_469_n N_VPWR_c_589_n 0.0119238f $X=6.675 $Y=2.99 $X2=0
+ $Y2=0
cc_412 N_A_27_368#_c_547_p N_VPWR_c_590_n 0.00751346f $X=2.08 $Y=2.365 $X2=0
+ $Y2=0
cc_413 N_A_27_368#_c_465_n N_VPWR_c_592_n 0.0124046f $X=0.28 $Y=2.435 $X2=0
+ $Y2=0
cc_414 N_A_27_368#_c_549_p N_VPWR_c_593_n 0.00712457f $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_415 N_A_27_368#_c_467_n N_VPWR_c_594_n 0.0144623f $X=3.03 $Y=2.815 $X2=0
+ $Y2=0
cc_416 N_A_27_368#_c_472_n N_VPWR_c_595_n 0.014549f $X=4.03 $Y=2.44 $X2=0 $Y2=0
cc_417 N_A_27_368#_c_521_n N_VPWR_c_596_n 0.0273216f $X=5.675 $Y=2.61 $X2=0
+ $Y2=0
cc_418 N_A_27_368#_c_468_n N_VPWR_c_597_n 0.0439895f $X=7.375 $Y=2.99 $X2=0
+ $Y2=0
cc_419 N_A_27_368#_c_469_n N_VPWR_c_597_n 0.0235512f $X=6.675 $Y=2.99 $X2=0
+ $Y2=0
cc_420 N_A_27_368#_c_470_n N_VPWR_c_597_n 0.0620536f $X=8.255 $Y=2.99 $X2=0
+ $Y2=0
cc_421 N_A_27_368#_c_473_n N_VPWR_c_597_n 0.0143373f $X=7.475 $Y=2.99 $X2=0
+ $Y2=0
cc_422 N_A_27_368#_c_465_n N_VPWR_c_583_n 0.0102675f $X=0.28 $Y=2.435 $X2=0
+ $Y2=0
cc_423 N_A_27_368#_c_549_p N_VPWR_c_583_n 0.00818839f $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_424 N_A_27_368#_c_547_p N_VPWR_c_583_n 0.00826681f $X=2.08 $Y=2.365 $X2=0
+ $Y2=0
cc_425 N_A_27_368#_c_467_n N_VPWR_c_583_n 0.0118344f $X=3.03 $Y=2.815 $X2=0
+ $Y2=0
cc_426 N_A_27_368#_c_468_n N_VPWR_c_583_n 0.0246728f $X=7.375 $Y=2.99 $X2=0
+ $Y2=0
cc_427 N_A_27_368#_c_469_n N_VPWR_c_583_n 0.0126924f $X=6.675 $Y=2.99 $X2=0
+ $Y2=0
cc_428 N_A_27_368#_c_470_n N_VPWR_c_583_n 0.0344172f $X=8.255 $Y=2.99 $X2=0
+ $Y2=0
cc_429 N_A_27_368#_c_472_n N_VPWR_c_583_n 0.0119743f $X=4.03 $Y=2.44 $X2=0 $Y2=0
cc_430 N_A_27_368#_c_521_n N_VPWR_c_583_n 0.0287492f $X=5.675 $Y=2.61 $X2=0
+ $Y2=0
cc_431 N_A_27_368#_c_473_n N_VPWR_c_583_n 0.00777554f $X=7.475 $Y=2.99 $X2=0
+ $Y2=0
cc_432 N_A_27_368#_c_468_n N_Y_M1001_d 0.00187091f $X=7.375 $Y=2.99 $X2=0 $Y2=0
cc_433 N_A_27_368#_c_470_n N_Y_M1007_d 0.00165831f $X=8.255 $Y=2.99 $X2=0 $Y2=0
cc_434 N_A_27_368#_M1006_d N_Y_c_712_n 0.0181255f $X=4.845 $Y=1.84 $X2=0 $Y2=0
cc_435 N_A_27_368#_M1018_d N_Y_c_712_n 0.00391812f $X=6.375 $Y=1.84 $X2=0 $Y2=0
cc_436 N_A_27_368#_c_512_n N_Y_c_712_n 0.0173758f $X=6.51 $Y=2.46 $X2=0 $Y2=0
cc_437 N_A_27_368#_c_518_n N_Y_c_712_n 0.106798f $X=4.865 $Y=2.61 $X2=0 $Y2=0
cc_438 N_A_27_368#_c_502_n N_Y_c_718_n 0.01102f $X=4.03 $Y=2.12 $X2=0 $Y2=0
cc_439 N_A_27_368#_c_518_n N_Y_c_718_n 0.0150788f $X=4.865 $Y=2.61 $X2=0 $Y2=0
cc_440 N_A_27_368#_M1004_s N_Y_c_749_n 0.00314376f $X=7.325 $Y=1.84 $X2=0 $Y2=0
cc_441 N_A_27_368#_c_576_p N_Y_c_749_n 0.0126919f $X=7.46 $Y=2.455 $X2=0 $Y2=0
cc_442 N_A_27_368#_c_512_n N_Y_c_733_n 0.0143399f $X=6.51 $Y=2.46 $X2=0 $Y2=0
cc_443 N_A_27_368#_c_513_n N_Y_c_733_n 0.0188059f $X=6.51 $Y=2.905 $X2=0 $Y2=0
cc_444 N_A_27_368#_c_468_n N_Y_c_733_n 0.0160291f $X=7.375 $Y=2.99 $X2=0 $Y2=0
cc_445 N_A_27_368#_c_470_n N_Y_c_762_n 0.0159318f $X=8.255 $Y=2.99 $X2=0 $Y2=0
cc_446 N_A_27_368#_c_466_n N_A_30_74#_c_814_n 0.00219923f $X=2.08 $Y=2.15 $X2=0
+ $Y2=0
cc_447 N_A_27_368#_c_466_n N_A_30_74#_c_818_n 0.00893125f $X=2.08 $Y=2.15 $X2=0
+ $Y2=0
cc_448 N_VPWR_M1017_s N_Y_c_712_n 0.00580794f $X=5.825 $Y=1.84 $X2=0 $Y2=0
cc_449 N_VPWR_M1002_s N_Y_c_718_n 0.00382469f $X=4.345 $Y=1.84 $X2=0 $Y2=0
cc_450 N_VPWR_M1002_s Y 0.00127105f $X=4.345 $Y=1.84 $X2=0 $Y2=0
cc_451 N_Y_c_699_n N_A_30_74#_c_815_n 0.0120611f $X=4.567 $Y=1.18 $X2=0 $Y2=0
cc_452 N_Y_c_699_n N_A_30_74#_c_816_n 0.0163927f $X=4.567 $Y=1.18 $X2=0 $Y2=0
cc_453 N_Y_c_697_n N_VGND_M1023_s 0.0146426f $X=8.195 $Y=1.095 $X2=0 $Y2=0
cc_454 N_Y_c_698_n N_VGND_c_889_n 0.0145639f $X=8.36 $Y=0.515 $X2=0 $Y2=0
cc_455 N_Y_c_696_n N_VGND_c_890_n 0.0119984f $X=6.675 $Y=0.515 $X2=0 $Y2=0
cc_456 N_Y_c_698_n N_VGND_c_890_n 0.0119984f $X=8.36 $Y=0.515 $X2=0 $Y2=0
cc_457 N_Y_c_696_n N_VGND_c_893_n 0.0145639f $X=6.675 $Y=0.515 $X2=0 $Y2=0
cc_458 N_Y_c_696_n N_VGND_c_894_n 0.0193213f $X=6.675 $Y=0.515 $X2=0 $Y2=0
cc_459 N_Y_c_697_n N_VGND_c_894_n 0.0802727f $X=8.195 $Y=1.095 $X2=0 $Y2=0
cc_460 N_Y_c_698_n N_VGND_c_894_n 0.0193213f $X=8.36 $Y=0.515 $X2=0 $Y2=0
cc_461 N_Y_c_694_n N_A_475_74#_M1000_s 0.00757665f $X=5.51 $Y=1.072 $X2=0 $Y2=0
cc_462 N_Y_c_695_n N_A_475_74#_M1024_s 0.00176461f $X=6.51 $Y=1.095 $X2=0 $Y2=0
cc_463 N_Y_M1000_d N_A_475_74#_c_969_n 0.00307175f $X=4.37 $Y=0.82 $X2=0 $Y2=0
cc_464 N_Y_c_694_n N_A_475_74#_c_969_n 0.00528925f $X=5.51 $Y=1.072 $X2=0 $Y2=0
cc_465 N_Y_c_699_n N_A_475_74#_c_969_n 0.0115653f $X=4.567 $Y=1.18 $X2=0 $Y2=0
cc_466 N_Y_c_694_n N_A_475_74#_c_980_n 0.0266194f $X=5.51 $Y=1.072 $X2=0 $Y2=0
cc_467 N_Y_c_720_n N_A_475_74#_c_980_n 0.0117291f $X=5.675 $Y=0.76 $X2=0 $Y2=0
cc_468 N_Y_c_699_n N_A_475_74#_c_980_n 0.00145033f $X=4.567 $Y=1.18 $X2=0 $Y2=0
cc_469 N_Y_M1005_d N_A_475_74#_c_970_n 0.00250873f $X=5.535 $Y=0.37 $X2=0 $Y2=0
cc_470 N_Y_c_694_n N_A_475_74#_c_970_n 0.00528925f $X=5.51 $Y=1.072 $X2=0 $Y2=0
cc_471 N_Y_c_720_n N_A_475_74#_c_970_n 0.0194097f $X=5.675 $Y=0.76 $X2=0 $Y2=0
cc_472 N_Y_c_695_n N_A_475_74#_c_970_n 0.00304353f $X=6.51 $Y=1.095 $X2=0 $Y2=0
cc_473 N_Y_c_696_n N_A_475_74#_c_970_n 0.00395312f $X=6.675 $Y=0.515 $X2=0 $Y2=0
cc_474 N_Y_c_695_n N_A_475_74#_c_985_n 0.0168694f $X=6.51 $Y=1.095 $X2=0 $Y2=0
cc_475 N_A_30_74#_c_809_n N_VGND_M1015_s 0.00176461f $X=1.07 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_476 N_A_30_74#_c_812_n N_VGND_M1028_s 0.00250873f $X=1.92 $Y=1.095 $X2=0
+ $Y2=0
cc_477 N_A_30_74#_c_808_n N_VGND_c_885_n 0.0182902f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_478 N_A_30_74#_c_809_n N_VGND_c_885_n 0.0170777f $X=1.07 $Y=1.095 $X2=0 $Y2=0
cc_479 N_A_30_74#_c_811_n N_VGND_c_885_n 0.0182488f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_480 N_A_30_74#_c_811_n N_VGND_c_886_n 0.0182488f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_481 N_A_30_74#_c_812_n N_VGND_c_886_n 0.0209867f $X=1.92 $Y=1.095 $X2=0 $Y2=0
cc_482 N_A_30_74#_c_813_n N_VGND_c_886_n 0.0199619f $X=2.085 $Y=0.495 $X2=0
+ $Y2=0
cc_483 N_A_30_74#_c_808_n N_VGND_c_887_n 0.011066f $X=0.295 $Y=0.515 $X2=0 $Y2=0
cc_484 N_A_30_74#_c_811_n N_VGND_c_888_n 0.00749631f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_485 N_A_30_74#_c_808_n N_VGND_c_890_n 0.00915947f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_486 N_A_30_74#_c_811_n N_VGND_c_890_n 0.0062048f $X=1.155 $Y=0.515 $X2=0
+ $Y2=0
cc_487 N_A_30_74#_c_813_n N_VGND_c_890_n 0.00915345f $X=2.085 $Y=0.495 $X2=0
+ $Y2=0
cc_488 N_A_30_74#_c_813_n N_VGND_c_893_n 0.0119552f $X=2.085 $Y=0.495 $X2=0
+ $Y2=0
cc_489 N_A_30_74#_c_814_n N_A_475_74#_M1003_d 0.00187091f $X=2.825 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_490 N_A_30_74#_c_815_n N_A_475_74#_M1022_d 0.00358162f $X=3.79 $Y=1.095 $X2=0
+ $Y2=0
cc_491 N_A_30_74#_c_814_n N_A_475_74#_c_974_n 0.0159089f $X=2.825 $Y=1.095 $X2=0
+ $Y2=0
cc_492 N_A_30_74#_M1012_s N_A_475_74#_c_967_n 0.00176461f $X=2.815 $Y=0.37 $X2=0
+ $Y2=0
cc_493 N_A_30_74#_c_814_n N_A_475_74#_c_967_n 0.0036669f $X=2.825 $Y=1.095 $X2=0
+ $Y2=0
cc_494 N_A_30_74#_c_842_n N_A_475_74#_c_967_n 0.014143f $X=2.955 $Y=0.76 $X2=0
+ $Y2=0
cc_495 N_A_30_74#_c_815_n N_A_475_74#_c_967_n 0.00304353f $X=3.79 $Y=1.095 $X2=0
+ $Y2=0
cc_496 N_A_30_74#_c_813_n N_A_475_74#_c_968_n 0.0053216f $X=2.085 $Y=0.495 $X2=0
+ $Y2=0
cc_497 N_A_30_74#_c_815_n N_A_475_74#_c_1011_n 0.0245926f $X=3.79 $Y=1.095 $X2=0
+ $Y2=0
cc_498 N_A_30_74#_M1026_s N_A_475_74#_c_969_n 0.00226085f $X=3.815 $Y=0.37 $X2=0
+ $Y2=0
cc_499 N_A_30_74#_c_815_n N_A_475_74#_c_969_n 0.00304353f $X=3.79 $Y=1.095 $X2=0
+ $Y2=0
cc_500 N_A_30_74#_c_816_n N_A_475_74#_c_969_n 0.0203911f $X=3.955 $Y=0.76 $X2=0
+ $Y2=0
cc_501 N_VGND_c_890_n N_A_475_74#_c_967_n 0.0225014f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_c_893_n N_A_475_74#_c_967_n 0.039974f $X=7.01 $Y=0.377 $X2=0 $Y2=0
cc_503 N_VGND_c_886_n N_A_475_74#_c_968_n 0.00238834f $X=1.585 $Y=0.675 $X2=0
+ $Y2=0
cc_504 N_VGND_c_890_n N_A_475_74#_c_968_n 0.0116972f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_505 N_VGND_c_893_n N_A_475_74#_c_968_n 0.0215329f $X=7.01 $Y=0.377 $X2=0
+ $Y2=0
cc_506 N_VGND_c_890_n N_A_475_74#_c_969_n 0.0480679f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_893_n N_A_475_74#_c_969_n 0.0837785f $X=7.01 $Y=0.377 $X2=0
+ $Y2=0
cc_508 N_VGND_c_890_n N_A_475_74#_c_970_n 0.0393024f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_893_n N_A_475_74#_c_970_n 0.0703543f $X=7.01 $Y=0.377 $X2=0
+ $Y2=0
cc_510 N_VGND_c_894_n N_A_475_74#_c_970_n 0.00292855f $X=8.025 $Y=0.377 $X2=0
+ $Y2=0
cc_511 N_VGND_c_890_n N_A_475_74#_c_971_n 0.0127797f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_893_n N_A_475_74#_c_971_n 0.023391f $X=7.01 $Y=0.377 $X2=0 $Y2=0
cc_513 N_VGND_c_890_n N_A_475_74#_c_972_n 0.0127537f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_893_n N_A_475_74#_c_972_n 0.0232521f $X=7.01 $Y=0.377 $X2=0
+ $Y2=0

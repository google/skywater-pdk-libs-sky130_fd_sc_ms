* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.016e+12p pd=1.704e+07u as=1.7584e+12p ps=1.21e+07u
M1001 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_709_74# A3 a_512_74# VNB nlowvt w=740000u l=150000u
+  ad=6.438e+11p pd=6.18e+06u as=4.144e+11p ps=4.08e+06u
M1005 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1008 VPWR A4 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_239_74# A2 a_512_74# VNB nlowvt w=740000u l=150000u
+  ad=6.808e+11p pd=6.28e+06u as=0p ps=0u
M1011 Y A1 a_239_74# VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1012 a_27_368# A4 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.069e+11p ps=4.33e+06u
M1014 a_709_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A4 a_709_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_512_74# A2 a_239_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_512_74# A3 a_709_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_239_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__dlclkp_2.pex.spice
* Created: Fri Aug 28 17:26:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%A_83_244# 1 2 9 13 15 16 18 19 21 23 24 26
+ 28 30 32 36 39
c90 36 0 1.23149e-19 $X=0.6 $Y=1.385
c91 18 0 5.08129e-20 $X=1.535 $Y=2.035
r92 36 40 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.385
+ $X2=0.59 $Y2=1.55
r93 36 39 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.385
+ $X2=0.59 $Y2=1.22
r94 35 37 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=1.385
+ $X2=0.61 $Y2=1.55
r95 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r96 32 35 6.25612 $w=3.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.61 $Y=1.195
+ $X2=0.61 $Y2=1.385
r97 28 30 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=1.705 $Y=2.715
+ $X2=2.24 $Y2=2.715
r98 24 26 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.56 $Y=0.785
+ $X2=1.985 $Y2=0.785
r99 23 28 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=2.55
+ $X2=1.705 $Y2=2.715
r100 22 23 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.55
r101 20 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=0.95
+ $X2=1.56 $Y2=0.785
r102 20 21 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.475 $Y=0.95
+ $X2=1.475 $Y2=1.11
r103 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.62 $Y2=2.12
r104 18 19 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=0.785 $Y2=2.035
r105 17 32 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.785 $Y=1.195
+ $X2=0.61 $Y2=1.195
r106 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.39 $Y=1.195
+ $X2=1.475 $Y2=1.11
r107 16 17 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.39 $Y=1.195
+ $X2=0.785 $Y2=1.195
r108 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.95
+ $X2=0.785 $Y2=2.035
r109 15 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.7 $Y=1.95 $X2=0.7
+ $Y2=1.55
r110 13 39 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.22
r111 9 40 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.55
r112 2 30 300 $w=1.7e-07 $l=9.67574e-07 $layer=licon1_PDIFF $count=2 $X=1.755
+ $Y=1.96 $X2=2.24 $Y2=2.715
r113 1 26 182 $w=1.7e-07 $l=5.29268e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.37 $X2=1.985 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%GATE 3 7 9 12
c39 9 0 1.23149e-19 $X=1.2 $Y=1.665
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.78
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.45
r42 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r43 7 14 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.26 $Y=0.69 $X2=1.26
+ $Y2=1.45
r44 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.245 $Y=2.46
+ $X2=1.245 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%A_315_48# 1 2 7 9 12 14 16 19 21 25 27 29
+ 30 33 36 45 46 51 52 53 55 60 62 64 66 67 77
c148 51 0 5.08129e-20 $X=2.39 $Y=2.215
c149 36 0 1.73462e-19 $X=4.43 $Y=0.74
c150 30 0 1.92985e-19 $X=3.155 $Y=2.135
c151 7 0 1.30966e-19 $X=1.65 $Y=1.12
r152 66 67 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=4.377 $Y=2.24
+ $X2=4.377 $Y2=2.075
r153 63 67 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=1.885
+ $X2=4.295 $Y2=2.075
r154 62 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.295 $Y=1.555
+ $X2=4.295 $Y2=1.275
r155 61 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.16 $Y=1.72 $X2=4.16
+ $Y2=1.63
r156 60 63 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.187 $Y=1.72
+ $X2=4.187 $Y2=1.885
r157 60 62 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.187 $Y=1.72
+ $X2=4.187 $Y2=1.555
r158 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.16
+ $Y=1.72 $X2=4.16 $Y2=1.72
r159 55 58 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=1.72
+ $X2=3.32 $Y2=1.885
r160 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.72 $X2=3.32 $Y2=1.72
r161 51 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=2.215
+ $X2=2.39 $Y2=2.38
r162 50 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.215
+ $X2=2.555 $Y2=2.215
r163 50 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.215
+ $X2=2.225 $Y2=2.215
r164 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=2.215 $X2=2.39 $Y2=2.215
r165 46 70 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.88 $Y=1.285
+ $X2=1.65 $Y2=1.285
r166 45 48 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.887 $Y=1.285
+ $X2=1.887 $Y2=1.45
r167 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.285 $X2=1.88 $Y2=1.285
r168 34 64 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=4.402 $Y=1.083
+ $X2=4.402 $Y2=1.275
r169 34 36 10.2672 $w=3.83e-07 $l=3.43e-07 $layer=LI1_cond $X=4.402 $Y=1.083
+ $X2=4.402 $Y2=0.74
r170 33 58 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=2.05
+ $X2=3.24 $Y2=1.885
r171 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.155 $Y=2.135
+ $X2=3.24 $Y2=2.05
r172 30 53 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.155 $Y=2.135
+ $X2=2.555 $Y2=2.135
r173 29 52 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.045 $Y=2.135
+ $X2=2.225 $Y2=2.135
r174 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.96 $Y=2.05
+ $X2=2.045 $Y2=2.135
r175 27 48 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.96 $Y=2.05 $X2=1.96
+ $Y2=1.45
r176 25 56 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.505 $Y=1.72
+ $X2=3.32 $Y2=1.72
r177 23 25 24.2346 $w=1.79e-07 $l=9e-08 $layer=POLY_cond $X=3.617 $Y=1.63
+ $X2=3.617 $Y2=1.72
r178 22 23 7.00825 $w=1.5e-07 $l=1.13e-07 $layer=POLY_cond $X=3.73 $Y=1.63
+ $X2=3.617 $Y2=1.63
r179 21 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.63
+ $X2=4.16 $Y2=1.63
r180 21 22 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.995 $Y=1.63
+ $X2=3.73 $Y2=1.63
r181 17 23 21.602 $w=1.79e-07 $l=9.20598e-08 $layer=POLY_cond $X=3.655 $Y=1.555
+ $X2=3.617 $Y2=1.63
r182 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.655 $Y=1.555
+ $X2=3.655 $Y2=0.995
r183 14 25 84.35 $w=1.8e-07 $l=3.25814e-07 $layer=POLY_cond $X=3.595 $Y=2.035
+ $X2=3.617 $Y2=1.72
r184 14 16 135.228 $w=1.8e-07 $l=5.05e-07 $layer=POLY_cond $X=3.595 $Y=2.035
+ $X2=3.595 $Y2=2.54
r185 12 76 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.465 $Y=2.75
+ $X2=2.465 $Y2=2.38
r186 7 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.12
+ $X2=1.65 $Y2=1.285
r187 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.65 $Y=1.12 $X2=1.65
+ $Y2=0.69
r188 2 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.235
+ $Y=2.095 $X2=4.38 $Y2=2.24
r189 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.285
+ $Y=0.595 $X2=4.43 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%A_315_338# 1 2 7 9 10 11 14 18 19 21 22 27
+ 31 33 34
c96 27 0 2.51472e-19 $X=3.82 $Y=2.265
c97 19 0 1.92985e-19 $X=2.42 $Y=1.675
r98 29 33 3.70735 $w=2.5e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.87 $Y=1.215
+ $X2=3.845 $Y2=1.3
r99 29 31 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.87 $Y=1.215
+ $X2=3.87 $Y2=0.77
r100 27 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=2.265
+ $X2=3.82 $Y2=2.1
r101 23 33 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.74 $Y=1.385
+ $X2=3.845 $Y2=1.3
r102 23 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.74 $Y=1.385
+ $X2=3.74 $Y2=2.1
r103 21 33 2.76166 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.655 $Y=1.3
+ $X2=3.845 $Y2=1.3
r104 21 22 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.655 $Y=1.3
+ $X2=2.585 $Y2=1.3
r105 19 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.42 $Y=1.675
+ $X2=2.42 $Y2=1.765
r106 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.675
+ $X2=2.42 $Y2=1.51
r107 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.675 $X2=2.42 $Y2=1.675
r108 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.42 $Y=1.385
+ $X2=2.585 $Y2=1.3
r109 16 18 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.42 $Y=1.385
+ $X2=2.42 $Y2=1.675
r110 14 36 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.395 $Y=0.8
+ $X2=2.395 $Y2=1.51
r111 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.765
+ $X2=2.42 $Y2=1.765
r112 10 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.255 $Y=1.765
+ $X2=1.755 $Y2=1.765
r113 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.665 $Y=1.84
+ $X2=1.755 $Y2=1.765
r114 7 9 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=1.665 $Y=1.84
+ $X2=1.665 $Y2=2.46
r115 2 27 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.685
+ $Y=2.12 $X2=3.82 $Y2=2.265
r116 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.73
+ $Y=0.625 $X2=3.87 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%CLK 3 5 7 10 12 14 15 24
c51 15 0 1.30706e-19 $X=5.04 $Y=1.665
c52 12 0 1.73462e-19 $X=5.145 $Y=1.445
r53 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.13 $Y=1.61
+ $X2=5.145 $Y2=1.61
r54 21 23 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=1.61
+ $X2=5.13 $Y2=1.61
r55 19 21 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=4.645 $Y=1.61
+ $X2=5.055 $Y2=1.61
r56 17 19 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.625 $Y=1.61
+ $X2=4.645 $Y2=1.61
r57 15 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.055
+ $Y=1.61 $X2=5.055 $Y2=1.61
r58 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.445
+ $X2=5.145 $Y2=1.61
r59 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.145 $Y=1.445
+ $X2=5.145 $Y2=0.965
r60 8 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.775
+ $X2=5.13 $Y2=1.61
r61 8 10 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.13 $Y=1.775
+ $X2=5.13 $Y2=2.435
r62 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.645 $Y=1.445
+ $X2=4.645 $Y2=1.61
r63 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.645 $Y=1.445
+ $X2=4.645 $Y2=0.965
r64 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.625 $Y=1.775
+ $X2=4.625 $Y2=1.61
r65 1 3 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=4.625 $Y=1.775
+ $X2=4.625 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%A_27_74# 1 2 10 11 13 15 20 23 27 30 36 38
+ 41 42 43 44 46 47 48 54
c127 38 0 1.30966e-19 $X=1.05 $Y=0.855
c128 27 0 1.30706e-19 $X=5.562 $Y=1.56
c129 13 0 1.86939e-19 $X=2.885 $Y=2.75
c130 11 0 6.45334e-20 $X=2.885 $Y=2.215
r131 52 57 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.977 $Y=0.42
+ $X2=2.977 $Y2=0.585
r132 52 54 37.9425 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=2.977 $Y=0.42
+ $X2=2.977 $Y2=0.18
r133 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=0.42 $X2=2.995 $Y2=0.42
r134 48 51 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.995 $Y=0.34
+ $X2=2.995 $Y2=0.42
r135 46 47 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=1.82
r136 42 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=0.34
+ $X2=2.995 $Y2=0.34
r137 42 43 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.83 $Y=0.34
+ $X2=1.22 $Y2=0.34
r138 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=0.425
+ $X2=1.22 $Y2=0.34
r139 40 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.135 $Y=0.425
+ $X2=1.135 $Y2=0.77
r140 39 44 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=0.855
+ $X2=0.23 $Y2=0.855
r141 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=0.855
+ $X2=1.135 $Y2=0.77
r142 38 39 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.05 $Y=0.855
+ $X2=0.365 $Y2=0.855
r143 34 46 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=1.985
r144 34 36 27.0001 $w=3.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=2.815
r145 32 44 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.18 $Y=0.94
+ $X2=0.23 $Y2=0.855
r146 32 47 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.18 $Y=0.94
+ $X2=0.18 $Y2=1.82
r147 28 44 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=0.77
+ $X2=0.23 $Y2=0.855
r148 28 30 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.23 $Y=0.77
+ $X2=0.23 $Y2=0.645
r149 26 27 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.562 $Y=1.41
+ $X2=5.562 $Y2=1.56
r150 23 27 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=5.605 $Y=2.435
+ $X2=5.605 $Y2=1.56
r151 20 26 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.505 $Y=0.965
+ $X2=5.505 $Y2=1.41
r152 17 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.505 $Y=0.255
+ $X2=5.505 $Y2=0.965
r153 16 54 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.16 $Y=0.18
+ $X2=2.977 $Y2=0.18
r154 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=5.505 $Y2=0.255
r155 15 16 1163.98 $w=1.5e-07 $l=2.27e-06 $layer=POLY_cond $X=5.43 $Y=0.18
+ $X2=3.16 $Y2=0.18
r156 11 25 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.885 $Y=2.215
+ $X2=2.885 $Y2=2.125
r157 11 13 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=2.885 $Y=2.215
+ $X2=2.885 $Y2=2.75
r158 10 25 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.87 $Y=0.905
+ $X2=2.87 $Y2=2.125
r159 10 57 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.87 $Y=0.905
+ $X2=2.87 $Y2=0.585
r160 2 46 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r161 2 36 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r162 1 30 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%A_1044_387# 1 2 7 8 11 15 17 21 23 25 27 28
+ 31 37 40 41 46 47
r70 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.14
+ $Y=1.105 $X2=6.14 $Y2=1.105
r71 44 46 7.49781 $w=6.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.72 $Y=1.275
+ $X2=6.14 $Y2=1.275
r72 42 44 4.37372 $w=6.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.475 $Y=1.275
+ $X2=5.72 $Y2=1.275
r73 40 41 7.81132 $w=3.43e-07 $l=1.45e-07 $layer=LI1_cond $X=5.387 $Y=2.095
+ $X2=5.387 $Y2=1.95
r74 35 44 4.89075 $w=3.3e-07 $l=3.35e-07 $layer=LI1_cond $X=5.72 $Y=0.94
+ $X2=5.72 $Y2=1.275
r75 35 37 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=5.72 $Y=0.94 $X2=5.72
+ $Y2=0.74
r76 33 42 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.475 $Y=1.61
+ $X2=5.475 $Y2=1.275
r77 33 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.475 $Y=1.61
+ $X2=5.475 $Y2=1.95
r78 29 40 0.901912 $w=3.43e-07 $l=2.7e-08 $layer=LI1_cond $X=5.387 $Y=2.122
+ $X2=5.387 $Y2=2.095
r79 29 31 22.9821 $w=3.43e-07 $l=6.88e-07 $layer=LI1_cond $X=5.387 $Y=2.122
+ $X2=5.387 $Y2=2.81
r80 26 47 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.14 $Y=1.37
+ $X2=6.14 $Y2=1.105
r81 23 28 27.536 $w=1.65e-07 $l=1.26491e-07 $layer=POLY_cond $X=7.185 $Y=1.31
+ $X2=7.085 $Y2=1.37
r82 23 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.185 $Y=1.31
+ $X2=7.185 $Y2=0.83
r83 19 28 27.536 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=7.175 $Y=1.61
+ $X2=7.085 $Y2=1.37
r84 19 21 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=7.175 $Y=1.61
+ $X2=7.175 $Y2=2.4
r85 18 27 7.86782 $w=2.4e-07 $l=9.8e-08 $layer=POLY_cond $X=6.83 $Y=1.49
+ $X2=6.732 $Y2=1.49
r86 17 28 0.138649 $w=2.4e-07 $l=1.2e-07 $layer=POLY_cond $X=7.085 $Y=1.49
+ $X2=7.085 $Y2=1.37
r87 17 18 65.9955 $w=2.4e-07 $l=2.55e-07 $layer=POLY_cond $X=7.085 $Y=1.49
+ $X2=6.83 $Y2=1.49
r88 13 27 16.8416 $w=1.5e-07 $l=1.30996e-07 $layer=POLY_cond $X=6.755 $Y=1.37
+ $X2=6.732 $Y2=1.49
r89 13 15 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.755 $Y=1.37
+ $X2=6.755 $Y2=0.83
r90 9 27 16.8416 $w=1.8e-07 $l=1.2345e-07 $layer=POLY_cond $X=6.725 $Y=1.61
+ $X2=6.732 $Y2=1.49
r91 9 11 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=6.725 $Y=1.61
+ $X2=6.725 $Y2=2.4
r92 8 26 27.8133 $w=2.4e-07 $l=2.16852e-07 $layer=POLY_cond $X=6.305 $Y=1.49
+ $X2=6.14 $Y2=1.37
r93 7 27 7.86782 $w=2.4e-07 $l=9.7e-08 $layer=POLY_cond $X=6.635 $Y=1.49
+ $X2=6.732 $Y2=1.49
r94 7 8 85.4059 $w=2.4e-07 $l=3.3e-07 $layer=POLY_cond $X=6.635 $Y=1.49
+ $X2=6.305 $Y2=1.49
r95 2 40 400 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.935 $X2=5.38 $Y2=2.095
r96 2 31 400 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.935 $X2=5.38 $Y2=2.81
r97 1 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.58
+ $Y=0.595 $X2=5.72 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%VPWR 1 2 3 4 5 20 24 28 32 36 38 43 44 45
+ 47 62 66 72 75 78 82
r83 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r84 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r85 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r86 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 70 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r88 70 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r90 67 78 15.5458 $w=1.7e-07 $l=4.53e-07 $layer=LI1_cond $X=6.635 $Y=3.33
+ $X2=6.182 $Y2=3.33
r91 67 69 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=3.33
+ $X2=6.96 $Y2=3.33
r92 66 81 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=7.497 $Y2=3.33
r93 66 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=6.96 $Y2=3.33
r94 65 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r95 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r96 62 78 15.5458 $w=1.7e-07 $l=4.52e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=6.182 $Y2=3.33
r97 62 64 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r99 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r100 58 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r102 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r103 55 75 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.215 $Y2=3.33
r104 55 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 54 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 51 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 48 72 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.88 $Y2=3.33
r112 48 50 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.2 $Y2=3.33
r113 47 75 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.215 $Y2=3.33
r114 47 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 45 61 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 45 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 43 60 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.88 $Y2=3.33
r119 42 64 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=4.88 $Y2=3.33
r121 38 41 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.44 $Y=1.985
+ $X2=7.44 $Y2=2.815
r122 36 81 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.497 $Y2=3.33
r123 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.44 $Y2=2.815
r124 32 35 9.36906 $w=9.03e-07 $l=6.95e-07 $layer=LI1_cond $X=6.182 $Y=2.115
+ $X2=6.182 $Y2=2.81
r125 30 78 3.35974 $w=9.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=3.33
r126 30 35 5.86409 $w=9.03e-07 $l=4.35e-07 $layer=LI1_cond $X=6.182 $Y=3.245
+ $X2=6.182 $Y2=2.81
r127 26 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=3.245
+ $X2=4.88 $Y2=3.33
r128 26 28 35.0971 $w=3.28e-07 $l=1.005e-06 $layer=LI1_cond $X=4.88 $Y=3.245
+ $X2=4.88 $Y2=2.24
r129 22 75 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=3.33
r130 22 24 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=3.215 $Y=3.245
+ $X2=3.215 $Y2=2.815
r131 18 72 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=3.33
r132 18 20 25.4128 $w=3.88e-07 $l=8.6e-07 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=2.385
r133 5 41 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.84 $X2=7.4 $Y2=2.815
r134 5 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.84 $X2=7.4 $Y2=1.985
r135 4 35 200 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=3 $X=5.695
+ $Y=1.935 $X2=5.835 $Y2=2.81
r136 4 32 200 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=3 $X=5.695
+ $Y=1.935 $X2=5.835 $Y2=2.115
r137 3 28 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=4.715
+ $Y=2.095 $X2=4.88 $Y2=2.24
r138 2 24 600 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_PDIFF $count=1 $X=2.975
+ $Y=2.54 $X2=3.215 $Y2=2.815
r139 1 20 300 $w=1.7e-07 $l=6.7257e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.88 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%GCLK 1 2 7 8 9 10 11 12 13
r19 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=2.405
+ $X2=6.97 $Y2=2.775
r20 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.97 $Y=1.985
+ $X2=6.97 $Y2=2.405
r21 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.97 $Y=1.665
+ $X2=6.97 $Y2=1.985
r22 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.665
r23 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=0.925 $X2=6.97
+ $Y2=1.295
r24 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.97 $Y=0.555 $X2=6.97
+ $Y2=0.925
r25 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.815
+ $Y=1.84 $X2=6.95 $Y2=2.815
r26 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.815
+ $Y=1.84 $X2=6.95 $Y2=1.985
r27 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.83
+ $Y=0.46 $X2=6.97 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_2%VGND 1 2 3 4 5 18 20 25 28 32 34 36 39 40
+ 43 45 57 64 69 75 78 81 85
r92 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r93 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r96 73 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r97 73 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r98 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r99 70 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.635 $Y=0 $X2=6.47
+ $Y2=0
r100 70 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=0
+ $X2=6.96 $Y2=0
r101 69 84 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.497 $Y2=0
r102 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=6.96 $Y2=0
r103 68 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r104 68 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r105 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r106 65 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=4.93
+ $Y2=0
r107 65 67 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=5.095 $Y=0 $X2=6
+ $Y2=0
r108 64 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6.47
+ $Y2=0
r109 64 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.305 $Y=0 $X2=6
+ $Y2=0
r110 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r111 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r112 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r113 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r114 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.93
+ $Y2=0
r115 57 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r116 56 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r117 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r118 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r119 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r121 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r122 50 75 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.712
+ $Y2=0
r123 50 52 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r124 48 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r125 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r126 45 75 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.712 $Y2=0
r127 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r128 43 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r129 43 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r130 39 55 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.12
+ $Y2=0
r131 39 40 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.437
+ $Y2=0
r132 38 59 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.6
+ $Y2=0
r133 38 40 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.437
+ $Y2=0
r134 34 84 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.497 $Y2=0
r135 34 36 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0.605
r136 30 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0
r137 30 32 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0.605
r138 26 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0
r139 26 28 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.93 $Y=0.085
+ $X2=4.93 $Y2=0.74
r140 25 42 3.91487 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=3.437 $Y=0.755
+ $X2=3.437 $Y2=0.88
r141 24 40 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.437 $Y2=0
r142 24 25 38.1072 $w=1.93e-07 $l=6.7e-07 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.437 $Y2=0.755
r143 20 42 3.03794 $w=2.5e-07 $l=9.7e-08 $layer=LI1_cond $X=3.34 $Y=0.88
+ $X2=3.437 $Y2=0.88
r144 20 22 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.34 $Y=0.88
+ $X2=3.085 $Y2=0.88
r145 16 75 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0
r146 16 18 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0.515
r147 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.26
+ $Y=0.46 $X2=7.4 $Y2=0.605
r148 4 32 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.46 $X2=6.47 $Y2=0.605
r149 3 28 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.72
+ $Y=0.595 $X2=4.93 $Y2=0.74
r150 2 42 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.695 $X2=3.44 $Y2=0.84
r151 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.695 $X2=3.085 $Y2=0.84
r152 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends


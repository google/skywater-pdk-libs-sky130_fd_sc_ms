* File: sky130_fd_sc_ms__a41oi_2.spice
* Created: Wed Sep  2 11:56:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a41oi_2.pex.spice"
.subckt sky130_fd_sc_ms__a41oi_2  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1013 N_Y_M1013_d N_B1_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A1_M1011_g N_A_239_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1011_d N_A1_M1018_g N_A_239_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_A_239_74#_M1018_s N_A2_M1010_g N_A_512_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_A_239_74#_M1016_d N_A2_M1016_g N_A_512_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_709_74#_M1004_d N_A3_M1004_g N_A_512_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_709_74#_M1017_d N_A3_M1017_g N_A_512_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_A_709_74#_M1017_d N_A4_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1015 N_A_709_74#_M1015_d N_A4_M1015_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2257 AS=0.1221 PD=2.09 PS=1.07 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_368#_M1007_d N_B1_M1007_g N_Y_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1009 N_A_27_368#_M1009_d N_B1_M1009_g N_Y_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1002 N_A_27_368#_M1009_d N_A1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.3136 PD=1.44 PS=1.68 NRD=0 NRS=24.625 M=1 R=6.22222 SA=90001.2
+ SB=90003.9 A=0.2016 P=2.6 MULT=1
MM1006 N_A_27_368#_M1006_d N_A1_M1006_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=1.68 NRD=0 NRS=24.625 M=1 R=6.22222 SA=90001.9
+ SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_27_368#_M1006_d N_A2_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.4
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1005 N_A_27_368#_M1005_d N_A2_M1005_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.9
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_27_368#_M1005_d N_A3_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.4
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1003 N_A_27_368#_M1003_d N_A3_M1003_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1988 AS=0.2072 PD=1.475 PS=1.49 NRD=1.7533 NRS=7.8997 M=1 R=6.22222
+ SA=90003.9 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A4_M1008_g N_A_27_368#_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1988 PD=1.39 PS=1.475 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90004.5
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1008_d N_A4_M1012_g N_A_27_368#_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3416 PD=1.39 PS=2.85 NRD=0 NRS=0.8668 M=1 R=6.22222 SA=90004.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX19_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__a41oi_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__and4b_2.spice
* Created: Fri Aug 28 17:14:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4b_2.pex.spice"
.subckt sky130_fd_sc_ms__and4b_2  VNB VPB A_N D C B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_N_M1010_g N_A_27_112#_M1010_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18.54 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.4 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1010_d N_A_186_48#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.144644 AS=0.1036 PD=1.26202 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_186_48#_M1013_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.23495 AS=0.1036 PD=1.375 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1000 A_459_74# N_D_M1000_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.23495 PD=0.98 PS=1.375 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1001 A_537_74# N_C_M1001_g A_459_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0888 PD=1.13 PS=0.98 NRD=22.692 NRS=10.536 M=1 R=4.93333 SA=75002.2
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1008 A_645_74# N_B_M1008_g A_537_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.1443 PD=1.13 PS=1.13 NRD=22.692 NRS=22.692 M=1 R=4.93333 SA=75002.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1012 N_A_186_48#_M1012_d N_A_27_112#_M1012_g A_645_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1443 PD=2.05 PS=1.13 NRD=0 NRS=22.692 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_112#_M1005_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1662 AS=0.2352 PD=1.27286 PS=2.24 NRD=33.49 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003.5 A=0.1512 P=2.04 MULT=1
MM1007 N_X_M1007_d N_A_186_48#_M1007_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2216 PD=1.39 PS=1.69714 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90000.6 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1007_d N_A_186_48#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.255592 PD=1.39 PS=1.6483 NRD=0 NRS=14.0658 M=1 R=6.22222
+ SA=90001.1 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1002 N_A_186_48#_M1002_d N_D_M1002_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.1475 AS=0.228208 PD=1.295 PS=1.4717 NRD=0.9653 NRS=16.7253 M=1 R=5.55556
+ SA=90001.7 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_A_186_48#_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.23305 AS=0.1475 PD=1.53 PS=1.295 NRD=16.7253 NRS=1.9503 M=1 R=5.55556
+ SA=90002.2 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1003 N_A_186_48#_M1003_d N_B_M1003_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.155 AS=0.23305 PD=1.31 PS=1.53 NRD=2.9353 NRS=16.7253 M=1 R=5.55556
+ SA=90002.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_27_112#_M1011_g N_A_186_48#_M1003_d VPB PSHORT L=0.18
+ W=1 AD=0.41835 AS=0.155 PD=2.96 PS=1.31 NRD=18.6953 NRS=2.9353 M=1 R=5.55556
+ SA=90003.3 SB=90000.3 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_43 VNB 0 1.93659e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__and4b_2.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__tap_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__tap_2 VGND VNB VPB VPWR
.ends


* File: sky130_fd_sc_ms__dfstp_4.pxi.spice
* Created: Wed Sep  2 12:03:49 2020
* 
x_PM_SKY130_FD_SC_MS__DFSTP_4%D N_D_c_274_n N_D_M1031_g N_D_M1032_g D D
+ N_D_c_276_n N_D_c_277_n N_D_c_281_n PM_SKY130_FD_SC_MS__DFSTP_4%D
x_PM_SKY130_FD_SC_MS__DFSTP_4%CLK N_CLK_M1035_g N_CLK_M1024_g CLK N_CLK_c_310_n
+ N_CLK_c_311_n PM_SKY130_FD_SC_MS__DFSTP_4%CLK
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_398_74# N_A_398_74#_M1018_d N_A_398_74#_M1027_d
+ N_A_398_74#_M1001_g N_A_398_74#_c_346_n N_A_398_74#_M1013_g
+ N_A_398_74#_M1006_g N_A_398_74#_M1036_g N_A_398_74#_c_348_n
+ N_A_398_74#_c_468_p N_A_398_74#_c_349_n N_A_398_74#_c_350_n
+ N_A_398_74#_c_367_n N_A_398_74#_c_368_n N_A_398_74#_c_351_n
+ N_A_398_74#_c_352_n N_A_398_74#_c_353_n N_A_398_74#_c_354_n
+ N_A_398_74#_c_373_n N_A_398_74#_c_374_n N_A_398_74#_c_375_n
+ N_A_398_74#_c_376_n N_A_398_74#_c_377_n N_A_398_74#_c_378_n
+ N_A_398_74#_c_379_n N_A_398_74#_c_380_n N_A_398_74#_c_355_n
+ N_A_398_74#_c_356_n N_A_398_74#_c_357_n N_A_398_74#_c_358_n
+ N_A_398_74#_c_382_n N_A_398_74#_c_359_n N_A_398_74#_c_360_n
+ N_A_398_74#_c_361_n N_A_398_74#_c_383_n N_A_398_74#_c_362_n
+ N_A_398_74#_c_363_n N_A_398_74#_c_385_n PM_SKY130_FD_SC_MS__DFSTP_4%A_398_74#
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_767_402# N_A_767_402#_M1026_s
+ N_A_767_402#_M1038_d N_A_767_402#_M1010_g N_A_767_402#_c_607_n
+ N_A_767_402#_M1003_g N_A_767_402#_c_608_n N_A_767_402#_c_609_n
+ N_A_767_402#_c_610_n N_A_767_402#_c_615_n N_A_767_402#_c_616_n
+ N_A_767_402#_c_617_n N_A_767_402#_c_611_n N_A_767_402#_c_618_n
+ N_A_767_402#_c_612_n PM_SKY130_FD_SC_MS__DFSTP_4%A_767_402#
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_612_74# N_A_612_74#_M1023_d N_A_612_74#_M1001_d
+ N_A_612_74#_M1038_g N_A_612_74#_c_693_n N_A_612_74#_M1026_g
+ N_A_612_74#_M1033_g N_A_612_74#_M1028_g N_A_612_74#_c_696_n
+ N_A_612_74#_c_697_n N_A_612_74#_c_698_n N_A_612_74#_c_699_n
+ N_A_612_74#_c_709_n N_A_612_74#_c_700_n N_A_612_74#_c_701_n
+ N_A_612_74#_c_702_n N_A_612_74#_c_703_n N_A_612_74#_c_704_n
+ N_A_612_74#_c_705_n N_A_612_74#_c_706_n PM_SKY130_FD_SC_MS__DFSTP_4%A_612_74#
x_PM_SKY130_FD_SC_MS__DFSTP_4%SET_B N_SET_B_M1011_g N_SET_B_M1016_g
+ N_SET_B_c_829_n N_SET_B_M1004_g N_SET_B_c_830_n N_SET_B_c_831_n
+ N_SET_B_M1019_g N_SET_B_c_832_n N_SET_B_c_833_n N_SET_B_c_834_n SET_B
+ N_SET_B_c_836_n N_SET_B_c_837_n N_SET_B_c_838_n
+ PM_SKY130_FD_SC_MS__DFSTP_4%SET_B
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_225_74# N_A_225_74#_M1035_s N_A_225_74#_M1024_s
+ N_A_225_74#_M1018_g N_A_225_74#_M1027_g N_A_225_74#_c_968_n
+ N_A_225_74#_c_956_n N_A_225_74#_c_969_n N_A_225_74#_c_970_n
+ N_A_225_74#_M1023_g N_A_225_74#_M1002_g N_A_225_74#_c_972_n
+ N_A_225_74#_M1025_g N_A_225_74#_c_958_n N_A_225_74#_c_959_n
+ N_A_225_74#_M1015_g N_A_225_74#_c_961_n N_A_225_74#_c_962_n
+ N_A_225_74#_c_963_n N_A_225_74#_c_979_n N_A_225_74#_c_964_n
+ N_A_225_74#_c_981_n N_A_225_74#_c_965_n N_A_225_74#_c_966_n
+ N_A_225_74#_c_983_n PM_SKY130_FD_SC_MS__DFSTP_4%A_225_74#
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_1484_62# N_A_1484_62#_M1005_d
+ N_A_1484_62#_M1012_d N_A_1484_62#_M1007_g N_A_1484_62#_M1014_g
+ N_A_1484_62#_c_1129_n N_A_1484_62#_c_1130_n N_A_1484_62#_c_1144_n
+ N_A_1484_62#_c_1131_n N_A_1484_62#_c_1132_n N_A_1484_62#_c_1136_n
+ N_A_1484_62#_c_1133_n N_A_1484_62#_c_1134_n
+ PM_SKY130_FD_SC_MS__DFSTP_4%A_1484_62#
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_1324_392# N_A_1324_392#_M1006_d
+ N_A_1324_392#_M1025_d N_A_1324_392#_M1019_d N_A_1324_392#_c_1210_n
+ N_A_1324_392#_M1005_g N_A_1324_392#_M1012_g N_A_1324_392#_c_1212_n
+ N_A_1324_392#_M1000_g N_A_1324_392#_c_1223_n N_A_1324_392#_M1020_g
+ N_A_1324_392#_c_1214_n N_A_1324_392#_c_1225_n N_A_1324_392#_M1021_g
+ N_A_1324_392#_c_1215_n N_A_1324_392#_c_1227_n N_A_1324_392#_c_1216_n
+ N_A_1324_392#_c_1228_n N_A_1324_392#_c_1229_n N_A_1324_392#_c_1230_n
+ N_A_1324_392#_c_1231_n N_A_1324_392#_c_1232_n N_A_1324_392#_c_1217_n
+ N_A_1324_392#_c_1218_n N_A_1324_392#_c_1233_n N_A_1324_392#_c_1219_n
+ N_A_1324_392#_c_1220_n N_A_1324_392#_c_1234_n N_A_1324_392#_c_1235_n
+ PM_SKY130_FD_SC_MS__DFSTP_4%A_1324_392#
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_1940_74# N_A_1940_74#_M1000_s
+ N_A_1940_74#_M1020_d N_A_1940_74#_c_1372_n N_A_1940_74#_M1008_g
+ N_A_1940_74#_c_1373_n N_A_1940_74#_c_1374_n N_A_1940_74#_c_1375_n
+ N_A_1940_74#_M1009_g N_A_1940_74#_M1022_g N_A_1940_74#_M1029_g
+ N_A_1940_74#_c_1378_n N_A_1940_74#_M1017_g N_A_1940_74#_M1030_g
+ N_A_1940_74#_c_1380_n N_A_1940_74#_M1034_g N_A_1940_74#_M1037_g
+ N_A_1940_74#_c_1383_n N_A_1940_74#_c_1384_n N_A_1940_74#_c_1385_n
+ N_A_1940_74#_c_1392_n N_A_1940_74#_c_1386_n N_A_1940_74#_c_1387_n
+ PM_SKY130_FD_SC_MS__DFSTP_4%A_1940_74#
x_PM_SKY130_FD_SC_MS__DFSTP_4%A_27_74# N_A_27_74#_M1032_s N_A_27_74#_M1023_s
+ N_A_27_74#_M1031_s N_A_27_74#_M1001_s N_A_27_74#_c_1489_n N_A_27_74#_c_1490_n
+ N_A_27_74#_c_1495_n N_A_27_74#_c_1496_n N_A_27_74#_c_1497_n
+ N_A_27_74#_c_1491_n N_A_27_74#_c_1492_n N_A_27_74#_c_1499_n
+ N_A_27_74#_c_1541_n N_A_27_74#_c_1493_n PM_SKY130_FD_SC_MS__DFSTP_4%A_27_74#
x_PM_SKY130_FD_SC_MS__DFSTP_4%VPWR N_VPWR_M1031_d N_VPWR_M1024_d N_VPWR_M1010_d
+ N_VPWR_M1011_d N_VPWR_M1014_d N_VPWR_M1012_s N_VPWR_M1020_s N_VPWR_M1021_s
+ N_VPWR_M1029_s N_VPWR_M1037_s N_VPWR_c_1559_n N_VPWR_c_1560_n N_VPWR_c_1561_n
+ N_VPWR_c_1562_n N_VPWR_c_1563_n N_VPWR_c_1564_n N_VPWR_c_1565_n
+ N_VPWR_c_1566_n N_VPWR_c_1567_n N_VPWR_c_1568_n N_VPWR_c_1569_n
+ N_VPWR_c_1570_n N_VPWR_c_1571_n N_VPWR_c_1572_n N_VPWR_c_1573_n VPWR
+ N_VPWR_c_1574_n N_VPWR_c_1575_n N_VPWR_c_1576_n N_VPWR_c_1577_n
+ N_VPWR_c_1578_n N_VPWR_c_1579_n N_VPWR_c_1580_n N_VPWR_c_1581_n
+ N_VPWR_c_1582_n N_VPWR_c_1583_n N_VPWR_c_1584_n N_VPWR_c_1585_n
+ N_VPWR_c_1586_n N_VPWR_c_1587_n N_VPWR_c_1588_n N_VPWR_c_1589_n
+ N_VPWR_c_1558_n PM_SKY130_FD_SC_MS__DFSTP_4%VPWR
x_PM_SKY130_FD_SC_MS__DFSTP_4%Q N_Q_M1008_d N_Q_M1017_d N_Q_M1022_d N_Q_M1030_d
+ N_Q_c_1738_n N_Q_c_1739_n N_Q_c_1740_n N_Q_c_1745_n N_Q_c_1746_n N_Q_c_1741_n
+ N_Q_c_1747_n N_Q_c_1742_n N_Q_c_1743_n Q Q Q N_Q_c_1750_n
+ PM_SKY130_FD_SC_MS__DFSTP_4%Q
x_PM_SKY130_FD_SC_MS__DFSTP_4%VGND N_VGND_M1032_d N_VGND_M1035_d N_VGND_M1003_d
+ N_VGND_M1016_d N_VGND_M1004_d N_VGND_M1000_d N_VGND_M1009_s N_VGND_M1034_s
+ N_VGND_c_1810_n N_VGND_c_1811_n N_VGND_c_1812_n N_VGND_c_1813_n
+ N_VGND_c_1814_n N_VGND_c_1815_n N_VGND_c_1816_n N_VGND_c_1817_n
+ N_VGND_c_1818_n N_VGND_c_1819_n N_VGND_c_1820_n VGND N_VGND_c_1821_n
+ N_VGND_c_1822_n N_VGND_c_1823_n N_VGND_c_1824_n N_VGND_c_1825_n
+ N_VGND_c_1826_n N_VGND_c_1827_n N_VGND_c_1828_n N_VGND_c_1829_n
+ N_VGND_c_1830_n N_VGND_c_1831_n N_VGND_c_1832_n N_VGND_c_1833_n
+ PM_SKY130_FD_SC_MS__DFSTP_4%VGND
cc_1 VNB N_D_c_274_n 0.0447809f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_2 VNB N_D_M1032_g 0.0283644f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_276_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_277_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_M1024_g 0.00712101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB CLK 0.00893055f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_7 VNB N_CLK_c_310_n 0.0322418f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_CLK_c_311_n 0.0199457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_398_74#_c_346_n 0.0227081f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A_398_74#_M1013_g 0.0525559f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_11 VNB N_A_398_74#_c_348_n 0.00169421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_398_74#_c_349_n 0.0153888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_398_74#_c_350_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_351_n 0.00190286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_352_n 0.0158101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_353_n 0.00125833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_354_n 0.0174283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_355_n 0.00185717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_356_n 0.00920071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_357_n 0.00225196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_358_n 0.00683192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_359_n 0.00505342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_360_n 0.03212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_361_n 0.00183894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_362_n 0.0136527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_398_74#_c_363_n 0.0192244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_767_402#_c_607_n 0.0191692f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_A_767_402#_c_608_n 0.0117603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_767_402#_c_609_n 0.00887451f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_30 VNB N_A_767_402#_c_610_n 0.0253986f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_31 VNB N_A_767_402#_c_611_n 0.0141708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_767_402#_c_612_n 0.0359736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_612_74#_M1038_g 0.0126793f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_34 VNB N_A_612_74#_c_693_n 0.0192259f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_35 VNB N_A_612_74#_M1033_g 0.00143836f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_36 VNB N_A_612_74#_M1028_g 0.0248687f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_37 VNB N_A_612_74#_c_696_n 0.00472968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_612_74#_c_697_n 0.0145886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_612_74#_c_698_n 0.00935088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_612_74#_c_699_n 0.0176834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_612_74#_c_700_n 0.00276658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_612_74#_c_701_n 0.00220525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_612_74#_c_702_n 0.00959991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_612_74#_c_703_n 0.00438751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_612_74#_c_704_n 0.00189138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_612_74#_c_705_n 0.0325974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_612_74#_c_706_n 0.0434133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_SET_B_M1016_g 0.0426396f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_49 VNB N_SET_B_c_829_n 0.0162437f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_50 VNB N_SET_B_c_830_n 0.0682954f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_51 VNB N_SET_B_c_831_n 0.0198191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SET_B_c_832_n 0.00103492f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_53 VNB N_SET_B_c_833_n 0.0123954f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_54 VNB N_SET_B_c_834_n 0.00109498f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_55 VNB SET_B 0.00124466f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_56 VNB N_SET_B_c_836_n 0.00324757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SET_B_c_837_n 0.00628056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_838_n 0.00233764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_225_74#_M1018_g 0.0251862f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_60 VNB N_A_225_74#_c_956_n 0.0336376f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_61 VNB N_A_225_74#_M1023_g 0.0294306f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_62 VNB N_A_225_74#_c_958_n 0.0103413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_225_74#_c_959_n 8.10579e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_225_74#_M1015_g 0.0515873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_225_74#_c_961_n 0.0124352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_225_74#_c_962_n 0.0269886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_225_74#_c_963_n 0.0195044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_225_74#_c_964_n 0.0115791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_225_74#_c_965_n 0.00374876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_225_74#_c_966_n 0.013166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1484_62#_M1007_g 0.0336842f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_72 VNB N_A_1484_62#_c_1129_n 0.00351864f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.145
cc_73 VNB N_A_1484_62#_c_1130_n 0.0138251f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_74 VNB N_A_1484_62#_c_1131_n 0.00682312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1484_62#_c_1132_n 0.00634625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1484_62#_c_1133_n 0.00805698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1484_62#_c_1134_n 0.0430611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1324_392#_c_1210_n 0.00412849f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_79 VNB N_A_1324_392#_M1005_g 0.0507006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1324_392#_c_1212_n 0.0686098f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.825
cc_81 VNB N_A_1324_392#_M1000_g 0.0297718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1324_392#_c_1214_n 0.0132882f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.825
cc_83 VNB N_A_1324_392#_c_1215_n 0.0141228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1324_392#_c_1216_n 0.00512183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1324_392#_c_1217_n 0.00272086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1324_392#_c_1218_n 0.0240576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1324_392#_c_1219_n 2.14136e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1324_392#_c_1220_n 0.00243428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1940_74#_c_1372_n 0.0181326f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_90 VNB N_A_1940_74#_c_1373_n 0.0145071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1940_74#_c_1374_n 0.00747839f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_92 VNB N_A_1940_74#_c_1375_n 0.0198904f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_93 VNB N_A_1940_74#_M1022_g 5.18122e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_94 VNB N_A_1940_74#_M1029_g 4.78866e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_95 VNB N_A_1940_74#_c_1378_n 0.0203684f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_96 VNB N_A_1940_74#_M1030_g 4.7855e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1940_74#_c_1380_n 0.109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1940_74#_M1034_g 0.0243152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1940_74#_M1037_g 5.20265e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1940_74#_c_1383_n 0.0146895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1940_74#_c_1384_n 0.00151156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1940_74#_c_1385_n 4.11739e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1940_74#_c_1386_n 0.00463811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1940_74#_c_1387_n 0.00402022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_27_74#_c_1489_n 0.0146704f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_106 VNB N_A_27_74#_c_1490_n 0.040185f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_107 VNB N_A_27_74#_c_1491_n 0.00677877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_27_74#_c_1492_n 0.00791533f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_109 VNB N_A_27_74#_c_1493_n 0.0065301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VPWR_c_1558_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_Q_c_1738_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_112 VNB N_Q_c_1739_n 0.00542399f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_113 VNB N_Q_c_1740_n 0.00228436f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_114 VNB N_Q_c_1741_n 0.00280896f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_115 VNB N_Q_c_1742_n 0.00893228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_Q_c_1743_n 0.00372816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB Q 0.0268698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1810_n 0.00766994f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_119 VNB N_VGND_c_1811_n 0.0223817f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_120 VNB N_VGND_c_1812_n 0.00555881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1813_n 0.0166819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1814_n 0.0172166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1815_n 0.00819684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1816_n 0.0118832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1817_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1818_n 0.0297496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1819_n 0.0376041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1820_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1821_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1822_n 0.0561972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1823_n 0.0341238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1824_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1825_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1826_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1827_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1828_n 0.00738258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1829_n 0.0511502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1830_n 0.0397556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1831_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1832_n 0.0127911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1833_n 0.714439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VPB N_D_c_274_n 0.0126446f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_143 VPB N_D_M1031_g 0.0599227f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.73
cc_144 VPB N_D_c_277_n 0.00226531f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_145 VPB N_D_c_281_n 0.0244074f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_146 VPB N_CLK_M1024_g 0.0243587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_398_74#_M1001_g 0.0226528f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_148 VPB N_A_398_74#_c_346_n 0.0166347f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_149 VPB N_A_398_74#_M1036_g 0.0261185f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_150 VPB N_A_398_74#_c_367_n 0.0206876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_398_74#_c_368_n 0.00246275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_398_74#_c_351_n 0.00198249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_398_74#_c_352_n 0.0371759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_398_74#_c_353_n 0.00593785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_398_74#_c_354_n 0.0185024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_398_74#_c_373_n 0.0027728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_398_74#_c_374_n 0.00885541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_398_74#_c_375_n 0.00434119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_398_74#_c_376_n 0.016715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_398_74#_c_377_n 0.00322702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_398_74#_c_378_n 0.00242579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_398_74#_c_379_n 0.00795467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_398_74#_c_380_n 5.72606e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_398_74#_c_355_n 0.00241745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_398_74#_c_382_n 0.00102518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_398_74#_c_383_n 8.45509e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_398_74#_c_362_n 0.00771009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_398_74#_c_385_n 0.039937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_767_402#_M1010_g 0.0207042f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_170 VPB N_A_767_402#_c_610_n 0.0023708f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_171 VPB N_A_767_402#_c_615_n 0.0132551f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_172 VPB N_A_767_402#_c_616_n 0.065417f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_173 VPB N_A_767_402#_c_617_n 0.00267421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_767_402#_c_618_n 0.00597358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_612_74#_M1038_g 0.0444077f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_176 VPB N_A_612_74#_M1033_g 0.0218971f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_177 VPB N_A_612_74#_c_709_n 0.00386855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_612_74#_c_700_n 0.00657325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_SET_B_M1011_g 0.02984f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.99
cc_180 VPB N_SET_B_M1016_g 0.00239435f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_181 VPB N_SET_B_M1019_g 0.0578308f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_182 VPB N_SET_B_c_832_n 0.0209448f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_183 VPB N_SET_B_c_833_n 0.0186138f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_184 VPB N_SET_B_c_834_n 0.0015583f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_185 VPB SET_B 0.00132511f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_186 VPB N_SET_B_c_836_n 0.00640286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_SET_B_c_837_n 0.0348872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_SET_B_c_838_n 0.00327236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_225_74#_M1027_g 0.0204871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_225_74#_c_968_n 0.0705799f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_191 VPB N_A_225_74#_c_969_n 0.0558158f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_192 VPB N_A_225_74#_c_970_n 0.0123683f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_193 VPB N_A_225_74#_M1002_g 0.0345512f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_194 VPB N_A_225_74#_c_972_n 0.227688f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_195 VPB N_A_225_74#_M1025_g 0.0169781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_225_74#_c_958_n 0.0386327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_225_74#_c_959_n 0.00703403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_225_74#_c_961_n 0.00169155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_225_74#_c_962_n 5.35904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_225_74#_c_963_n 0.00573612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_225_74#_c_979_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_225_74#_c_964_n 0.00180372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_225_74#_c_981_n 0.0047582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_225_74#_c_965_n 2.33575e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_225_74#_c_983_n 0.0138824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1484_62#_M1014_g 0.061553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1484_62#_c_1136_n 0.00738766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1484_62#_c_1133_n 0.0181569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1324_392#_c_1210_n 0.0473246f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_210 VPB N_A_1324_392#_M1012_g 0.0262214f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_211 VPB N_A_1324_392#_c_1223_n 0.0175515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1324_392#_c_1214_n 0.0099104f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_213 VPB N_A_1324_392#_c_1225_n 0.0169447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1324_392#_c_1215_n 0.00568743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1324_392#_c_1227_n 0.00276818f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1324_392#_c_1228_n 0.00457775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1324_392#_c_1229_n 0.00959247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1324_392#_c_1230_n 0.00760636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1324_392#_c_1231_n 0.00835114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1324_392#_c_1232_n 0.0133368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1324_392#_c_1233_n 0.0325225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1324_392#_c_1234_n 0.00300345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1324_392#_c_1235_n 0.00509406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1940_74#_M1022_g 0.0238147f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_225 VPB N_A_1940_74#_M1029_g 0.021629f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_226 VPB N_A_1940_74#_M1030_g 0.0216045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1940_74#_M1037_g 0.0246636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1940_74#_c_1392_n 0.0035517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_27_74#_c_1490_n 0.0275147f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_230 VPB N_A_27_74#_c_1495_n 0.02407f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_231 VPB N_A_27_74#_c_1496_n 0.0258928f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_232 VPB N_A_27_74#_c_1497_n 0.0153732f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_233 VPB N_A_27_74#_c_1491_n 0.00245721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_27_74#_c_1499_n 0.0109181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1559_n 0.0136412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1560_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1561_n 0.00595966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1562_n 0.00636858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1563_n 0.00803143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1564_n 0.0122991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1565_n 0.0350016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1566_n 0.0213734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1567_n 0.0211536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1568_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1569_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1570_n 0.0346609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1571_n 0.00180198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1572_n 0.036062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1573_n 0.0034365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1574_n 0.0182335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1575_n 0.0214173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1576_n 0.0487365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1577_n 0.0536763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1578_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1579_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1580_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1581_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1582_n 0.00628274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1583_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1584_n 0.00223746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1585_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1586_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1587_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1588_n 0.00535984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1589_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1558_n 0.123252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_Q_c_1745_n 0.00205506f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_268 VPB N_Q_c_1746_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_269 VPB N_Q_c_1747_n 0.00233077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB Q 0.00844788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB Q 0.0182893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_Q_c_1750_n 0.00267489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 N_D_c_274_n N_CLK_M1024_g 0.00441433f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_274 N_D_c_274_n N_CLK_c_310_n 0.00572583f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_275 N_D_c_276_n N_CLK_c_311_n 0.00232413f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_276 N_D_c_274_n N_A_225_74#_c_964_n 0.0035771f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_277 N_D_M1032_g N_A_225_74#_c_966_n 0.00621603f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_278 N_D_c_276_n N_A_225_74#_c_966_n 0.0035771f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_279 N_D_c_277_n N_A_225_74#_c_966_n 0.0557245f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_280 N_D_c_274_n N_A_225_74#_c_983_n 0.00296994f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_281 N_D_M1031_g N_A_225_74#_c_983_n 0.00249516f $X=0.505 $Y=2.73 $X2=0 $Y2=0
cc_282 N_D_c_277_n N_A_225_74#_c_983_n 0.02241f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_283 N_D_M1032_g N_A_27_74#_c_1489_n 0.00146243f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_284 N_D_M1032_g N_A_27_74#_c_1490_n 0.00600966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_285 N_D_c_276_n N_A_27_74#_c_1490_n 0.0338681f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_286 N_D_c_277_n N_A_27_74#_c_1490_n 0.0697394f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_287 N_D_M1031_g N_A_27_74#_c_1495_n 0.00561317f $X=0.505 $Y=2.73 $X2=0 $Y2=0
cc_288 N_D_M1031_g N_A_27_74#_c_1496_n 0.0218542f $X=0.505 $Y=2.73 $X2=0 $Y2=0
cc_289 N_D_c_277_n N_A_27_74#_c_1496_n 0.019138f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_290 N_D_c_281_n N_A_27_74#_c_1496_n 0.00134301f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_291 N_D_M1031_g N_VPWR_c_1559_n 0.0135514f $X=0.505 $Y=2.73 $X2=0 $Y2=0
cc_292 N_D_M1031_g N_VPWR_c_1574_n 0.00562069f $X=0.505 $Y=2.73 $X2=0 $Y2=0
cc_293 N_D_M1031_g N_VPWR_c_1558_n 0.0054305f $X=0.505 $Y=2.73 $X2=0 $Y2=0
cc_294 N_D_M1032_g N_VGND_c_1810_n 0.0137856f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_295 N_D_c_276_n N_VGND_c_1810_n 0.00175174f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_296 N_D_c_277_n N_VGND_c_1810_n 0.0220022f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_297 N_D_M1032_g N_VGND_c_1821_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_298 N_D_M1032_g N_VGND_c_1833_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_299 CLK N_A_225_74#_M1018_g 0.00400177f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_300 N_CLK_c_310_n N_A_225_74#_M1018_g 0.0206752f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_301 N_CLK_c_311_n N_A_225_74#_M1018_g 0.0131399f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_302 N_CLK_M1024_g N_A_225_74#_M1027_g 0.0472331f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_303 N_CLK_M1024_g N_A_225_74#_c_961_n 0.00781426f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_304 N_CLK_M1024_g N_A_225_74#_c_964_n 0.00356278f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_305 CLK N_A_225_74#_c_964_n 0.0286813f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_306 N_CLK_c_310_n N_A_225_74#_c_964_n 0.00297156f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_307 N_CLK_c_311_n N_A_225_74#_c_964_n 0.00330079f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_308 N_CLK_M1024_g N_A_225_74#_c_981_n 0.00932745f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_309 N_CLK_c_310_n N_A_225_74#_c_981_n 5.60514e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_310 N_CLK_M1024_g N_A_225_74#_c_965_n 8.97049e-19 $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_311 CLK N_A_225_74#_c_965_n 0.0162505f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_312 CLK N_A_225_74#_c_966_n 0.00763035f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_313 N_CLK_c_310_n N_A_225_74#_c_966_n 0.00114664f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_314 N_CLK_c_311_n N_A_225_74#_c_966_n 0.00811931f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_315 N_CLK_M1024_g N_A_225_74#_c_983_n 0.00699187f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_316 CLK N_A_225_74#_c_983_n 0.0353752f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_317 N_CLK_c_310_n N_A_225_74#_c_983_n 0.00317947f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_318 N_CLK_M1024_g N_A_27_74#_c_1496_n 0.018001f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_319 CLK N_A_27_74#_c_1491_n 0.00460396f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_320 N_CLK_M1024_g N_VPWR_c_1559_n 0.0131823f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_321 N_CLK_M1024_g N_VPWR_c_1560_n 0.0251708f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_322 N_CLK_M1024_g N_VPWR_c_1575_n 0.00460063f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_323 N_CLK_M1024_g N_VPWR_c_1558_n 0.00913687f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_324 N_CLK_c_311_n N_VGND_c_1810_n 0.00280144f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_325 N_CLK_c_311_n N_VGND_c_1811_n 0.00434054f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_326 CLK N_VGND_c_1812_n 0.013855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_327 N_CLK_c_311_n N_VGND_c_1812_n 0.0027655f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_328 N_CLK_c_311_n N_VGND_c_1833_n 0.0082522f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_329 N_A_398_74#_c_373_n N_A_767_402#_M1010_g 0.0025182f $X=3.71 $Y=2.905
+ $X2=0 $Y2=0
cc_330 N_A_398_74#_c_374_n N_A_767_402#_M1010_g 0.0200606f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_331 N_A_398_74#_c_375_n N_A_767_402#_M1010_g 0.00368728f $X=4.6 $Y=2.905
+ $X2=0 $Y2=0
cc_332 N_A_398_74#_M1013_g N_A_767_402#_c_607_n 0.0422629f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_333 N_A_398_74#_c_353_n N_A_767_402#_c_610_n 6.69553e-19 $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_354_n N_A_767_402#_c_610_n 0.00851627f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_335 N_A_398_74#_c_353_n N_A_767_402#_c_615_n 0.0123371f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_c_354_n N_A_767_402#_c_615_n 2.62742e-19 $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_337 N_A_398_74#_c_374_n N_A_767_402#_c_615_n 0.0444853f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_338 N_A_398_74#_c_352_n N_A_767_402#_c_616_n 0.00106832f $X=2.95 $Y=1.62
+ $X2=0 $Y2=0
cc_339 N_A_398_74#_c_353_n N_A_767_402#_c_616_n 0.00758688f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_340 N_A_398_74#_c_354_n N_A_767_402#_c_616_n 0.00891788f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_341 N_A_398_74#_c_374_n N_A_767_402#_c_616_n 0.0129825f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_342 N_A_398_74#_c_374_n N_A_767_402#_c_617_n 0.0104876f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_c_378_n N_A_767_402#_c_617_n 0.00133539f $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_344 N_A_398_74#_c_380_n N_A_767_402#_c_617_n 0.00853861f $X=5.51 $Y=2.18
+ $X2=0 $Y2=0
cc_345 N_A_398_74#_M1013_g N_A_767_402#_c_611_n 8.22539e-19 $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_346 N_A_398_74#_c_374_n N_A_767_402#_c_618_n 0.0032594f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_c_375_n N_A_767_402#_c_618_n 0.0294669f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_348 N_A_398_74#_c_376_n N_A_767_402#_c_618_n 0.020903f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_349 N_A_398_74#_c_378_n N_A_767_402#_c_618_n 0.0156619f $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_350 N_A_398_74#_M1013_g N_A_767_402#_c_612_n 0.00603499f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_351 N_A_398_74#_c_374_n N_A_612_74#_M1038_g 0.00391134f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_352 N_A_398_74#_c_375_n N_A_612_74#_M1038_g 0.0123464f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_353 N_A_398_74#_c_376_n N_A_612_74#_M1038_g 0.00283539f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_354 N_A_398_74#_c_378_n N_A_612_74#_M1038_g 6.03531e-19 $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_355 N_A_398_74#_c_378_n N_A_612_74#_M1033_g 0.00346038f $X=5.425 $Y=2.905
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_c_379_n N_A_612_74#_M1033_g 0.02026f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_357 N_A_398_74#_c_355_n N_A_612_74#_M1033_g 0.00914775f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_358 N_A_398_74#_c_357_n N_A_612_74#_M1028_g 0.00161751f $X=6.475 $Y=0.34
+ $X2=0 $Y2=0
cc_359 N_A_398_74#_c_360_n N_A_612_74#_M1028_g 0.00397266f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_360 N_A_398_74#_c_361_n N_A_612_74#_M1028_g 0.00869284f $X=6.5 $Y=1.12 $X2=0
+ $Y2=0
cc_361 N_A_398_74#_c_363_n N_A_612_74#_M1028_g 0.0195997f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_M1013_g N_A_612_74#_c_696_n 0.0187196f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_363 N_A_398_74#_c_349_n N_A_612_74#_c_696_n 0.00381334f $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_364 N_A_398_74#_c_358_n N_A_612_74#_c_696_n 0.0403355f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_M1013_g N_A_612_74#_c_697_n 0.0142826f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_366 N_A_398_74#_c_353_n N_A_612_74#_c_697_n 0.0132987f $X=3.71 $Y=1.635 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_c_354_n N_A_612_74#_c_697_n 0.0039875f $X=3.71 $Y=1.635 $X2=0
+ $Y2=0
cc_368 N_A_398_74#_M1001_g N_A_612_74#_c_709_n 3.31415e-19 $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_369 N_A_398_74#_c_346_n N_A_612_74#_c_709_n 0.00503148f $X=3.51 $Y=1.635
+ $X2=0 $Y2=0
cc_370 N_A_398_74#_c_367_n N_A_612_74#_c_709_n 0.0219188f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_M1001_g N_A_612_74#_c_700_n 0.00259065f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_372 N_A_398_74#_c_346_n N_A_612_74#_c_700_n 0.0221174f $X=3.51 $Y=1.635 $X2=0
+ $Y2=0
cc_373 N_A_398_74#_M1013_g N_A_612_74#_c_700_n 0.00425975f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_374 N_A_398_74#_c_352_n N_A_612_74#_c_700_n 0.00608023f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_375 N_A_398_74#_c_353_n N_A_612_74#_c_700_n 0.0498141f $X=3.71 $Y=1.635 $X2=0
+ $Y2=0
cc_376 N_A_398_74#_c_358_n N_A_612_74#_c_700_n 0.0606779f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_377 N_A_398_74#_c_382_n N_A_612_74#_c_700_n 0.0129295f $X=3.71 $Y=2.25 $X2=0
+ $Y2=0
cc_378 N_A_398_74#_c_346_n N_A_612_74#_c_701_n 0.00242402f $X=3.51 $Y=1.635
+ $X2=0 $Y2=0
cc_379 N_A_398_74#_M1013_g N_A_612_74#_c_701_n 0.00427915f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_380 N_A_398_74#_c_358_n N_A_612_74#_c_701_n 0.0143568f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_381 N_A_398_74#_M1013_g N_A_612_74#_c_702_n 0.00178188f $X=3.585 $Y=0.58
+ $X2=0 $Y2=0
cc_382 N_A_398_74#_c_353_n N_A_612_74#_c_702_n 0.00715168f $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_383 N_A_398_74#_c_354_n N_A_612_74#_c_702_n 9.47085e-19 $X=3.71 $Y=1.635
+ $X2=0 $Y2=0
cc_384 N_A_398_74#_c_374_n N_A_612_74#_c_702_n 0.00485285f $X=4.515 $Y=2.25
+ $X2=0 $Y2=0
cc_385 N_A_398_74#_c_379_n N_A_612_74#_c_704_n 0.00295832f $X=6.305 $Y=2.18
+ $X2=0 $Y2=0
cc_386 N_A_398_74#_c_359_n N_A_612_74#_c_704_n 0.0230196f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_387 N_A_398_74#_c_360_n N_A_612_74#_c_704_n 2.80493e-19 $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_388 N_A_398_74#_c_379_n N_A_612_74#_c_705_n 0.00199466f $X=6.305 $Y=2.18
+ $X2=0 $Y2=0
cc_389 N_A_398_74#_c_359_n N_A_612_74#_c_705_n 0.00389788f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_390 N_A_398_74#_c_360_n N_A_612_74#_c_705_n 0.0139138f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_391 N_A_398_74#_c_376_n N_SET_B_M1011_g 0.00295426f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_392 N_A_398_74#_c_378_n N_SET_B_M1011_g 0.0164116f $X=5.425 $Y=2.905 $X2=0
+ $Y2=0
cc_393 N_A_398_74#_c_380_n N_SET_B_M1011_g 0.00680112f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_394 N_A_398_74#_c_379_n N_SET_B_c_833_n 0.0190347f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_395 N_A_398_74#_c_355_n N_SET_B_c_833_n 0.0222258f $X=6.39 $Y=2.095 $X2=0
+ $Y2=0
cc_396 N_A_398_74#_c_359_n N_SET_B_c_833_n 0.00959624f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_c_383_n N_SET_B_c_833_n 0.00572674f $X=7.21 $Y=2.185 $X2=0
+ $Y2=0
cc_398 N_A_398_74#_c_362_n N_SET_B_c_833_n 0.0208316f $X=7.21 $Y=2.02 $X2=0
+ $Y2=0
cc_399 N_A_398_74#_c_385_n N_SET_B_c_833_n 0.00108214f $X=7.325 $Y=2.185 $X2=0
+ $Y2=0
cc_400 N_A_398_74#_c_379_n N_SET_B_c_834_n 0.00190675f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_401 N_A_398_74#_c_380_n N_SET_B_c_834_n 8.05363e-19 $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_402 N_A_398_74#_c_379_n N_SET_B_c_836_n 0.00913037f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_403 N_A_398_74#_c_380_n N_SET_B_c_836_n 0.0133873f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_355_n N_SET_B_c_836_n 0.00814397f $X=6.39 $Y=2.095 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_379_n N_SET_B_c_837_n 0.00156156f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_380_n N_SET_B_c_837_n 0.00317486f $X=5.51 $Y=2.18 $X2=0
+ $Y2=0
cc_407 N_A_398_74#_c_348_n N_A_225_74#_M1018_g 0.00164183f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_408 N_A_398_74#_c_350_n N_A_225_74#_M1018_g 0.00266901f $X=2.215 $Y=0.34
+ $X2=0 $Y2=0
cc_409 N_A_398_74#_c_368_n N_A_225_74#_M1027_g 0.00144344f $X=2.275 $Y=2.99
+ $X2=0 $Y2=0
cc_410 N_A_398_74#_M1001_g N_A_225_74#_c_968_n 0.0181106f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_411 N_A_398_74#_c_468_p N_A_225_74#_c_968_n 0.00598552f $X=2.19 $Y=2.575
+ $X2=0 $Y2=0
cc_412 N_A_398_74#_c_367_n N_A_225_74#_c_968_n 0.0101668f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_413 N_A_398_74#_c_351_n N_A_225_74#_c_968_n 3.80136e-19 $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_414 N_A_398_74#_c_349_n N_A_225_74#_c_956_n 0.00237694f $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_415 N_A_398_74#_c_351_n N_A_225_74#_c_956_n 0.00105733f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_416 N_A_398_74#_c_352_n N_A_225_74#_c_956_n 0.0147005f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_417 N_A_398_74#_c_358_n N_A_225_74#_c_956_n 0.00695648f $X=2.95 $Y=1.455
+ $X2=0 $Y2=0
cc_418 N_A_398_74#_M1001_g N_A_225_74#_c_969_n 0.0105864f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_419 N_A_398_74#_c_367_n N_A_225_74#_c_969_n 0.0128457f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_420 N_A_398_74#_M1013_g N_A_225_74#_M1023_g 0.0179618f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_421 N_A_398_74#_c_348_n N_A_225_74#_M1023_g 0.00395905f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_349_n N_A_225_74#_M1023_g 0.010044f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_423 N_A_398_74#_c_358_n N_A_225_74#_M1023_g 0.0216123f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_424 N_A_398_74#_M1001_g N_A_225_74#_M1002_g 0.0108932f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_346_n N_A_225_74#_M1002_g 0.00779081f $X=3.51 $Y=1.635
+ $X2=0 $Y2=0
cc_426 N_A_398_74#_c_367_n N_A_225_74#_M1002_g 0.0183218f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_427 N_A_398_74#_c_373_n N_A_225_74#_M1002_g 0.0063525f $X=3.71 $Y=2.905 $X2=0
+ $Y2=0
cc_428 N_A_398_74#_c_382_n N_A_225_74#_M1002_g 0.00113129f $X=3.71 $Y=2.25 $X2=0
+ $Y2=0
cc_429 N_A_398_74#_c_367_n N_A_225_74#_c_972_n 0.00410612f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_430 N_A_398_74#_c_376_n N_A_225_74#_c_972_n 0.0135663f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_431 N_A_398_74#_c_377_n N_A_225_74#_c_972_n 0.00420304f $X=4.685 $Y=2.99
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_M1036_g N_A_225_74#_M1025_g 0.00476377f $X=7.325 $Y=2.75
+ $X2=0 $Y2=0
cc_433 N_A_398_74#_c_379_n N_A_225_74#_M1025_g 0.00613584f $X=6.305 $Y=2.18
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_c_355_n N_A_225_74#_M1025_g 0.00587557f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_383_n N_A_225_74#_c_958_n 0.00103484f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_436 N_A_398_74#_c_385_n N_A_225_74#_c_958_n 0.00901519f $X=7.325 $Y=2.185
+ $X2=0 $Y2=0
cc_437 N_A_398_74#_c_355_n N_A_225_74#_c_959_n 0.00373037f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_438 N_A_398_74#_c_359_n N_A_225_74#_c_959_n 0.001254f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_439 N_A_398_74#_c_360_n N_A_225_74#_c_959_n 0.0172301f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_440 N_A_398_74#_c_355_n N_A_225_74#_M1015_g 8.38958e-19 $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_441 N_A_398_74#_c_356_n N_A_225_74#_M1015_g 0.0127652f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_442 N_A_398_74#_c_359_n N_A_225_74#_M1015_g 3.27596e-19 $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_360_n N_A_225_74#_M1015_g 0.0110658f $X=6.53 $Y=1.285 $X2=0
+ $Y2=0
cc_444 N_A_398_74#_c_362_n N_A_225_74#_M1015_g 0.00923424f $X=7.21 $Y=2.02 $X2=0
+ $Y2=0
cc_445 N_A_398_74#_c_363_n N_A_225_74#_M1015_g 0.0190732f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_446 N_A_398_74#_c_348_n N_A_225_74#_c_962_n 5.90715e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_c_349_n N_A_225_74#_c_962_n 9.09485e-19 $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_448 N_A_398_74#_c_351_n N_A_225_74#_c_962_n 3.80136e-19 $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_449 N_A_398_74#_c_352_n N_A_225_74#_c_962_n 0.0394012f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_450 N_A_398_74#_c_358_n N_A_225_74#_c_962_n 8.19775e-19 $X=2.95 $Y=1.455
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_348_n N_A_225_74#_c_963_n 0.00102206f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_M1027_d N_A_225_74#_c_981_n 0.00231044f $X=2.055 $Y=1.84
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_348_n N_A_225_74#_c_965_n 0.0120964f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_454 N_A_398_74#_c_356_n N_A_1484_62#_M1007_g 0.00169096f $X=7.205 $Y=0.34
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_362_n N_A_1484_62#_M1007_g 0.00722371f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_456 N_A_398_74#_c_383_n N_A_1484_62#_M1014_g 0.00174361f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_457 N_A_398_74#_c_362_n N_A_1484_62#_M1014_g 0.00915762f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_458 N_A_398_74#_c_385_n N_A_1484_62#_M1014_g 0.0575918f $X=7.325 $Y=2.185
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_362_n N_A_1484_62#_c_1129_n 0.0479592f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_362_n N_A_1484_62#_c_1144_n 0.0127905f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_461 N_A_398_74#_c_356_n N_A_1324_392#_M1006_d 0.00205663f $X=7.205 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_462 N_A_398_74#_M1036_g N_A_1324_392#_c_1227_n 0.00234858f $X=7.325 $Y=2.75
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_355_n N_A_1324_392#_c_1227_n 0.0148971f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_383_n N_A_1324_392#_c_1227_n 0.0185355f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_362_n N_A_1324_392#_c_1227_n 0.0100217f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_466 N_A_398_74#_c_385_n N_A_1324_392#_c_1227_n 0.00319533f $X=7.325 $Y=2.185
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_c_355_n N_A_1324_392#_c_1216_n 0.00689075f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_359_n N_A_1324_392#_c_1216_n 0.0251223f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_c_360_n N_A_1324_392#_c_1216_n 0.00226999f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_361_n N_A_1324_392#_c_1216_n 0.00627822f $X=6.5 $Y=1.12
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_362_n N_A_1324_392#_c_1216_n 0.0496067f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_472 N_A_398_74#_c_363_n N_A_1324_392#_c_1216_n 0.00150671f $X=6.53 $Y=1.12
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_M1036_g N_A_1324_392#_c_1228_n 0.00995194f $X=7.325 $Y=2.75
+ $X2=0 $Y2=0
cc_474 N_A_398_74#_c_383_n N_A_1324_392#_c_1228_n 0.00826905f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_M1036_g N_A_1324_392#_c_1229_n 0.0107571f $X=7.325 $Y=2.75
+ $X2=0 $Y2=0
cc_476 N_A_398_74#_c_383_n N_A_1324_392#_c_1229_n 0.0181124f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_477 N_A_398_74#_c_385_n N_A_1324_392#_c_1229_n 0.00461229f $X=7.325 $Y=2.185
+ $X2=0 $Y2=0
cc_478 N_A_398_74#_c_356_n N_A_1324_392#_c_1219_n 0.0218291f $X=7.205 $Y=0.34
+ $X2=0 $Y2=0
cc_479 N_A_398_74#_c_359_n N_A_1324_392#_c_1219_n 0.00246577f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_362_n N_A_1324_392#_c_1219_n 0.0150761f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_481 N_A_398_74#_c_363_n N_A_1324_392#_c_1219_n 0.00408225f $X=6.53 $Y=1.12
+ $X2=0 $Y2=0
cc_482 N_A_398_74#_c_355_n N_A_1324_392#_c_1220_n 0.0101597f $X=6.39 $Y=2.095
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_359_n N_A_1324_392#_c_1220_n 0.00157906f $X=6.53 $Y=1.285
+ $X2=0 $Y2=0
cc_484 N_A_398_74#_c_362_n N_A_1324_392#_c_1220_n 0.0119049f $X=7.21 $Y=2.02
+ $X2=0 $Y2=0
cc_485 N_A_398_74#_c_385_n N_A_1324_392#_c_1234_n 0.00367764f $X=7.325 $Y=2.185
+ $X2=0 $Y2=0
cc_486 N_A_398_74#_c_349_n N_A_27_74#_M1023_s 0.00416589f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_487 N_A_398_74#_M1027_d N_A_27_74#_c_1497_n 0.00574218f $X=2.055 $Y=1.84
+ $X2=0 $Y2=0
cc_488 N_A_398_74#_M1001_g N_A_27_74#_c_1497_n 0.00813468f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_489 N_A_398_74#_c_468_p N_A_27_74#_c_1497_n 0.0380749f $X=2.19 $Y=2.575 $X2=0
+ $Y2=0
cc_490 N_A_398_74#_c_367_n N_A_27_74#_c_1497_n 0.0395555f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_491 N_A_398_74#_c_351_n N_A_27_74#_c_1497_n 0.0181995f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_492 N_A_398_74#_c_352_n N_A_27_74#_c_1497_n 0.00131676f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_493 N_A_398_74#_c_348_n N_A_27_74#_c_1491_n 0.0119813f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_494 N_A_398_74#_c_351_n N_A_27_74#_c_1491_n 0.0461461f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_495 N_A_398_74#_c_352_n N_A_27_74#_c_1491_n 0.00357538f $X=2.95 $Y=1.62 $X2=0
+ $Y2=0
cc_496 N_A_398_74#_c_358_n N_A_27_74#_c_1491_n 0.023467f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_497 N_A_398_74#_c_348_n N_A_27_74#_c_1493_n 0.0206593f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_498 N_A_398_74#_c_349_n N_A_27_74#_c_1493_n 0.0239262f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_499 N_A_398_74#_c_358_n N_A_27_74#_c_1493_n 0.0244211f $X=2.95 $Y=1.455 $X2=0
+ $Y2=0
cc_500 N_A_398_74#_c_374_n N_VPWR_M1010_d 0.0100399f $X=4.515 $Y=2.25 $X2=0
+ $Y2=0
cc_501 N_A_398_74#_c_375_n N_VPWR_M1010_d 0.0115414f $X=4.6 $Y=2.905 $X2=0 $Y2=0
cc_502 N_A_398_74#_c_378_n N_VPWR_M1011_d 0.0044983f $X=5.425 $Y=2.905 $X2=0
+ $Y2=0
cc_503 N_A_398_74#_c_379_n N_VPWR_M1011_d 0.00568979f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_504 N_A_398_74#_c_368_n N_VPWR_c_1560_n 0.0103602f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_367_n N_VPWR_c_1561_n 0.0132711f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_373_n N_VPWR_c_1561_n 0.00998696f $X=3.71 $Y=2.905 $X2=0
+ $Y2=0
cc_507 N_A_398_74#_c_375_n N_VPWR_c_1561_n 0.00670097f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_508 N_A_398_74#_c_377_n N_VPWR_c_1561_n 0.00852847f $X=4.685 $Y=2.99 $X2=0
+ $Y2=0
cc_509 N_A_398_74#_c_376_n N_VPWR_c_1562_n 0.0147865f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_c_378_n N_VPWR_c_1562_n 0.0356944f $X=5.425 $Y=2.905 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_379_n N_VPWR_c_1562_n 0.0162955f $X=6.305 $Y=2.18 $X2=0
+ $Y2=0
cc_512 N_A_398_74#_c_373_n N_VPWR_c_1571_n 0.00929866f $X=3.71 $Y=2.905 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_374_n N_VPWR_c_1571_n 0.0224779f $X=4.515 $Y=2.25 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_375_n N_VPWR_c_1571_n 0.0192298f $X=4.6 $Y=2.905 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_376_n N_VPWR_c_1572_n 0.0537108f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_377_n N_VPWR_c_1572_n 0.0115893f $X=4.685 $Y=2.99 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_367_n N_VPWR_c_1576_n 0.0975205f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_368_n N_VPWR_c_1576_n 0.0121664f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_M1036_g N_VPWR_c_1577_n 0.00389275f $X=7.325 $Y=2.75 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_M1036_g N_VPWR_c_1558_n 0.0049743f $X=7.325 $Y=2.75 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_367_n N_VPWR_c_1558_n 0.0514634f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_368_n N_VPWR_c_1558_n 0.00660537f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_376_n N_VPWR_c_1558_n 0.0278398f $X=5.34 $Y=2.99 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_377_n N_VPWR_c_1558_n 0.00583135f $X=4.685 $Y=2.99 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_373_n A_719_463# 0.00150957f $X=3.71 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_526 N_A_398_74#_c_379_n A_1223_347# 0.0106143f $X=6.305 $Y=2.18 $X2=-0.19
+ $Y2=-0.245
cc_527 N_A_398_74#_c_355_n A_1223_347# 0.00481312f $X=6.39 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_528 N_A_398_74#_c_350_n N_VGND_c_1812_n 0.0109685f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_529 N_A_398_74#_M1013_g N_VGND_c_1813_n 0.00126697f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_530 N_A_398_74#_c_357_n N_VGND_c_1814_n 0.00917417f $X=6.475 $Y=0.34 $X2=0
+ $Y2=0
cc_531 N_A_398_74#_c_361_n N_VGND_c_1814_n 0.0285193f $X=6.5 $Y=1.12 $X2=0 $Y2=0
cc_532 N_A_398_74#_c_363_n N_VGND_c_1814_n 4.42772e-19 $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_533 N_A_398_74#_M1013_g N_VGND_c_1822_n 0.00434272f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_534 N_A_398_74#_c_349_n N_VGND_c_1822_n 0.0586507f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_535 N_A_398_74#_c_350_n N_VGND_c_1822_n 0.0121867f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_536 N_A_398_74#_c_356_n N_VGND_c_1829_n 0.0587172f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_537 N_A_398_74#_c_357_n N_VGND_c_1829_n 0.0121867f $X=6.475 $Y=0.34 $X2=0
+ $Y2=0
cc_538 N_A_398_74#_c_363_n N_VGND_c_1829_n 0.00278271f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_539 N_A_398_74#_c_356_n N_VGND_c_1830_n 0.00636506f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_540 N_A_398_74#_c_362_n N_VGND_c_1830_n 0.00405322f $X=7.21 $Y=2.02 $X2=0
+ $Y2=0
cc_541 N_A_398_74#_M1013_g N_VGND_c_1833_n 0.00822443f $X=3.585 $Y=0.58 $X2=0
+ $Y2=0
cc_542 N_A_398_74#_c_349_n N_VGND_c_1833_n 0.0333627f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_543 N_A_398_74#_c_350_n N_VGND_c_1833_n 0.00660921f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_544 N_A_398_74#_c_356_n N_VGND_c_1833_n 0.033365f $X=7.205 $Y=0.34 $X2=0
+ $Y2=0
cc_545 N_A_398_74#_c_357_n N_VGND_c_1833_n 0.00660921f $X=6.475 $Y=0.34 $X2=0
+ $Y2=0
cc_546 N_A_398_74#_c_363_n N_VGND_c_1833_n 0.00359494f $X=6.53 $Y=1.12 $X2=0
+ $Y2=0
cc_547 N_A_398_74#_c_357_n A_1225_74# 7.18263e-19 $X=6.475 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_548 N_A_398_74#_c_361_n A_1225_74# 0.00947773f $X=6.5 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_549 N_A_398_74#_c_362_n A_1436_88# 0.00181261f $X=7.21 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_550 N_A_767_402#_c_615_n N_A_612_74#_M1038_g 0.0151251f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_551 N_A_767_402#_c_616_n N_A_612_74#_M1038_g 0.0185659f $X=4.28 $Y=1.865
+ $X2=0 $Y2=0
cc_552 N_A_767_402#_c_617_n N_A_612_74#_M1038_g 0.00831739f $X=4.94 $Y=2.295
+ $X2=0 $Y2=0
cc_553 N_A_767_402#_c_618_n N_A_612_74#_M1038_g 0.00856245f $X=5.085 $Y=2.515
+ $X2=0 $Y2=0
cc_554 N_A_767_402#_c_611_n N_A_612_74#_c_693_n 0.00995281f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_555 N_A_767_402#_c_612_n N_A_612_74#_c_693_n 0.00382576f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_556 N_A_767_402#_c_607_n N_A_612_74#_c_696_n 0.00306844f $X=3.975 $Y=0.9
+ $X2=0 $Y2=0
cc_557 N_A_767_402#_c_612_n N_A_612_74#_c_696_n 3.7427e-19 $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_558 N_A_767_402#_c_609_n N_A_612_74#_c_697_n 0.00297558f $X=4.05 $Y=0.975
+ $X2=0 $Y2=0
cc_559 N_A_767_402#_c_608_n N_A_612_74#_c_698_n 0.00182267f $X=4.23 $Y=0.975
+ $X2=0 $Y2=0
cc_560 N_A_767_402#_c_610_n N_A_612_74#_c_698_n 0.0126255f $X=4.305 $Y=1.7 $X2=0
+ $Y2=0
cc_561 N_A_767_402#_c_615_n N_A_612_74#_c_698_n 0.0475354f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_562 N_A_767_402#_c_616_n N_A_612_74#_c_698_n 0.00174649f $X=4.28 $Y=1.865
+ $X2=0 $Y2=0
cc_563 N_A_767_402#_c_611_n N_A_612_74#_c_698_n 0.0290223f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_564 N_A_767_402#_c_612_n N_A_612_74#_c_698_n 0.00105029f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_565 N_A_767_402#_c_611_n N_A_612_74#_c_699_n 0.00128907f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_566 N_A_767_402#_M1010_g N_A_612_74#_c_700_n 4.34548e-19 $X=3.925 $Y=2.525
+ $X2=0 $Y2=0
cc_567 N_A_767_402#_c_609_n N_A_612_74#_c_702_n 0.0059641f $X=4.05 $Y=0.975
+ $X2=0 $Y2=0
cc_568 N_A_767_402#_c_610_n N_A_612_74#_c_702_n 3.58867e-19 $X=4.305 $Y=1.7
+ $X2=0 $Y2=0
cc_569 N_A_767_402#_c_615_n N_A_612_74#_c_702_n 0.00151836f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_570 N_A_767_402#_c_616_n N_A_612_74#_c_702_n 0.00315033f $X=4.28 $Y=1.865
+ $X2=0 $Y2=0
cc_571 N_A_767_402#_c_611_n N_A_612_74#_c_702_n 0.00746874f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_572 N_A_767_402#_c_612_n N_A_612_74#_c_702_n 0.00363451f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_573 N_A_767_402#_c_610_n N_A_612_74#_c_703_n 7.77514e-19 $X=4.305 $Y=1.7
+ $X2=0 $Y2=0
cc_574 N_A_767_402#_c_615_n N_A_612_74#_c_703_n 0.0206269f $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_575 N_A_767_402#_c_611_n N_A_612_74#_c_703_n 0.0261626f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_576 N_A_767_402#_c_610_n N_A_612_74#_c_706_n 0.0148476f $X=4.305 $Y=1.7 $X2=0
+ $Y2=0
cc_577 N_A_767_402#_c_615_n N_A_612_74#_c_706_n 4.25161e-19 $X=4.855 $Y=1.867
+ $X2=0 $Y2=0
cc_578 N_A_767_402#_c_611_n N_A_612_74#_c_706_n 0.00234761f $X=4.395 $Y=1.065
+ $X2=0 $Y2=0
cc_579 N_A_767_402#_c_612_n N_A_612_74#_c_706_n 0.00699025f $X=4.395 $Y=0.975
+ $X2=0 $Y2=0
cc_580 N_A_767_402#_c_617_n N_SET_B_M1011_g 0.00336143f $X=4.94 $Y=2.295 $X2=0
+ $Y2=0
cc_581 N_A_767_402#_c_618_n N_SET_B_M1011_g 2.64649e-19 $X=5.085 $Y=2.515 $X2=0
+ $Y2=0
cc_582 N_A_767_402#_c_611_n N_SET_B_M1016_g 9.88858e-19 $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_583 N_A_767_402#_c_615_n N_SET_B_c_834_n 2.23271e-19 $X=4.855 $Y=1.867 $X2=0
+ $Y2=0
cc_584 N_A_767_402#_c_615_n N_SET_B_c_836_n 0.0156891f $X=4.855 $Y=1.867 $X2=0
+ $Y2=0
cc_585 N_A_767_402#_c_615_n N_SET_B_c_837_n 0.00255214f $X=4.855 $Y=1.867 $X2=0
+ $Y2=0
cc_586 N_A_767_402#_M1010_g N_A_225_74#_M1002_g 0.0310264f $X=3.925 $Y=2.525
+ $X2=0 $Y2=0
cc_587 N_A_767_402#_M1010_g N_A_225_74#_c_972_n 0.0123711f $X=3.925 $Y=2.525
+ $X2=0 $Y2=0
cc_588 N_A_767_402#_M1010_g N_VPWR_c_1561_n 0.00352584f $X=3.925 $Y=2.525 $X2=0
+ $Y2=0
cc_589 N_A_767_402#_M1010_g N_VPWR_c_1571_n 0.00374568f $X=3.925 $Y=2.525 $X2=0
+ $Y2=0
cc_590 N_A_767_402#_M1010_g N_VPWR_c_1558_n 9.455e-19 $X=3.925 $Y=2.525 $X2=0
+ $Y2=0
cc_591 N_A_767_402#_c_611_n N_VGND_M1003_d 0.00118908f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_592 N_A_767_402#_c_607_n N_VGND_c_1813_n 0.0098944f $X=3.975 $Y=0.9 $X2=0
+ $Y2=0
cc_593 N_A_767_402#_c_608_n N_VGND_c_1813_n 0.0079331f $X=4.23 $Y=0.975 $X2=0
+ $Y2=0
cc_594 N_A_767_402#_c_611_n N_VGND_c_1813_n 0.00929432f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_595 N_A_767_402#_c_612_n N_VGND_c_1813_n 6.63116e-19 $X=4.395 $Y=0.975 $X2=0
+ $Y2=0
cc_596 N_A_767_402#_c_611_n N_VGND_c_1814_n 0.00958081f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_597 N_A_767_402#_c_611_n N_VGND_c_1819_n 0.00824154f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_598 N_A_767_402#_c_607_n N_VGND_c_1822_n 0.00383152f $X=3.975 $Y=0.9 $X2=0
+ $Y2=0
cc_599 N_A_767_402#_c_607_n N_VGND_c_1833_n 0.0075725f $X=3.975 $Y=0.9 $X2=0
+ $Y2=0
cc_600 N_A_767_402#_c_611_n N_VGND_c_1833_n 0.0209055f $X=4.395 $Y=1.065 $X2=0
+ $Y2=0
cc_601 N_A_612_74#_M1038_g N_SET_B_M1011_g 0.021147f $X=4.86 $Y=2.525 $X2=0
+ $Y2=0
cc_602 N_A_612_74#_M1033_g N_SET_B_M1011_g 0.0133015f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_603 N_A_612_74#_M1038_g N_SET_B_M1016_g 0.00427675f $X=4.86 $Y=2.525 $X2=0
+ $Y2=0
cc_604 N_A_612_74#_c_693_n N_SET_B_M1016_g 0.0531748f $X=5.1 $Y=1.12 $X2=0 $Y2=0
cc_605 N_A_612_74#_M1033_g N_SET_B_M1016_g 0.0151427f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_606 N_A_612_74#_M1028_g N_SET_B_M1016_g 0.0120624f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_607 N_A_612_74#_c_699_n N_SET_B_M1016_g 0.0144612f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_608 N_A_612_74#_c_703_n N_SET_B_M1016_g 0.00275571f $X=4.935 $Y=1.285 $X2=0
+ $Y2=0
cc_609 N_A_612_74#_c_704_n N_SET_B_M1016_g 8.93876e-19 $X=5.97 $Y=1.285 $X2=0
+ $Y2=0
cc_610 N_A_612_74#_c_705_n N_SET_B_M1016_g 0.0185109f $X=5.97 $Y=1.365 $X2=0
+ $Y2=0
cc_611 N_A_612_74#_M1033_g N_SET_B_c_833_n 0.00732598f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_612 N_A_612_74#_c_699_n N_SET_B_c_833_n 0.00599672f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_613 N_A_612_74#_c_704_n N_SET_B_c_833_n 0.010239f $X=5.97 $Y=1.285 $X2=0
+ $Y2=0
cc_614 N_A_612_74#_c_705_n N_SET_B_c_833_n 0.00389225f $X=5.97 $Y=1.365 $X2=0
+ $Y2=0
cc_615 N_A_612_74#_M1033_g N_SET_B_c_834_n 0.00133736f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_616 N_A_612_74#_c_699_n N_SET_B_c_834_n 0.00787805f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_617 N_A_612_74#_M1038_g N_SET_B_c_836_n 0.00301198f $X=4.86 $Y=2.525 $X2=0
+ $Y2=0
cc_618 N_A_612_74#_M1033_g N_SET_B_c_836_n 0.00322608f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_619 N_A_612_74#_c_699_n N_SET_B_c_836_n 0.0292376f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_620 N_A_612_74#_c_703_n N_SET_B_c_836_n 0.00150495f $X=4.935 $Y=1.285 $X2=0
+ $Y2=0
cc_621 N_A_612_74#_M1038_g N_SET_B_c_837_n 0.0172323f $X=4.86 $Y=2.525 $X2=0
+ $Y2=0
cc_622 N_A_612_74#_c_699_n N_SET_B_c_837_n 0.00115559f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_623 N_A_612_74#_c_701_n N_A_225_74#_c_956_n 3.27724e-19 $X=3.41 $Y=1.215
+ $X2=0 $Y2=0
cc_624 N_A_612_74#_c_696_n N_A_225_74#_M1023_g 0.00260688f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_625 N_A_612_74#_c_709_n N_A_225_74#_M1002_g 0.00631895f $X=3.28 $Y=2.515
+ $X2=0 $Y2=0
cc_626 N_A_612_74#_c_700_n N_A_225_74#_M1002_g 0.00274132f $X=3.285 $Y=2.295
+ $X2=0 $Y2=0
cc_627 N_A_612_74#_M1038_g N_A_225_74#_c_972_n 0.0105864f $X=4.86 $Y=2.525 $X2=0
+ $Y2=0
cc_628 N_A_612_74#_M1033_g N_A_225_74#_c_972_n 0.0124851f $X=6.025 $Y=2.235
+ $X2=0 $Y2=0
cc_629 N_A_612_74#_M1033_g N_A_225_74#_c_959_n 0.0439011f $X=6.025 $Y=2.235
+ $X2=0 $Y2=0
cc_630 N_A_612_74#_M1033_g N_A_1324_392#_c_1229_n 6.56447e-19 $X=6.025 $Y=2.235
+ $X2=0 $Y2=0
cc_631 N_A_612_74#_c_709_n N_A_27_74#_c_1497_n 0.0184847f $X=3.28 $Y=2.515 $X2=0
+ $Y2=0
cc_632 N_A_612_74#_c_700_n N_A_27_74#_c_1497_n 0.00522751f $X=3.285 $Y=2.295
+ $X2=0 $Y2=0
cc_633 N_A_612_74#_M1033_g N_VPWR_c_1562_n 0.00969538f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_634 N_A_612_74#_M1033_g N_VPWR_c_1558_n 0.00110204f $X=6.025 $Y=2.235 $X2=0
+ $Y2=0
cc_635 N_A_612_74#_c_693_n N_VGND_c_1813_n 0.00327534f $X=5.1 $Y=1.12 $X2=0
+ $Y2=0
cc_636 N_A_612_74#_c_696_n N_VGND_c_1813_n 0.00786568f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_637 N_A_612_74#_c_702_n N_VGND_c_1813_n 0.00302077f $X=4.05 $Y=1.215 $X2=0
+ $Y2=0
cc_638 N_A_612_74#_M1028_g N_VGND_c_1814_n 0.0144111f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_639 N_A_612_74#_c_699_n N_VGND_c_1814_n 0.010974f $X=5.805 $Y=1.285 $X2=0
+ $Y2=0
cc_640 N_A_612_74#_c_704_n N_VGND_c_1814_n 0.0156226f $X=5.97 $Y=1.285 $X2=0
+ $Y2=0
cc_641 N_A_612_74#_c_705_n N_VGND_c_1814_n 0.00133381f $X=5.97 $Y=1.365 $X2=0
+ $Y2=0
cc_642 N_A_612_74#_c_693_n N_VGND_c_1819_n 0.00417521f $X=5.1 $Y=1.12 $X2=0
+ $Y2=0
cc_643 N_A_612_74#_c_696_n N_VGND_c_1822_n 0.0109942f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_644 N_A_612_74#_M1028_g N_VGND_c_1829_n 0.00383152f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_645 N_A_612_74#_c_693_n N_VGND_c_1833_n 0.00479212f $X=5.1 $Y=1.12 $X2=0
+ $Y2=0
cc_646 N_A_612_74#_M1028_g N_VGND_c_1833_n 0.00758607f $X=6.05 $Y=0.69 $X2=0
+ $Y2=0
cc_647 N_A_612_74#_c_696_n N_VGND_c_1833_n 0.00904371f $X=3.37 $Y=0.58 $X2=0
+ $Y2=0
cc_648 N_SET_B_M1011_g N_A_225_74#_c_972_n 0.0109545f $X=5.31 $Y=2.525 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_833_n N_A_225_74#_c_958_n 0.00400315f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_833_n N_A_225_74#_c_959_n 0.00599883f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_651 N_SET_B_c_833_n N_A_225_74#_M1015_g 0.00633119f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_829_n N_A_1484_62#_M1007_g 0.040286f $X=7.885 $Y=0.935 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_830_n N_A_1484_62#_M1007_g 0.00387759f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_832_n N_A_1484_62#_M1014_g 0.0541219f $X=8.31 $Y=1.85 $X2=0
+ $Y2=0
cc_655 N_SET_B_c_833_n N_A_1484_62#_M1014_g 0.00374132f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_838_n N_A_1484_62#_M1014_g 0.00130941f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_830_n N_A_1484_62#_c_1129_n 0.0102598f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_833_n N_A_1484_62#_c_1129_n 0.0238932f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_659 SET_B N_A_1484_62#_c_1129_n 2.66384e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_660 N_SET_B_c_838_n N_A_1484_62#_c_1129_n 0.0214964f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_661 N_SET_B_c_829_n N_A_1484_62#_c_1130_n 0.0046649f $X=7.885 $Y=0.935 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_830_n N_A_1484_62#_c_1130_n 0.018828f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_833_n N_A_1484_62#_c_1130_n 0.00842616f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_664 SET_B N_A_1484_62#_c_1130_n 0.001949f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_665 N_SET_B_c_838_n N_A_1484_62#_c_1130_n 0.0251801f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_829_n N_A_1484_62#_c_1144_n 0.00326479f $X=7.885 $Y=0.935 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_830_n N_A_1484_62#_c_1144_n 0.00123586f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_830_n N_A_1484_62#_c_1134_n 0.0230148f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_833_n N_A_1484_62#_c_1134_n 0.00840235f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_838_n N_A_1484_62#_c_1134_n 0.00111154f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_831_n N_A_1324_392#_c_1210_n 0.0121016f $X=8.31 $Y=1.645 $X2=0
+ $Y2=0
cc_672 N_SET_B_M1019_g N_A_1324_392#_c_1210_n 0.0141535f $X=8.195 $Y=2.75 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_830_n N_A_1324_392#_M1005_g 0.0053109f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_838_n N_A_1324_392#_M1005_g 0.00102865f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_833_n N_A_1324_392#_c_1227_n 0.00168835f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_676 N_SET_B_c_833_n N_A_1324_392#_c_1216_n 0.0101492f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_677 N_SET_B_M1019_g N_A_1324_392#_c_1230_n 0.01124f $X=8.195 $Y=2.75 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_833_n N_A_1324_392#_c_1230_n 0.012116f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_838_n N_A_1324_392#_c_1230_n 0.00197365f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_680 N_SET_B_M1019_g N_A_1324_392#_c_1231_n 0.00956346f $X=8.195 $Y=2.75 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_830_n N_A_1324_392#_c_1217_n 0.00165128f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_682 N_SET_B_M1019_g N_A_1324_392#_c_1217_n 0.00252386f $X=8.195 $Y=2.75 $X2=0
+ $Y2=0
cc_683 SET_B N_A_1324_392#_c_1217_n 0.00699971f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_684 N_SET_B_c_838_n N_A_1324_392#_c_1217_n 0.0218297f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_830_n N_A_1324_392#_c_1218_n 0.0121016f $X=8.31 $Y=1.385 $X2=0
+ $Y2=0
cc_686 SET_B N_A_1324_392#_c_1218_n 0.00410251f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_687 N_SET_B_c_838_n N_A_1324_392#_c_1218_n 0.0022247f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_833_n N_A_1324_392#_c_1220_n 0.020282f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_689 N_SET_B_M1019_g N_A_1324_392#_c_1234_n 5.38189e-19 $X=8.195 $Y=2.75 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_833_n N_A_1324_392#_c_1234_n 0.00323313f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_691 N_SET_B_M1019_g N_A_1324_392#_c_1235_n 0.00484387f $X=8.195 $Y=2.75 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_832_n N_A_1324_392#_c_1235_n 0.00153883f $X=8.31 $Y=1.85 $X2=0
+ $Y2=0
cc_693 SET_B N_A_1324_392#_c_1235_n 0.00301214f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_694 N_SET_B_c_838_n N_A_1324_392#_c_1235_n 0.00864852f $X=8.35 $Y=1.345 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_833_n N_VPWR_M1011_d 0.00248692f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_696 N_SET_B_M1011_g N_VPWR_c_1562_n 0.00133144f $X=5.31 $Y=2.525 $X2=0 $Y2=0
cc_697 N_SET_B_M1019_g N_VPWR_c_1563_n 0.0027763f $X=8.195 $Y=2.75 $X2=0 $Y2=0
cc_698 N_SET_B_M1019_g N_VPWR_c_1564_n 0.00338437f $X=8.195 $Y=2.75 $X2=0 $Y2=0
cc_699 N_SET_B_M1019_g N_VPWR_c_1578_n 0.005209f $X=8.195 $Y=2.75 $X2=0 $Y2=0
cc_700 N_SET_B_M1019_g N_VPWR_c_1558_n 0.00540654f $X=8.195 $Y=2.75 $X2=0 $Y2=0
cc_701 N_SET_B_c_833_n A_1223_347# 0.00189006f $X=8.255 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_702 N_SET_B_M1016_g N_VGND_c_1814_n 0.0111202f $X=5.49 $Y=0.8 $X2=0 $Y2=0
cc_703 N_SET_B_c_833_n N_VGND_c_1814_n 6.575e-19 $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_704 N_SET_B_M1016_g N_VGND_c_1819_n 0.00434252f $X=5.49 $Y=0.8 $X2=0 $Y2=0
cc_705 N_SET_B_c_829_n N_VGND_c_1829_n 0.00438299f $X=7.885 $Y=0.935 $X2=0 $Y2=0
cc_706 N_SET_B_c_829_n N_VGND_c_1830_n 0.0103808f $X=7.885 $Y=0.935 $X2=0 $Y2=0
cc_707 N_SET_B_c_830_n N_VGND_c_1830_n 0.00175578f $X=8.31 $Y=1.385 $X2=0 $Y2=0
cc_708 N_SET_B_M1016_g N_VGND_c_1833_n 0.00479212f $X=5.49 $Y=0.8 $X2=0 $Y2=0
cc_709 N_SET_B_c_829_n N_VGND_c_1833_n 0.00436392f $X=7.885 $Y=0.935 $X2=0 $Y2=0
cc_710 N_A_225_74#_M1015_g N_A_1484_62#_M1007_g 0.0609879f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_711 N_A_225_74#_M1015_g N_A_1484_62#_M1014_g 0.00359614f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_712 N_A_225_74#_M1025_g N_A_1324_392#_c_1227_n 0.00346582f $X=6.53 $Y=2.46
+ $X2=0 $Y2=0
cc_713 N_A_225_74#_c_958_n N_A_1324_392#_c_1227_n 0.00551143f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_714 N_A_225_74#_c_958_n N_A_1324_392#_c_1216_n 0.00171411f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_715 N_A_225_74#_M1015_g N_A_1324_392#_c_1216_n 0.0138144f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_716 N_A_225_74#_M1025_g N_A_1324_392#_c_1229_n 0.00924668f $X=6.53 $Y=2.46
+ $X2=0 $Y2=0
cc_717 N_A_225_74#_c_958_n N_A_1324_392#_c_1229_n 0.00485374f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_718 N_A_225_74#_M1015_g N_A_1324_392#_c_1219_n 0.00761503f $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_719 N_A_225_74#_c_958_n N_A_1324_392#_c_1220_n 0.0193936f $X=7.03 $Y=1.735
+ $X2=0 $Y2=0
cc_720 N_A_225_74#_M1015_g N_A_1324_392#_c_1220_n 9.78128e-19 $X=7.105 $Y=0.65
+ $X2=0 $Y2=0
cc_721 N_A_225_74#_M1024_s N_A_27_74#_c_1496_n 0.0117665f $X=1.145 $Y=1.84 $X2=0
+ $Y2=0
cc_722 N_A_225_74#_c_981_n N_A_27_74#_c_1496_n 0.00567797f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_723 N_A_225_74#_c_983_n N_A_27_74#_c_1496_n 0.0326558f $X=1.455 $Y=1.895
+ $X2=0 $Y2=0
cc_724 N_A_225_74#_M1027_g N_A_27_74#_c_1497_n 0.0165411f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_725 N_A_225_74#_c_968_n N_A_27_74#_c_1497_n 0.0259855f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_726 N_A_225_74#_c_963_n N_A_27_74#_c_1497_n 0.00191316f $X=2.41 $Y=1.515
+ $X2=0 $Y2=0
cc_727 N_A_225_74#_c_981_n N_A_27_74#_c_1497_n 0.0263833f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_728 N_A_225_74#_M1018_g N_A_27_74#_c_1491_n 9.17507e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_729 N_A_225_74#_M1027_g N_A_27_74#_c_1491_n 0.00121124f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_730 N_A_225_74#_c_968_n N_A_27_74#_c_1491_n 0.00915392f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_731 N_A_225_74#_c_956_n N_A_27_74#_c_1491_n 0.00588052f $X=2.91 $Y=1.14 $X2=0
+ $Y2=0
cc_732 N_A_225_74#_M1023_g N_A_27_74#_c_1491_n 0.00249586f $X=2.985 $Y=0.58
+ $X2=0 $Y2=0
cc_733 N_A_225_74#_c_962_n N_A_27_74#_c_1491_n 0.0199619f $X=2.485 $Y=1.14 $X2=0
+ $Y2=0
cc_734 N_A_225_74#_c_981_n N_A_27_74#_c_1491_n 0.0136281f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_735 N_A_225_74#_c_965_n N_A_27_74#_c_1491_n 0.0265108f $X=2.11 $Y=1.515 $X2=0
+ $Y2=0
cc_736 N_A_225_74#_M1027_g N_A_27_74#_c_1541_n 0.00236708f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_737 N_A_225_74#_c_981_n N_A_27_74#_c_1541_n 0.00973529f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_738 N_A_225_74#_c_956_n N_A_27_74#_c_1493_n 0.00616968f $X=2.91 $Y=1.14 $X2=0
+ $Y2=0
cc_739 N_A_225_74#_M1023_g N_A_27_74#_c_1493_n 0.0066603f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_740 N_A_225_74#_c_962_n N_A_27_74#_c_1493_n 9.04452e-19 $X=2.485 $Y=1.14
+ $X2=0 $Y2=0
cc_741 N_A_225_74#_c_981_n N_VPWR_M1024_d 0.00168828f $X=1.945 $Y=1.805 $X2=0
+ $Y2=0
cc_742 N_A_225_74#_M1027_g N_VPWR_c_1560_n 0.00921044f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_743 N_A_225_74#_c_970_n N_VPWR_c_1560_n 0.00241896f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_744 N_A_225_74#_M1002_g N_VPWR_c_1561_n 8.25145e-19 $X=3.505 $Y=2.525 $X2=0
+ $Y2=0
cc_745 N_A_225_74#_c_972_n N_VPWR_c_1561_n 0.016146f $X=6.44 $Y=3.15 $X2=0 $Y2=0
cc_746 N_A_225_74#_c_972_n N_VPWR_c_1562_n 0.0218775f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_747 N_A_225_74#_M1025_g N_VPWR_c_1562_n 0.00598235f $X=6.53 $Y=2.46 $X2=0
+ $Y2=0
cc_748 N_A_225_74#_c_972_n N_VPWR_c_1571_n 0.00411927f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_749 N_A_225_74#_c_972_n N_VPWR_c_1572_n 0.0365645f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_750 N_A_225_74#_M1027_g N_VPWR_c_1576_n 0.00460063f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_751 N_A_225_74#_c_970_n N_VPWR_c_1576_n 0.0367413f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_752 N_A_225_74#_c_972_n N_VPWR_c_1577_n 0.0245531f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_753 N_A_225_74#_M1027_g N_VPWR_c_1558_n 0.00909358f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_754 N_A_225_74#_c_969_n N_VPWR_c_1558_n 0.0201297f $X=3.415 $Y=3.15 $X2=0
+ $Y2=0
cc_755 N_A_225_74#_c_970_n N_VPWR_c_1558_n 0.00599933f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_756 N_A_225_74#_c_972_n N_VPWR_c_1558_n 0.0938983f $X=6.44 $Y=3.15 $X2=0
+ $Y2=0
cc_757 N_A_225_74#_c_979_n N_VPWR_c_1558_n 0.00445015f $X=3.505 $Y=3.15 $X2=0
+ $Y2=0
cc_758 N_A_225_74#_c_966_n N_VGND_c_1810_n 0.0371671f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_759 N_A_225_74#_c_966_n N_VGND_c_1811_n 0.0212023f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_760 N_A_225_74#_M1018_g N_VGND_c_1812_n 0.0115741f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_761 N_A_225_74#_c_966_n N_VGND_c_1812_n 0.0263763f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_762 N_A_225_74#_M1018_g N_VGND_c_1822_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_763 N_A_225_74#_M1023_g N_VGND_c_1822_n 0.00278159f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_764 N_A_225_74#_M1015_g N_VGND_c_1829_n 8.27887e-19 $X=7.105 $Y=0.65 $X2=0
+ $Y2=0
cc_765 N_A_225_74#_M1018_g N_VGND_c_1833_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_766 N_A_225_74#_M1023_g N_VGND_c_1833_n 0.00359882f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_767 N_A_225_74#_c_966_n N_VGND_c_1833_n 0.0168959f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_768 N_A_1484_62#_c_1133_n N_A_1324_392#_c_1210_n 0.0285604f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_769 N_A_1484_62#_c_1130_n N_A_1324_392#_M1005_g 0.0116315f $X=9.12 $Y=0.925
+ $X2=0 $Y2=0
cc_770 N_A_1484_62#_c_1131_n N_A_1324_392#_M1005_g 0.0110008f $X=9.285 $Y=0.65
+ $X2=0 $Y2=0
cc_771 N_A_1484_62#_c_1132_n N_A_1324_392#_M1005_g 0.00495915f $X=9.285 $Y=0.925
+ $X2=0 $Y2=0
cc_772 N_A_1484_62#_c_1133_n N_A_1324_392#_M1005_g 0.0127661f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_773 N_A_1484_62#_c_1136_n N_A_1324_392#_M1012_g 0.00614026f $X=9.395 $Y=2.815
+ $X2=0 $Y2=0
cc_774 N_A_1484_62#_c_1133_n N_A_1324_392#_c_1212_n 0.0212496f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_775 N_A_1484_62#_c_1133_n N_A_1324_392#_M1000_g 5.80505e-19 $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_776 N_A_1484_62#_c_1133_n N_A_1324_392#_c_1215_n 0.00653497f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_777 N_A_1484_62#_M1014_g N_A_1324_392#_c_1229_n 9.64533e-19 $X=7.745 $Y=2.75
+ $X2=0 $Y2=0
cc_778 N_A_1484_62#_M1014_g N_A_1324_392#_c_1230_n 0.0104411f $X=7.745 $Y=2.75
+ $X2=0 $Y2=0
cc_779 N_A_1484_62#_c_1129_n N_A_1324_392#_c_1230_n 0.00172307f $X=7.71 $Y=1.49
+ $X2=0 $Y2=0
cc_780 N_A_1484_62#_M1014_g N_A_1324_392#_c_1231_n 5.30739e-19 $X=7.745 $Y=2.75
+ $X2=0 $Y2=0
cc_781 N_A_1484_62#_c_1133_n N_A_1324_392#_c_1232_n 0.0135416f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_782 N_A_1484_62#_c_1130_n N_A_1324_392#_c_1217_n 0.0144687f $X=9.12 $Y=0.925
+ $X2=0 $Y2=0
cc_783 N_A_1484_62#_c_1133_n N_A_1324_392#_c_1217_n 0.0696093f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_784 N_A_1484_62#_c_1130_n N_A_1324_392#_c_1218_n 0.00126969f $X=9.12 $Y=0.925
+ $X2=0 $Y2=0
cc_785 N_A_1484_62#_c_1132_n N_A_1324_392#_c_1218_n 0.00171994f $X=9.285
+ $Y=0.925 $X2=0 $Y2=0
cc_786 N_A_1484_62#_M1014_g N_A_1324_392#_c_1234_n 0.00986239f $X=7.745 $Y=2.75
+ $X2=0 $Y2=0
cc_787 N_A_1484_62#_c_1129_n N_A_1324_392#_c_1234_n 0.00209394f $X=7.71 $Y=1.49
+ $X2=0 $Y2=0
cc_788 N_A_1484_62#_c_1134_n N_A_1324_392#_c_1234_n 5.89701e-19 $X=7.745 $Y=1.49
+ $X2=0 $Y2=0
cc_789 N_A_1484_62#_c_1131_n N_A_1940_74#_c_1383_n 0.0282823f $X=9.285 $Y=0.65
+ $X2=0 $Y2=0
cc_790 N_A_1484_62#_c_1132_n N_A_1940_74#_c_1383_n 0.0121618f $X=9.285 $Y=0.925
+ $X2=0 $Y2=0
cc_791 N_A_1484_62#_c_1133_n N_A_1940_74#_c_1383_n 0.0198356f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_792 N_A_1484_62#_c_1133_n N_A_1940_74#_c_1385_n 0.0105853f $X=9.395 $Y=2.65
+ $X2=0 $Y2=0
cc_793 N_A_1484_62#_M1014_g N_VPWR_c_1563_n 0.00287402f $X=7.745 $Y=2.75 $X2=0
+ $Y2=0
cc_794 N_A_1484_62#_c_1136_n N_VPWR_c_1564_n 0.011548f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_795 N_A_1484_62#_c_1136_n N_VPWR_c_1565_n 0.0244397f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_796 N_A_1484_62#_c_1133_n N_VPWR_c_1565_n 0.042748f $X=9.395 $Y=2.65 $X2=0
+ $Y2=0
cc_797 N_A_1484_62#_M1014_g N_VPWR_c_1577_n 0.00502389f $X=7.745 $Y=2.75 $X2=0
+ $Y2=0
cc_798 N_A_1484_62#_c_1136_n N_VPWR_c_1579_n 0.0142041f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_799 N_A_1484_62#_M1014_g N_VPWR_c_1558_n 0.00539457f $X=7.745 $Y=2.75 $X2=0
+ $Y2=0
cc_800 N_A_1484_62#_c_1136_n N_VPWR_c_1558_n 0.0118403f $X=9.395 $Y=2.815 $X2=0
+ $Y2=0
cc_801 N_A_1484_62#_c_1130_n N_VGND_M1004_d 0.0100699f $X=9.12 $Y=0.925 $X2=0
+ $Y2=0
cc_802 N_A_1484_62#_c_1131_n N_VGND_c_1823_n 0.0112889f $X=9.285 $Y=0.65 $X2=0
+ $Y2=0
cc_803 N_A_1484_62#_M1007_g N_VGND_c_1829_n 0.00527445f $X=7.495 $Y=0.65 $X2=0
+ $Y2=0
cc_804 N_A_1484_62#_M1007_g N_VGND_c_1830_n 0.00104583f $X=7.495 $Y=0.65 $X2=0
+ $Y2=0
cc_805 N_A_1484_62#_c_1130_n N_VGND_c_1830_n 0.0747503f $X=9.12 $Y=0.925 $X2=0
+ $Y2=0
cc_806 N_A_1484_62#_c_1131_n N_VGND_c_1830_n 0.0102732f $X=9.285 $Y=0.65 $X2=0
+ $Y2=0
cc_807 N_A_1484_62#_M1007_g N_VGND_c_1833_n 0.00523671f $X=7.495 $Y=0.65 $X2=0
+ $Y2=0
cc_808 N_A_1484_62#_c_1130_n N_VGND_c_1833_n 0.010553f $X=9.12 $Y=0.925 $X2=0
+ $Y2=0
cc_809 N_A_1484_62#_c_1144_n N_VGND_c_1833_n 0.0126596f $X=7.875 $Y=0.925 $X2=0
+ $Y2=0
cc_810 N_A_1484_62#_c_1131_n N_VGND_c_1833_n 0.0115369f $X=9.285 $Y=0.65 $X2=0
+ $Y2=0
cc_811 N_A_1484_62#_c_1144_n A_1514_88# 0.00299242f $X=7.875 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_812 N_A_1324_392#_M1000_g N_A_1940_74#_c_1372_n 0.0119421f $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_813 N_A_1324_392#_c_1214_n N_A_1940_74#_c_1374_n 0.0072081f $X=10.505 $Y=1.69
+ $X2=0 $Y2=0
cc_814 N_A_1324_392#_c_1215_n N_A_1940_74#_c_1374_n 0.0119421f $X=10.055 $Y=1.37
+ $X2=0 $Y2=0
cc_815 N_A_1324_392#_c_1214_n N_A_1940_74#_M1022_g 0.0213464f $X=10.505 $Y=1.69
+ $X2=0 $Y2=0
cc_816 N_A_1324_392#_c_1214_n N_A_1940_74#_c_1380_n 0.00148303f $X=10.505
+ $Y=1.69 $X2=0 $Y2=0
cc_817 N_A_1324_392#_M1005_g N_A_1940_74#_c_1383_n 0.00323395f $X=9.07 $Y=0.65
+ $X2=0 $Y2=0
cc_818 N_A_1324_392#_M1000_g N_A_1940_74#_c_1383_n 0.0230336f $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_819 N_A_1324_392#_c_1212_n N_A_1940_74#_c_1384_n 0.00238371f $X=10.055
+ $Y=1.492 $X2=0 $Y2=0
cc_820 N_A_1324_392#_M1000_g N_A_1940_74#_c_1384_n 0.00759579f $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_821 N_A_1324_392#_c_1215_n N_A_1940_74#_c_1384_n 0.00825982f $X=10.055
+ $Y=1.37 $X2=0 $Y2=0
cc_822 N_A_1324_392#_c_1212_n N_A_1940_74#_c_1385_n 0.0198827f $X=10.055
+ $Y=1.492 $X2=0 $Y2=0
cc_823 N_A_1324_392#_c_1223_n N_A_1940_74#_c_1392_n 0.0168202f $X=10.145
+ $Y=1.765 $X2=0 $Y2=0
cc_824 N_A_1324_392#_c_1214_n N_A_1940_74#_c_1392_n 0.00735076f $X=10.505
+ $Y=1.69 $X2=0 $Y2=0
cc_825 N_A_1324_392#_c_1225_n N_A_1940_74#_c_1392_n 0.0148637f $X=10.595
+ $Y=1.765 $X2=0 $Y2=0
cc_826 N_A_1324_392#_c_1215_n N_A_1940_74#_c_1392_n 0.00504166f $X=10.055
+ $Y=1.37 $X2=0 $Y2=0
cc_827 N_A_1324_392#_c_1214_n N_A_1940_74#_c_1386_n 0.00975883f $X=10.505
+ $Y=1.69 $X2=0 $Y2=0
cc_828 N_A_1324_392#_M1000_g N_A_1940_74#_c_1387_n 6.82259e-19 $X=10.13 $Y=0.74
+ $X2=0 $Y2=0
cc_829 N_A_1324_392#_c_1214_n N_A_1940_74#_c_1387_n 0.00687641f $X=10.505
+ $Y=1.69 $X2=0 $Y2=0
cc_830 N_A_1324_392#_c_1215_n N_A_1940_74#_c_1387_n 0.0148745f $X=10.055 $Y=1.37
+ $X2=0 $Y2=0
cc_831 N_A_1324_392#_c_1229_n N_VPWR_c_1562_n 0.0088797f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_832 N_A_1324_392#_c_1229_n N_VPWR_c_1563_n 0.0050121f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_833 N_A_1324_392#_c_1230_n N_VPWR_c_1563_n 0.0130545f $X=8.255 $Y=2.395 $X2=0
+ $Y2=0
cc_834 N_A_1324_392#_c_1231_n N_VPWR_c_1563_n 0.0115095f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_835 N_A_1324_392#_M1012_g N_VPWR_c_1564_n 0.00501904f $X=9.17 $Y=2.75 $X2=0
+ $Y2=0
cc_836 N_A_1324_392#_c_1231_n N_VPWR_c_1564_n 0.0244395f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_837 N_A_1324_392#_c_1232_n N_VPWR_c_1564_n 0.0220489f $X=8.78 $Y=2.395 $X2=0
+ $Y2=0
cc_838 N_A_1324_392#_c_1233_n N_VPWR_c_1564_n 0.00149279f $X=8.945 $Y=2.215
+ $X2=0 $Y2=0
cc_839 N_A_1324_392#_M1012_g N_VPWR_c_1565_n 0.00334936f $X=9.17 $Y=2.75 $X2=0
+ $Y2=0
cc_840 N_A_1324_392#_c_1212_n N_VPWR_c_1565_n 0.0048892f $X=10.055 $Y=1.492
+ $X2=0 $Y2=0
cc_841 N_A_1324_392#_c_1223_n N_VPWR_c_1565_n 0.00873579f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_842 N_A_1324_392#_c_1223_n N_VPWR_c_1566_n 0.00465228f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_843 N_A_1324_392#_c_1225_n N_VPWR_c_1566_n 0.00465228f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_844 N_A_1324_392#_c_1225_n N_VPWR_c_1567_n 0.00790409f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_845 N_A_1324_392#_c_1228_n N_VPWR_c_1577_n 0.00385839f $X=7.545 $Y=2.565
+ $X2=0 $Y2=0
cc_846 N_A_1324_392#_c_1229_n N_VPWR_c_1577_n 0.0293565f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_847 N_A_1324_392#_c_1234_n N_VPWR_c_1577_n 0.00227646f $X=7.63 $Y=2.395 $X2=0
+ $Y2=0
cc_848 N_A_1324_392#_c_1231_n N_VPWR_c_1578_n 0.0145333f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_849 N_A_1324_392#_M1012_g N_VPWR_c_1579_n 0.005209f $X=9.17 $Y=2.75 $X2=0
+ $Y2=0
cc_850 N_A_1324_392#_M1012_g N_VPWR_c_1558_n 0.00904034f $X=9.17 $Y=2.75 $X2=0
+ $Y2=0
cc_851 N_A_1324_392#_c_1223_n N_VPWR_c_1558_n 0.00555093f $X=10.145 $Y=1.765
+ $X2=0 $Y2=0
cc_852 N_A_1324_392#_c_1225_n N_VPWR_c_1558_n 0.00555093f $X=10.595 $Y=1.765
+ $X2=0 $Y2=0
cc_853 N_A_1324_392#_c_1228_n N_VPWR_c_1558_n 0.00697082f $X=7.545 $Y=2.565
+ $X2=0 $Y2=0
cc_854 N_A_1324_392#_c_1229_n N_VPWR_c_1558_n 0.0244131f $X=7.265 $Y=2.565 $X2=0
+ $Y2=0
cc_855 N_A_1324_392#_c_1230_n N_VPWR_c_1558_n 0.0113321f $X=8.255 $Y=2.395 $X2=0
+ $Y2=0
cc_856 N_A_1324_392#_c_1231_n N_VPWR_c_1558_n 0.0119681f $X=8.42 $Y=2.75 $X2=0
+ $Y2=0
cc_857 N_A_1324_392#_c_1232_n N_VPWR_c_1558_n 0.010474f $X=8.78 $Y=2.395 $X2=0
+ $Y2=0
cc_858 N_A_1324_392#_c_1234_n N_VPWR_c_1558_n 0.00447679f $X=7.63 $Y=2.395 $X2=0
+ $Y2=0
cc_859 N_A_1324_392#_c_1228_n A_1483_508# 0.00159568f $X=7.545 $Y=2.565
+ $X2=-0.19 $Y2=-0.245
cc_860 N_A_1324_392#_c_1234_n A_1483_508# 0.00123523f $X=7.63 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_861 N_A_1324_392#_M1000_g N_VGND_c_1815_n 0.0163444f $X=10.13 $Y=0.74 $X2=0
+ $Y2=0
cc_862 N_A_1324_392#_c_1215_n N_VGND_c_1815_n 0.00127334f $X=10.055 $Y=1.37
+ $X2=0 $Y2=0
cc_863 N_A_1324_392#_M1005_g N_VGND_c_1823_n 0.00504315f $X=9.07 $Y=0.65 $X2=0
+ $Y2=0
cc_864 N_A_1324_392#_M1000_g N_VGND_c_1823_n 0.00383152f $X=10.13 $Y=0.74 $X2=0
+ $Y2=0
cc_865 N_A_1324_392#_M1005_g N_VGND_c_1830_n 0.0100857f $X=9.07 $Y=0.65 $X2=0
+ $Y2=0
cc_866 N_A_1324_392#_M1005_g N_VGND_c_1833_n 0.00523671f $X=9.07 $Y=0.65 $X2=0
+ $Y2=0
cc_867 N_A_1324_392#_M1000_g N_VGND_c_1833_n 0.00762539f $X=10.13 $Y=0.74 $X2=0
+ $Y2=0
cc_868 N_A_1940_74#_c_1385_n N_VPWR_c_1565_n 0.013441f $X=10.01 $Y=1.405 $X2=0
+ $Y2=0
cc_869 N_A_1940_74#_c_1392_n N_VPWR_c_1565_n 0.030344f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_870 N_A_1940_74#_c_1392_n N_VPWR_c_1566_n 0.00657675f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_871 N_A_1940_74#_c_1373_n N_VPWR_c_1567_n 0.00111964f $X=10.985 $Y=1.3 $X2=0
+ $Y2=0
cc_872 N_A_1940_74#_M1022_g N_VPWR_c_1567_n 0.00429323f $X=11.115 $Y=2.4 $X2=0
+ $Y2=0
cc_873 N_A_1940_74#_c_1380_n N_VPWR_c_1567_n 5.17557e-19 $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_874 N_A_1940_74#_c_1392_n N_VPWR_c_1567_n 0.0316306f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_875 N_A_1940_74#_c_1386_n N_VPWR_c_1567_n 0.0245135f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_876 N_A_1940_74#_M1022_g N_VPWR_c_1568_n 5.53279e-19 $X=11.115 $Y=2.4 $X2=0
+ $Y2=0
cc_877 N_A_1940_74#_M1029_g N_VPWR_c_1568_n 0.0138856f $X=11.565 $Y=2.4 $X2=0
+ $Y2=0
cc_878 N_A_1940_74#_M1030_g N_VPWR_c_1568_n 0.0138034f $X=12.015 $Y=2.4 $X2=0
+ $Y2=0
cc_879 N_A_1940_74#_M1037_g N_VPWR_c_1568_n 5.21408e-19 $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_880 N_A_1940_74#_M1030_g N_VPWR_c_1570_n 5.02386e-19 $X=12.015 $Y=2.4 $X2=0
+ $Y2=0
cc_881 N_A_1940_74#_M1037_g N_VPWR_c_1570_n 0.0134762f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_882 N_A_1940_74#_M1022_g N_VPWR_c_1580_n 0.005209f $X=11.115 $Y=2.4 $X2=0
+ $Y2=0
cc_883 N_A_1940_74#_M1029_g N_VPWR_c_1580_n 0.00460063f $X=11.565 $Y=2.4 $X2=0
+ $Y2=0
cc_884 N_A_1940_74#_M1030_g N_VPWR_c_1581_n 0.00460063f $X=12.015 $Y=2.4 $X2=0
+ $Y2=0
cc_885 N_A_1940_74#_M1037_g N_VPWR_c_1581_n 0.00460063f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_886 N_A_1940_74#_M1022_g N_VPWR_c_1558_n 0.00986727f $X=11.115 $Y=2.4 $X2=0
+ $Y2=0
cc_887 N_A_1940_74#_M1029_g N_VPWR_c_1558_n 0.00908554f $X=11.565 $Y=2.4 $X2=0
+ $Y2=0
cc_888 N_A_1940_74#_M1030_g N_VPWR_c_1558_n 0.00908554f $X=12.015 $Y=2.4 $X2=0
+ $Y2=0
cc_889 N_A_1940_74#_M1037_g N_VPWR_c_1558_n 0.00908554f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_890 N_A_1940_74#_c_1392_n N_VPWR_c_1558_n 0.00992028f $X=10.37 $Y=1.985 $X2=0
+ $Y2=0
cc_891 N_A_1940_74#_c_1372_n N_Q_c_1738_n 0.00761489f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_892 N_A_1940_74#_c_1375_n N_Q_c_1738_n 0.0137392f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_893 N_A_1940_74#_c_1375_n N_Q_c_1739_n 0.0127216f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_894 N_A_1940_74#_c_1378_n N_Q_c_1739_n 0.0150954f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_895 N_A_1940_74#_c_1380_n N_Q_c_1739_n 0.0153125f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_896 N_A_1940_74#_c_1386_n N_Q_c_1739_n 0.072964f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_897 N_A_1940_74#_c_1372_n N_Q_c_1740_n 0.00276819f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_898 N_A_1940_74#_c_1373_n N_Q_c_1740_n 0.00224597f $X=10.985 $Y=1.3 $X2=0
+ $Y2=0
cc_899 N_A_1940_74#_c_1375_n N_Q_c_1740_n 0.00121617f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_900 N_A_1940_74#_c_1383_n N_Q_c_1740_n 5.79493e-19 $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_901 N_A_1940_74#_c_1386_n N_Q_c_1740_n 0.0275317f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_902 N_A_1940_74#_M1022_g N_Q_c_1745_n 0.0036068f $X=11.115 $Y=2.4 $X2=0 $Y2=0
cc_903 N_A_1940_74#_c_1380_n N_Q_c_1745_n 0.00220488f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_904 N_A_1940_74#_c_1386_n N_Q_c_1745_n 0.0234813f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_905 N_A_1940_74#_M1022_g N_Q_c_1746_n 0.0111678f $X=11.115 $Y=2.4 $X2=0 $Y2=0
cc_906 N_A_1940_74#_M1029_g N_Q_c_1746_n 3.83863e-19 $X=11.565 $Y=2.4 $X2=0
+ $Y2=0
cc_907 N_A_1940_74#_c_1378_n N_Q_c_1741_n 4.78514e-19 $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_908 N_A_1940_74#_M1034_g N_Q_c_1741_n 0.0133757f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_909 N_A_1940_74#_M1030_g N_Q_c_1747_n 3.8104e-19 $X=12.015 $Y=2.4 $X2=0 $Y2=0
cc_910 N_A_1940_74#_M1037_g N_Q_c_1747_n 3.8104e-19 $X=12.465 $Y=2.4 $X2=0 $Y2=0
cc_911 N_A_1940_74#_c_1380_n N_Q_c_1742_n 0.00213685f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_912 N_A_1940_74#_M1034_g N_Q_c_1742_n 0.0145085f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_913 N_A_1940_74#_c_1380_n N_Q_c_1743_n 0.00480942f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_914 N_A_1940_74#_M1034_g N_Q_c_1743_n 0.00162456f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_915 N_A_1940_74#_c_1380_n Q 0.0124746f $X=12.395 $Y=1.32 $X2=0 $Y2=0
cc_916 N_A_1940_74#_M1034_g Q 0.0121215f $X=12.395 $Y=0.74 $X2=0 $Y2=0
cc_917 N_A_1940_74#_c_1386_n Q 0.0100186f $X=11.83 $Y=1.485 $X2=0 $Y2=0
cc_918 N_A_1940_74#_c_1380_n Q 0.00278253f $X=12.395 $Y=1.32 $X2=0 $Y2=0
cc_919 N_A_1940_74#_M1037_g Q 0.0245319f $X=12.465 $Y=2.4 $X2=0 $Y2=0
cc_920 N_A_1940_74#_M1029_g N_Q_c_1750_n 0.0174262f $X=11.565 $Y=2.4 $X2=0 $Y2=0
cc_921 N_A_1940_74#_M1030_g N_Q_c_1750_n 0.0189673f $X=12.015 $Y=2.4 $X2=0 $Y2=0
cc_922 N_A_1940_74#_c_1380_n N_Q_c_1750_n 0.00236536f $X=12.395 $Y=1.32 $X2=0
+ $Y2=0
cc_923 N_A_1940_74#_c_1386_n N_Q_c_1750_n 0.0409106f $X=11.83 $Y=1.485 $X2=0
+ $Y2=0
cc_924 N_A_1940_74#_c_1372_n N_VGND_c_1815_n 0.00590268f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_925 N_A_1940_74#_c_1383_n N_VGND_c_1815_n 0.0308485f $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_926 N_A_1940_74#_c_1384_n N_VGND_c_1815_n 0.00164036f $X=10.205 $Y=1.405
+ $X2=0 $Y2=0
cc_927 N_A_1940_74#_c_1387_n N_VGND_c_1815_n 0.0263154f $X=10.37 $Y=1.485 $X2=0
+ $Y2=0
cc_928 N_A_1940_74#_c_1375_n N_VGND_c_1816_n 0.00322722f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_929 N_A_1940_74#_c_1378_n N_VGND_c_1816_n 0.00352244f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_930 N_A_1940_74#_M1034_g N_VGND_c_1818_n 0.0122304f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_931 N_A_1940_74#_c_1383_n N_VGND_c_1823_n 0.0146357f $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_932 N_A_1940_74#_c_1372_n N_VGND_c_1824_n 0.00434272f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_933 N_A_1940_74#_c_1375_n N_VGND_c_1824_n 0.00434272f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_934 N_A_1940_74#_c_1378_n N_VGND_c_1825_n 0.00460063f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_935 N_A_1940_74#_M1034_g N_VGND_c_1825_n 0.00434272f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_936 N_A_1940_74#_c_1372_n N_VGND_c_1833_n 0.00820772f $X=10.63 $Y=1.225 $X2=0
+ $Y2=0
cc_937 N_A_1940_74#_c_1375_n N_VGND_c_1833_n 0.00823001f $X=11.06 $Y=1.225 $X2=0
+ $Y2=0
cc_938 N_A_1940_74#_c_1378_n N_VGND_c_1833_n 0.00910475f $X=11.92 $Y=1.225 $X2=0
+ $Y2=0
cc_939 N_A_1940_74#_M1034_g N_VGND_c_1833_n 0.00824368f $X=12.395 $Y=0.74 $X2=0
+ $Y2=0
cc_940 N_A_1940_74#_c_1383_n N_VGND_c_1833_n 0.0121141f $X=9.845 $Y=0.515 $X2=0
+ $Y2=0
cc_941 N_A_27_74#_c_1497_n N_VPWR_M1024_d 9.98109e-19 $X=2.445 $Y=2.155 $X2=0
+ $Y2=0
cc_942 N_A_27_74#_c_1541_n N_VPWR_M1024_d 0.00557716f $X=1.71 $Y=2.155 $X2=0
+ $Y2=0
cc_943 N_A_27_74#_c_1495_n N_VPWR_c_1559_n 0.0131953f $X=0.28 $Y=2.73 $X2=0
+ $Y2=0
cc_944 N_A_27_74#_c_1496_n N_VPWR_c_1559_n 0.0243665f $X=1.625 $Y=2.325 $X2=0
+ $Y2=0
cc_945 N_A_27_74#_c_1496_n N_VPWR_c_1560_n 0.00216696f $X=1.625 $Y=2.325 $X2=0
+ $Y2=0
cc_946 N_A_27_74#_c_1497_n N_VPWR_c_1560_n 0.00236221f $X=2.445 $Y=2.155 $X2=0
+ $Y2=0
cc_947 N_A_27_74#_c_1541_n N_VPWR_c_1560_n 0.01132f $X=1.71 $Y=2.155 $X2=0 $Y2=0
cc_948 N_A_27_74#_c_1495_n N_VPWR_c_1574_n 0.0102563f $X=0.28 $Y=2.73 $X2=0
+ $Y2=0
cc_949 N_A_27_74#_c_1495_n N_VPWR_c_1558_n 0.0090542f $X=0.28 $Y=2.73 $X2=0
+ $Y2=0
cc_950 N_A_27_74#_c_1489_n N_VGND_c_1810_n 0.0172562f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_951 N_A_27_74#_c_1489_n N_VGND_c_1821_n 0.0109681f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_952 N_A_27_74#_c_1489_n N_VGND_c_1833_n 0.00912188f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_953 N_VPWR_c_1567_n N_Q_c_1745_n 0.0117266f $X=10.89 $Y=1.985 $X2=0 $Y2=0
cc_954 N_VPWR_c_1567_n N_Q_c_1746_n 0.0336653f $X=10.89 $Y=1.985 $X2=0 $Y2=0
cc_955 N_VPWR_c_1568_n N_Q_c_1746_n 0.0281624f $X=11.79 $Y=2.335 $X2=0 $Y2=0
cc_956 N_VPWR_c_1580_n N_Q_c_1746_n 0.0123179f $X=11.625 $Y=3.33 $X2=0 $Y2=0
cc_957 N_VPWR_c_1558_n N_Q_c_1746_n 0.0101276f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_958 N_VPWR_c_1568_n N_Q_c_1747_n 0.0281397f $X=11.79 $Y=2.335 $X2=0 $Y2=0
cc_959 N_VPWR_c_1570_n N_Q_c_1747_n 0.0255132f $X=12.69 $Y=2.405 $X2=0 $Y2=0
cc_960 N_VPWR_c_1581_n N_Q_c_1747_n 0.0101736f $X=12.525 $Y=3.33 $X2=0 $Y2=0
cc_961 N_VPWR_c_1558_n N_Q_c_1747_n 0.0084208f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_962 N_VPWR_M1037_s Q 0.00385022f $X=12.555 $Y=1.84 $X2=0 $Y2=0
cc_963 N_VPWR_c_1570_n Q 0.0212555f $X=12.69 $Y=2.405 $X2=0 $Y2=0
cc_964 N_VPWR_M1029_s N_Q_c_1750_n 0.00168016f $X=11.655 $Y=1.84 $X2=0 $Y2=0
cc_965 N_VPWR_c_1568_n N_Q_c_1750_n 0.0175329f $X=11.79 $Y=2.335 $X2=0 $Y2=0
cc_966 N_Q_c_1739_n N_VGND_M1009_s 0.0089885f $X=12.015 $Y=1.065 $X2=0 $Y2=0
cc_967 N_Q_c_1742_n N_VGND_M1034_s 0.00451232f $X=12.605 $Y=1.065 $X2=0 $Y2=0
cc_968 N_Q_c_1738_n N_VGND_c_1815_n 0.0243921f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_969 N_Q_c_1740_n N_VGND_c_1815_n 0.00711243f $X=11.01 $Y=1.065 $X2=0 $Y2=0
cc_970 N_Q_c_1738_n N_VGND_c_1816_n 0.0177638f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_971 N_Q_c_1739_n N_VGND_c_1816_n 0.0464602f $X=12.015 $Y=1.065 $X2=0 $Y2=0
cc_972 N_Q_c_1741_n N_VGND_c_1816_n 0.0183183f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_973 N_Q_c_1741_n N_VGND_c_1818_n 0.0180508f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_974 N_Q_c_1742_n N_VGND_c_1818_n 0.0270821f $X=12.605 $Y=1.065 $X2=0 $Y2=0
cc_975 N_Q_c_1738_n N_VGND_c_1824_n 0.0144922f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_976 N_Q_c_1741_n N_VGND_c_1825_n 0.0145639f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_977 N_Q_c_1738_n N_VGND_c_1833_n 0.0118826f $X=10.845 $Y=0.515 $X2=0 $Y2=0
cc_978 N_Q_c_1741_n N_VGND_c_1833_n 0.0119984f $X=12.18 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__fah_4.spice
* Created: Wed Sep  2 12:09:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fah_4.pex.spice"
.subckt sky130_fd_sc_ms__fah_4  VNB VPB A B CI VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1037 N_VGND_M1037_d N_A_M1037_g N_A_27_74#_M1037_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1038 N_A_200_74#_M1038_d N_A_M1038_g N_VGND_M1037_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_430_362#_M1007_d N_A_27_74#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.124942 AS=0.418 PD=1.14217 PS=2.8 NRD=7.296 NRS=34.86 M=1
+ R=4.93333 SA=75000.4 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1018 N_A_536_114#_M1018_d N_B_M1018_g N_A_430_362#_M1007_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.108058 PD=0.92 PS=0.987826 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1030 N_A_200_74#_M1030_d N_A_586_257#_M1030_g N_A_536_114#_M1018_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1222 AS=0.0896 PD=1.08 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1027 N_A_531_362#_M1027_d N_B_M1027_g N_A_200_74#_M1030_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1024 AS=0.1222 PD=0.96 PS=1.08 NRD=7.488 NRS=14.988 M=1 R=4.26667
+ SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1035 N_A_430_362#_M1035_d N_A_586_257#_M1035_g N_A_531_362#_M1027_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1024 PD=1.81 PS=0.96 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1025 N_A_586_257#_M1025_d N_B_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.27675 PD=2.05 PS=2.42 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_A_1278_102#_M1021_d N_A_531_362#_M1021_g N_A_1183_102#_M1021_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.122062 AS=0.208 PD=1.105 PS=1.93 NRD=1.872 NRS=9.372
+ M=1 R=4.26667 SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1040 N_A_1378_125#_M1040_d N_A_536_114#_M1040_g N_A_1278_102#_M1021_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.0896 AS=0.122062 PD=0.92 PS=1.105 NRD=0 NRS=12.18
+ M=1 R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1041 N_A_1268_379#_M1041_d N_A_531_362#_M1041_g N_A_1378_125#_M1040_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.118425 AS=0.0896 PD=1.09 PS=0.92 NRD=11.244 NRS=0
+ M=1 R=4.26667 SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1026 N_A_586_257#_M1026_d N_A_536_114#_M1026_g N_A_1268_379#_M1041_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.356425 AS=0.118425 PD=3.14 PS=1.09 NRD=94.104 NRS=0
+ M=1 R=4.26667 SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A_1378_125#_M1020_g N_A_1183_102#_M1020_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.307107 AS=0.23505 PD=1.76232 PS=2.02 NRD=79.656 NRS=14.988
+ M=1 R=4.26667 SA=75000.3 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1009 N_COUT_M1009_d N_A_1268_379#_M1009_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.355093 PD=1.02 PS=2.03768 NRD=0 NRS=68.892 M=1 R=4.93333
+ SA=75001.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1011 N_COUT_M1009_d N_A_1268_379#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.18675 PD=1.02 PS=1.45 NRD=0 NRS=32.004 M=1 R=4.93333
+ SA=75001.6 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1014 N_COUT_M1014_d N_A_1268_379#_M1014_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.18675 PD=1.02 PS=1.45 NRD=0 NRS=32.004 M=1 R=4.93333
+ SA=75002.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1022 N_COUT_M1014_d N_A_1268_379#_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.36 PD=1.02 PS=2.83 NRD=0 NRS=69.96 M=1 R=4.93333
+ SA=75002.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_CI_M1017_g N_A_1378_125#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.194087 AS=0.1824 PD=1.3913 PS=1.85 NRD=46.548 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1017_d N_A_1278_102#_M1002_g N_SUM_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.224413 AS=0.1036 PD=1.6087 PS=1.02 NRD=40.248 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_A_1278_102#_M1028_g N_SUM_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1028_d N_A_1278_102#_M1031_g N_SUM_M1031_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1042 N_VGND_M1042_d N_A_1278_102#_M1042_g N_SUM_M1031_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_27_74#_M1005_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_A_200_74#_M1006_d N_A_M1006_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_A_430_362#_M1003_d N_A_27_74#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.196 AS=0.4995 PD=1.65143 PS=3.52 NRD=8.7862 NRS=68.753 M=1
+ R=6.22222 SA=90000.3 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1033 N_A_531_362#_M1033_d N_B_M1033_g N_A_430_362#_M1003_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1155 AS=0.147 PD=1.115 PS=1.23857 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.8 SB=90001.7 A=0.1512 P=2.04 MULT=1
MM1019 N_A_200_74#_M1019_d N_A_586_257#_M1019_g N_A_531_362#_M1033_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.22685 AS=0.1155 PD=1.57 PS=1.115 NRD=50.432 NRS=0 M=1
+ R=4.66667 SA=90001.2 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1023 N_A_536_114#_M1023_d N_B_M1023_g N_A_200_74#_M1019_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.22685 PD=1.11 PS=1.57 NRD=0 NRS=50.432 M=1 R=4.66667
+ SA=90001.9 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1029 N_A_430_362#_M1029_d N_A_586_257#_M1029_g N_A_536_114#_M1023_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.1134 PD=2.24 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90002.3 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1010 N_A_586_257#_M1010_d N_B_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.214257 AS=0.3136 PD=1.68571 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1000 N_A_1268_379#_M1000_d N_A_531_362#_M1000_g N_A_586_257#_M1010_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.1743 AS=0.160693 PD=1.255 PS=1.26429 NRD=32.8202
+ NRS=18.7544 M=1 R=4.66667 SA=90000.7 SB=90004.4 A=0.1512 P=2.04 MULT=1
MM1004 N_A_1378_125#_M1004_d N_A_536_114#_M1004_g N_A_1268_379#_M1000_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.21245 AS=0.1743 PD=1.52 PS=1.255 NRD=46.4132 NRS=0
+ M=1 R=4.66667 SA=90001.3 SB=90003.8 A=0.1512 P=2.04 MULT=1
MM1043 N_A_1278_102#_M1043_d N_A_531_362#_M1043_g N_A_1378_125#_M1004_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.3234 AS=0.21245 PD=1.61 PS=1.52 NRD=116.072
+ NRS=11.7215 M=1 R=4.66667 SA=90001.5 SB=90004 A=0.1512 P=2.04 MULT=1
MM1001 N_A_1183_102#_M1001_d N_A_536_114#_M1001_g N_A_1278_102#_M1043_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.165774 AS=0.3234 PD=1.34217 PS=1.61 NRD=33.3718
+ NRS=0 M=1 R=4.66667 SA=90002.5 SB=90003 A=0.1512 P=2.04 MULT=1
MM1016 N_VPWR_M1016_d N_A_1378_125#_M1016_g N_A_1183_102#_M1001_d VPB PSHORT
+ L=0.18 W=1 AD=0.41 AS=0.197351 PD=1.90566 PS=1.59783 NRD=69.9153 NRS=0 M=1
+ R=5.55556 SA=90002.4 SB=90003 A=0.18 P=2.36 MULT=1
MM1008 N_COUT_M1008_d N_A_1268_379#_M1008_g N_VPWR_M1016_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.4592 PD=1.39 PS=2.13434 NRD=0 NRS=62.4293 M=1 R=6.22222
+ SA=90002.9 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1024 N_COUT_M1008_d N_A_1268_379#_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.280475 PD=1.39 PS=1.795 NRD=0 NRS=34.3568 M=1 R=6.22222
+ SA=90003.4 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1036 N_COUT_M1036_d N_A_1268_379#_M1036_g N_VPWR_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.280475 PD=1.39 PS=1.795 NRD=0 NRS=34.3568 M=1 R=6.22222
+ SA=90004 SB=90001 A=0.2016 P=2.6 MULT=1
MM1039 N_COUT_M1036_d N_A_1268_379#_M1039_g N_VPWR_M1039_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.8746 PD=1.39 PS=4.01 NRD=0 NRS=127.676 M=1 R=6.22222
+ SA=90004.5 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1034 N_VPWR_M1034_d N_CI_M1034_g N_A_1378_125#_M1034_s VPB PSHORT L=0.18 W=1
+ AD=0.209717 AS=0.28 PD=1.43868 PS=2.56 NRD=16.0752 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1012 N_SUM_M1012_d N_A_1278_102#_M1012_g N_VPWR_M1034_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.234883 PD=1.39 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.7 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1013 N_SUM_M1012_d N_A_1278_102#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.2 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1015 N_SUM_M1015_d N_A_1278_102#_M1015_g N_VPWR_M1013_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1568 AS=0.2016 PD=1.4 PS=1.48 NRD=0.8668 NRS=6.1464 M=1 R=6.22222
+ SA=90001.7 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1032 N_SUM_M1015_d N_A_1278_102#_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1568 AS=0.3136 PD=1.4 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX44_noxref VNB VPB NWDIODE A=29.3716 P=35.37
c_164 VNB 0 3.55461e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__fah_4.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__nand3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand3b_4 A_N B C VGND VNB VPB VPWR Y
M1000 VGND A_N a_89_172# VNB nlowvt w=740000u l=150000u
+  ad=1.1492e+12p pd=8.02e+06u as=1.9515e+11p ps=2.05e+06u
M1001 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=4.8426e+12p pd=1.966e+07u as=1.3328e+12p ps=9.1e+06u
M1002 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_744_74# B a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=1.0672e+12p pd=1.036e+07u as=8.806e+11p ps=8.3e+06u
M1004 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_744_74# a_89_172# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1006 a_297_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_744_74# B a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_89_172# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_89_172# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_297_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_89_172# a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_89_172# a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_297_82# B a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_297_82# B a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_89_172# A_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1018 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_744_74# a_89_172# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A_N a_89_172# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


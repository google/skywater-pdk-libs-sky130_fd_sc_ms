* File: sky130_fd_sc_ms__dlclkp_4.pxi.spice
* Created: Wed Sep  2 12:04:50 2020
* 
x_PM_SKY130_FD_SC_MS__DLCLKP_4%A_84_48# N_A_84_48#_M1018_d N_A_84_48#_M1000_d
+ N_A_84_48#_c_150_n N_A_84_48#_M1020_g N_A_84_48#_M1003_g N_A_84_48#_c_152_n
+ N_A_84_48#_c_153_n N_A_84_48#_c_162_p N_A_84_48#_c_222_p N_A_84_48#_c_154_n
+ N_A_84_48#_c_190_p N_A_84_48#_c_209_p N_A_84_48#_c_177_p N_A_84_48#_c_227_p
+ N_A_84_48#_c_159_n N_A_84_48#_c_155_n N_A_84_48#_c_156_n
+ PM_SKY130_FD_SC_MS__DLCLKP_4%A_84_48#
x_PM_SKY130_FD_SC_MS__DLCLKP_4%GATE N_GATE_M1023_g N_GATE_M1017_g GATE
+ N_GATE_c_244_n PM_SKY130_FD_SC_MS__DLCLKP_4%GATE
x_PM_SKY130_FD_SC_MS__DLCLKP_4%A_334_54# N_A_334_54#_M1019_s N_A_334_54#_M1012_s
+ N_A_334_54#_c_278_n N_A_334_54#_M1018_g N_A_334_54#_M1024_g
+ N_A_334_54#_M1015_g N_A_334_54#_M1025_g N_A_334_54#_c_280_n
+ N_A_334_54#_c_281_n N_A_334_54#_c_290_n N_A_334_54#_c_308_n
+ N_A_334_54#_c_291_n N_A_334_54#_c_282_n N_A_334_54#_c_356_p
+ N_A_334_54#_c_293_n N_A_334_54#_c_357_p N_A_334_54#_c_283_n
+ N_A_334_54#_c_284_n N_A_334_54#_c_294_n N_A_334_54#_c_285_n
+ N_A_334_54#_c_286_n PM_SKY130_FD_SC_MS__DLCLKP_4%A_334_54#
x_PM_SKY130_FD_SC_MS__DLCLKP_4%A_334_338# N_A_334_338#_M1025_d
+ N_A_334_338#_M1015_d N_A_334_338#_c_409_n N_A_334_338#_M1000_g
+ N_A_334_338#_c_402_n N_A_334_338#_c_411_n N_A_334_338#_M1011_g
+ N_A_334_338#_c_404_n N_A_334_338#_c_405_n N_A_334_338#_c_406_n
+ N_A_334_338#_c_414_n N_A_334_338#_c_407_n N_A_334_338#_c_408_n
+ PM_SKY130_FD_SC_MS__DLCLKP_4%A_334_338#
x_PM_SKY130_FD_SC_MS__DLCLKP_4%A_27_74# N_A_27_74#_M1020_s N_A_27_74#_M1003_s
+ N_A_27_74#_c_481_n N_A_27_74#_M1002_g N_A_27_74#_M1001_g N_A_27_74#_M1021_g
+ N_A_27_74#_M1014_g N_A_27_74#_c_486_n N_A_27_74#_c_498_n N_A_27_74#_c_505_n
+ N_A_27_74#_c_509_n N_A_27_74#_c_487_n N_A_27_74#_c_488_n N_A_27_74#_c_489_n
+ N_A_27_74#_c_490_n N_A_27_74#_c_491_n N_A_27_74#_c_549_n N_A_27_74#_c_492_n
+ N_A_27_74#_c_499_n N_A_27_74#_c_493_n N_A_27_74#_c_494_n N_A_27_74#_c_495_n
+ PM_SKY130_FD_SC_MS__DLCLKP_4%A_27_74#
x_PM_SKY130_FD_SC_MS__DLCLKP_4%CLK N_CLK_M1012_g N_CLK_M1019_g N_CLK_M1008_g
+ N_CLK_M1005_g CLK N_CLK_c_625_n N_CLK_c_626_n PM_SKY130_FD_SC_MS__DLCLKP_4%CLK
x_PM_SKY130_FD_SC_MS__DLCLKP_4%A_1047_368# N_A_1047_368#_M1021_d
+ N_A_1047_368#_M1008_d N_A_1047_368#_c_668_n N_A_1047_368#_M1004_g
+ N_A_1047_368#_M1006_g N_A_1047_368#_M1007_g N_A_1047_368#_M1009_g
+ N_A_1047_368#_c_671_n N_A_1047_368#_c_672_n N_A_1047_368#_M1010_g
+ N_A_1047_368#_M1013_g N_A_1047_368#_M1022_g N_A_1047_368#_M1016_g
+ N_A_1047_368#_c_675_n N_A_1047_368#_c_688_n N_A_1047_368#_c_689_n
+ N_A_1047_368#_c_690_n N_A_1047_368#_c_676_n N_A_1047_368#_c_677_n
+ N_A_1047_368#_c_678_n N_A_1047_368#_c_679_n
+ PM_SKY130_FD_SC_MS__DLCLKP_4%A_1047_368#
x_PM_SKY130_FD_SC_MS__DLCLKP_4%VPWR N_VPWR_M1003_d N_VPWR_M1002_d N_VPWR_M1012_d
+ N_VPWR_M1014_d N_VPWR_M1007_s N_VPWR_M1022_s N_VPWR_c_796_n N_VPWR_c_797_n
+ N_VPWR_c_798_n N_VPWR_c_799_n N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_802_n
+ N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_805_n N_VPWR_c_806_n VPWR
+ N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n
+ N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_795_n PM_SKY130_FD_SC_MS__DLCLKP_4%VPWR
x_PM_SKY130_FD_SC_MS__DLCLKP_4%GCLK N_GCLK_M1006_d N_GCLK_M1013_d N_GCLK_M1004_d
+ N_GCLK_M1010_d N_GCLK_c_908_n N_GCLK_c_901_n N_GCLK_c_909_n N_GCLK_c_929_n
+ N_GCLK_c_902_n N_GCLK_c_903_n N_GCLK_c_910_n N_GCLK_c_904_n N_GCLK_c_905_n
+ N_GCLK_c_906_n GCLK GCLK PM_SKY130_FD_SC_MS__DLCLKP_4%GCLK
x_PM_SKY130_FD_SC_MS__DLCLKP_4%VGND N_VGND_M1020_d N_VGND_M1001_d N_VGND_M1019_d
+ N_VGND_M1006_s N_VGND_M1009_s N_VGND_M1016_s N_VGND_c_976_n N_VGND_c_977_n
+ N_VGND_c_978_n N_VGND_c_979_n N_VGND_c_980_n N_VGND_c_981_n VGND
+ N_VGND_c_982_n N_VGND_c_983_n N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n
+ N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n N_VGND_c_991_n
+ N_VGND_c_992_n PM_SKY130_FD_SC_MS__DLCLKP_4%VGND
cc_1 VNB N_A_84_48#_c_150_n 0.0230635f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_84_48#_M1003_g 0.00704416f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.4
cc_3 VNB N_A_84_48#_c_152_n 0.00150907f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.97
cc_4 VNB N_A_84_48#_c_153_n 0.01229f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.275
cc_5 VNB N_A_84_48#_c_154_n 0.00256251f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_6 VNB N_A_84_48#_c_155_n 0.00621205f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.275
cc_7 VNB N_A_84_48#_c_156_n 0.0443355f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_8 VNB N_GATE_M1017_g 0.0348671f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_9 VNB GATE 0.00265138f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_GATE_c_244_n 0.0194668f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.4
cc_11 VNB N_A_334_54#_c_278_n 0.0179936f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_12 VNB N_A_334_54#_M1025_g 0.0241088f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_13 VNB N_A_334_54#_c_280_n 0.00525847f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=0.815
cc_14 VNB N_A_334_54#_c_281_n 0.0373992f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_15 VNB N_A_334_54#_c_282_n 0.00268632f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.275
cc_16 VNB N_A_334_54#_c_283_n 0.00716059f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_17 VNB N_A_334_54#_c_284_n 0.0618249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_334_54#_c_285_n 0.00537146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_334_54#_c_286_n 0.0330284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_334_338#_c_402_n 0.00433237f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.55
cc_21 VNB N_A_334_338#_M1011_g 0.0377623f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.55
cc_22 VNB N_A_334_338#_c_404_n 0.00766943f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.055
cc_23 VNB N_A_334_338#_c_405_n 0.00409063f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.98
cc_24 VNB N_A_334_338#_c_406_n 0.0223667f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=0.815
cc_25 VNB N_A_334_338#_c_407_n 0.0113424f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.275
cc_26 VNB N_A_334_338#_c_408_n 0.00929218f $X=-0.19 $Y=-0.245 $X2=0.707
+ $Y2=1.385
cc_27 VNB N_A_27_74#_c_481_n 0.00576023f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_28 VNB N_A_27_74#_M1002_g 0.0106067f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_29 VNB N_A_27_74#_M1001_g 0.0266169f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.55
cc_30 VNB N_A_27_74#_M1021_g 0.023672f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.275
cc_31 VNB N_A_27_74#_M1014_g 0.00171287f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_32 VNB N_A_27_74#_c_486_n 0.0207357f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_33 VNB N_A_27_74#_c_487_n 0.0309217f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_34 VNB N_A_27_74#_c_488_n 0.00233902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_489_n 0.00122215f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_36 VNB N_A_27_74#_c_490_n 0.00767704f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_37 VNB N_A_27_74#_c_491_n 0.0354209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_492_n 0.00704942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_493_n 0.0312479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_494_n 0.0460418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_495_n 0.02825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_CLK_M1019_g 0.0293985f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_43 VNB N_CLK_M1005_g 0.0222599f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.97
cc_44 VNB N_CLK_c_625_n 0.00487367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_CLK_c_626_n 0.0519309f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.685
cc_46 VNB N_A_1047_368#_c_668_n 0.0171186f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_47 VNB N_A_1047_368#_M1006_g 0.0265413f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.97
cc_48 VNB N_A_1047_368#_M1009_g 0.025436f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.52
cc_49 VNB N_A_1047_368#_c_671_n 0.0122982f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_50 VNB N_A_1047_368#_c_672_n 0.0201218f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_51 VNB N_A_1047_368#_M1013_g 0.0254487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1047_368#_M1016_g 0.036104f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_53 VNB N_A_1047_368#_c_675_n 0.0317946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1047_368#_c_676_n 0.0281117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1047_368#_c_677_n 0.00409086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1047_368#_c_678_n 0.0599216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1047_368#_c_679_n 0.01192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_795_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_GCLK_c_901_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_60 VNB N_GCLK_c_902_n 0.00766134f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_61 VNB N_GCLK_c_903_n 0.00158543f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_62 VNB N_GCLK_c_904_n 0.00316097f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_63 VNB N_GCLK_c_905_n 3.53034e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_64 VNB N_GCLK_c_906_n 0.00194448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB GCLK 0.00915128f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_66 VNB N_VGND_c_976_n 0.00727256f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_67 VNB N_VGND_c_977_n 0.00972604f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_68 VNB N_VGND_c_978_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.685
cc_69 VNB N_VGND_c_979_n 0.00807502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_980_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_71 VNB N_VGND_c_981_n 0.0353267f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.55
cc_72 VNB N_VGND_c_982_n 0.01755f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_73 VNB N_VGND_c_983_n 0.0565077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_984_n 0.0277574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_985_n 0.0549955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_986_n 0.0190448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_987_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_988_n 0.0070281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_989_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_990_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_991_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_992_n 0.467177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VPB N_A_84_48#_M1003_g 0.0296879f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_84 VPB N_A_84_48#_c_152_n 0.00329282f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.97
cc_85 VPB N_A_84_48#_c_159_n 0.00258331f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_86 VPB N_GATE_M1023_g 0.0246086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB GATE 0.00239443f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_88 VPB N_GATE_c_244_n 0.0131315f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_89 VPB N_A_334_54#_M1024_g 0.0250486f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_90 VPB N_A_334_54#_M1015_g 0.028097f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.275
cc_91 VPB N_A_334_54#_c_280_n 0.00486805f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=0.815
cc_92 VPB N_A_334_54#_c_290_n 0.0246311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_334_54#_c_291_n 0.0311256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_334_54#_c_282_n 0.00270934f $X=-0.19 $Y=1.66 $X2=0.707 $Y2=1.275
cc_95 VPB N_A_334_54#_c_293_n 0.019332f $X=-0.19 $Y=1.66 $X2=0.707 $Y2=1.385
cc_96 VPB N_A_334_54#_c_294_n 0.0136411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_334_54#_c_286_n 0.0099419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_334_338#_c_409_n 0.0224247f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_99 VPB N_A_334_338#_c_402_n 0.0278659f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.55
cc_100 VPB N_A_334_338#_c_411_n 0.00817298f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_101 VPB N_A_334_338#_c_404_n 0.00538878f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=2.055
cc_102 VPB N_A_334_338#_c_406_n 0.0127529f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=0.815
cc_103 VPB N_A_334_338#_c_414_n 0.00202688f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_104 VPB N_A_27_74#_M1002_g 0.0663643f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_105 VPB N_A_27_74#_M1014_g 0.0251205f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.19
cc_106 VPB N_A_27_74#_c_498_n 0.04385f $X=-0.19 $Y=1.66 $X2=0.707 $Y2=1.275
cc_107 VPB N_A_27_74#_c_499_n 0.0124642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_74#_c_493_n 0.00819868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_CLK_M1012_g 0.0447498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_CLK_M1008_g 0.0225005f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_111 VPB N_CLK_c_625_n 0.00619808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_CLK_c_626_n 0.00831757f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_113 VPB N_A_1047_368#_c_668_n 0.00997041f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_114 VPB N_A_1047_368#_M1004_g 0.022724f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_115 VPB N_A_1047_368#_M1007_g 0.0210234f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=2.055
cc_116 VPB N_A_1047_368#_c_671_n 0.00421806f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_117 VPB N_A_1047_368#_c_672_n 0.00436988f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_118 VPB N_A_1047_368#_M1010_g 0.0208406f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_119 VPB N_A_1047_368#_M1022_g 0.0253255f $X=-0.19 $Y=1.66 $X2=0.707 $Y2=1.55
cc_120 VPB N_A_1047_368#_c_675_n 0.00448104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_1047_368#_c_688_n 0.00312943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_1047_368#_c_689_n 0.00275612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_1047_368#_c_690_n 0.00652416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_1047_368#_c_677_n 0.00307504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_1047_368#_c_679_n 0.0103718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_796_n 0.0104796f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.19
cc_127 VPB N_VPWR_c_797_n 0.00772962f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_128 VPB N_VPWR_c_798_n 0.00663805f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_129 VPB N_VPWR_c_799_n 0.014133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_800_n 0.00749022f $X=-0.19 $Y=1.66 $X2=0.707 $Y2=1.55
cc_131 VPB N_VPWR_c_801_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.385
cc_132 VPB N_VPWR_c_802_n 0.0481756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_803_n 0.0238191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_804_n 0.00718714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_805_n 0.0354159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_806_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_807_n 0.0556468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_808_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_809_n 0.0186436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_810_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_811_n 0.00631473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_812_n 0.0169969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_813_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_795_n 0.102501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_GCLK_c_908_n 0.0024448f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.97
cc_146 VPB N_GCLK_c_909_n 0.00423197f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.52
cc_147 VPB N_GCLK_c_910_n 0.00257518f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_148 VPB GCLK 8.14549e-19 $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_149 VPB GCLK 0.00903753f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.385
cc_150 N_A_84_48#_M1003_g N_GATE_M1023_g 0.019037f $X=0.6 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_84_48#_c_152_n N_GATE_M1023_g 0.0031117f $X=0.795 $Y=1.97 $X2=0 $Y2=0
cc_152 N_A_84_48#_c_162_p N_GATE_M1023_g 0.017501f $X=1.435 $Y=2.055 $X2=0 $Y2=0
cc_153 N_A_84_48#_c_150_n N_GATE_M1017_g 0.00900631f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_154 N_A_84_48#_c_153_n N_GATE_M1017_g 0.0148109f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_155 N_A_84_48#_c_154_n N_GATE_M1017_g 0.00393105f $X=1.52 $Y=1.19 $X2=0 $Y2=0
cc_156 N_A_84_48#_c_155_n N_GATE_M1017_g 0.00224326f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_157 N_A_84_48#_c_156_n N_GATE_M1017_g 0.00628804f $X=0.695 $Y=1.385 $X2=0
+ $Y2=0
cc_158 N_A_84_48#_c_153_n GATE 0.0250347f $X=1.435 $Y=1.275 $X2=0 $Y2=0
cc_159 N_A_84_48#_c_162_p GATE 0.0226356f $X=1.435 $Y=2.055 $X2=0 $Y2=0
cc_160 N_A_84_48#_c_155_n GATE 0.0188052f $X=0.707 $Y=1.275 $X2=0 $Y2=0
cc_161 N_A_84_48#_M1003_g N_GATE_c_244_n 0.00587708f $X=0.6 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_84_48#_c_153_n N_GATE_c_244_n 0.00445796f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_163 N_A_84_48#_c_162_p N_GATE_c_244_n 0.00323803f $X=1.435 $Y=2.055 $X2=0
+ $Y2=0
cc_164 N_A_84_48#_c_155_n N_GATE_c_244_n 0.00229548f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_165 N_A_84_48#_c_156_n N_GATE_c_244_n 0.00429519f $X=0.695 $Y=1.385 $X2=0
+ $Y2=0
cc_166 N_A_84_48#_c_154_n N_A_334_54#_c_278_n 0.00417838f $X=1.52 $Y=1.19 $X2=0
+ $Y2=0
cc_167 N_A_84_48#_c_177_p N_A_334_54#_c_278_n 0.0208157f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_168 N_A_84_48#_c_159_n N_A_334_54#_M1024_g 0.0139011f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_169 N_A_84_48#_M1000_d N_A_334_54#_c_280_n 0.00367686f $X=1.85 $Y=1.96 $X2=0
+ $Y2=0
cc_170 N_A_84_48#_c_153_n N_A_334_54#_c_280_n 0.0142091f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_171 N_A_84_48#_c_162_p N_A_334_54#_c_280_n 0.00651026f $X=1.435 $Y=2.055
+ $X2=0 $Y2=0
cc_172 N_A_84_48#_c_154_n N_A_334_54#_c_280_n 0.00293885f $X=1.52 $Y=1.19 $X2=0
+ $Y2=0
cc_173 N_A_84_48#_c_177_p N_A_334_54#_c_280_n 0.021323f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_174 N_A_84_48#_c_153_n N_A_334_54#_c_281_n 0.00140598f $X=1.435 $Y=1.275
+ $X2=0 $Y2=0
cc_175 N_A_84_48#_c_177_p N_A_334_54#_c_281_n 0.00166298f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_176 N_A_84_48#_M1000_d N_A_334_54#_c_290_n 0.00136409f $X=1.85 $Y=1.96 $X2=0
+ $Y2=0
cc_177 N_A_84_48#_c_159_n N_A_334_54#_c_290_n 0.03372f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_178 N_A_84_48#_M1000_d N_A_334_54#_c_308_n 0.00232285f $X=1.85 $Y=1.96 $X2=0
+ $Y2=0
cc_179 N_A_84_48#_c_162_p N_A_334_54#_c_308_n 0.00786627f $X=1.435 $Y=2.055
+ $X2=0 $Y2=0
cc_180 N_A_84_48#_c_190_p N_A_334_54#_c_308_n 0.0164691f $X=1.52 $Y=2.52 $X2=0
+ $Y2=0
cc_181 N_A_84_48#_c_159_n N_A_334_54#_c_308_n 0.0193557f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_182 N_A_84_48#_c_159_n N_A_334_54#_c_291_n 0.00354136f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_183 N_A_84_48#_c_162_p N_A_334_338#_c_409_n 0.00127882f $X=1.435 $Y=2.055
+ $X2=0 $Y2=0
cc_184 N_A_84_48#_c_190_p N_A_334_338#_c_409_n 0.00527479f $X=1.52 $Y=2.52 $X2=0
+ $Y2=0
cc_185 N_A_84_48#_c_159_n N_A_334_338#_c_409_n 0.0235437f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_186 N_A_84_48#_c_159_n N_A_334_338#_c_402_n 7.89305e-19 $X=2.15 $Y=2.685
+ $X2=0 $Y2=0
cc_187 N_A_84_48#_c_177_p N_A_334_338#_M1011_g 0.0121963f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_188 N_A_84_48#_c_177_p N_A_334_338#_c_405_n 9.67748e-19 $X=2.06 $Y=0.815
+ $X2=0 $Y2=0
cc_189 N_A_84_48#_c_159_n N_A_27_74#_M1002_g 0.00156106f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_190 N_A_84_48#_c_177_p N_A_27_74#_M1001_g 3.05797e-19 $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_191 N_A_84_48#_c_150_n N_A_27_74#_c_486_n 0.00159473f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_192 N_A_84_48#_M1003_g N_A_27_74#_c_498_n 0.0199149f $X=0.6 $Y=2.4 $X2=0
+ $Y2=0
cc_193 N_A_84_48#_c_150_n N_A_27_74#_c_505_n 0.0144795f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_194 N_A_84_48#_c_153_n N_A_27_74#_c_505_n 0.0280388f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_195 N_A_84_48#_c_155_n N_A_27_74#_c_505_n 0.0254697f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_196 N_A_84_48#_c_156_n N_A_27_74#_c_505_n 0.0017501f $X=0.695 $Y=1.385 $X2=0
+ $Y2=0
cc_197 N_A_84_48#_c_150_n N_A_27_74#_c_509_n 0.00257528f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_198 N_A_84_48#_M1018_d N_A_27_74#_c_487_n 0.00241797f $X=1.82 $Y=0.4 $X2=0
+ $Y2=0
cc_199 N_A_84_48#_c_209_p N_A_27_74#_c_487_n 0.00707909f $X=1.605 $Y=0.815 $X2=0
+ $Y2=0
cc_200 N_A_84_48#_c_177_p N_A_27_74#_c_487_n 0.0325781f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_201 N_A_84_48#_c_150_n N_A_27_74#_c_488_n 3.78932e-19 $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_202 N_A_84_48#_c_177_p N_A_27_74#_c_490_n 0.012421f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_203 N_A_84_48#_M1003_g N_A_27_74#_c_499_n 0.00440232f $X=0.6 $Y=2.4 $X2=0
+ $Y2=0
cc_204 N_A_84_48#_c_152_n N_A_27_74#_c_499_n 0.00656531f $X=0.795 $Y=1.97 $X2=0
+ $Y2=0
cc_205 N_A_84_48#_c_156_n N_A_27_74#_c_499_n 0.00391223f $X=0.695 $Y=1.385 $X2=0
+ $Y2=0
cc_206 N_A_84_48#_c_150_n N_A_27_74#_c_493_n 0.0129583f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_207 N_A_84_48#_M1003_g N_A_27_74#_c_493_n 0.00614644f $X=0.6 $Y=2.4 $X2=0
+ $Y2=0
cc_208 N_A_84_48#_c_152_n N_A_27_74#_c_493_n 0.0127446f $X=0.795 $Y=1.97 $X2=0
+ $Y2=0
cc_209 N_A_84_48#_c_155_n N_A_27_74#_c_493_n 0.027924f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_210 N_A_84_48#_c_152_n N_VPWR_M1003_d 0.00270963f $X=0.795 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_211 N_A_84_48#_c_162_p N_VPWR_M1003_d 0.0107381f $X=1.435 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A_84_48#_c_222_p N_VPWR_M1003_d 0.00403994f $X=0.88 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_84_48#_M1003_g N_VPWR_c_796_n 0.0109471f $X=0.6 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_84_48#_c_162_p N_VPWR_c_796_n 0.0226626f $X=1.435 $Y=2.055 $X2=0
+ $Y2=0
cc_215 N_A_84_48#_c_222_p N_VPWR_c_796_n 0.00843013f $X=0.88 $Y=2.055 $X2=0
+ $Y2=0
cc_216 N_A_84_48#_M1003_g N_VPWR_c_803_n 0.005209f $X=0.6 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A_84_48#_c_227_p N_VPWR_c_807_n 0.00409999f $X=1.605 $Y=2.685 $X2=0
+ $Y2=0
cc_218 N_A_84_48#_c_159_n N_VPWR_c_807_n 0.0211957f $X=2.15 $Y=2.685 $X2=0 $Y2=0
cc_219 N_A_84_48#_M1003_g N_VPWR_c_795_n 0.00989564f $X=0.6 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_84_48#_c_227_p N_VPWR_c_795_n 0.00576021f $X=1.605 $Y=2.685 $X2=0
+ $Y2=0
cc_221 N_A_84_48#_c_159_n N_VPWR_c_795_n 0.0279392f $X=2.15 $Y=2.685 $X2=0 $Y2=0
cc_222 N_A_84_48#_c_162_p A_286_392# 0.00365807f $X=1.435 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_84_48#_c_190_p A_286_392# 0.00372192f $X=1.52 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_224 N_A_84_48#_c_227_p A_286_392# 0.00180109f $X=1.605 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A_84_48#_c_159_n A_286_392# 3.90667e-19 $X=2.15 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_84_48#_c_150_n N_VGND_c_976_n 0.0112574f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_227 N_A_84_48#_c_150_n N_VGND_c_982_n 0.00398535f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_228 N_A_84_48#_c_150_n N_VGND_c_992_n 0.00404969f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_229 N_A_84_48#_c_154_n A_286_80# 6.49906e-19 $X=1.52 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_230 N_A_84_48#_c_209_p A_286_80# 0.00147622f $X=1.605 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_84_48#_c_177_p A_286_80# 3.7187e-19 $X=2.06 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_232 N_GATE_M1017_g N_A_334_54#_c_278_n 0.0308885f $X=1.355 $Y=0.72 $X2=0
+ $Y2=0
cc_233 N_GATE_M1017_g N_A_334_54#_c_280_n 7.74843e-19 $X=1.355 $Y=0.72 $X2=0
+ $Y2=0
cc_234 GATE N_A_334_54#_c_280_n 0.0120209f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_235 N_GATE_c_244_n N_A_334_54#_c_280_n 0.00372683f $X=1.265 $Y=1.635 $X2=0
+ $Y2=0
cc_236 N_GATE_c_244_n N_A_334_54#_c_281_n 0.0308885f $X=1.265 $Y=1.635 $X2=0
+ $Y2=0
cc_237 N_GATE_M1023_g N_A_334_338#_c_409_n 0.0355123f $X=1.34 $Y=2.46 $X2=0
+ $Y2=0
cc_238 GATE N_A_334_338#_c_411_n 4.93257e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_239 N_GATE_c_244_n N_A_334_338#_c_411_n 0.0355123f $X=1.265 $Y=1.635 $X2=0
+ $Y2=0
cc_240 N_GATE_M1017_g N_A_27_74#_c_487_n 0.0147887f $X=1.355 $Y=0.72 $X2=0 $Y2=0
cc_241 N_GATE_M1023_g N_VPWR_c_796_n 0.0136797f $X=1.34 $Y=2.46 $X2=0 $Y2=0
cc_242 N_GATE_M1023_g N_VPWR_c_807_n 0.00553757f $X=1.34 $Y=2.46 $X2=0 $Y2=0
cc_243 N_GATE_M1023_g N_VPWR_c_795_n 0.0109163f $X=1.34 $Y=2.46 $X2=0 $Y2=0
cc_244 N_GATE_M1017_g N_VGND_c_976_n 9.39772e-19 $X=1.355 $Y=0.72 $X2=0 $Y2=0
cc_245 N_GATE_M1017_g N_VGND_c_983_n 9.29978e-19 $X=1.355 $Y=0.72 $X2=0 $Y2=0
cc_246 N_A_334_54#_c_293_n N_A_334_338#_M1015_d 0.00717307f $X=4.205 $Y=2.605
+ $X2=0 $Y2=0
cc_247 N_A_334_54#_M1024_g N_A_334_338#_c_409_n 0.0141534f $X=2.545 $Y=2.75
+ $X2=0 $Y2=0
cc_248 N_A_334_54#_c_280_n N_A_334_338#_c_409_n 0.00782653f $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_249 N_A_334_54#_c_308_n N_A_334_338#_c_409_n 0.0103724f $X=2.065 $Y=2.2 $X2=0
+ $Y2=0
cc_250 N_A_334_54#_c_291_n N_A_334_338#_c_409_n 0.00787863f $X=2.47 $Y=2.215
+ $X2=0 $Y2=0
cc_251 N_A_334_54#_c_280_n N_A_334_338#_c_402_n 0.0132375f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_252 N_A_334_54#_c_290_n N_A_334_338#_c_402_n 0.00839201f $X=3.305 $Y=2.2
+ $X2=0 $Y2=0
cc_253 N_A_334_54#_c_280_n N_A_334_338#_c_411_n 0.00355197f $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_254 N_A_334_54#_c_281_n N_A_334_338#_c_411_n 0.0275626f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_255 N_A_334_54#_c_278_n N_A_334_338#_M1011_g 0.016863f $X=1.745 $Y=1.15 $X2=0
+ $Y2=0
cc_256 N_A_334_54#_c_280_n N_A_334_338#_M1011_g 0.00174539f $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_257 N_A_334_54#_c_281_n N_A_334_338#_M1011_g 0.0178648f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_258 N_A_334_54#_M1015_g N_A_334_338#_c_404_n 0.0038186f $X=3.585 $Y=2.54
+ $X2=0 $Y2=0
cc_259 N_A_334_54#_M1025_g N_A_334_338#_c_404_n 0.0100418f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_260 N_A_334_54#_c_282_n N_A_334_338#_c_404_n 0.0286547f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_261 N_A_334_54#_c_294_n N_A_334_338#_c_404_n 0.00615349f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_262 N_A_334_54#_c_280_n N_A_334_338#_c_405_n 0.0259472f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_263 N_A_334_54#_c_281_n N_A_334_338#_c_405_n 4.56399e-19 $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_264 N_A_334_54#_c_290_n N_A_334_338#_c_405_n 0.018746f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_265 N_A_334_54#_c_291_n N_A_334_338#_c_405_n 0.00117723f $X=2.47 $Y=2.215
+ $X2=0 $Y2=0
cc_266 N_A_334_54#_c_282_n N_A_334_338#_c_405_n 0.0029232f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_267 N_A_334_54#_c_280_n N_A_334_338#_c_406_n 0.0045632f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_268 N_A_334_54#_c_290_n N_A_334_338#_c_406_n 0.00128281f $X=3.305 $Y=2.2
+ $X2=0 $Y2=0
cc_269 N_A_334_54#_c_291_n N_A_334_338#_c_406_n 0.0215977f $X=2.47 $Y=2.215
+ $X2=0 $Y2=0
cc_270 N_A_334_54#_M1015_g N_A_334_338#_c_414_n 0.00300921f $X=3.585 $Y=2.54
+ $X2=0 $Y2=0
cc_271 N_A_334_54#_c_282_n N_A_334_338#_c_414_n 5.72571e-19 $X=3.39 $Y=2.35
+ $X2=0 $Y2=0
cc_272 N_A_334_54#_c_293_n N_A_334_338#_c_414_n 0.0211711f $X=4.205 $Y=2.605
+ $X2=0 $Y2=0
cc_273 N_A_334_54#_c_294_n N_A_334_338#_c_414_n 0.0121633f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_274 N_A_334_54#_c_286_n N_A_334_338#_c_414_n 0.00241703f $X=3.695 $Y=1.795
+ $X2=0 $Y2=0
cc_275 N_A_334_54#_M1025_g N_A_334_338#_c_407_n 0.0138783f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_276 N_A_334_54#_c_290_n N_A_334_338#_c_407_n 0.0228749f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_277 N_A_334_54#_c_282_n N_A_334_338#_c_407_n 0.0268965f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_278 N_A_334_54#_c_286_n N_A_334_338#_c_407_n 0.00771188f $X=3.695 $Y=1.795
+ $X2=0 $Y2=0
cc_279 N_A_334_54#_M1025_g N_A_334_338#_c_408_n 0.002462f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_280 N_A_334_54#_M1015_g N_A_27_74#_M1002_g 0.0250706f $X=3.585 $Y=2.54 $X2=0
+ $Y2=0
cc_281 N_A_334_54#_c_290_n N_A_27_74#_M1002_g 0.0258066f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_282 N_A_334_54#_c_291_n N_A_27_74#_M1002_g 0.0576075f $X=2.47 $Y=2.215 $X2=0
+ $Y2=0
cc_283 N_A_334_54#_c_282_n N_A_27_74#_M1002_g 0.00627566f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_284 N_A_334_54#_c_356_p N_A_27_74#_M1002_g 0.00342789f $X=3.39 $Y=2.52 $X2=0
+ $Y2=0
cc_285 N_A_334_54#_c_357_p N_A_27_74#_M1002_g 0.00453023f $X=3.475 $Y=2.605
+ $X2=0 $Y2=0
cc_286 N_A_334_54#_c_286_n N_A_27_74#_M1002_g 0.0152868f $X=3.695 $Y=1.795 $X2=0
+ $Y2=0
cc_287 N_A_334_54#_M1025_g N_A_27_74#_M1001_g 0.0171519f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_334_54#_c_278_n N_A_27_74#_c_487_n 0.0119481f $X=1.745 $Y=1.15 $X2=0
+ $Y2=0
cc_289 N_A_334_54#_M1025_g N_A_27_74#_c_490_n 0.00318939f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_290 N_A_334_54#_M1019_s N_A_27_74#_c_491_n 0.00239646f $X=4.3 $Y=0.37 $X2=0
+ $Y2=0
cc_291 N_A_334_54#_M1025_g N_A_27_74#_c_491_n 0.0175247f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_334_54#_c_283_n N_A_27_74#_c_491_n 0.0151779f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_293 N_A_334_54#_c_284_n N_A_27_74#_c_491_n 0.00634638f $X=3.98 $Y=0.35 $X2=0
+ $Y2=0
cc_294 N_A_334_54#_c_285_n N_A_27_74#_c_491_n 0.0258904f $X=4.445 $Y=0.685 $X2=0
+ $Y2=0
cc_295 N_A_334_54#_c_284_n N_A_27_74#_c_494_n 0.00690617f $X=3.98 $Y=0.35 $X2=0
+ $Y2=0
cc_296 N_A_334_54#_c_293_n N_CLK_M1012_g 0.00837497f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_297 N_A_334_54#_c_294_n N_CLK_M1012_g 0.00758617f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_298 N_A_334_54#_c_283_n N_CLK_M1019_g 0.0023f $X=4.28 $Y=0.385 $X2=0 $Y2=0
cc_299 N_A_334_54#_c_284_n N_CLK_M1019_g 0.00464769f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_300 N_A_334_54#_c_294_n N_CLK_c_625_n 0.00767395f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_301 N_A_334_54#_M1025_g N_CLK_c_626_n 0.00408582f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_334_54#_c_294_n N_CLK_c_626_n 6.37339e-19 $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_303 N_A_334_54#_c_290_n N_VPWR_M1002_d 0.00177961f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_304 N_A_334_54#_c_282_n N_VPWR_M1002_d 0.00148466f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_305 N_A_334_54#_c_356_p N_VPWR_M1002_d 0.00215336f $X=3.39 $Y=2.52 $X2=0
+ $Y2=0
cc_306 N_A_334_54#_c_357_p N_VPWR_M1002_d 0.00398396f $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_307 N_A_334_54#_M1015_g N_VPWR_c_797_n 0.00440778f $X=3.585 $Y=2.54 $X2=0
+ $Y2=0
cc_308 N_A_334_54#_c_290_n N_VPWR_c_797_n 0.00732173f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_309 N_A_334_54#_c_357_p N_VPWR_c_797_n 0.0112162f $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_310 N_A_334_54#_c_293_n N_VPWR_c_798_n 0.0159435f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_311 N_A_334_54#_c_294_n N_VPWR_c_798_n 0.0145507f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_312 N_A_334_54#_M1015_g N_VPWR_c_805_n 0.00392086f $X=3.585 $Y=2.54 $X2=0
+ $Y2=0
cc_313 N_A_334_54#_c_293_n N_VPWR_c_805_n 0.0260715f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_314 N_A_334_54#_M1024_g N_VPWR_c_807_n 0.00523141f $X=2.545 $Y=2.75 $X2=0
+ $Y2=0
cc_315 N_A_334_54#_M1024_g N_VPWR_c_795_n 0.00986058f $X=2.545 $Y=2.75 $X2=0
+ $Y2=0
cc_316 N_A_334_54#_M1015_g N_VPWR_c_795_n 0.00502116f $X=3.585 $Y=2.54 $X2=0
+ $Y2=0
cc_317 N_A_334_54#_c_293_n N_VPWR_c_795_n 0.0319548f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_318 N_A_334_54#_c_357_p N_VPWR_c_795_n 0.00178054f $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_319 N_A_334_54#_M1025_g N_VGND_c_977_n 0.00921355f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_320 N_A_334_54#_c_283_n N_VGND_c_977_n 0.0205948f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_321 N_A_334_54#_c_284_n N_VGND_c_977_n 0.0115834f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_322 N_A_334_54#_c_285_n N_VGND_c_977_n 0.00972897f $X=4.445 $Y=0.685 $X2=0
+ $Y2=0
cc_323 N_A_334_54#_c_283_n N_VGND_c_978_n 0.0151168f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_324 N_A_334_54#_c_284_n N_VGND_c_978_n 9.77729e-19 $X=3.98 $Y=0.35 $X2=0
+ $Y2=0
cc_325 N_A_334_54#_c_278_n N_VGND_c_983_n 9.29978e-19 $X=1.745 $Y=1.15 $X2=0
+ $Y2=0
cc_326 N_A_334_54#_c_283_n N_VGND_c_984_n 0.0532296f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_327 N_A_334_54#_c_284_n N_VGND_c_984_n 0.0118937f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_328 N_A_334_54#_c_283_n N_VGND_c_992_n 0.0289216f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_329 N_A_334_54#_c_284_n N_VGND_c_992_n 0.0190295f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_330 N_A_334_338#_M1011_g N_A_27_74#_c_481_n 8.86417e-19 $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_331 N_A_334_338#_c_405_n N_A_27_74#_c_481_n 0.00163581f $X=2.47 $Y=1.445
+ $X2=0 $Y2=0
cc_332 N_A_334_338#_c_406_n N_A_27_74#_c_481_n 0.0209296f $X=2.47 $Y=1.64 $X2=0
+ $Y2=0
cc_333 N_A_334_338#_c_407_n N_A_27_74#_c_481_n 0.00918689f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_334 N_A_334_338#_M1011_g N_A_27_74#_M1001_g 0.0213372f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_335 N_A_334_338#_c_407_n N_A_27_74#_M1001_g 0.00564586f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_336 N_A_334_338#_M1011_g N_A_27_74#_c_487_n 0.00658236f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_337 N_A_334_338#_M1011_g N_A_27_74#_c_490_n 0.00591925f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_338 N_A_334_338#_M1025_d N_A_27_74#_c_491_n 0.0056672f $X=3.77 $Y=0.625 $X2=0
+ $Y2=0
cc_339 N_A_334_338#_c_407_n N_A_27_74#_c_491_n 0.0652325f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_340 N_A_334_338#_M1011_g N_A_27_74#_c_549_n 0.00396757f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_341 N_A_334_338#_c_407_n N_A_27_74#_c_549_n 0.0167062f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_342 N_A_334_338#_M1011_g N_A_27_74#_c_494_n 0.00202272f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_343 N_A_334_338#_c_404_n N_CLK_M1012_g 0.00826661f $X=3.91 $Y=2.18 $X2=0
+ $Y2=0
cc_344 N_A_334_338#_c_404_n N_CLK_c_625_n 0.00747805f $X=3.91 $Y=2.18 $X2=0
+ $Y2=0
cc_345 N_A_334_338#_c_408_n N_CLK_c_625_n 0.0164788f $X=3.99 $Y=1.445 $X2=0
+ $Y2=0
cc_346 N_A_334_338#_c_404_n N_CLK_c_626_n 2.7829e-19 $X=3.91 $Y=2.18 $X2=0 $Y2=0
cc_347 N_A_334_338#_c_408_n N_CLK_c_626_n 0.00121403f $X=3.99 $Y=1.445 $X2=0
+ $Y2=0
cc_348 N_A_334_338#_c_409_n N_VPWR_c_807_n 0.00370063f $X=1.76 $Y=1.84 $X2=0
+ $Y2=0
cc_349 N_A_334_338#_c_409_n N_VPWR_c_795_n 0.00455969f $X=1.76 $Y=1.84 $X2=0
+ $Y2=0
cc_350 N_A_334_338#_c_407_n N_VGND_M1001_d 0.00483981f $X=3.825 $Y=1.485 $X2=0
+ $Y2=0
cc_351 N_A_334_338#_c_405_n A_491_124# 0.00338728f $X=2.47 $Y=1.445 $X2=-0.19
+ $Y2=-0.245
cc_352 N_A_334_338#_c_407_n A_491_124# 0.00720817f $X=3.825 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_27_74#_c_491_n N_CLK_M1019_g 0.0163338f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_354 N_A_27_74#_M1021_g N_CLK_M1005_g 0.0350457f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_491_n N_CLK_M1005_g 0.0253727f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_356 N_A_27_74#_M1014_g N_CLK_c_625_n 6.72627e-19 $X=5.63 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_491_n N_CLK_c_625_n 0.0723728f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_358 N_A_27_74#_M1014_g N_CLK_c_626_n 0.0162011f $X=5.63 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_491_n N_CLK_c_626_n 0.00876998f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_495_n N_CLK_c_626_n 0.0350457f $X=5.64 $Y=1.465 $X2=0 $Y2=0
cc_361 N_A_27_74#_M1014_g N_A_1047_368#_c_688_n 0.00113429f $X=5.63 $Y=2.4 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_491_n N_A_1047_368#_c_688_n 0.0262166f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_363 N_A_27_74#_c_495_n N_A_1047_368#_c_688_n 5.01421e-19 $X=5.64 $Y=1.465
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_M1014_g N_A_1047_368#_c_689_n 0.0181361f $X=5.63 $Y=2.4 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_M1014_g N_A_1047_368#_c_690_n 0.0150412f $X=5.63 $Y=2.4 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_491_n N_A_1047_368#_c_690_n 0.0157153f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_367 N_A_27_74#_c_495_n N_A_1047_368#_c_690_n 5.84989e-19 $X=5.64 $Y=1.465
+ $X2=0 $Y2=0
cc_368 N_A_27_74#_M1021_g N_A_1047_368#_c_676_n 0.0148811f $X=5.55 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_491_n N_A_1047_368#_c_676_n 0.0228054f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_370 N_A_27_74#_c_495_n N_A_1047_368#_c_676_n 0.00141568f $X=5.64 $Y=1.465
+ $X2=0 $Y2=0
cc_371 N_A_27_74#_M1021_g N_A_1047_368#_c_677_n 0.00143549f $X=5.55 $Y=0.74
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_M1014_g N_A_1047_368#_c_677_n 0.00599397f $X=5.63 $Y=2.4 $X2=0
+ $Y2=0
cc_373 N_A_27_74#_c_491_n N_A_1047_368#_c_677_n 0.0337495f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_374 N_A_27_74#_c_495_n N_A_1047_368#_c_677_n 0.00111362f $X=5.64 $Y=1.465
+ $X2=0 $Y2=0
cc_375 N_A_27_74#_M1021_g N_A_1047_368#_c_678_n 0.0121306f $X=5.55 $Y=0.74 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_491_n N_A_1047_368#_c_678_n 3.72912e-19 $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_377 N_A_27_74#_c_495_n N_A_1047_368#_c_678_n 0.0208223f $X=5.64 $Y=1.465
+ $X2=0 $Y2=0
cc_378 N_A_27_74#_M1014_g N_A_1047_368#_c_679_n 0.00190646f $X=5.63 $Y=2.4 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_c_498_n N_VPWR_c_796_n 0.0404605f $X=0.375 $Y=2.815 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_M1002_g N_VPWR_c_797_n 0.00440778f $X=2.965 $Y=2.75 $X2=0
+ $Y2=0
cc_381 N_A_27_74#_M1014_g N_VPWR_c_798_n 5.70732e-19 $X=5.63 $Y=2.4 $X2=0 $Y2=0
cc_382 N_A_27_74#_M1014_g N_VPWR_c_799_n 0.00761722f $X=5.63 $Y=2.4 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_498_n N_VPWR_c_803_n 0.018788f $X=0.375 $Y=2.815 $X2=0 $Y2=0
cc_384 N_A_27_74#_M1002_g N_VPWR_c_807_n 0.00553757f $X=2.965 $Y=2.75 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_M1014_g N_VPWR_c_808_n 0.005209f $X=5.63 $Y=2.4 $X2=0 $Y2=0
cc_386 N_A_27_74#_M1002_g N_VPWR_c_795_n 0.0109009f $X=2.965 $Y=2.75 $X2=0 $Y2=0
cc_387 N_A_27_74#_M1014_g N_VPWR_c_795_n 0.00987161f $X=5.63 $Y=2.4 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_498_n N_VPWR_c_795_n 0.0154829f $X=0.375 $Y=2.815 $X2=0
+ $Y2=0
cc_389 N_A_27_74#_c_505_n N_VGND_M1020_d 0.0166022f $X=1.095 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_390 N_A_27_74#_c_509_n N_VGND_M1020_d 0.00684638f $X=1.18 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_391 N_A_27_74#_c_488_n N_VGND_M1020_d 2.48347e-19 $X=1.265 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_392 N_A_27_74#_c_490_n N_VGND_M1001_d 0.00120802f $X=2.98 $Y=1.02 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_491_n N_VGND_M1001_d 0.015135f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_394 N_A_27_74#_c_549_n N_VGND_M1001_d 3.54991e-19 $X=3.145 $Y=1.105 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_491_n N_VGND_M1019_d 0.00176461f $X=5.26 $Y=1.105 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_486_n N_VGND_c_976_n 0.0125137f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_397 N_A_27_74#_c_505_n N_VGND_c_976_n 0.0250287f $X=1.095 $Y=0.935 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_509_n N_VGND_c_976_n 0.0196481f $X=1.18 $Y=0.85 $X2=0 $Y2=0
cc_399 N_A_27_74#_c_488_n N_VGND_c_976_n 0.0150932f $X=1.265 $Y=0.34 $X2=0 $Y2=0
cc_400 N_A_27_74#_M1001_g N_VGND_c_977_n 0.00104285f $X=2.98 $Y=1.155 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_489_n N_VGND_c_977_n 0.0142656f $X=2.98 $Y=0.425 $X2=0 $Y2=0
cc_402 N_A_27_74#_c_490_n N_VGND_c_977_n 0.0348535f $X=2.98 $Y=1.02 $X2=0 $Y2=0
cc_403 N_A_27_74#_c_491_n N_VGND_c_977_n 0.0219153f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_404 N_A_27_74#_c_494_n N_VGND_c_977_n 0.00260146f $X=2.98 $Y=0.38 $X2=0 $Y2=0
cc_405 N_A_27_74#_M1021_g N_VGND_c_978_n 0.00197566f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_27_74#_c_491_n N_VGND_c_978_n 0.0170777f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_407 N_A_27_74#_c_486_n N_VGND_c_982_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_408 N_A_27_74#_c_487_n N_VGND_c_983_n 0.0997901f $X=2.815 $Y=0.34 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_488_n N_VGND_c_983_n 0.0121867f $X=1.265 $Y=0.34 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_489_n N_VGND_c_983_n 0.0224969f $X=2.98 $Y=0.425 $X2=0 $Y2=0
cc_411 N_A_27_74#_c_494_n N_VGND_c_983_n 0.00612073f $X=2.98 $Y=0.38 $X2=0 $Y2=0
cc_412 N_A_27_74#_M1021_g N_VGND_c_985_n 0.00748462f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_413 N_A_27_74#_M1021_g N_VGND_c_992_n 0.0082231f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_414 N_A_27_74#_c_486_n N_VGND_c_992_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_415 N_A_27_74#_c_505_n N_VGND_c_992_n 0.0124076f $X=1.095 $Y=0.935 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_487_n N_VGND_c_992_n 0.0582686f $X=2.815 $Y=0.34 $X2=0 $Y2=0
cc_417 N_A_27_74#_c_488_n N_VGND_c_992_n 0.00660921f $X=1.265 $Y=0.34 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_489_n N_VGND_c_992_n 0.0113197f $X=2.98 $Y=0.425 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_494_n N_VGND_c_992_n 0.00853275f $X=2.98 $Y=0.38 $X2=0 $Y2=0
cc_420 N_A_27_74#_c_487_n A_286_80# 0.00150293f $X=2.815 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_421 N_A_27_74#_c_490_n A_491_124# 0.00107962f $X=2.98 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_422 N_A_27_74#_c_549_n A_491_124# 0.00308074f $X=3.145 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_423 N_A_27_74#_c_491_n A_1047_74# 0.0056254f $X=5.26 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_424 N_CLK_M1008_g N_A_1047_368#_c_688_n 6.55893e-19 $X=5.145 $Y=2.4 $X2=0
+ $Y2=0
cc_425 N_CLK_M1008_g N_A_1047_368#_c_689_n 4.35897e-19 $X=5.145 $Y=2.4 $X2=0
+ $Y2=0
cc_426 N_CLK_M1005_g N_A_1047_368#_c_676_n 0.00233225f $X=5.16 $Y=0.74 $X2=0
+ $Y2=0
cc_427 N_CLK_M1012_g N_VPWR_c_798_n 0.00819006f $X=4.595 $Y=2.53 $X2=0 $Y2=0
cc_428 N_CLK_M1008_g N_VPWR_c_798_n 0.0156325f $X=5.145 $Y=2.4 $X2=0 $Y2=0
cc_429 N_CLK_c_625_n N_VPWR_c_798_n 0.0170757f $X=4.905 $Y=1.515 $X2=0 $Y2=0
cc_430 N_CLK_c_626_n N_VPWR_c_798_n 0.00114703f $X=5.16 $Y=1.515 $X2=0 $Y2=0
cc_431 N_CLK_M1012_g N_VPWR_c_805_n 0.0065193f $X=4.595 $Y=2.53 $X2=0 $Y2=0
cc_432 N_CLK_M1008_g N_VPWR_c_808_n 0.0050621f $X=5.145 $Y=2.4 $X2=0 $Y2=0
cc_433 N_CLK_M1012_g N_VPWR_c_795_n 0.00651205f $X=4.595 $Y=2.53 $X2=0 $Y2=0
cc_434 N_CLK_M1008_g N_VPWR_c_795_n 0.00999308f $X=5.145 $Y=2.4 $X2=0 $Y2=0
cc_435 N_CLK_M1019_g N_VGND_c_978_n 0.0104121f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_436 N_CLK_M1005_g N_VGND_c_978_n 0.0140817f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_437 N_CLK_M1019_g N_VGND_c_984_n 0.00383152f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_438 N_CLK_M1005_g N_VGND_c_985_n 0.00383152f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_439 N_CLK_M1019_g N_VGND_c_992_n 0.00759393f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_440 N_CLK_M1005_g N_VGND_c_992_n 0.0075725f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_441 N_A_1047_368#_c_690_n N_VPWR_M1014_d 0.0115435f $X=5.975 $Y=1.905 $X2=0
+ $Y2=0
cc_442 N_A_1047_368#_c_689_n N_VPWR_c_798_n 0.0341854f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_443 N_A_1047_368#_M1004_g N_VPWR_c_799_n 0.00761722f $X=6.735 $Y=2.4 $X2=0
+ $Y2=0
cc_444 N_A_1047_368#_c_689_n N_VPWR_c_799_n 0.0316504f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_445 N_A_1047_368#_c_690_n N_VPWR_c_799_n 0.0498832f $X=5.975 $Y=1.905 $X2=0
+ $Y2=0
cc_446 N_A_1047_368#_c_679_n N_VPWR_c_799_n 0.00965925f $X=6.185 $Y=1.4 $X2=0
+ $Y2=0
cc_447 N_A_1047_368#_M1007_g N_VPWR_c_800_n 0.00190234f $X=7.2 $Y=2.4 $X2=0
+ $Y2=0
cc_448 N_A_1047_368#_c_671_n N_VPWR_c_800_n 8.91722e-19 $X=7.595 $Y=1.54 $X2=0
+ $Y2=0
cc_449 N_A_1047_368#_M1010_g N_VPWR_c_800_n 0.00172337f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_450 N_A_1047_368#_M1010_g N_VPWR_c_802_n 6.88684e-19 $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_451 N_A_1047_368#_M1022_g N_VPWR_c_802_n 0.017993f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_452 N_A_1047_368#_c_689_n N_VPWR_c_808_n 0.014549f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_453 N_A_1047_368#_M1004_g N_VPWR_c_809_n 0.005209f $X=6.735 $Y=2.4 $X2=0
+ $Y2=0
cc_454 N_A_1047_368#_M1007_g N_VPWR_c_809_n 0.00537895f $X=7.2 $Y=2.4 $X2=0
+ $Y2=0
cc_455 N_A_1047_368#_M1010_g N_VPWR_c_810_n 0.005209f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_456 N_A_1047_368#_M1022_g N_VPWR_c_810_n 0.00460063f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_457 N_A_1047_368#_M1004_g N_VPWR_c_795_n 0.00986878f $X=6.735 $Y=2.4 $X2=0
+ $Y2=0
cc_458 N_A_1047_368#_M1007_g N_VPWR_c_795_n 0.0103679f $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_459 N_A_1047_368#_M1010_g N_VPWR_c_795_n 0.00982612f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_460 N_A_1047_368#_M1022_g N_VPWR_c_795_n 0.00908554f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_461 N_A_1047_368#_c_689_n N_VPWR_c_795_n 0.0119743f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_462 N_A_1047_368#_M1004_g N_GCLK_c_908_n 0.0247138f $X=6.735 $Y=2.4 $X2=0
+ $Y2=0
cc_463 N_A_1047_368#_M1007_g N_GCLK_c_908_n 0.0167554f $X=7.2 $Y=2.4 $X2=0 $Y2=0
cc_464 N_A_1047_368#_M1010_g N_GCLK_c_908_n 6.92718e-19 $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_465 N_A_1047_368#_c_690_n N_GCLK_c_908_n 0.00670758f $X=5.975 $Y=1.905 $X2=0
+ $Y2=0
cc_466 N_A_1047_368#_c_677_n N_GCLK_c_908_n 0.00385961f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_467 N_A_1047_368#_M1006_g N_GCLK_c_901_n 0.0205429f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_468 N_A_1047_368#_M1009_g N_GCLK_c_901_n 0.0126177f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_469 N_A_1047_368#_M1013_g N_GCLK_c_901_n 6.13796e-19 $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_470 N_A_1047_368#_c_676_n N_GCLK_c_901_n 0.015596f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_471 N_A_1047_368#_c_677_n N_GCLK_c_901_n 0.00255045f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_472 N_A_1047_368#_c_678_n N_GCLK_c_901_n 7.55566e-19 $X=6.185 $Y=0.835 $X2=0
+ $Y2=0
cc_473 N_A_1047_368#_M1007_g N_GCLK_c_909_n 0.00832805f $X=7.2 $Y=2.4 $X2=0
+ $Y2=0
cc_474 N_A_1047_368#_c_671_n N_GCLK_c_909_n 0.00864502f $X=7.595 $Y=1.54 $X2=0
+ $Y2=0
cc_475 N_A_1047_368#_c_672_n N_GCLK_c_909_n 0.00392988f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_476 N_A_1047_368#_M1010_g N_GCLK_c_909_n 0.00761093f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_477 N_A_1047_368#_c_675_n N_GCLK_c_909_n 0.00357204f $X=8.135 $Y=1.54 $X2=0
+ $Y2=0
cc_478 N_A_1047_368#_M1004_g N_GCLK_c_929_n 0.00120554f $X=6.735 $Y=2.4 $X2=0
+ $Y2=0
cc_479 N_A_1047_368#_M1007_g N_GCLK_c_929_n 5.28008e-19 $X=7.2 $Y=2.4 $X2=0
+ $Y2=0
cc_480 N_A_1047_368#_c_672_n N_GCLK_c_929_n 0.0150556f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_481 N_A_1047_368#_c_677_n N_GCLK_c_929_n 0.00641561f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_482 N_A_1047_368#_M1009_g N_GCLK_c_902_n 0.0113124f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_483 N_A_1047_368#_c_671_n N_GCLK_c_902_n 0.00465995f $X=7.595 $Y=1.54 $X2=0
+ $Y2=0
cc_484 N_A_1047_368#_M1013_g N_GCLK_c_902_n 0.0113115f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_485 N_A_1047_368#_M1006_g N_GCLK_c_903_n 0.00524345f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_1047_368#_M1009_g N_GCLK_c_903_n 0.00272521f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_1047_368#_c_672_n N_GCLK_c_903_n 0.00287768f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_488 N_A_1047_368#_c_677_n N_GCLK_c_903_n 0.00581761f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_489 N_A_1047_368#_c_678_n N_GCLK_c_903_n 5.80746e-19 $X=6.185 $Y=0.835 $X2=0
+ $Y2=0
cc_490 N_A_1047_368#_M1007_g N_GCLK_c_910_n 5.81657e-19 $X=7.2 $Y=2.4 $X2=0
+ $Y2=0
cc_491 N_A_1047_368#_M1010_g N_GCLK_c_910_n 0.0166159f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_492 N_A_1047_368#_M1022_g N_GCLK_c_910_n 0.00187859f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_493 N_A_1047_368#_M1009_g N_GCLK_c_904_n 6.95109e-19 $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A_1047_368#_M1013_g N_GCLK_c_904_n 0.0122683f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A_1047_368#_M1016_g N_GCLK_c_904_n 0.00292368f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A_1047_368#_M1013_g N_GCLK_c_905_n 4.96773e-19 $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_497 N_A_1047_368#_M1016_g N_GCLK_c_905_n 4.72088e-19 $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A_1047_368#_c_675_n N_GCLK_c_905_n 0.0181007f $X=8.135 $Y=1.54 $X2=0
+ $Y2=0
cc_499 N_A_1047_368#_M1013_g N_GCLK_c_906_n 0.00223615f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_1047_368#_M1016_g N_GCLK_c_906_n 0.0053794f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_1047_368#_M1010_g GCLK 0.00247135f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_502 N_A_1047_368#_c_675_n GCLK 0.00622489f $X=8.135 $Y=1.54 $X2=0 $Y2=0
cc_503 N_A_1047_368#_M1022_g GCLK 0.0120697f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_504 N_A_1047_368#_c_675_n GCLK 0.014038f $X=8.135 $Y=1.54 $X2=0 $Y2=0
cc_505 N_A_1047_368#_c_676_n N_VGND_c_978_n 0.0163082f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_506 N_A_1047_368#_M1009_g N_VGND_c_979_n 0.00659576f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_1047_368#_M1013_g N_VGND_c_979_n 0.00170206f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A_1047_368#_M1013_g N_VGND_c_981_n 5.78878e-19 $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_509 N_A_1047_368#_M1016_g N_VGND_c_981_n 0.0128863f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_1047_368#_M1006_g N_VGND_c_985_n 0.00777188f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_1047_368#_c_676_n N_VGND_c_985_n 0.0480661f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_512 N_A_1047_368#_c_678_n N_VGND_c_985_n 0.00197975f $X=6.185 $Y=0.835 $X2=0
+ $Y2=0
cc_513 N_A_1047_368#_M1006_g N_VGND_c_986_n 0.00434272f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_514 N_A_1047_368#_M1009_g N_VGND_c_986_n 0.00434272f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_1047_368#_M1013_g N_VGND_c_987_n 0.00434272f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_516 N_A_1047_368#_M1016_g N_VGND_c_987_n 0.00383152f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_1047_368#_M1006_g N_VGND_c_992_n 0.00825283f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_518 N_A_1047_368#_M1009_g N_VGND_c_992_n 0.00820718f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_519 N_A_1047_368#_M1013_g N_VGND_c_992_n 0.00820942f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_520 N_A_1047_368#_M1016_g N_VGND_c_992_n 0.0075754f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_1047_368#_c_676_n N_VGND_c_992_n 0.0198939f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_799_n N_GCLK_c_908_n 0.0316504f $X=6.46 $Y=2.26 $X2=0 $Y2=0
cc_523 N_VPWR_c_800_n N_GCLK_c_908_n 0.0416573f $X=7.46 $Y=2.055 $X2=0 $Y2=0
cc_524 N_VPWR_c_809_n N_GCLK_c_908_n 0.0145071f $X=7.295 $Y=3.33 $X2=0 $Y2=0
cc_525 N_VPWR_c_795_n N_GCLK_c_908_n 0.0119067f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_800_n N_GCLK_c_909_n 0.0179486f $X=7.46 $Y=2.055 $X2=0 $Y2=0
cc_527 N_VPWR_c_800_n N_GCLK_c_910_n 0.0350907f $X=7.46 $Y=2.055 $X2=0 $Y2=0
cc_528 N_VPWR_c_802_n N_GCLK_c_910_n 0.0346097f $X=8.36 $Y=2.035 $X2=0 $Y2=0
cc_529 N_VPWR_c_810_n N_GCLK_c_910_n 0.0109793f $X=8.195 $Y=3.33 $X2=0 $Y2=0
cc_530 N_VPWR_c_795_n N_GCLK_c_910_n 0.00901959f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_531 N_VPWR_c_802_n GCLK 0.0241685f $X=8.36 $Y=2.035 $X2=0 $Y2=0
cc_532 N_GCLK_c_901_n N_VGND_c_979_n 0.0266484f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_533 N_GCLK_c_902_n N_VGND_c_979_n 0.0199684f $X=7.765 $Y=1.295 $X2=0 $Y2=0
cc_534 N_GCLK_c_904_n N_VGND_c_979_n 0.0244284f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_535 N_GCLK_c_904_n N_VGND_c_981_n 0.0254585f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_536 GCLK N_VGND_c_981_n 0.0109035f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_537 N_GCLK_c_901_n N_VGND_c_985_n 0.00618339f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_538 N_GCLK_c_901_n N_VGND_c_986_n 0.0144922f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_539 N_GCLK_c_904_n N_VGND_c_987_n 0.0109942f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_540 N_GCLK_c_901_n N_VGND_c_992_n 0.0118826f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_541 N_GCLK_c_904_n N_VGND_c_992_n 0.00904371f $X=7.93 $Y=0.515 $X2=0 $Y2=0

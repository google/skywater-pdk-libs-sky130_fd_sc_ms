* File: sky130_fd_sc_ms__a211oi_2.pex.spice
* Created: Fri Aug 28 16:57:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A211OI_2%A1 3 5 7 10 12 14 15 24
c47 12 0 2.33874e-19 $X=0.96 $Y=1.22
r48 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.945 $Y=1.385
+ $X2=0.96 $Y2=1.385
r49 22 23 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=0.53 $Y=1.385
+ $X2=0.945 $Y2=1.385
r50 21 22 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.53 $Y2=1.385
r51 18 21 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.325 $Y=1.385
+ $X2=0.495 $Y2=1.385
r52 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.325
+ $Y=1.385 $X2=0.325 $Y2=1.385
r53 15 19 2.92169 $w=3.53e-07 $l=9e-08 $layer=LI1_cond $X=0.302 $Y=1.295
+ $X2=0.302 $Y2=1.385
r54 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.22
+ $X2=0.96 $Y2=1.385
r55 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.96 $Y=1.22 $X2=0.96
+ $Y2=0.74
r56 8 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.55
+ $X2=0.945 $Y2=1.385
r57 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.945 $Y=1.55
+ $X2=0.945 $Y2=2.4
r58 5 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.22
+ $X2=0.53 $Y2=1.385
r59 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.53 $Y=1.22 $X2=0.53
+ $Y2=0.74
r60 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=1.385
r61 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%A2 3 7 11 15 17 18 19 30
r55 29 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.845 $Y=1.515
+ $X2=1.86 $Y2=1.515
r56 27 29 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.77 $Y=1.515
+ $X2=1.845 $Y2=1.515
r57 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=1.515 $X2=1.77 $Y2=1.515
r58 25 27 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.395 $Y=1.515
+ $X2=1.77 $Y2=1.515
r59 23 25 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.39 $Y=1.515
+ $X2=1.395 $Y2=1.515
r60 19 28 12.8415 $w=3.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=1.77 $Y2=1.605
r61 18 28 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.605 $X2=1.77
+ $Y2=1.605
r62 17 18 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=1.68 $Y2=1.605
r63 13 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=1.515
r64 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=0.74
r65 9 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.68
+ $X2=1.845 $Y2=1.515
r66 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.845 $Y=1.68
+ $X2=1.845 $Y2=2.4
r67 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=1.515
r68 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.39 $Y=1.35 $X2=1.39
+ $Y2=0.74
r69 1 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.68
+ $X2=1.395 $Y2=1.515
r70 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.395 $Y=1.68
+ $X2=1.395 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%B1 1 3 6 10 12 13 22
c46 22 0 1.71329e-19 $X=3.305 $Y=1.385
r47 20 22 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.26 $Y=1.385
+ $X2=3.305 $Y2=1.385
r48 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.385 $X2=3.26 $Y2=1.385
r49 18 20 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=2.855 $Y=1.385
+ $X2=3.26 $Y2=1.385
r50 16 18 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.84 $Y=1.385
+ $X2=2.855 $Y2=1.385
r51 13 21 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.26
+ $Y2=1.365
r52 12 21 4.3606 $w=3.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.26 $Y2=1.365
r53 8 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.55
+ $X2=3.305 $Y2=1.385
r54 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.305 $Y=1.55
+ $X2=3.305 $Y2=2.4
r55 4 18 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.55
+ $X2=2.855 $Y2=1.385
r56 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.855 $Y=1.55
+ $X2=2.855 $Y2=2.4
r57 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.22
+ $X2=2.84 $Y2=1.385
r58 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.84 $Y=1.22 $X2=2.84
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%C1 1 3 6 10 12 13 22
c33 13 0 1.71329e-19 $X=4.56 $Y=1.295
r34 20 22 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.13 $Y=1.385
+ $X2=4.205 $Y2=1.385
r35 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.385 $X2=4.13 $Y2=1.385
r36 18 20 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.755 $Y=1.385
+ $X2=4.13 $Y2=1.385
r37 16 18 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.71 $Y=1.385
+ $X2=3.755 $Y2=1.385
r38 13 21 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.365
+ $X2=4.13 $Y2=1.365
r39 12 21 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.365 $X2=4.13
+ $Y2=1.365
r40 8 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.205 $Y=1.55
+ $X2=4.205 $Y2=1.385
r41 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.205 $Y=1.55
+ $X2=4.205 $Y2=2.4
r42 4 18 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.55
+ $X2=3.755 $Y2=1.385
r43 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.755 $Y=1.55
+ $X2=3.755 $Y2=2.4
r44 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.22
+ $X2=3.71 $Y2=1.385
r45 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.71 $Y=1.22 $X2=3.71
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%VPWR 1 2 3 10 12 18 22 24 26 31 38 39 45 48
r60 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.07 $Y2=3.33
r65 36 38 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=4.56 $Y2=3.33
r66 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r67 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r70 32 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.07 $Y2=3.33
r72 31 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r74 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 27 42 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r77 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r79 26 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 24 39 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 24 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=3.33
r83 20 22 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=2.485
r84 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r85 16 18 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.375
r86 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.23 $Y=1.985
+ $X2=0.23 $Y2=2.815
r87 10 42 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r88 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.815
r89 3 22 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.485
r90 2 18 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=2.375
r91 1 15 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r92 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%A_117_368# 1 2 3 10 12 14 18 20 22 24 26 31
+ 32
r47 24 34 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=2.23
+ $X2=3.105 $Y2=2.145
r48 24 26 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.105 $Y=2.23
+ $X2=3.105 $Y2=2.57
r49 22 34 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.965 $Y=2.145
+ $X2=3.105 $Y2=2.145
r50 22 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.965 $Y=2.145
+ $X2=2.355 $Y2=2.145
r51 21 31 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.09
+ $X2=1.62 $Y2=2.09
r52 20 32 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.215 $Y=2.09
+ $X2=2.355 $Y2=2.09
r53 20 21 20.9909 $w=2.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.215 $Y=2.09
+ $X2=1.705 $Y2=2.09
r54 16 31 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.62 $Y=2.23 $X2=1.62
+ $Y2=2.09
r55 16 18 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.62 $Y=2.23
+ $X2=1.62 $Y2=2.44
r56 15 29 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.68 $Y2=1.97
r57 14 31 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.62 $Y2=2.09
r58 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=0.805 $Y2=2.035
r59 10 29 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.68 $Y=2.12 $X2=0.68
+ $Y2=1.97
r60 10 12 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.68 $Y=2.12
+ $X2=0.68 $Y2=2.4
r61 3 34 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.145
r62 3 26 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.57
r63 2 31 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=2.035
r64 2 18 300 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=2.44
r65 1 29 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
r66 1 12 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%A_497_368# 1 2 3 12 14 15 18 20 24 28
r37 24 27 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.47 $Y=1.985
+ $X2=4.47 $Y2=2.815
r38 22 27 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.47 $Y=2.905 $X2=4.47
+ $Y2=2.815
r39 21 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=2.99
+ $X2=3.53 $Y2=2.99
r40 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.345 $Y=2.99
+ $X2=4.47 $Y2=2.905
r41 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.345 $Y=2.99
+ $X2=3.615 $Y2=2.99
r42 16 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=2.905
+ $X2=3.53 $Y2=2.99
r43 16 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.53 $Y=2.905
+ $X2=3.53 $Y2=2.225
r44 14 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=2.99
+ $X2=3.53 $Y2=2.99
r45 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.445 $Y=2.99
+ $X2=2.795 $Y2=2.99
r46 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.63 $Y=2.905
+ $X2=2.795 $Y2=2.99
r47 10 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.63 $Y=2.905
+ $X2=2.63 $Y2=2.485
r48 3 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.295
+ $Y=1.84 $X2=4.43 $Y2=2.815
r49 3 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.295
+ $Y=1.84 $X2=4.43 $Y2=1.985
r50 2 18 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=1.84 $X2=3.53 $Y2=2.225
r51 1 12 300 $w=1.7e-07 $l=7.13828e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.84 $X2=2.63 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%Y 1 2 3 12 14 15 16 18 22 27 31 32 37 38 40
+ 44
r75 45 46 15.7216 $w=1.94e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=0.925
+ $X2=2.64 $Y2=1.175
r76 38 44 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.64 $Y=1.72
+ $X2=2.64 $Y2=1.665
r77 37 40 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.64 $Y=1.26
+ $X2=2.64 $Y2=1.295
r78 32 38 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.805 $X2=2.64
+ $Y2=1.72
r79 32 44 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=1.65
+ $X2=2.64 $Y2=1.665
r80 31 37 1.66045 $w=2.3e-07 $l=2.5e-08 $layer=LI1_cond $X=2.64 $Y=1.235
+ $X2=2.64 $Y2=1.26
r81 31 46 3.7732 $w=1.94e-07 $l=6e-08 $layer=LI1_cond $X=2.64 $Y=1.235 $X2=2.64
+ $Y2=1.175
r82 31 32 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.64 $Y=1.32
+ $X2=2.64 $Y2=1.65
r83 31 40 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.64 $Y=1.32
+ $X2=2.64 $Y2=1.295
r84 27 29 8.16371 $w=6.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.275 $Y=0.495
+ $X2=3.275 $Y2=0.925
r85 22 24 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.98 $Y=1.97
+ $X2=3.98 $Y2=2.65
r86 20 22 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.98 $Y=1.89 $X2=3.98
+ $Y2=1.97
r87 19 32 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=1.805
+ $X2=2.64 $Y2=1.805
r88 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.815 $Y=1.805
+ $X2=3.98 $Y2=1.89
r89 18 19 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.815 $Y=1.805
+ $X2=2.755 $Y2=1.805
r90 17 45 1.50975 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=0.925
+ $X2=2.64 $Y2=0.925
r91 16 29 8.63246 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=2.96 $Y=0.925
+ $X2=3.275 $Y2=0.925
r92 16 17 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.96 $Y=0.925
+ $X2=2.755 $Y2=0.925
r93 14 46 1.50975 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.525 $Y=1.175
+ $X2=2.64 $Y2=1.175
r94 14 15 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=2.525 $Y=1.175
+ $X2=0.83 $Y2=1.175
r95 10 15 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.74 $Y=1.09
+ $X2=0.83 $Y2=1.175
r96 10 12 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.74 $Y=1.09
+ $X2=0.74 $Y2=0.8
r97 3 24 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.84 $X2=3.98 $Y2=2.65
r98 3 22 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.84 $X2=3.98 $Y2=1.97
r99 2 27 45.5 $w=1.7e-07 $l=5.69078e-07 $layer=licon1_NDIFF $count=4 $X=2.915
+ $Y=0.37 $X2=3.425 $Y2=0.495
r100 1 12 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%A_38_74# 1 2 3 12 14 15 17 19 20 22 24
r45 22 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=0.75
+ $X2=2.115 $Y2=0.835
r46 22 24 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.115 $Y=0.75
+ $X2=2.115 $Y2=0.495
r47 21 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.26 $Y=0.835
+ $X2=1.135 $Y2=0.835
r48 20 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.99 $Y=0.835
+ $X2=2.115 $Y2=0.835
r49 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.99 $Y=0.835
+ $X2=1.26 $Y2=0.835
r50 17 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.75
+ $X2=1.135 $Y2=0.835
r51 17 19 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.135 $Y=0.75
+ $X2=1.135 $Y2=0.495
r52 16 19 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=1.135 $Y=0.425
+ $X2=1.135 $Y2=0.495
r53 14 16 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.01 $Y=0.34
+ $X2=1.135 $Y2=0.425
r54 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.01 $Y=0.34
+ $X2=0.48 $Y2=0.34
r55 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.315 $Y=0.425
+ $X2=0.48 $Y2=0.34
r56 10 12 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.315 $Y=0.425
+ $X2=0.315 $Y2=0.535
r57 3 29 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.37 $X2=2.075 $Y2=0.835
r58 3 24 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.37 $X2=2.075 $Y2=0.495
r59 2 27 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.835
r60 2 19 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.495
r61 1 12 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.19
+ $Y=0.37 $X2=0.315 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_2%VGND 1 2 3 11 14 18 21 22 26 29 30 31 40 49
+ 50 53
c60 26 0 9.12126e-20 $X=1.625 $Y=0.495
c61 11 0 1.42661e-19 $X=1.525 $Y=0.33
r62 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r64 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r65 47 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r66 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r67 44 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.625
+ $Y2=0
r68 44 46 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=3.6
+ $Y2=0
r69 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 40 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.625
+ $Y2=0
r71 40 42 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.16
+ $Y2=0
r72 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r73 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r74 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r75 34 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r76 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 31 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r78 31 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r79 29 46 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.6
+ $Y2=0
r80 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.925
+ $Y2=0
r81 28 49 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.56
+ $Y2=0
r82 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.925
+ $Y2=0
r83 23 26 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=1.525 $Y=0.455
+ $X2=1.625 $Y2=0.455
r84 21 38 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r85 21 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.525
+ $Y2=0
r86 20 42 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.16
+ $Y2=0
r87 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.525
+ $Y2=0
r88 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r89 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.515
r90 12 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0
r91 12 14 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0.55
r92 11 23 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.525 $Y=0.33
+ $X2=1.525 $Y2=0.455
r93 10 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=0.085
+ $X2=1.525 $Y2=0
r94 10 11 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.525 $Y=0.085
+ $X2=1.525 $Y2=0.33
r95 3 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.785
+ $Y=0.37 $X2=3.925 $Y2=0.515
r96 2 14 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.37 $X2=2.625 $Y2=0.55
r97 1 26 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.625 $Y2=0.495
.ends


* NGSPICE file created from sky130_fd_sc_ms__o21a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_219_387# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=5.64e+11p pd=4.92e+06u as=1.9384e+12p ps=1.45e+07u
M1001 VGND a_219_387# X VNB nlowvt w=740000u l=150000u
+  ad=1.1573e+12p pd=1.034e+07u as=4.144e+11p ps=4.08e+06u
M1002 X a_219_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=7.744e+11p pd=7.54e+06u as=0p ps=0u
M1004 VGND A2 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_219_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_219_387# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_219_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1008 VPWR B1 a_219_387# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_219_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_125# B1 a_219_387# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 a_219_387# A2 a_119_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.4e+11p ps=5.28e+06u
M1012 VPWR a_219_387# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_119_387# A2 a_219_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A1 a_119_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_119_387# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_219_387# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_219_387# B1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.413400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.905000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.835000 1.410000 ;
        RECT 0.615000 0.350000 0.945000 0.960000 ;
        RECT 0.615000 0.960000 1.945000 1.130000 ;
        RECT 0.615000 1.130000 0.835000 1.180000 ;
        RECT 0.660000 1.410000 0.835000 1.800000 ;
        RECT 0.660000 1.800000 1.730000 1.970000 ;
        RECT 0.660000 1.970000 0.835000 2.980000 ;
        RECT 1.560000 1.970000 1.730000 2.980000 ;
        RECT 1.615000 0.350000 1.945000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.010000 ;
      RECT 0.130000  1.820000 0.460000 3.245000 ;
      RECT 1.030000  2.140000 1.360000 3.245000 ;
      RECT 1.060000  1.300000 2.285000 1.630000 ;
      RECT 1.115000  0.085000 1.445000 0.790000 ;
      RECT 1.930000  1.820000 2.260000 3.245000 ;
      RECT 2.115000  0.085000 2.745000 0.680000 ;
      RECT 2.115000  0.960000 3.245000 1.130000 ;
      RECT 2.115000  1.130000 2.285000 1.300000 ;
      RECT 2.465000  1.950000 3.245000 2.200000 ;
      RECT 2.915000  0.350000 3.245000 0.960000 ;
      RECT 2.915000  2.370000 3.245000 3.245000 ;
      RECT 3.075000  1.130000 3.245000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ms__buf_4
END LIBRARY

* File: sky130_fd_sc_ms__a22oi_2.pex.spice
* Created: Wed Sep  2 11:53:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A22OI_2%A1 3 7 11 15 17 18 19 20 23 26 27 32 39 41
c91 39 0 1.71862e-19 $X=2.34 $Y=1.515
c92 15 0 7.10839e-20 $X=2.34 $Y=2.4
c93 11 0 1.09905e-19 $X=2.025 $Y=0.74
r94 32 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.515
+ $X2=0.605 $Y2=1.68
r95 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.515
+ $X2=0.605 $Y2=1.35
r96 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.515 $X2=0.605 $Y2=1.515
r97 27 41 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=1.605
+ $X2=0.71 $Y2=1.605
r98 27 41 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.672 $Y=1.605
+ $X2=0.71 $Y2=1.605
r99 27 33 2.20611 $w=3.48e-07 $l=6.7e-08 $layer=LI1_cond $X=0.672 $Y=1.605
+ $X2=0.605 $Y2=1.605
r100 26 33 12.0183 $w=3.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=1.605
+ $X2=0.605 $Y2=1.605
r101 24 39 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=2.045 $Y=1.515
+ $X2=2.34 $Y2=1.515
r102 24 36 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.045 $Y=1.515
+ $X2=2.025 $Y2=1.515
r103 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.045
+ $Y=1.515 $X2=2.045 $Y2=1.515
r104 21 23 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.045 $Y=1.95
+ $X2=2.045 $Y2=1.515
r105 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.88 $Y=2.035
+ $X2=2.045 $Y2=1.95
r106 19 20 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.88 $Y=2.035
+ $X2=0.88 $Y2=2.035
r107 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.795 $Y=1.95
+ $X2=0.88 $Y2=2.035
r108 17 27 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.795 $Y=1.78
+ $X2=0.795 $Y2=1.605
r109 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.795 $Y=1.78
+ $X2=0.795 $Y2=1.95
r110 13 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.68
+ $X2=2.34 $Y2=1.515
r111 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.34 $Y=1.68
+ $X2=2.34 $Y2=2.4
r112 9 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=1.35
+ $X2=2.025 $Y2=1.515
r113 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.025 $Y=1.35
+ $X2=2.025 $Y2=0.74
r114 7 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.68 $Y=2.4 $X2=0.68
+ $Y2=1.68
r115 3 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.665 $Y=0.74
+ $X2=0.665 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%A2 3 7 11 15 17 24 26
r52 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.595 $Y2=1.515
r53 23 25 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.215 $Y=1.515
+ $X2=1.58 $Y2=1.515
r54 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.515 $X2=1.215 $Y2=1.515
r55 21 23 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.215 $Y2=1.515
r56 19 21 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.095 $Y=1.515
+ $X2=1.13 $Y2=1.515
r57 17 24 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.235 $Y=1.665
+ $X2=1.235 $Y2=1.515
r58 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.35
+ $X2=1.595 $Y2=1.515
r59 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.595 $Y=1.35
+ $X2=1.595 $Y2=0.74
r60 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.68
+ $X2=1.58 $Y2=1.515
r61 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.58 $Y=1.68 $X2=1.58
+ $Y2=2.4
r62 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.68
+ $X2=1.13 $Y2=1.515
r63 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.13 $Y=1.68 $X2=1.13
+ $Y2=2.4
r64 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.095 $Y2=1.515
r65 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.095 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%B1 3 6 10 14 16 21 22 25 27 36
c79 36 0 2.81767e-19 $X=3.235 $Y=1.32
c80 25 0 6.84215e-20 $X=2.805 $Y=1.385
c81 21 0 1.74224e-19 $X=4.205 $Y=1.465
r82 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.385
+ $X2=2.805 $Y2=1.55
r83 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.385
+ $X2=2.805 $Y2=1.22
r84 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.385 $X2=2.805 $Y2=1.385
r85 22 36 7.98002 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.32
+ $X2=3.235 $Y2=1.32
r86 22 26 8.19054 $w=4.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.12 $Y=1.32
+ $X2=2.805 $Y2=1.32
r87 21 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.205 $Y=1.465
+ $X2=4.205 $Y2=1.63
r88 21 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.205 $Y=1.465
+ $X2=4.205 $Y2=1.3
r89 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.465 $X2=4.205 $Y2=1.465
r90 16 20 10.1086 $w=3.5e-07 $l=3.89076e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=4.137 $Y2=1.465
r91 16 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=3.235 $Y2=1.175
r92 14 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.17 $Y=2.4 $X2=4.17
+ $Y2=1.63
r93 10 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.115 $Y=0.74
+ $X2=4.115 $Y2=1.3
r94 6 28 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.79 $Y=2.4 $X2=2.79
+ $Y2=1.55
r95 3 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.715 $Y=0.74
+ $X2=2.715 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%B2 3 7 11 15 17 24 26
c51 24 0 2.42645e-19 $X=3.57 $Y=1.515
r52 25 26 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.685 $Y=1.515
+ $X2=3.72 $Y2=1.515
r53 23 25 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.57 $Y=1.515
+ $X2=3.685 $Y2=1.515
r54 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.515 $X2=3.57 $Y2=1.515
r55 21 23 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=3.27 $Y=1.515 $X2=3.57
+ $Y2=1.515
r56 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.255 $Y=1.515
+ $X2=3.27 $Y2=1.515
r57 17 24 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.515
r58 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.68
+ $X2=3.72 $Y2=1.515
r59 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.72 $Y=1.68
+ $X2=3.72 $Y2=2.4
r60 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=1.35
+ $X2=3.685 $Y2=1.515
r61 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.685 $Y=1.35
+ $X2=3.685 $Y2=0.74
r62 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.68
+ $X2=3.27 $Y2=1.515
r63 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.27 $Y=1.68 $X2=3.27
+ $Y2=2.4
r64 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=1.515
r65 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%A_66_368# 1 2 3 4 5 18 22 24 28 33 34 35 38
+ 40 44 46 48 50 53
r78 50 52 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.565 $Y=2.15
+ $X2=2.565 $Y2=2.375
r79 42 44 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.395 $Y=2.905
+ $X2=4.395 $Y2=2.385
r80 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=2.99
+ $X2=3.495 $Y2=2.99
r81 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.23 $Y=2.99
+ $X2=4.395 $Y2=2.905
r82 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.23 $Y=2.99
+ $X2=3.66 $Y2=2.99
r83 36 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.905
+ $X2=3.495 $Y2=2.99
r84 36 38 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.495 $Y=2.905
+ $X2=3.495 $Y2=2.385
r85 34 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=2.99
+ $X2=3.495 $Y2=2.99
r86 34 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.33 $Y=2.99 $X2=2.73
+ $Y2=2.99
r87 31 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.565 $Y=2.905
+ $X2=2.73 $Y2=2.99
r88 31 33 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.565 $Y=2.905
+ $X2=2.565 $Y2=2.83
r89 30 52 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2.46
+ $X2=2.565 $Y2=2.375
r90 30 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.565 $Y=2.46
+ $X2=2.565 $Y2=2.83
r91 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=2.375
+ $X2=1.355 $Y2=2.375
r92 28 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=2.375
+ $X2=2.565 $Y2=2.375
r93 28 29 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.4 $Y=2.375
+ $X2=1.52 $Y2=2.375
r94 25 46 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.54 $Y=2.375
+ $X2=0.415 $Y2=2.375
r95 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=2.375
+ $X2=1.355 $Y2=2.375
r96 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.19 $Y=2.375
+ $X2=0.54 $Y2=2.375
r97 20 46 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=2.46
+ $X2=0.415 $Y2=2.375
r98 20 22 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.415 $Y=2.46
+ $X2=0.415 $Y2=2.465
r99 16 46 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=2.29
+ $X2=0.415 $Y2=2.375
r100 16 18 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.415 $Y=2.29
+ $X2=0.415 $Y2=2.115
r101 5 44 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=4.26
+ $Y=1.84 $X2=4.395 $Y2=2.385
r102 4 38 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.84 $X2=3.495 $Y2=2.385
r103 3 50 400 $w=1.7e-07 $l=3.71416e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.565 $Y2=2.15
r104 3 33 400 $w=1.7e-07 $l=1.05534e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.565 $Y2=2.83
r105 2 48 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.84 $X2=1.355 $Y2=2.375
r106 1 22 300 $w=1.7e-07 $l=6.84653e-07 $layer=licon1_PDIFF $count=2 $X=0.33
+ $Y=1.84 $X2=0.455 $Y2=2.465
r107 1 18 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.84 $X2=0.455 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%VPWR 1 2 9 13 16 17 18 24 30 31 34
r54 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 28 34 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.23 $Y=3.33 $X2=1.96
+ $Y2=3.33
r57 28 30 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=2.23 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 24 34 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.69 $Y=3.33 $X2=1.96
+ $Y2=3.33
r61 24 26 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=3.33 $X2=1.68
+ $Y2=3.33
r62 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 18 31 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.56 $Y2=3.33
r65 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 16 21 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=3.33 $X2=0.72
+ $Y2=3.33
r67 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=0.865 $Y2=3.33
r68 15 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.68
+ $Y2=3.33
r69 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.865 $Y2=3.33
r70 11 34 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=3.33
r71 11 13 9.74582 $w=5.38e-07 $l=4.4e-07 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=2.805
r72 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r73 7 9 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.805
r74 2 13 600 $w=1.7e-07 $l=1.10049e-06 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.84 $X2=1.96 $Y2=2.805
r75 1 9 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.84 $X2=0.905 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%Y 1 2 3 4 5 18 20 21 24 27 28 29 32 34 38 40
+ 44 47 48 54 55 56
c98 48 0 7.10839e-20 $X=3.03 $Y=1.805
r99 63 64 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=1.175
+ $X2=2.295 $Y2=1.26
r100 62 63 4.92503 $w=5.08e-07 $l=2.1e-07 $layer=LI1_cond $X=2.295 $Y=0.965
+ $X2=2.295 $Y2=1.175
r101 56 62 0.938101 $w=5.08e-07 $l=4e-08 $layer=LI1_cond $X=2.295 $Y=0.925
+ $X2=2.295 $Y2=0.965
r102 56 59 3.23794 $w=5.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.295 $Y=0.925
+ $X2=2.295 $Y2=0.81
r103 51 52 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=3.03 $Y=1.985
+ $X2=3.03 $Y2=2.035
r104 48 51 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=3.03 $Y=1.805
+ $X2=3.03 $Y2=1.985
r105 47 55 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=4.625 $Y=1.95
+ $X2=4.625 $Y2=1.13
r106 42 55 11.032 $w=4.63e-07 $l=2.32e-07 $layer=LI1_cond $X=4.477 $Y=0.898
+ $X2=4.477 $Y2=1.13
r107 42 44 9.85157 $w=4.63e-07 $l=3.83e-07 $layer=LI1_cond $X=4.477 $Y=0.898
+ $X2=4.477 $Y2=0.515
r108 41 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.035
+ $X2=3.945 $Y2=2.035
r109 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.54 $Y=2.035
+ $X2=4.625 $Y2=1.95
r110 40 41 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.54 $Y=2.035
+ $X2=4.03 $Y2=2.035
r111 36 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=2.12
+ $X2=3.945 $Y2=2.035
r112 36 38 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.945 $Y=2.12
+ $X2=3.945 $Y2=2.57
r113 35 52 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.13 $Y=2.035 $X2=3.03
+ $Y2=2.035
r114 34 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=2.035
+ $X2=3.945 $Y2=2.035
r115 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.86 $Y=2.035
+ $X2=3.13 $Y2=2.035
r116 30 52 4.71364 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.12
+ $X2=3.03 $Y2=2.035
r117 30 32 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=3.03 $Y=2.12
+ $X2=3.03 $Y2=2.57
r118 28 48 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.93 $Y=1.805 $X2=3.03
+ $Y2=1.805
r119 28 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.93 $Y=1.805
+ $X2=2.55 $Y2=1.805
r120 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=1.72
+ $X2=2.55 $Y2=1.805
r121 27 64 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.465 $Y=1.72
+ $X2=2.465 $Y2=1.26
r122 24 59 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=2.347 $Y=0.515
+ $X2=2.347 $Y2=0.81
r123 20 63 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.04 $Y=1.175
+ $X2=2.295 $Y2=1.175
r124 20 21 98.1872 $w=1.68e-07 $l=1.505e-06 $layer=LI1_cond $X=2.04 $Y=1.175
+ $X2=0.535 $Y2=1.175
r125 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.41 $Y=1.09
+ $X2=0.535 $Y2=1.175
r126 16 18 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=0.41 $Y=1.09
+ $X2=0.41 $Y2=0.515
r127 5 54 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.84 $X2=3.945 $Y2=2.035
r128 5 38 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.84 $X2=3.945 $Y2=2.57
r129 4 51 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=1.985
r130 4 32 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=2.57
r131 3 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.19
+ $Y=0.37 $X2=4.33 $Y2=0.515
r132 2 62 182 $w=1.7e-07 $l=7.06965e-07 $layer=licon1_NDIFF $count=1 $X=2.1
+ $Y=0.37 $X2=2.345 $Y2=0.965
r133 2 24 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=2.1
+ $Y=0.37 $X2=2.345 $Y2=0.515
r134 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.325
+ $Y=0.37 $X2=0.45 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%A_148_74# 1 2 7 9 11 16
r29 16 17 14.5817 $w=2.51e-07 $l=3e-07 $layer=LI1_cond $X=1.81 $Y=0.535 $X2=1.81
+ $Y2=0.835
r30 12 14 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.965 $Y=0.835
+ $X2=0.84 $Y2=0.835
r31 11 17 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0.835
+ $X2=1.81 $Y2=0.835
r32 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.645 $Y=0.835
+ $X2=0.965 $Y2=0.835
r33 7 14 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0.75 $X2=0.84
+ $Y2=0.835
r34 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.84 $Y=0.75 $X2=0.84
+ $Y2=0.495
r35 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.37 $X2=1.81 $Y2=0.535
r36 1 14 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.37 $X2=0.88 $Y2=0.835
r37 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.37 $X2=0.88 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r62 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r63 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r64 33 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r65 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.47
+ $Y2=0
r67 30 32 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=4.56
+ $Y2=0
r68 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r71 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r72 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.31
+ $Y2=0
r74 23 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.68
+ $Y2=0
r75 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.47
+ $Y2=0
r76 22 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.12
+ $Y2=0
r77 20 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r78 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r79 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=1.31
+ $Y2=0
r80 17 19 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=0.24
+ $Y2=0
r81 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r82 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r83 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=0.085
+ $X2=3.47 $Y2=0
r84 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.47 $Y=0.085
+ $X2=3.47 $Y2=0.495
r85 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085 $X2=1.31
+ $Y2=0
r86 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.31 $Y=0.085 $X2=1.31
+ $Y2=0.495
r87 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.37 $X2=3.47 $Y2=0.495
r88 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.17
+ $Y=0.37 $X2=1.31 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_2%A_558_74# 1 2 7 9 11 13 15
r28 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.94 $Y=0.75 $X2=3.94
+ $Y2=0.835
r29 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.94 $Y=0.75
+ $X2=3.94 $Y2=0.495
r30 12 18 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.135 $Y=0.835
+ $X2=2.985 $Y2=0.835
r31 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.815 $Y=0.835
+ $X2=3.94 $Y2=0.835
r32 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.815 $Y=0.835
+ $X2=3.135 $Y2=0.835
r33 7 18 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.75 $X2=2.985
+ $Y2=0.835
r34 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.985 $Y=0.75
+ $X2=2.985 $Y2=0.495
r35 2 20 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.37 $X2=3.9 $Y2=0.835
r36 2 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.37 $X2=3.9 $Y2=0.495
r37 1 18 182 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=3 $Y2=0.835
r38 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=3 $Y2=0.495
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR SCE a_310_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X1 a_27_79# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VGND a_852_119# a_1025_119# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_2006_373# a_1790_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X4 a_2158_74# a_1790_74# a_2006_373# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 a_388_79# a_1025_119# a_1223_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X6 VGND a_2607_392# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_388_79# a_852_119# a_1223_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X8 a_310_464# D a_388_79# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X9 a_1223_119# a_852_119# a_1328_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X10 a_223_79# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_223_79# a_27_79# a_310_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 a_388_79# SCE a_547_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_1401_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 VPWR a_2607_392# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_852_119# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 VPWR RESET_B a_388_79# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X17 a_852_119# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR a_1790_74# a_2607_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X19 VGND RESET_B a_2158_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VGND a_1790_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 Q a_2607_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VPWR a_852_119# a_1025_119# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 a_1328_457# a_1370_290# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X24 a_1958_471# a_2006_373# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X25 a_1223_119# a_1025_119# a_1323_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 VGND a_1790_74# a_2607_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 a_27_79# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X28 a_541_483# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X29 a_1370_290# a_852_119# a_1790_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X30 VPWR a_1790_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 a_2000_74# a_2006_373# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_1790_74# a_1025_119# a_1958_471# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X33 VPWR RESET_B a_2006_373# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X34 a_1790_74# a_852_119# a_2000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 VGND a_1223_119# a_1370_290# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X36 a_388_79# a_27_79# a_541_483# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X37 a_310_79# D a_388_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 Q a_2607_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X39 VPWR a_1223_119# a_1370_290# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X40 a_547_79# SCD a_223_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X41 VPWR RESET_B a_1223_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X42 a_1323_119# a_1370_290# a_1401_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X43 Q_N a_1790_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X44 a_1370_290# a_1025_119# a_1790_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X45 Q_N a_1790_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

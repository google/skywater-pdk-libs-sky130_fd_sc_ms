* File: sky130_fd_sc_ms__dlrbp_2.pxi.spice
* Created: Fri Aug 28 17:27:20 2020
* 
x_PM_SKY130_FD_SC_MS__DLRBP_2%D N_D_M1000_g N_D_M1015_g D N_D_c_180_n
+ PM_SKY130_FD_SC_MS__DLRBP_2%D
x_PM_SKY130_FD_SC_MS__DLRBP_2%GATE N_GATE_M1013_g N_GATE_M1017_g GATE
+ N_GATE_c_219_n N_GATE_c_220_n PM_SKY130_FD_SC_MS__DLRBP_2%GATE
x_PM_SKY130_FD_SC_MS__DLRBP_2%A_230_74# N_A_230_74#_M1013_d N_A_230_74#_M1017_d
+ N_A_230_74#_c_255_n N_A_230_74#_c_256_n N_A_230_74#_M1001_g
+ N_A_230_74#_c_258_n N_A_230_74#_M1002_g N_A_230_74#_c_269_n
+ N_A_230_74#_M1014_g N_A_230_74#_c_270_n N_A_230_74#_c_271_n
+ N_A_230_74#_M1003_g N_A_230_74#_c_273_n N_A_230_74#_c_260_n
+ N_A_230_74#_c_261_n N_A_230_74#_c_262_n N_A_230_74#_c_263_n
+ N_A_230_74#_c_264_n N_A_230_74#_c_274_n N_A_230_74#_c_265_n
+ N_A_230_74#_c_266_n N_A_230_74#_c_267_n PM_SKY130_FD_SC_MS__DLRBP_2%A_230_74#
x_PM_SKY130_FD_SC_MS__DLRBP_2%A_27_112# N_A_27_112#_M1015_s N_A_27_112#_M1000_s
+ N_A_27_112#_M1010_g N_A_27_112#_M1004_g N_A_27_112#_c_393_n
+ N_A_27_112#_c_399_n N_A_27_112#_c_400_n N_A_27_112#_c_401_n
+ N_A_27_112#_c_394_n N_A_27_112#_c_395_n N_A_27_112#_c_396_n
+ N_A_27_112#_c_404_n N_A_27_112#_c_397_n PM_SKY130_FD_SC_MS__DLRBP_2%A_27_112#
x_PM_SKY130_FD_SC_MS__DLRBP_2%A_363_82# N_A_363_82#_M1002_s N_A_363_82#_M1001_s
+ N_A_363_82#_M1023_g N_A_363_82#_M1020_g N_A_363_82#_c_477_n
+ N_A_363_82#_c_478_n N_A_363_82#_c_479_n N_A_363_82#_c_480_n
+ N_A_363_82#_c_487_n N_A_363_82#_c_488_n N_A_363_82#_c_489_n
+ N_A_363_82#_c_490_n N_A_363_82#_c_491_n N_A_363_82#_c_481_n
+ N_A_363_82#_c_482_n N_A_363_82#_c_483_n PM_SKY130_FD_SC_MS__DLRBP_2%A_363_82#
x_PM_SKY130_FD_SC_MS__DLRBP_2%A_821_98# N_A_821_98#_M1016_s N_A_821_98#_M1027_d
+ N_A_821_98#_c_596_n N_A_821_98#_M1018_g N_A_821_98#_M1007_g
+ N_A_821_98#_M1024_g N_A_821_98#_M1021_g N_A_821_98#_M1025_g
+ N_A_821_98#_M1022_g N_A_821_98#_c_601_n N_A_821_98#_c_602_n
+ N_A_821_98#_M1012_g N_A_821_98#_M1006_g N_A_821_98#_c_605_n
+ N_A_821_98#_c_606_n N_A_821_98#_c_616_n N_A_821_98#_c_617_n
+ N_A_821_98#_c_607_n N_A_821_98#_c_618_n N_A_821_98#_c_619_n
+ N_A_821_98#_c_608_n N_A_821_98#_c_726_p N_A_821_98#_c_609_n
+ N_A_821_98#_c_621_n N_A_821_98#_c_610_n N_A_821_98#_c_611_n
+ PM_SKY130_FD_SC_MS__DLRBP_2%A_821_98#
x_PM_SKY130_FD_SC_MS__DLRBP_2%A_641_80# N_A_641_80#_M1023_d N_A_641_80#_M1014_d
+ N_A_641_80#_M1027_g N_A_641_80#_M1016_g N_A_641_80#_c_765_n
+ N_A_641_80#_c_766_n N_A_641_80#_c_779_n N_A_641_80#_c_774_n
+ N_A_641_80#_c_767_n N_A_641_80#_c_768_n N_A_641_80#_c_769_n
+ N_A_641_80#_c_770_n PM_SKY130_FD_SC_MS__DLRBP_2%A_641_80#
x_PM_SKY130_FD_SC_MS__DLRBP_2%RESET_B N_RESET_B_M1009_g N_RESET_B_M1026_g
+ RESET_B N_RESET_B_c_851_n N_RESET_B_c_852_n N_RESET_B_c_853_n
+ PM_SKY130_FD_SC_MS__DLRBP_2%RESET_B
x_PM_SKY130_FD_SC_MS__DLRBP_2%A_1449_368# N_A_1449_368#_M1006_s
+ N_A_1449_368#_M1012_s N_A_1449_368#_M1005_g N_A_1449_368#_M1011_g
+ N_A_1449_368#_M1008_g N_A_1449_368#_M1019_g N_A_1449_368#_c_894_n
+ N_A_1449_368#_c_895_n N_A_1449_368#_c_896_n N_A_1449_368#_c_897_n
+ N_A_1449_368#_c_898_n N_A_1449_368#_c_912_n N_A_1449_368#_c_899_n
+ PM_SKY130_FD_SC_MS__DLRBP_2%A_1449_368#
x_PM_SKY130_FD_SC_MS__DLRBP_2%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1007_d
+ N_VPWR_M1026_d N_VPWR_M1022_s N_VPWR_M1012_d N_VPWR_M1008_s N_VPWR_c_962_n
+ N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n N_VPWR_c_966_n N_VPWR_c_967_n
+ N_VPWR_c_968_n N_VPWR_c_969_n N_VPWR_c_970_n N_VPWR_c_971_n N_VPWR_c_972_n
+ VPWR N_VPWR_c_973_n N_VPWR_c_974_n N_VPWR_c_975_n N_VPWR_c_976_n
+ N_VPWR_c_977_n N_VPWR_c_978_n N_VPWR_c_979_n N_VPWR_c_980_n N_VPWR_c_961_n
+ PM_SKY130_FD_SC_MS__DLRBP_2%VPWR
x_PM_SKY130_FD_SC_MS__DLRBP_2%Q N_Q_M1024_d N_Q_M1021_d N_Q_c_1076_n
+ N_Q_c_1080_n N_Q_c_1081_n N_Q_c_1082_n N_Q_c_1077_n N_Q_c_1078_n Q
+ PM_SKY130_FD_SC_MS__DLRBP_2%Q
x_PM_SKY130_FD_SC_MS__DLRBP_2%Q_N N_Q_N_M1011_d N_Q_N_M1005_d N_Q_N_c_1129_n
+ N_Q_N_c_1130_n Q_N Q_N N_Q_N_c_1131_n PM_SKY130_FD_SC_MS__DLRBP_2%Q_N
x_PM_SKY130_FD_SC_MS__DLRBP_2%VGND N_VGND_M1015_d N_VGND_M1002_d N_VGND_M1018_d
+ N_VGND_M1009_d N_VGND_M1025_s N_VGND_M1006_d N_VGND_M1019_s N_VGND_c_1160_n
+ N_VGND_c_1161_n N_VGND_c_1162_n N_VGND_c_1163_n N_VGND_c_1164_n
+ N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n N_VGND_c_1168_n
+ N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n N_VGND_c_1172_n
+ N_VGND_c_1173_n VGND N_VGND_c_1174_n N_VGND_c_1175_n N_VGND_c_1176_n
+ N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n
+ PM_SKY130_FD_SC_MS__DLRBP_2%VGND
cc_1 VNB N_D_M1015_g 0.0375151f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB D 0.00242107f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_c_180_n 0.0220003f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_4 VNB N_GATE_M1017_g 0.00639429f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_5 VNB GATE 0.0061593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_GATE_c_219_n 0.0351695f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.615
cc_7 VNB N_GATE_c_220_n 0.0226366f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_8 VNB N_A_230_74#_c_255_n 0.0153485f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_9 VNB N_A_230_74#_c_256_n 0.0150744f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A_230_74#_M1001_g 0.00785243f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.615
cc_11 VNB N_A_230_74#_c_258_n 0.0187611f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_12 VNB N_A_230_74#_M1003_g 0.0417255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_230_74#_c_260_n 0.00580127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_230_74#_c_261_n 0.00163151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_230_74#_c_262_n 0.00874055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_230_74#_c_263_n 0.0446354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_230_74#_c_264_n 0.0163502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_230_74#_c_265_n 0.00543595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_230_74#_c_266_n 0.00643839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_230_74#_c_267_n 0.0272613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_112#_M1004_g 0.0326722f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_22 VNB N_A_27_112#_c_393_n 0.0201039f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.78
cc_23 VNB N_A_27_112#_c_394_n 0.00196261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_112#_c_395_n 0.0208665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_112#_c_396_n 0.013652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_112#_c_397_n 0.0253939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_363_82#_c_477_n 0.00623344f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.45
cc_28 VNB N_A_363_82#_c_478_n 0.00153466f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.78
cc_29 VNB N_A_363_82#_c_479_n 0.0177304f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_30 VNB N_A_363_82#_c_480_n 0.00287888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_363_82#_c_481_n 0.00746834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_363_82#_c_482_n 0.0308969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_363_82#_c_483_n 0.0159056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_821_98#_c_596_n 0.0171346f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_35 VNB N_A_821_98#_M1024_g 0.0223246f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_36 VNB N_A_821_98#_M1021_g 0.00151147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_821_98#_M1025_g 0.0227941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_821_98#_M1022_g 0.00169796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_821_98#_c_601_n 0.0762963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_821_98#_c_602_n 0.0334681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_821_98#_M1012_g 0.0020378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_821_98#_M1006_g 0.0259366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_821_98#_c_605_n 0.0198739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_821_98#_c_606_n 0.00991002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_821_98#_c_607_n 0.00813778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_821_98#_c_608_n 0.00536874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_821_98#_c_609_n 0.00577602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_821_98#_c_610_n 0.00387127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_821_98#_c_611_n 0.0227549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_641_80#_M1016_g 0.0266521f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_51 VNB N_A_641_80#_c_765_n 0.0311649f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.78
cc_52 VNB N_A_641_80#_c_766_n 0.0126002f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_53 VNB N_A_641_80#_c_767_n 0.00574196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_641_80#_c_768_n 0.0140086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_641_80#_c_769_n 0.007314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_641_80#_c_770_n 0.00856244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_M1026_g 0.00653808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_58 VNB N_RESET_B_c_851_n 0.0276452f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.615
cc_59 VNB N_RESET_B_c_852_n 0.00860315f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_60 VNB N_RESET_B_c_853_n 0.0172008f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_61 VNB N_A_1449_368#_M1005_g 0.00169308f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_62 VNB N_A_1449_368#_M1011_g 0.0229007f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_63 VNB N_A_1449_368#_M1008_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1449_368#_M1019_g 0.0260184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1449_368#_c_894_n 0.00924021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1449_368#_c_895_n 0.00129392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1449_368#_c_896_n 2.15008e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1449_368#_c_897_n 0.00569931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1449_368#_c_898_n 0.00140993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1449_368#_c_899_n 0.0651793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VPWR_c_961_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_Q_c_1076_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_73 VNB N_Q_c_1077_n 0.00849508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_Q_c_1078_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB Q 0.00348326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_Q_N_c_1129_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_77 VNB N_Q_N_c_1130_n 0.00429087f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_78 VNB N_Q_N_c_1131_n 0.00141953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1160_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1161_n 0.0219756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1162_n 0.00650187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1163_n 0.0171896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1164_n 0.0166669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1165_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1166_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1167_n 0.0514319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1168_n 0.0393212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1169_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1170_n 0.0294964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1171_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1172_n 0.0199677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1173_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1174_n 0.020108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1175_n 0.0221748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1176_n 0.0189349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1177_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1178_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1179_n 0.519539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VPB N_D_M1000_g 0.0298218f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_100 VPB D 0.00201744f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_101 VPB N_D_c_180_n 0.0139774f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_102 VPB N_GATE_M1017_g 0.0366343f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_103 VPB N_A_230_74#_M1001_g 0.036851f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.615
cc_104 VPB N_A_230_74#_c_269_n 0.0185141f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_105 VPB N_A_230_74#_c_270_n 0.0407751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_230_74#_c_271_n 0.00723652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_230_74#_M1003_g 0.00178447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_230_74#_c_273_n 0.00637912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_230_74#_c_274_n 0.0103231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_230_74#_c_265_n 0.007206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_230_74#_c_267_n 0.0100279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_112#_M1010_g 0.0228445f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_113 VPB N_A_27_112#_c_399_n 0.00900146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_112#_c_400_n 0.0094938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_112#_c_401_n 0.0224391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_112#_c_394_n 0.0011621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_112#_c_395_n 0.0154774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_112#_c_404_n 0.0136598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_112#_c_397_n 0.0137381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_363_82#_M1020_g 0.0228867f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_121 VPB N_A_363_82#_c_478_n 0.0037823f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.78
cc_122 VPB N_A_363_82#_c_480_n 0.00199465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_363_82#_c_487_n 0.00545495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_363_82#_c_488_n 0.00161412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_363_82#_c_489_n 0.00462548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_363_82#_c_490_n 0.0419973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_363_82#_c_491_n 0.00514446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_821_98#_M1007_g 0.0300701f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.45
cc_129 VPB N_A_821_98#_M1021_g 0.0228447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_821_98#_M1022_g 0.0248245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_821_98#_M1012_g 0.026758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_821_98#_c_616_n 0.0085437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_821_98#_c_617_n 0.031649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_821_98#_c_618_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_821_98#_c_619_n 0.00648423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_821_98#_c_608_n 8.45725e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_821_98#_c_621_n 0.00760266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_821_98#_c_610_n 6.12609e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_821_98#_c_611_n 0.0239464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_641_80#_M1027_g 0.0237964f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_141 VPB N_A_641_80#_c_765_n 0.013129f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.78
cc_142 VPB N_A_641_80#_c_766_n 6.79367e-19 $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_143 VPB N_A_641_80#_c_774_n 0.00481065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_641_80#_c_768_n 0.0101806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_641_80#_c_769_n 2.16397e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_641_80#_c_770_n 0.00406649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_M1026_g 0.0235049f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_148 VPB N_A_1449_368#_M1005_g 0.0239816f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_149 VPB N_A_1449_368#_M1008_g 0.0274013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_1449_368#_c_896_n 0.00459592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_962_n 0.0212529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_963_n 0.0128974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_964_n 0.00823421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_965_n 0.0172466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_966_n 0.0176566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_967_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_968_n 0.0644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_969_n 0.0185677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_970_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_971_n 0.0175592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_972_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_973_n 0.0428961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_974_n 0.0443808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_975_n 0.0212658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_976_n 0.0194151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_977_n 0.0270908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_978_n 0.00680249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_979_n 0.0176638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_980_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_961_n 0.120264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_Q_c_1080_n 0.00180133f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_172 VPB N_Q_c_1081_n 0.00769988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_Q_c_1082_n 0.00156994f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_174 VPB Q 0.00234304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB Q_N 0.00447264f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.45
cc_176 VPB Q_N 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_Q_N_c_1131_n 0.0010488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 N_D_M1000_g N_GATE_M1017_g 0.0301116f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_179 D N_GATE_M1017_g 0.00243125f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_180 N_D_c_180_n N_GATE_M1017_g 0.00959987f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_181 N_D_M1015_g GATE 0.00204708f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_182 D GATE 0.00792655f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_183 N_D_M1015_g N_GATE_c_219_n 0.00769876f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_184 D N_GATE_c_219_n 5.77592e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_185 N_D_c_180_n N_GATE_c_219_n 0.0062543f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_186 N_D_M1015_g N_GATE_c_220_n 0.0167806f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_187 N_D_M1000_g N_A_230_74#_c_274_n 0.00109847f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_188 D N_A_230_74#_c_265_n 0.00736576f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_189 N_D_M1015_g N_A_27_112#_c_393_n 0.00673958f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_190 N_D_M1000_g N_A_27_112#_c_399_n 0.00599381f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_191 N_D_M1000_g N_A_27_112#_c_400_n 0.0123041f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_192 D N_A_27_112#_c_400_n 0.00917545f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_193 N_D_c_180_n N_A_27_112#_c_400_n 0.00243769f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_194 N_D_M1000_g N_A_27_112#_c_401_n 0.00854305f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_195 N_D_M1015_g N_A_27_112#_c_396_n 0.00583243f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_196 D N_A_27_112#_c_396_n 9.01811e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_197 N_D_c_180_n N_A_27_112#_c_396_n 2.01578e-19 $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_198 N_D_M1000_g N_A_27_112#_c_404_n 0.004898f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_199 D N_A_27_112#_c_404_n 0.00151667f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_200 N_D_M1015_g N_A_27_112#_c_397_n 0.00927701f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_201 D N_A_27_112#_c_397_n 0.0250412f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_202 N_D_c_180_n N_A_27_112#_c_397_n 0.011781f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_203 N_D_M1000_g N_VPWR_c_962_n 0.00407412f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_204 N_D_M1000_g N_VPWR_c_977_n 0.00539235f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_205 N_D_M1000_g N_VPWR_c_961_n 0.00595788f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_206 N_D_M1015_g N_VGND_c_1160_n 0.00610345f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_207 D N_VGND_c_1160_n 0.00727791f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_208 N_D_c_180_n N_VGND_c_1160_n 0.00252403f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_209 N_D_M1015_g N_VGND_c_1174_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_210 N_D_M1015_g N_VGND_c_1179_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_211 GATE N_A_230_74#_c_264_n 0.0110796f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_212 N_GATE_c_219_n N_A_230_74#_c_264_n 0.00124546f $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_213 N_GATE_c_220_n N_A_230_74#_c_264_n 0.0080587f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_214 N_GATE_M1017_g N_A_230_74#_c_274_n 0.00700445f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_215 GATE N_A_230_74#_c_274_n 0.00405092f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_216 N_GATE_c_219_n N_A_230_74#_c_274_n 7.65906e-19 $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_217 N_GATE_M1017_g N_A_230_74#_c_265_n 0.00897006f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_218 GATE N_A_230_74#_c_266_n 0.0289292f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_219 N_GATE_c_219_n N_A_230_74#_c_266_n 0.00404058f $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_220 N_GATE_c_220_n N_A_230_74#_c_266_n 0.00376199f $X=1.13 $Y=1.22 $X2=0
+ $Y2=0
cc_221 N_GATE_M1017_g N_A_230_74#_c_267_n 0.00418042f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_222 GATE N_A_230_74#_c_267_n 2.22836e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_223 N_GATE_c_219_n N_A_230_74#_c_267_n 0.0110794f $X=1.13 $Y=1.385 $X2=0
+ $Y2=0
cc_224 N_GATE_c_220_n N_A_27_112#_c_393_n 6.40098e-19 $X=1.13 $Y=1.22 $X2=0
+ $Y2=0
cc_225 N_GATE_M1017_g N_A_27_112#_c_400_n 0.0205793f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_226 N_GATE_M1017_g N_A_27_112#_c_401_n 7.80168e-19 $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_227 N_GATE_M1017_g N_A_27_112#_c_404_n 0.00181332f $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_228 N_GATE_M1017_g N_A_363_82#_c_491_n 3.52257e-19 $X=1.125 $Y=2.38 $X2=0
+ $Y2=0
cc_229 N_GATE_M1017_g N_VPWR_c_962_n 0.00443659f $X=1.125 $Y=2.38 $X2=0 $Y2=0
cc_230 N_GATE_M1017_g N_VPWR_c_973_n 0.00562877f $X=1.125 $Y=2.38 $X2=0 $Y2=0
cc_231 N_GATE_M1017_g N_VPWR_c_961_n 0.00595788f $X=1.125 $Y=2.38 $X2=0 $Y2=0
cc_232 N_GATE_c_220_n N_VGND_c_1160_n 0.00984417f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_233 N_GATE_c_220_n N_VGND_c_1167_n 0.00434272f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_234 N_GATE_c_220_n N_VGND_c_1179_n 0.00830058f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_235 N_A_230_74#_M1001_g N_A_27_112#_M1010_g 0.026453f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_236 N_A_230_74#_c_269_n N_A_27_112#_M1010_g 0.0352008f $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_237 N_A_230_74#_c_256_n N_A_27_112#_M1004_g 0.00760431f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_238 N_A_230_74#_c_258_n N_A_27_112#_M1004_g 0.0247978f $X=2.175 $Y=1.225
+ $X2=0 $Y2=0
cc_239 N_A_230_74#_c_260_n N_A_27_112#_M1004_g 0.00971882f $X=2.81 $Y=0.665
+ $X2=0 $Y2=0
cc_240 N_A_230_74#_c_261_n N_A_27_112#_M1004_g 0.00982733f $X=2.98 $Y=0.382
+ $X2=0 $Y2=0
cc_241 N_A_230_74#_c_262_n N_A_27_112#_M1004_g 2.18501e-19 $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_242 N_A_230_74#_M1017_d N_A_27_112#_c_400_n 0.0095968f $X=1.215 $Y=1.96 $X2=0
+ $Y2=0
cc_243 N_A_230_74#_M1001_g N_A_27_112#_c_400_n 0.0179132f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_244 N_A_230_74#_c_274_n N_A_27_112#_c_400_n 0.0286837f $X=1.54 $Y=2.065 $X2=0
+ $Y2=0
cc_245 N_A_230_74#_c_267_n N_A_27_112#_c_400_n 0.00207455f $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_246 N_A_230_74#_c_256_n N_A_27_112#_c_394_n 0.0011064f $X=2.185 $Y=1.49 $X2=0
+ $Y2=0
cc_247 N_A_230_74#_M1001_g N_A_27_112#_c_394_n 0.00712986f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_248 N_A_230_74#_c_271_n N_A_27_112#_c_394_n 6.49375e-19 $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_249 N_A_230_74#_c_256_n N_A_27_112#_c_395_n 0.019726f $X=2.185 $Y=1.49 $X2=0
+ $Y2=0
cc_250 N_A_230_74#_c_271_n N_A_27_112#_c_395_n 0.0352008f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_251 N_A_230_74#_c_260_n N_A_363_82#_M1002_s 0.00689956f $X=2.81 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_252 N_A_230_74#_c_256_n N_A_363_82#_c_477_n 0.00189668f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_253 N_A_230_74#_c_258_n N_A_363_82#_c_477_n 0.00934554f $X=2.175 $Y=1.225
+ $X2=0 $Y2=0
cc_254 N_A_230_74#_c_260_n N_A_363_82#_c_477_n 0.0267031f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_255 N_A_230_74#_c_264_n N_A_363_82#_c_477_n 0.0209634f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_256 N_A_230_74#_c_265_n N_A_363_82#_c_477_n 0.00539606f $X=1.7 $Y=1.505 $X2=0
+ $Y2=0
cc_257 N_A_230_74#_c_266_n N_A_363_82#_c_477_n 0.00596096f $X=1.66 $Y=1.34 $X2=0
+ $Y2=0
cc_258 N_A_230_74#_c_267_n N_A_363_82#_c_477_n 0.00663024f $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_259 N_A_230_74#_c_255_n N_A_363_82#_c_478_n 0.00541098f $X=2.095 $Y=1.415
+ $X2=0 $Y2=0
cc_260 N_A_230_74#_c_256_n N_A_363_82#_c_478_n 0.00546978f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_261 N_A_230_74#_M1001_g N_A_363_82#_c_478_n 0.0137143f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_262 N_A_230_74#_c_273_n N_A_363_82#_c_478_n 0.0110443f $X=1.54 $Y=1.94 $X2=0
+ $Y2=0
cc_263 N_A_230_74#_c_265_n N_A_363_82#_c_478_n 0.0246582f $X=1.7 $Y=1.505 $X2=0
+ $Y2=0
cc_264 N_A_230_74#_c_266_n N_A_363_82#_c_478_n 0.00159827f $X=1.66 $Y=1.34 $X2=0
+ $Y2=0
cc_265 N_A_230_74#_c_267_n N_A_363_82#_c_478_n 9.9735e-19 $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_266 N_A_230_74#_c_256_n N_A_363_82#_c_479_n 0.00510753f $X=2.185 $Y=1.49
+ $X2=0 $Y2=0
cc_267 N_A_230_74#_c_258_n N_A_363_82#_c_479_n 0.00284581f $X=2.175 $Y=1.225
+ $X2=0 $Y2=0
cc_268 N_A_230_74#_c_260_n N_A_363_82#_c_479_n 0.0204051f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_269 N_A_230_74#_c_261_n N_A_363_82#_c_479_n 0.005856f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_270 N_A_230_74#_c_269_n N_A_363_82#_c_480_n 0.0215112f $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_271 N_A_230_74#_c_271_n N_A_363_82#_c_480_n 0.00421618f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_272 N_A_230_74#_M1003_g N_A_363_82#_c_480_n 8.84971e-19 $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_273 N_A_230_74#_c_269_n N_A_363_82#_c_487_n 0.0101099f $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_274 N_A_230_74#_c_269_n N_A_363_82#_c_488_n 0.00217084f $X=3.175 $Y=1.84
+ $X2=0 $Y2=0
cc_275 N_A_230_74#_c_269_n N_A_363_82#_c_489_n 7.18546e-19 $X=3.175 $Y=1.84
+ $X2=0 $Y2=0
cc_276 N_A_230_74#_c_270_n N_A_363_82#_c_489_n 6.37973e-19 $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_277 N_A_230_74#_c_269_n N_A_363_82#_c_490_n 0.0213756f $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_278 N_A_230_74#_c_270_n N_A_363_82#_c_490_n 0.0163458f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_279 N_A_230_74#_c_255_n N_A_363_82#_c_491_n 0.00469925f $X=2.095 $Y=1.415
+ $X2=0 $Y2=0
cc_280 N_A_230_74#_M1001_g N_A_363_82#_c_491_n 0.0070225f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_281 N_A_230_74#_c_274_n N_A_363_82#_c_491_n 0.0216496f $X=1.54 $Y=2.065 $X2=0
+ $Y2=0
cc_282 N_A_230_74#_c_265_n N_A_363_82#_c_491_n 0.00379671f $X=1.7 $Y=1.505 $X2=0
+ $Y2=0
cc_283 N_A_230_74#_c_267_n N_A_363_82#_c_491_n 4.58946e-19 $X=1.7 $Y=1.415 $X2=0
+ $Y2=0
cc_284 N_A_230_74#_c_271_n N_A_363_82#_c_481_n 0.00125576f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_285 N_A_230_74#_M1003_g N_A_363_82#_c_481_n 4.00544e-19 $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_286 N_A_230_74#_c_262_n N_A_363_82#_c_481_n 0.00497076f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_287 N_A_230_74#_c_271_n N_A_363_82#_c_482_n 0.0194307f $X=3.265 $Y=1.765
+ $X2=0 $Y2=0
cc_288 N_A_230_74#_M1003_g N_A_363_82#_c_482_n 0.0113395f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_289 N_A_230_74#_M1003_g N_A_363_82#_c_483_n 0.0147384f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_290 N_A_230_74#_c_261_n N_A_363_82#_c_483_n 0.00569577f $X=2.98 $Y=0.382
+ $X2=0 $Y2=0
cc_291 N_A_230_74#_c_262_n N_A_363_82#_c_483_n 0.0137397f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_292 N_A_230_74#_c_263_n N_A_363_82#_c_483_n 0.00778027f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_293 N_A_230_74#_M1003_g N_A_821_98#_c_596_n 0.0393303f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_294 N_A_230_74#_c_263_n N_A_821_98#_c_596_n 0.00120024f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_295 N_A_230_74#_M1003_g N_A_821_98#_c_611_n 0.0188158f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_296 N_A_230_74#_c_262_n N_A_641_80#_M1023_d 0.0024671f $X=3.73 $Y=0.345
+ $X2=-0.19 $Y2=-0.245
cc_297 N_A_230_74#_M1003_g N_A_641_80#_c_779_n 0.00630606f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_298 N_A_230_74#_c_262_n N_A_641_80#_c_779_n 0.0227491f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_299 N_A_230_74#_c_263_n N_A_641_80#_c_779_n 0.00305359f $X=3.73 $Y=0.345
+ $X2=0 $Y2=0
cc_300 N_A_230_74#_c_269_n N_A_641_80#_c_774_n 0.00310466f $X=3.175 $Y=1.84
+ $X2=0 $Y2=0
cc_301 N_A_230_74#_c_270_n N_A_641_80#_c_774_n 0.00595711f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_302 N_A_230_74#_c_270_n N_A_641_80#_c_767_n 0.00150476f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_303 N_A_230_74#_M1003_g N_A_641_80#_c_767_n 0.0202191f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_304 N_A_230_74#_c_270_n N_A_641_80#_c_768_n 0.00422622f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_305 N_A_230_74#_M1003_g N_A_641_80#_c_768_n 0.00648948f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_306 N_A_230_74#_c_270_n N_A_641_80#_c_769_n 0.0187322f $X=3.715 $Y=1.765
+ $X2=0 $Y2=0
cc_307 N_A_230_74#_M1003_g N_A_641_80#_c_769_n 9.81799e-19 $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_308 N_A_230_74#_M1001_g N_VPWR_c_963_n 0.00436483f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_309 N_A_230_74#_c_269_n N_VPWR_c_963_n 4.16264e-19 $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_310 N_A_230_74#_M1001_g N_VPWR_c_973_n 0.00562877f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_311 N_A_230_74#_c_269_n N_VPWR_c_974_n 0.00333867f $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_312 N_A_230_74#_M1001_g N_VPWR_c_961_n 0.00595788f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_313 N_A_230_74#_c_269_n N_VPWR_c_961_n 0.00423361f $X=3.175 $Y=1.84 $X2=0
+ $Y2=0
cc_314 N_A_230_74#_c_260_n N_VGND_M1002_d 0.00930264f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_315 N_A_230_74#_c_264_n N_VGND_c_1160_n 0.02718f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_316 N_A_230_74#_M1003_g N_VGND_c_1161_n 0.00214993f $X=3.79 $Y=0.83 $X2=0
+ $Y2=0
cc_317 N_A_230_74#_c_262_n N_VGND_c_1161_n 0.01269f $X=3.73 $Y=0.345 $X2=0 $Y2=0
cc_318 N_A_230_74#_c_263_n N_VGND_c_1161_n 0.00337434f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_319 N_A_230_74#_c_258_n N_VGND_c_1167_n 0.00794823f $X=2.175 $Y=1.225 $X2=0
+ $Y2=0
cc_320 N_A_230_74#_c_260_n N_VGND_c_1167_n 0.037305f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_321 N_A_230_74#_c_261_n N_VGND_c_1167_n 0.0113147f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_322 N_A_230_74#_c_264_n N_VGND_c_1167_n 0.0221178f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_323 N_A_230_74#_c_260_n N_VGND_c_1168_n 0.00276577f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_324 N_A_230_74#_c_261_n N_VGND_c_1168_n 0.0117598f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_325 N_A_230_74#_c_262_n N_VGND_c_1168_n 0.0596213f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_326 N_A_230_74#_c_263_n N_VGND_c_1168_n 0.00653686f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_327 N_A_230_74#_c_258_n N_VGND_c_1179_n 0.00533081f $X=2.175 $Y=1.225 $X2=0
+ $Y2=0
cc_328 N_A_230_74#_c_260_n N_VGND_c_1179_n 0.0268131f $X=2.81 $Y=0.665 $X2=0
+ $Y2=0
cc_329 N_A_230_74#_c_261_n N_VGND_c_1179_n 0.00647831f $X=2.98 $Y=0.382 $X2=0
+ $Y2=0
cc_330 N_A_230_74#_c_262_n N_VGND_c_1179_n 0.0332028f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_331 N_A_230_74#_c_263_n N_VGND_c_1179_n 0.0102677f $X=3.73 $Y=0.345 $X2=0
+ $Y2=0
cc_332 N_A_230_74#_c_264_n N_VGND_c_1179_n 0.0182647f $X=1.29 $Y=0.515 $X2=0
+ $Y2=0
cc_333 N_A_230_74#_c_261_n A_569_80# 0.00410008f $X=2.98 $Y=0.382 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_230_74#_c_262_n A_569_80# 6.30424e-19 $X=3.73 $Y=0.345 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_27_112#_c_400_n N_A_363_82#_M1001_s 0.00757931f $X=2.485 $Y=2.445
+ $X2=0 $Y2=0
cc_336 N_A_27_112#_M1004_g N_A_363_82#_c_477_n 0.00107979f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_337 N_A_27_112#_M1004_g N_A_363_82#_c_478_n 8.52697e-19 $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_338 N_A_27_112#_c_394_n N_A_363_82#_c_478_n 0.0230359f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_339 N_A_27_112#_c_395_n N_A_363_82#_c_478_n 0.00105459f $X=2.65 $Y=1.635
+ $X2=0 $Y2=0
cc_340 N_A_27_112#_M1004_g N_A_363_82#_c_479_n 0.0124182f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_341 N_A_27_112#_c_394_n N_A_363_82#_c_479_n 0.0250055f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_342 N_A_27_112#_c_395_n N_A_363_82#_c_479_n 0.00147052f $X=2.65 $Y=1.635
+ $X2=0 $Y2=0
cc_343 N_A_27_112#_c_400_n N_A_363_82#_c_480_n 0.0133618f $X=2.485 $Y=2.445
+ $X2=0 $Y2=0
cc_344 N_A_27_112#_c_395_n N_A_363_82#_c_480_n 0.00961468f $X=2.65 $Y=1.635
+ $X2=0 $Y2=0
cc_345 N_A_27_112#_M1010_g N_A_363_82#_c_488_n 0.0014421f $X=2.755 $Y=2.46 $X2=0
+ $Y2=0
cc_346 N_A_27_112#_M1010_g N_A_363_82#_c_491_n 2.27089e-19 $X=2.755 $Y=2.46
+ $X2=0 $Y2=0
cc_347 N_A_27_112#_c_400_n N_A_363_82#_c_491_n 0.0258418f $X=2.485 $Y=2.445
+ $X2=0 $Y2=0
cc_348 N_A_27_112#_c_394_n N_A_363_82#_c_491_n 0.0133851f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_349 N_A_27_112#_M1004_g N_A_363_82#_c_481_n 0.00977096f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_350 N_A_27_112#_c_394_n N_A_363_82#_c_481_n 0.066144f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_351 N_A_27_112#_c_395_n N_A_363_82#_c_482_n 0.0376213f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_352 N_A_27_112#_M1004_g N_A_363_82#_c_483_n 0.0376213f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_353 N_A_27_112#_M1004_g N_A_641_80#_c_779_n 8.37329e-19 $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_354 N_A_27_112#_c_400_n N_VPWR_M1000_d 0.0134589f $X=2.485 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_27_112#_c_400_n N_VPWR_M1001_d 0.00898525f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_356 N_A_27_112#_c_394_n N_VPWR_M1001_d 0.00461397f $X=2.65 $Y=1.635 $X2=0
+ $Y2=0
cc_357 N_A_27_112#_c_400_n N_VPWR_c_962_n 0.025956f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_358 N_A_27_112#_c_401_n N_VPWR_c_962_n 0.00464231f $X=0.445 $Y=2.445 $X2=0
+ $Y2=0
cc_359 N_A_27_112#_M1010_g N_VPWR_c_963_n 0.00907098f $X=2.755 $Y=2.46 $X2=0
+ $Y2=0
cc_360 N_A_27_112#_c_400_n N_VPWR_c_963_n 0.0252777f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_361 N_A_27_112#_M1010_g N_VPWR_c_974_n 0.00460063f $X=2.755 $Y=2.46 $X2=0
+ $Y2=0
cc_362 N_A_27_112#_c_401_n N_VPWR_c_977_n 0.00961497f $X=0.445 $Y=2.445 $X2=0
+ $Y2=0
cc_363 N_A_27_112#_M1010_g N_VPWR_c_961_n 0.00571695f $X=2.755 $Y=2.46 $X2=0
+ $Y2=0
cc_364 N_A_27_112#_c_400_n N_VPWR_c_961_n 0.0601041f $X=2.485 $Y=2.445 $X2=0
+ $Y2=0
cc_365 N_A_27_112#_c_401_n N_VPWR_c_961_n 0.0119199f $X=0.445 $Y=2.445 $X2=0
+ $Y2=0
cc_366 N_A_27_112#_c_393_n N_VGND_c_1160_n 0.0177942f $X=0.265 $Y=0.95 $X2=0
+ $Y2=0
cc_367 N_A_27_112#_M1004_g N_VGND_c_1167_n 0.00142194f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_368 N_A_27_112#_M1004_g N_VGND_c_1168_n 0.00347067f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_369 N_A_27_112#_c_393_n N_VGND_c_1174_n 0.00885135f $X=0.265 $Y=0.95 $X2=0
+ $Y2=0
cc_370 N_A_27_112#_M1004_g N_VGND_c_1179_n 0.00414706f $X=2.77 $Y=0.72 $X2=0
+ $Y2=0
cc_371 N_A_27_112#_c_393_n N_VGND_c_1179_n 0.0115776f $X=0.265 $Y=0.95 $X2=0
+ $Y2=0
cc_372 N_A_363_82#_M1020_g N_A_821_98#_M1007_g 0.0137938f $X=3.71 $Y=2.75 $X2=0
+ $Y2=0
cc_373 N_A_363_82#_c_487_n N_A_821_98#_M1007_g 0.00177596f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_374 N_A_363_82#_c_489_n N_A_821_98#_M1007_g 0.00917517f $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_375 N_A_363_82#_c_490_n N_A_821_98#_M1007_g 0.00343718f $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_376 N_A_363_82#_c_489_n N_A_821_98#_c_616_n 0.0181165f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_377 N_A_363_82#_c_490_n N_A_821_98#_c_616_n 9.76153e-19 $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_378 N_A_363_82#_c_489_n N_A_821_98#_c_617_n 3.39771e-19 $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_379 N_A_363_82#_c_490_n N_A_821_98#_c_617_n 0.0172854f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_380 N_A_363_82#_c_487_n N_A_641_80#_M1014_d 0.00473638f $X=3.705 $Y=2.99
+ $X2=0 $Y2=0
cc_381 N_A_363_82#_c_481_n N_A_641_80#_c_779_n 0.0138103f $X=3.18 $Y=1.215 $X2=0
+ $Y2=0
cc_382 N_A_363_82#_c_482_n N_A_641_80#_c_779_n 0.00107163f $X=3.22 $Y=1.315
+ $X2=0 $Y2=0
cc_383 N_A_363_82#_c_483_n N_A_641_80#_c_779_n 0.00686671f $X=3.22 $Y=1.15 $X2=0
+ $Y2=0
cc_384 N_A_363_82#_c_480_n N_A_641_80#_c_774_n 0.0361307f $X=3.06 $Y=2.905 $X2=0
+ $Y2=0
cc_385 N_A_363_82#_c_487_n N_A_641_80#_c_774_n 0.0123303f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_386 N_A_363_82#_c_489_n N_A_641_80#_c_774_n 0.0414419f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_387 N_A_363_82#_c_490_n N_A_641_80#_c_774_n 0.00550019f $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_388 N_A_363_82#_c_480_n N_A_641_80#_c_767_n 0.00677684f $X=3.06 $Y=2.905
+ $X2=0 $Y2=0
cc_389 N_A_363_82#_c_481_n N_A_641_80#_c_767_n 0.0251828f $X=3.18 $Y=1.215 $X2=0
+ $Y2=0
cc_390 N_A_363_82#_c_482_n N_A_641_80#_c_767_n 0.00224196f $X=3.22 $Y=1.315
+ $X2=0 $Y2=0
cc_391 N_A_363_82#_c_483_n N_A_641_80#_c_767_n 0.00309916f $X=3.22 $Y=1.15 $X2=0
+ $Y2=0
cc_392 N_A_363_82#_c_490_n N_A_641_80#_c_768_n 0.00111766f $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_393 N_A_363_82#_c_480_n N_A_641_80#_c_769_n 0.0131205f $X=3.06 $Y=2.905 $X2=0
+ $Y2=0
cc_394 N_A_363_82#_c_489_n N_A_641_80#_c_769_n 0.0201952f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_395 N_A_363_82#_c_490_n N_A_641_80#_c_769_n 8.29613e-19 $X=3.87 $Y=2.215
+ $X2=0 $Y2=0
cc_396 N_A_363_82#_c_481_n N_A_641_80#_c_769_n 0.00523479f $X=3.18 $Y=1.215
+ $X2=0 $Y2=0
cc_397 N_A_363_82#_c_482_n N_A_641_80#_c_769_n 2.01687e-19 $X=3.22 $Y=1.315
+ $X2=0 $Y2=0
cc_398 N_A_363_82#_c_480_n N_VPWR_c_963_n 0.0103728f $X=3.06 $Y=2.905 $X2=0
+ $Y2=0
cc_399 N_A_363_82#_c_488_n N_VPWR_c_963_n 0.00984682f $X=3.145 $Y=2.99 $X2=0
+ $Y2=0
cc_400 N_A_363_82#_M1020_g N_VPWR_c_974_n 0.00333833f $X=3.71 $Y=2.75 $X2=0
+ $Y2=0
cc_401 N_A_363_82#_c_487_n N_VPWR_c_974_n 0.0587151f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_402 N_A_363_82#_c_488_n N_VPWR_c_974_n 0.011907f $X=3.145 $Y=2.99 $X2=0 $Y2=0
cc_403 N_A_363_82#_M1020_g N_VPWR_c_979_n 4.05858e-19 $X=3.71 $Y=2.75 $X2=0
+ $Y2=0
cc_404 N_A_363_82#_c_487_n N_VPWR_c_979_n 0.00796896f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_405 N_A_363_82#_c_489_n N_VPWR_c_979_n 0.0109521f $X=3.87 $Y=2.215 $X2=0
+ $Y2=0
cc_406 N_A_363_82#_M1020_g N_VPWR_c_961_n 0.00425285f $X=3.71 $Y=2.75 $X2=0
+ $Y2=0
cc_407 N_A_363_82#_c_487_n N_VPWR_c_961_n 0.0325052f $X=3.705 $Y=2.99 $X2=0
+ $Y2=0
cc_408 N_A_363_82#_c_488_n N_VPWR_c_961_n 0.0063247f $X=3.145 $Y=2.99 $X2=0
+ $Y2=0
cc_409 N_A_363_82#_c_480_n A_569_392# 0.00869394f $X=3.06 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_410 N_A_363_82#_c_488_n A_569_392# 5.7967e-19 $X=3.145 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_411 N_A_363_82#_c_487_n A_760_508# 8.66307e-19 $X=3.705 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_412 N_A_363_82#_c_489_n A_760_508# 0.00564058f $X=3.87 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_413 N_A_363_82#_c_479_n N_VGND_M1002_d 0.00306155f $X=2.975 $Y=1.215 $X2=0
+ $Y2=0
cc_414 N_A_363_82#_c_483_n N_VGND_c_1168_n 9.29978e-19 $X=3.22 $Y=1.15 $X2=0
+ $Y2=0
cc_415 N_A_821_98#_M1007_g N_A_641_80#_M1027_g 0.0152228f $X=4.365 $Y=2.75 $X2=0
+ $Y2=0
cc_416 N_A_821_98#_c_616_n N_A_641_80#_M1027_g 0.0131759f $X=5.095 $Y=2.155
+ $X2=0 $Y2=0
cc_417 N_A_821_98#_c_617_n N_A_641_80#_M1027_g 0.00737988f $X=4.41 $Y=2.155
+ $X2=0 $Y2=0
cc_418 N_A_821_98#_c_618_n N_A_641_80#_M1027_g 3.04814e-19 $X=5.4 $Y=2.4 $X2=0
+ $Y2=0
cc_419 N_A_821_98#_c_621_n N_A_641_80#_M1027_g 0.0235234f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_420 N_A_821_98#_c_610_n N_A_641_80#_M1027_g 8.86568e-19 $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_421 N_A_821_98#_c_611_n N_A_641_80#_M1027_g 0.00559257f $X=4.41 $Y=1.99 $X2=0
+ $Y2=0
cc_422 N_A_821_98#_c_605_n N_A_641_80#_M1016_g 0.00506044f $X=4.32 $Y=1.19 $X2=0
+ $Y2=0
cc_423 N_A_821_98#_c_607_n N_A_641_80#_M1016_g 0.0120602f $X=4.955 $Y=0.515
+ $X2=0 $Y2=0
cc_424 N_A_821_98#_c_609_n N_A_641_80#_M1016_g 0.00418289f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_425 N_A_821_98#_c_610_n N_A_641_80#_M1016_g 0.0114535f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_426 N_A_821_98#_c_616_n N_A_641_80#_c_765_n 0.00452694f $X=5.095 $Y=2.155
+ $X2=0 $Y2=0
cc_427 N_A_821_98#_c_609_n N_A_641_80#_c_765_n 0.00842608f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_428 N_A_821_98#_c_611_n N_A_641_80#_c_765_n 0.0223372f $X=4.41 $Y=1.99 $X2=0
+ $Y2=0
cc_429 N_A_821_98#_c_610_n N_A_641_80#_c_766_n 0.0105381f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_430 N_A_821_98#_c_596_n N_A_641_80#_c_779_n 4.80093e-19 $X=4.18 $Y=1.115
+ $X2=0 $Y2=0
cc_431 N_A_821_98#_c_596_n N_A_641_80#_c_767_n 0.00135697f $X=4.18 $Y=1.115
+ $X2=0 $Y2=0
cc_432 N_A_821_98#_c_611_n N_A_641_80#_c_767_n 0.00180539f $X=4.41 $Y=1.99 $X2=0
+ $Y2=0
cc_433 N_A_821_98#_c_605_n N_A_641_80#_c_768_n 0.00449484f $X=4.32 $Y=1.19 $X2=0
+ $Y2=0
cc_434 N_A_821_98#_c_616_n N_A_641_80#_c_768_n 0.0266186f $X=5.095 $Y=2.155
+ $X2=0 $Y2=0
cc_435 N_A_821_98#_c_617_n N_A_641_80#_c_768_n 0.00427209f $X=4.41 $Y=2.155
+ $X2=0 $Y2=0
cc_436 N_A_821_98#_c_611_n N_A_641_80#_c_768_n 0.0129419f $X=4.41 $Y=1.99 $X2=0
+ $Y2=0
cc_437 N_A_821_98#_c_616_n N_A_641_80#_c_770_n 0.027116f $X=5.095 $Y=2.155 $X2=0
+ $Y2=0
cc_438 N_A_821_98#_c_609_n N_A_641_80#_c_770_n 0.00950973f $X=5.027 $Y=1.13
+ $X2=0 $Y2=0
cc_439 N_A_821_98#_c_610_n N_A_641_80#_c_770_n 0.034555f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_440 N_A_821_98#_c_611_n N_A_641_80#_c_770_n 0.00226185f $X=4.41 $Y=1.99 $X2=0
+ $Y2=0
cc_441 N_A_821_98#_M1021_g N_RESET_B_M1026_g 0.0138422f $X=6.155 $Y=2.4 $X2=0
+ $Y2=0
cc_442 N_A_821_98#_c_602_n N_RESET_B_M1026_g 0.00291797f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_443 N_A_821_98#_c_618_n N_RESET_B_M1026_g 0.008244f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_444 N_A_821_98#_c_619_n N_RESET_B_M1026_g 0.013393f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_445 N_A_821_98#_c_608_n N_RESET_B_M1026_g 0.00349399f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_446 N_A_821_98#_c_621_n N_RESET_B_M1026_g 0.00979138f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_447 N_A_821_98#_c_610_n N_RESET_B_M1026_g 0.00318065f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_448 N_A_821_98#_M1024_g N_RESET_B_c_851_n 0.0178261f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_449 N_A_821_98#_c_619_n N_RESET_B_c_851_n 0.00156944f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_450 N_A_821_98#_c_608_n N_RESET_B_c_851_n 7.51785e-19 $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_451 N_A_821_98#_c_621_n N_RESET_B_c_851_n 0.00206086f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_452 N_A_821_98#_c_610_n N_RESET_B_c_851_n 9.18528e-19 $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_453 N_A_821_98#_M1024_g N_RESET_B_c_852_n 0.00141176f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_454 N_A_821_98#_c_602_n N_RESET_B_c_852_n 2.72691e-19 $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_455 N_A_821_98#_c_619_n N_RESET_B_c_852_n 0.0161187f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_456 N_A_821_98#_c_608_n N_RESET_B_c_852_n 0.0188908f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_457 N_A_821_98#_c_621_n N_RESET_B_c_852_n 0.010918f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_458 N_A_821_98#_c_610_n N_RESET_B_c_852_n 0.0294391f $X=5.33 $Y=1.72 $X2=0
+ $Y2=0
cc_459 N_A_821_98#_M1024_g N_RESET_B_c_853_n 0.0158216f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_460 N_A_821_98#_c_607_n N_RESET_B_c_853_n 0.00349897f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_461 N_A_821_98#_M1012_g N_A_1449_368#_M1005_g 0.00965813f $X=7.615 $Y=2.34
+ $X2=0 $Y2=0
cc_462 N_A_821_98#_M1006_g N_A_1449_368#_M1011_g 0.0200925f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_463 N_A_821_98#_M1025_g N_A_1449_368#_c_894_n 0.00494994f $X=6.53 $Y=0.74
+ $X2=0 $Y2=0
cc_464 N_A_821_98#_M1006_g N_A_1449_368#_c_894_n 0.005981f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_465 N_A_821_98#_M1006_g N_A_1449_368#_c_895_n 0.00655853f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_466 N_A_821_98#_M1022_g N_A_1449_368#_c_896_n 0.00629436f $X=6.605 $Y=2.4
+ $X2=0 $Y2=0
cc_467 N_A_821_98#_M1012_g N_A_1449_368#_c_896_n 0.0205493f $X=7.615 $Y=2.34
+ $X2=0 $Y2=0
cc_468 N_A_821_98#_c_606_n N_A_1449_368#_c_897_n 0.0211541f $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_469 N_A_821_98#_M1006_g N_A_1449_368#_c_898_n 0.00231106f $X=7.625 $Y=0.79
+ $X2=0 $Y2=0
cc_470 N_A_821_98#_c_601_n N_A_1449_368#_c_912_n 0.023405f $X=7.525 $Y=1.465
+ $X2=0 $Y2=0
cc_471 N_A_821_98#_c_606_n N_A_1449_368#_c_912_n 9.32228e-19 $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_472 N_A_821_98#_c_606_n N_A_1449_368#_c_899_n 0.0216214f $X=7.615 $Y=1.465
+ $X2=0 $Y2=0
cc_473 N_A_821_98#_c_616_n N_VPWR_M1007_d 0.00613881f $X=5.095 $Y=2.155 $X2=0
+ $Y2=0
cc_474 N_A_821_98#_c_619_n N_VPWR_M1026_d 0.00206187f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_475 N_A_821_98#_c_608_n N_VPWR_M1026_d 6.9418e-19 $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_476 N_A_821_98#_M1021_g N_VPWR_c_964_n 0.0020069f $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A_821_98#_c_619_n N_VPWR_c_964_n 0.0148886f $X=5.955 $Y=1.805 $X2=0
+ $Y2=0
cc_478 N_A_821_98#_c_608_n N_VPWR_c_964_n 0.00463957f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_479 N_A_821_98#_c_621_n N_VPWR_c_964_n 0.0358158f $X=5.33 $Y=1.805 $X2=0
+ $Y2=0
cc_480 N_A_821_98#_M1021_g N_VPWR_c_965_n 5.92659e-19 $X=6.155 $Y=2.4 $X2=0
+ $Y2=0
cc_481 N_A_821_98#_M1022_g N_VPWR_c_965_n 0.0181408f $X=6.605 $Y=2.4 $X2=0 $Y2=0
cc_482 N_A_821_98#_c_601_n N_VPWR_c_965_n 6.85105e-19 $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_483 N_A_821_98#_M1012_g N_VPWR_c_965_n 0.00426005f $X=7.615 $Y=2.34 $X2=0
+ $Y2=0
cc_484 N_A_821_98#_M1012_g N_VPWR_c_966_n 0.00365f $X=7.615 $Y=2.34 $X2=0 $Y2=0
cc_485 N_A_821_98#_c_618_n N_VPWR_c_969_n 0.014549f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_486 N_A_821_98#_M1021_g N_VPWR_c_971_n 0.00552356f $X=6.155 $Y=2.4 $X2=0
+ $Y2=0
cc_487 N_A_821_98#_M1022_g N_VPWR_c_971_n 0.00460063f $X=6.605 $Y=2.4 $X2=0
+ $Y2=0
cc_488 N_A_821_98#_M1007_g N_VPWR_c_974_n 0.00461464f $X=4.365 $Y=2.75 $X2=0
+ $Y2=0
cc_489 N_A_821_98#_M1012_g N_VPWR_c_975_n 0.00567889f $X=7.615 $Y=2.34 $X2=0
+ $Y2=0
cc_490 N_A_821_98#_M1007_g N_VPWR_c_979_n 0.0170354f $X=4.365 $Y=2.75 $X2=0
+ $Y2=0
cc_491 N_A_821_98#_c_616_n N_VPWR_c_979_n 0.0284872f $X=5.095 $Y=2.155 $X2=0
+ $Y2=0
cc_492 N_A_821_98#_c_617_n N_VPWR_c_979_n 0.00230817f $X=4.41 $Y=2.155 $X2=0
+ $Y2=0
cc_493 N_A_821_98#_c_618_n N_VPWR_c_979_n 0.0144922f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_494 N_A_821_98#_M1007_g N_VPWR_c_961_n 0.00910297f $X=4.365 $Y=2.75 $X2=0
+ $Y2=0
cc_495 N_A_821_98#_M1021_g N_VPWR_c_961_n 0.0108836f $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_496 N_A_821_98#_M1022_g N_VPWR_c_961_n 0.00908554f $X=6.605 $Y=2.4 $X2=0
+ $Y2=0
cc_497 N_A_821_98#_M1012_g N_VPWR_c_961_n 0.00610055f $X=7.615 $Y=2.34 $X2=0
+ $Y2=0
cc_498 N_A_821_98#_c_618_n N_VPWR_c_961_n 0.0119743f $X=5.4 $Y=2.4 $X2=0 $Y2=0
cc_499 N_A_821_98#_M1024_g N_Q_c_1076_n 0.00802514f $X=6.1 $Y=0.74 $X2=0 $Y2=0
cc_500 N_A_821_98#_M1025_g N_Q_c_1076_n 0.0131993f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A_821_98#_M1021_g N_Q_c_1080_n 3.70642e-19 $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_502 N_A_821_98#_M1022_g N_Q_c_1080_n 3.62369e-19 $X=6.605 $Y=2.4 $X2=0 $Y2=0
cc_503 N_A_821_98#_M1022_g N_Q_c_1081_n 0.0168943f $X=6.605 $Y=2.4 $X2=0 $Y2=0
cc_504 N_A_821_98#_c_601_n N_Q_c_1081_n 0.00163358f $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_505 N_A_821_98#_M1012_g N_Q_c_1081_n 4.08485e-19 $X=7.615 $Y=2.34 $X2=0 $Y2=0
cc_506 N_A_821_98#_c_726_p N_Q_c_1081_n 0.0133617f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_507 N_A_821_98#_M1021_g N_Q_c_1082_n 3.24225e-19 $X=6.155 $Y=2.4 $X2=0 $Y2=0
cc_508 N_A_821_98#_c_602_n N_Q_c_1082_n 0.00233326f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_509 N_A_821_98#_c_608_n N_Q_c_1082_n 0.00488278f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_510 N_A_821_98#_c_726_p N_Q_c_1082_n 0.0143383f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_511 N_A_821_98#_M1025_g N_Q_c_1077_n 0.0128805f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_512 N_A_821_98#_c_601_n N_Q_c_1077_n 0.00442505f $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_513 N_A_821_98#_M1006_g N_Q_c_1077_n 3.42629e-19 $X=7.625 $Y=0.79 $X2=0 $Y2=0
cc_514 N_A_821_98#_c_726_p N_Q_c_1077_n 0.0122755f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_515 N_A_821_98#_M1024_g N_Q_c_1078_n 0.00374068f $X=6.1 $Y=0.74 $X2=0 $Y2=0
cc_516 N_A_821_98#_M1025_g N_Q_c_1078_n 9.7541e-19 $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_517 N_A_821_98#_c_602_n N_Q_c_1078_n 0.00260566f $X=6.695 $Y=1.465 $X2=0
+ $Y2=0
cc_518 N_A_821_98#_c_726_p N_Q_c_1078_n 0.0276081f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_519 N_A_821_98#_M1025_g Q 0.00556303f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A_821_98#_M1022_g Q 0.00625258f $X=6.605 $Y=2.4 $X2=0 $Y2=0
cc_521 N_A_821_98#_c_601_n Q 0.0259674f $X=7.525 $Y=1.465 $X2=0 $Y2=0
cc_522 N_A_821_98#_M1012_g Q 6.63467e-19 $X=7.615 $Y=2.34 $X2=0 $Y2=0
cc_523 N_A_821_98#_M1006_g Q 6.46089e-19 $X=7.625 $Y=0.79 $X2=0 $Y2=0
cc_524 N_A_821_98#_c_726_p Q 0.0223699f $X=6.53 $Y=1.465 $X2=0 $Y2=0
cc_525 N_A_821_98#_c_596_n N_VGND_c_1161_n 0.0144666f $X=4.18 $Y=1.115 $X2=0
+ $Y2=0
cc_526 N_A_821_98#_c_605_n N_VGND_c_1161_n 0.00540622f $X=4.32 $Y=1.19 $X2=0
+ $Y2=0
cc_527 N_A_821_98#_c_607_n N_VGND_c_1161_n 0.0491859f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_528 N_A_821_98#_M1024_g N_VGND_c_1162_n 0.00889628f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_529 N_A_821_98#_c_607_n N_VGND_c_1162_n 0.0145513f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_530 N_A_821_98#_M1025_g N_VGND_c_1163_n 0.013225f $X=6.53 $Y=0.74 $X2=0 $Y2=0
cc_531 N_A_821_98#_c_601_n N_VGND_c_1163_n 7.73684e-19 $X=7.525 $Y=1.465 $X2=0
+ $Y2=0
cc_532 N_A_821_98#_M1006_g N_VGND_c_1163_n 0.00336635f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_533 N_A_821_98#_M1006_g N_VGND_c_1164_n 0.0074703f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_534 N_A_821_98#_c_596_n N_VGND_c_1168_n 0.00347405f $X=4.18 $Y=1.115 $X2=0
+ $Y2=0
cc_535 N_A_821_98#_c_607_n N_VGND_c_1170_n 0.0206573f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_536 N_A_821_98#_M1024_g N_VGND_c_1172_n 0.00434272f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_537 N_A_821_98#_M1025_g N_VGND_c_1172_n 0.00434272f $X=6.53 $Y=0.74 $X2=0
+ $Y2=0
cc_538 N_A_821_98#_M1006_g N_VGND_c_1175_n 0.00485498f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_539 N_A_821_98#_c_596_n N_VGND_c_1179_n 0.00395485f $X=4.18 $Y=1.115 $X2=0
+ $Y2=0
cc_540 N_A_821_98#_M1024_g N_VGND_c_1179_n 0.00821985f $X=6.1 $Y=0.74 $X2=0
+ $Y2=0
cc_541 N_A_821_98#_M1025_g N_VGND_c_1179_n 0.00825059f $X=6.53 $Y=0.74 $X2=0
+ $Y2=0
cc_542 N_A_821_98#_M1006_g N_VGND_c_1179_n 0.00514438f $X=7.625 $Y=0.79 $X2=0
+ $Y2=0
cc_543 N_A_821_98#_c_607_n N_VGND_c_1179_n 0.016746f $X=4.955 $Y=0.515 $X2=0
+ $Y2=0
cc_544 N_A_641_80#_c_766_n N_RESET_B_M1026_g 0.0170261f $X=5.035 $Y=1.35 $X2=0
+ $Y2=0
cc_545 N_A_641_80#_M1016_g N_RESET_B_c_851_n 0.0181352f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_A_641_80#_c_766_n N_RESET_B_c_851_n 0.00276431f $X=5.035 $Y=1.35 $X2=0
+ $Y2=0
cc_547 N_A_641_80#_M1016_g N_RESET_B_c_852_n 0.00101423f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_548 N_A_641_80#_M1016_g N_RESET_B_c_853_n 0.0496133f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_549 N_A_641_80#_M1027_g N_VPWR_c_969_n 0.00461464f $X=5.125 $Y=2.4 $X2=0
+ $Y2=0
cc_550 N_A_641_80#_M1027_g N_VPWR_c_979_n 0.0156218f $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_551 N_A_641_80#_M1027_g N_VPWR_c_961_n 0.00909121f $X=5.125 $Y=2.4 $X2=0
+ $Y2=0
cc_552 N_A_641_80#_M1016_g N_VGND_c_1161_n 0.00414178f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_553 N_A_641_80#_c_779_n N_VGND_c_1161_n 0.00562511f $X=3.57 $Y=0.875 $X2=0
+ $Y2=0
cc_554 N_A_641_80#_c_767_n N_VGND_c_1161_n 0.00300042f $X=3.655 $Y=1.65 $X2=0
+ $Y2=0
cc_555 N_A_641_80#_c_768_n N_VGND_c_1161_n 0.0109219f $X=4.605 $Y=1.735 $X2=0
+ $Y2=0
cc_556 N_A_641_80#_M1016_g N_VGND_c_1162_n 0.00125099f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_557 N_A_641_80#_M1016_g N_VGND_c_1170_n 0.00291513f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_558 N_A_641_80#_M1016_g N_VGND_c_1179_n 0.00363725f $X=5.17 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_RESET_B_M1026_g N_VPWR_c_964_n 0.00200449f $X=5.625 $Y=2.4 $X2=0 $Y2=0
cc_560 N_RESET_B_M1026_g N_VPWR_c_969_n 0.005209f $X=5.625 $Y=2.4 $X2=0 $Y2=0
cc_561 N_RESET_B_M1026_g N_VPWR_c_979_n 4.25103e-19 $X=5.625 $Y=2.4 $X2=0 $Y2=0
cc_562 N_RESET_B_M1026_g N_VPWR_c_961_n 0.00982981f $X=5.625 $Y=2.4 $X2=0 $Y2=0
cc_563 N_RESET_B_c_853_n N_Q_c_1078_n 3.46348e-19 $X=5.62 $Y=1.22 $X2=0 $Y2=0
cc_564 N_RESET_B_c_851_n N_VGND_c_1162_n 9.00259e-19 $X=5.62 $Y=1.385 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_852_n N_VGND_c_1162_n 0.0124443f $X=5.62 $Y=1.385 $X2=0 $Y2=0
cc_566 N_RESET_B_c_853_n N_VGND_c_1162_n 0.0136038f $X=5.62 $Y=1.22 $X2=0 $Y2=0
cc_567 N_RESET_B_c_853_n N_VGND_c_1170_n 0.00383152f $X=5.62 $Y=1.22 $X2=0 $Y2=0
cc_568 N_RESET_B_c_853_n N_VGND_c_1179_n 0.0075725f $X=5.62 $Y=1.22 $X2=0 $Y2=0
cc_569 N_A_1449_368#_c_896_n N_VPWR_c_965_n 0.0444755f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_570 N_A_1449_368#_M1005_g N_VPWR_c_966_n 0.00580407f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_571 N_A_1449_368#_c_896_n N_VPWR_c_966_n 0.0402324f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_572 N_A_1449_368#_c_897_n N_VPWR_c_966_n 0.026236f $X=8.08 $Y=1.465 $X2=0
+ $Y2=0
cc_573 N_A_1449_368#_c_899_n N_VPWR_c_966_n 0.00320573f $X=8.625 $Y=1.465 $X2=0
+ $Y2=0
cc_574 N_A_1449_368#_M1008_g N_VPWR_c_968_n 0.00647357f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_575 N_A_1449_368#_c_896_n N_VPWR_c_975_n 0.00915997f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_A_1449_368#_M1005_g N_VPWR_c_976_n 0.005209f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_577 N_A_1449_368#_M1008_g N_VPWR_c_976_n 0.0048691f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_578 N_A_1449_368#_M1005_g N_VPWR_c_961_n 0.00986727f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_579 N_A_1449_368#_M1008_g N_VPWR_c_961_n 0.00875947f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_580 N_A_1449_368#_c_896_n N_VPWR_c_961_n 0.0104921f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_581 N_A_1449_368#_c_896_n N_Q_c_1081_n 0.0147753f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_582 N_A_1449_368#_c_894_n N_Q_c_1077_n 0.0149965f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_583 N_A_1449_368#_c_895_n Q 0.0135906f $X=7.4 $Y=1.3 $X2=0 $Y2=0
cc_584 N_A_1449_368#_c_896_n Q 0.0136317f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_585 N_A_1449_368#_c_912_n Q 0.0256724f $X=7.4 $Y=1.465 $X2=0 $Y2=0
cc_586 N_A_1449_368#_M1011_g N_Q_N_c_1129_n 0.00746865f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_587 N_A_1449_368#_M1019_g N_Q_N_c_1129_n 0.0081896f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_588 N_A_1449_368#_M1011_g N_Q_N_c_1130_n 0.00322812f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_589 N_A_1449_368#_M1019_g N_Q_N_c_1130_n 0.00215589f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_590 N_A_1449_368#_c_899_n N_Q_N_c_1130_n 0.00244427f $X=8.625 $Y=1.465 $X2=0
+ $Y2=0
cc_591 N_A_1449_368#_M1005_g Q_N 0.00307491f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_592 N_A_1449_368#_M1008_g Q_N 0.00270934f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_593 N_A_1449_368#_c_897_n Q_N 0.00138666f $X=8.08 $Y=1.465 $X2=0 $Y2=0
cc_594 N_A_1449_368#_c_899_n Q_N 0.00310238f $X=8.625 $Y=1.465 $X2=0 $Y2=0
cc_595 N_A_1449_368#_M1005_g Q_N 0.0122016f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_596 N_A_1449_368#_M1008_g Q_N 0.0149161f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_597 N_A_1449_368#_M1005_g N_Q_N_c_1131_n 0.00293165f $X=8.165 $Y=2.4 $X2=0
+ $Y2=0
cc_598 N_A_1449_368#_M1011_g N_Q_N_c_1131_n 0.0025553f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_599 N_A_1449_368#_M1008_g N_Q_N_c_1131_n 0.00994275f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_600 N_A_1449_368#_M1019_g N_Q_N_c_1131_n 0.00866774f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_601 N_A_1449_368#_c_897_n N_Q_N_c_1131_n 0.0249855f $X=8.08 $Y=1.465 $X2=0
+ $Y2=0
cc_602 N_A_1449_368#_c_899_n N_Q_N_c_1131_n 0.0238138f $X=8.625 $Y=1.465 $X2=0
+ $Y2=0
cc_603 N_A_1449_368#_c_894_n N_VGND_c_1163_n 0.0207909f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_604 N_A_1449_368#_M1011_g N_VGND_c_1164_n 0.0093706f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_605 N_A_1449_368#_c_894_n N_VGND_c_1164_n 0.0270587f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_606 N_A_1449_368#_c_897_n N_VGND_c_1164_n 0.028359f $X=8.08 $Y=1.465 $X2=0
+ $Y2=0
cc_607 N_A_1449_368#_c_899_n N_VGND_c_1164_n 0.00370401f $X=8.625 $Y=1.465 $X2=0
+ $Y2=0
cc_608 N_A_1449_368#_M1019_g N_VGND_c_1166_n 0.00646793f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_609 N_A_1449_368#_c_894_n N_VGND_c_1175_n 0.0103491f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_610 N_A_1449_368#_M1011_g N_VGND_c_1176_n 0.00434272f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_611 N_A_1449_368#_M1019_g N_VGND_c_1176_n 0.00422942f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_612 N_A_1449_368#_M1011_g N_VGND_c_1179_n 0.00825059f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_613 N_A_1449_368#_M1019_g N_VGND_c_1179_n 0.00787255f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_614 N_A_1449_368#_c_894_n N_VGND_c_1179_n 0.0113354f $X=7.41 $Y=0.615 $X2=0
+ $Y2=0
cc_615 N_VPWR_c_964_n N_Q_c_1080_n 0.0315118f $X=5.9 $Y=2.145 $X2=0 $Y2=0
cc_616 N_VPWR_c_965_n N_Q_c_1080_n 0.0283117f $X=6.83 $Y=2.305 $X2=0 $Y2=0
cc_617 N_VPWR_c_971_n N_Q_c_1080_n 0.00749631f $X=6.665 $Y=3.33 $X2=0 $Y2=0
cc_618 N_VPWR_c_961_n N_Q_c_1080_n 0.0062048f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_619 N_VPWR_M1022_s N_Q_c_1081_n 0.00313614f $X=6.695 $Y=1.84 $X2=0 $Y2=0
cc_620 N_VPWR_c_965_n N_Q_c_1081_n 0.0231981f $X=6.83 $Y=2.305 $X2=0 $Y2=0
cc_621 N_VPWR_c_966_n Q_N 0.0456524f $X=7.89 $Y=1.985 $X2=0 $Y2=0
cc_622 N_VPWR_c_968_n Q_N 0.0455874f $X=8.84 $Y=1.985 $X2=0 $Y2=0
cc_623 N_VPWR_c_976_n Q_N 0.0157112f $X=8.755 $Y=3.33 $X2=0 $Y2=0
cc_624 N_VPWR_c_961_n Q_N 0.0127977f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_625 N_Q_c_1077_n N_VGND_M1025_s 0.00464869f $X=6.845 $Y=1.045 $X2=0 $Y2=0
cc_626 N_Q_c_1076_n N_VGND_c_1162_n 0.0402483f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_627 N_Q_c_1078_n N_VGND_c_1162_n 0.00349775f $X=6.48 $Y=1.045 $X2=0 $Y2=0
cc_628 N_Q_c_1076_n N_VGND_c_1163_n 0.0173003f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_629 N_Q_c_1077_n N_VGND_c_1163_n 0.027001f $X=6.845 $Y=1.045 $X2=0 $Y2=0
cc_630 N_Q_c_1076_n N_VGND_c_1172_n 0.0144922f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_631 N_Q_c_1076_n N_VGND_c_1179_n 0.0118826f $X=6.315 $Y=0.515 $X2=0 $Y2=0
cc_632 N_Q_N_c_1129_n N_VGND_c_1164_n 0.0309448f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_633 N_Q_N_c_1129_n N_VGND_c_1166_n 0.0308798f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_634 N_Q_N_c_1129_n N_VGND_c_1176_n 0.0149085f $X=8.41 $Y=0.515 $X2=0 $Y2=0
cc_635 N_Q_N_c_1129_n N_VGND_c_1179_n 0.0122037f $X=8.41 $Y=0.515 $X2=0 $Y2=0

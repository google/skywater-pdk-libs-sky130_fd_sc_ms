* File: sky130_fd_sc_ms__o21bai_2.pxi.spice
* Created: Wed Sep  2 12:22:36 2020
* 
x_PM_SKY130_FD_SC_MS__O21BAI_2%B1_N N_B1_N_M1011_g N_B1_N_M1000_g B1_N
+ N_B1_N_c_81_n N_B1_N_c_82_n PM_SKY130_FD_SC_MS__O21BAI_2%B1_N
x_PM_SKY130_FD_SC_MS__O21BAI_2%A_27_74# N_A_27_74#_M1011_s N_A_27_74#_M1000_s
+ N_A_27_74#_M1008_g N_A_27_74#_c_114_n N_A_27_74#_M1007_g N_A_27_74#_M1009_g
+ N_A_27_74#_c_116_n N_A_27_74#_M1013_g N_A_27_74#_c_117_n N_A_27_74#_c_118_n
+ N_A_27_74#_c_119_n N_A_27_74#_c_126_n N_A_27_74#_c_120_n N_A_27_74#_c_121_n
+ N_A_27_74#_c_122_n N_A_27_74#_c_127_n N_A_27_74#_c_123_n
+ PM_SKY130_FD_SC_MS__O21BAI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O21BAI_2%A1 N_A1_M1004_g N_A1_M1001_g N_A1_M1012_g
+ N_A1_M1006_g N_A1_c_202_n N_A1_c_203_n N_A1_c_220_p N_A1_c_217_n A1
+ N_A1_c_204_n N_A1_c_205_n A1 PM_SKY130_FD_SC_MS__O21BAI_2%A1
x_PM_SKY130_FD_SC_MS__O21BAI_2%A2 N_A2_M1002_g N_A2_M1005_g N_A2_M1003_g
+ N_A2_M1010_g A2 N_A2_c_286_n N_A2_c_287_n PM_SKY130_FD_SC_MS__O21BAI_2%A2
x_PM_SKY130_FD_SC_MS__O21BAI_2%VPWR N_VPWR_M1000_d N_VPWR_M1009_s N_VPWR_M1012_s
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n VPWR
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n
+ N_VPWR_c_339_n PM_SKY130_FD_SC_MS__O21BAI_2%VPWR
x_PM_SKY130_FD_SC_MS__O21BAI_2%Y N_Y_M1007_s N_Y_M1008_d N_Y_M1002_d N_Y_c_397_n
+ N_Y_c_395_n N_Y_c_403_n N_Y_c_433_p N_Y_c_404_n Y Y Y Y
+ PM_SKY130_FD_SC_MS__O21BAI_2%Y
x_PM_SKY130_FD_SC_MS__O21BAI_2%A_510_368# N_A_510_368#_M1001_d
+ N_A_510_368#_M1003_s N_A_510_368#_c_438_n N_A_510_368#_c_444_n
+ N_A_510_368#_c_439_n PM_SKY130_FD_SC_MS__O21BAI_2%A_510_368#
x_PM_SKY130_FD_SC_MS__O21BAI_2%VGND N_VGND_M1011_d N_VGND_M1004_s N_VGND_M1010_s
+ N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n VGND N_VGND_c_468_n
+ N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n
+ N_VGND_c_474_n N_VGND_c_475_n PM_SKY130_FD_SC_MS__O21BAI_2%VGND
x_PM_SKY130_FD_SC_MS__O21BAI_2%A_225_74# N_A_225_74#_M1007_d N_A_225_74#_M1013_d
+ N_A_225_74#_M1005_d N_A_225_74#_M1006_d N_A_225_74#_c_519_n
+ N_A_225_74#_c_520_n N_A_225_74#_c_521_n N_A_225_74#_c_540_n
+ N_A_225_74#_c_522_n N_A_225_74#_c_523_n N_A_225_74#_c_524_n
+ N_A_225_74#_c_525_n N_A_225_74#_c_526_n N_A_225_74#_c_527_n
+ PM_SKY130_FD_SC_MS__O21BAI_2%A_225_74#
cc_1 VNB N_B1_N_M1011_g 0.0392908f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_B1_N_c_81_n 0.00536388f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_3 VNB N_B1_N_c_82_n 0.0306368f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.515
cc_4 VNB N_A_27_74#_M1008_g 0.00662559f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_5 VNB N_A_27_74#_c_114_n 0.0184105f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_6 VNB N_A_27_74#_M1009_g 0.00663413f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.515
cc_7 VNB N_A_27_74#_c_116_n 0.016529f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.515
cc_8 VNB N_A_27_74#_c_117_n 0.0396459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_118_n 0.0344881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_119_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_120_n 0.0243345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_121_n 0.00511234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_122_n 0.0109678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_123_n 0.022547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1004_g 0.025715f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_16 VNB N_A1_M1012_g 7.72232e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_17 VNB N_A1_M1006_g 0.030416f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_18 VNB N_A1_c_202_n 0.00166985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_203_n 0.0270502f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.665
cc_20 VNB N_A1_c_204_n 0.0346418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_205_n 0.0191473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A1 8.32086e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1005_g 0.024925f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.34
cc_24 VNB N_A2_M1010_g 0.0230333f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_25 VNB N_A2_c_286_n 0.00138642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_287_n 0.036618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_339_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_395_n 4.51115e-19 $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.515
cc_29 VNB Y 0.00224001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_465_n 0.0107462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_466_n 0.00842841f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.515
cc_32 VNB N_VGND_c_467_n 0.00327765f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.665
cc_33 VNB N_VGND_c_468_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_469_n 0.0405043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_470_n 0.0162351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_471_n 0.0180274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_472_n 0.262471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_473_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_474_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_475_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_225_74#_c_519_n 0.00379275f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_42 VNB N_A_225_74#_c_520_n 0.00452721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_225_74#_c_521_n 0.00417961f $X=-0.19 $Y=-0.245 $X2=0.647 $Y2=1.515
cc_44 VNB N_A_225_74#_c_522_n 0.00968069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_225_74#_c_523_n 0.0100176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_225_74#_c_524_n 0.00179461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_225_74#_c_525_n 0.015761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_225_74#_c_526_n 0.0255089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_225_74#_c_527_n 0.00193677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_B1_N_M1000_g 0.0282787f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.34
cc_51 VPB N_B1_N_c_81_n 0.00578639f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.515
cc_52 VPB N_B1_N_c_82_n 0.0071055f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.515
cc_53 VPB N_A_27_74#_M1008_g 0.0245385f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_54 VPB N_A_27_74#_M1009_g 0.022286f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.515
cc_55 VPB N_A_27_74#_c_126_n 0.0356507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_74#_c_127_n 0.0137373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_74#_c_123_n 0.0143228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A1_M1001_g 0.0207467f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.34
cc_59 VPB N_A1_M1012_g 0.0281549f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_60 VPB N_A1_c_202_n 0.00269395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A1_c_203_n 0.00564567f $X=-0.19 $Y=1.66 $X2=0.647 $Y2=1.665
cc_62 VPB A1 0.00323722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A2_M1002_g 0.0203281f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.69
cc_64 VPB N_A2_M1003_g 0.0207479f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_65 VPB N_A2_c_286_n 0.00284416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A2_c_287_n 0.00466114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_340_n 0.0155971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_341_n 0.00579614f $X=-0.19 $Y=1.66 $X2=0.647 $Y2=1.515
cc_69 VPB N_VPWR_c_342_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.647 $Y2=1.665
cc_70 VPB N_VPWR_c_343_n 0.0576944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_344_n 0.030897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_345_n 0.0183662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_346_n 0.0388892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_347_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_348_n 0.00689346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_339_n 0.0760481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_Y_c_397_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_510_368#_c_438_n 0.00392434f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.34
cc_79 VPB N_A_510_368#_c_439_n 0.00195131f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.515
cc_80 N_B1_N_c_81_n N_A_27_74#_M1008_g 0.00401955f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B1_N_c_82_n N_A_27_74#_M1008_g 0.0178034f $X=0.7 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B1_N_M1011_g N_A_27_74#_c_117_n 0.0040089f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_83 N_B1_N_c_81_n N_A_27_74#_c_117_n 0.00135338f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_84 N_B1_N_c_82_n N_A_27_74#_c_117_n 0.0111951f $X=0.7 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B1_N_M1011_g N_A_27_74#_c_119_n 4.43891e-19 $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_86 N_B1_N_M1000_g N_A_27_74#_c_126_n 0.0116287f $X=0.7 $Y=2.34 $X2=0 $Y2=0
cc_87 N_B1_N_M1011_g N_A_27_74#_c_120_n 0.0189149f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_88 N_B1_N_c_81_n N_A_27_74#_c_120_n 0.0285306f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B1_N_c_82_n N_A_27_74#_c_120_n 0.00153394f $X=0.7 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B1_N_M1011_g N_A_27_74#_c_121_n 0.00179141f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_91 N_B1_N_c_81_n N_A_27_74#_c_121_n 0.014429f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B1_N_c_82_n N_A_27_74#_c_121_n 2.33686e-19 $X=0.7 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B1_N_M1000_g N_A_27_74#_c_127_n 0.00479039f $X=0.7 $Y=2.34 $X2=0 $Y2=0
cc_94 N_B1_N_c_81_n N_A_27_74#_c_127_n 0.0129929f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_95 N_B1_N_c_82_n N_A_27_74#_c_127_n 0.00254876f $X=0.7 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B1_N_M1011_g N_A_27_74#_c_123_n 0.0139236f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_97 N_B1_N_M1000_g N_A_27_74#_c_123_n 0.00386959f $X=0.7 $Y=2.34 $X2=0 $Y2=0
cc_98 N_B1_N_c_81_n N_A_27_74#_c_123_n 0.0323502f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_99 N_B1_N_M1000_g N_VPWR_c_340_n 0.0157737f $X=0.7 $Y=2.34 $X2=0 $Y2=0
cc_100 N_B1_N_M1000_g N_VPWR_c_344_n 0.00567889f $X=0.7 $Y=2.34 $X2=0 $Y2=0
cc_101 N_B1_N_M1000_g N_VPWR_c_339_n 0.00610055f $X=0.7 $Y=2.34 $X2=0 $Y2=0
cc_102 N_B1_N_M1011_g N_VGND_c_465_n 0.0156976f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_103 N_B1_N_M1011_g N_VGND_c_468_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_104 N_B1_N_M1011_g N_VGND_c_472_n 0.00761198f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_105 N_B1_N_M1011_g N_A_225_74#_c_519_n 8.38994e-19 $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_106 N_B1_N_M1011_g N_A_225_74#_c_521_n 7.24903e-19 $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_107 N_A_27_74#_c_116_n N_A1_M1004_g 0.0238637f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A_27_74#_M1009_g N_A1_M1001_g 0.0386604f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_27_74#_M1009_g N_A1_c_202_n 0.00227635f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_118_n N_A1_c_202_n 0.0013665f $X=1.915 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_118_n N_A1_c_203_n 0.0177085f $X=1.915 $Y=1.385 $X2=0 $Y2=0
cc_112 N_A_27_74#_M1009_g N_A1_c_217_n 0.00159214f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_27_74#_M1008_g N_VPWR_c_340_n 0.0131925f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_27_74#_c_117_n N_VPWR_c_340_n 0.00226699f $X=1.38 $Y=1.385 $X2=0
+ $Y2=0
cc_115 N_A_27_74#_c_120_n N_VPWR_c_340_n 7.87179e-19 $X=1.03 $Y=1.095 $X2=0
+ $Y2=0
cc_116 N_A_27_74#_c_121_n N_VPWR_c_340_n 0.0187766f $X=1.195 $Y=1.385 $X2=0
+ $Y2=0
cc_117 N_A_27_74#_c_127_n N_VPWR_c_340_n 0.0406188f $X=0.475 $Y=2.035 $X2=0
+ $Y2=0
cc_118 N_A_27_74#_M1008_g N_VPWR_c_341_n 4.45232e-19 $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_27_74#_M1009_g N_VPWR_c_341_n 0.00880347f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_126_n N_VPWR_c_344_n 0.0156062f $X=0.475 $Y=2.715 $X2=0
+ $Y2=0
cc_121 N_A_27_74#_M1008_g N_VPWR_c_345_n 0.005209f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_27_74#_M1009_g N_VPWR_c_345_n 0.00460063f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_27_74#_M1008_g N_VPWR_c_339_n 0.00987287f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_27_74#_M1009_g N_VPWR_c_339_n 0.00908554f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_27_74#_c_126_n N_VPWR_c_339_n 0.0178368f $X=0.475 $Y=2.715 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_M1008_g N_Y_c_397_n 0.00710505f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_27_74#_M1009_g N_Y_c_397_n 2.60789e-19 $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_27_74#_c_114_n N_Y_c_395_n 0.00107507f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_116_n N_Y_c_395_n 0.00779056f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_27_74#_c_120_n N_Y_c_395_n 0.00446815f $X=1.03 $Y=1.095 $X2=0 $Y2=0
cc_131 N_A_27_74#_M1009_g N_Y_c_403_n 0.0163663f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_27_74#_M1008_g N_Y_c_404_n 0.00211414f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_27_74#_M1009_g N_Y_c_404_n 0.00218557f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A_27_74#_M1008_g Y 0.0213544f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_27_74#_c_114_n Y 0.00240384f $X=1.485 $Y=1.22 $X2=0 $Y2=0
cc_136 N_A_27_74#_M1009_g Y 0.0172218f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_27_74#_c_116_n Y 0.0012234f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_138 N_A_27_74#_c_118_n Y 0.0235171f $X=1.915 $Y=1.385 $X2=0 $Y2=0
cc_139 N_A_27_74#_c_121_n Y 0.0278451f $X=1.195 $Y=1.385 $X2=0 $Y2=0
cc_140 N_A_27_74#_c_114_n N_VGND_c_465_n 0.00184366f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_141 N_A_27_74#_c_119_n N_VGND_c_465_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_120_n N_VGND_c_465_n 0.0243991f $X=1.03 $Y=1.095 $X2=0 $Y2=0
cc_143 N_A_27_74#_c_119_n N_VGND_c_468_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_144 N_A_27_74#_c_114_n N_VGND_c_469_n 0.00278247f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_145 N_A_27_74#_c_116_n N_VGND_c_469_n 0.00278271f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_146 N_A_27_74#_c_114_n N_VGND_c_472_n 0.00358425f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_147 N_A_27_74#_c_116_n N_VGND_c_472_n 0.0035414f $X=1.915 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A_27_74#_c_119_n N_VGND_c_472_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_c_120_n N_A_225_74#_M1007_d 0.00281428f $X=1.03 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_150 N_A_27_74#_c_114_n N_A_225_74#_c_519_n 0.00809982f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_151 N_A_27_74#_c_116_n N_A_225_74#_c_519_n 5.5293e-19 $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_152 N_A_27_74#_c_117_n N_A_225_74#_c_519_n 0.00120271f $X=1.38 $Y=1.385 $X2=0
+ $Y2=0
cc_153 N_A_27_74#_c_120_n N_A_225_74#_c_519_n 0.0217145f $X=1.03 $Y=1.095 $X2=0
+ $Y2=0
cc_154 N_A_27_74#_c_114_n N_A_225_74#_c_520_n 0.0100711f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_155 N_A_27_74#_c_116_n N_A_225_74#_c_520_n 0.0133867f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_156 N_A_27_74#_c_114_n N_A_225_74#_c_521_n 0.00395315f $X=1.485 $Y=1.22 $X2=0
+ $Y2=0
cc_157 N_A_27_74#_c_116_n N_A_225_74#_c_523_n 0.00116009f $X=1.915 $Y=1.22 $X2=0
+ $Y2=0
cc_158 N_A1_M1001_g N_A2_M1002_g 0.0506622f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A1_c_202_n N_A2_M1002_g 0.00220334f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A1_c_220_p N_A2_M1002_g 0.0115514f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_161 N_A1_M1004_g N_A2_M1005_g 0.0254412f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A1_c_220_p N_A2_M1003_g 0.0214565f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_163 N_A1_M1006_g N_A2_M1010_g 0.0314638f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_c_204_n N_A2_M1010_g 0.0221478f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_165 N_A1_c_205_n N_A2_M1010_g 0.0043055f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_166 N_A1_c_202_n N_A2_c_286_n 0.0253277f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A1_c_203_n N_A2_c_286_n 0.00121367f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A1_c_220_p N_A2_c_286_n 0.0290075f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_169 N_A1_c_204_n N_A2_c_286_n 2.15819e-19 $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_170 N_A1_c_205_n N_A2_c_286_n 0.0189163f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_171 A1 N_A2_c_286_n 0.00805575f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_172 N_A1_M1012_g N_A2_c_287_n 0.0221478f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_c_202_n N_A2_c_287_n 0.00137425f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A1_c_203_n N_A2_c_287_n 0.0179603f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_175 N_A1_c_220_p N_A2_c_287_n 4.88468e-19 $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_176 A1 N_A2_c_287_n 0.00323361f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_177 N_A1_c_202_n N_VPWR_M1009_s 0.00134673f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A1_c_217_n N_VPWR_M1009_s 0.00283555f $X=2.58 $Y=2.035 $X2=0 $Y2=0
cc_179 N_A1_M1001_g N_VPWR_c_341_n 0.00332485f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A1_M1012_g N_VPWR_c_343_n 0.00478817f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A1_c_204_n N_VPWR_c_343_n 0.00230627f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_182 N_A1_c_205_n N_VPWR_c_343_n 0.008349f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_183 A1 N_VPWR_c_343_n 0.00118327f $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_184 N_A1_M1001_g N_VPWR_c_346_n 0.00518311f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_M1012_g N_VPWR_c_346_n 0.00517089f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1001_g N_VPWR_c_339_n 0.00981524f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1012_g N_VPWR_c_339_n 0.00981377f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_c_220_p N_Y_M1002_d 0.00314031f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_189 N_A1_M1001_g N_Y_c_403_n 0.0164405f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A1_c_203_n N_Y_c_403_n 2.85826e-19 $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A1_c_220_p N_Y_c_403_n 0.0357287f $X=3.485 $Y=2.035 $X2=0 $Y2=0
cc_192 N_A1_c_217_n N_Y_c_403_n 0.0187923f $X=2.58 $Y=2.035 $X2=0 $Y2=0
cc_193 N_A1_M1004_g Y 7.96105e-19 $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1001_g Y 0.00118541f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A1_c_202_n Y 0.0242551f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A1_c_203_n Y 9.77722e-19 $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_197 N_A1_c_217_n Y 0.00748773f $X=2.58 $Y=2.035 $X2=0 $Y2=0
cc_198 N_A1_c_220_p N_A_510_368#_M1001_d 0.00761462f $X=3.485 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A1_c_220_p N_A_510_368#_M1003_s 0.00209824f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_200 A1 N_A_510_368#_M1003_s 2.29261e-19 $X=3.6 $Y=1.665 $X2=0 $Y2=0
cc_201 N_A1_M1012_g N_A_510_368#_c_438_n 0.00360372f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A1_M1012_g N_A_510_368#_c_444_n 0.00911188f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A1_c_220_p N_A_510_368#_c_444_n 0.0162961f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_204 N_A1_c_205_n N_A_510_368#_c_444_n 9.50316e-19 $X=3.89 $Y=1.485 $X2=0
+ $Y2=0
cc_205 N_A1_M1001_g N_A_510_368#_c_439_n 0.00705822f $X=2.46 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A1_M1004_g N_VGND_c_466_n 0.00404801f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A1_M1006_g N_VGND_c_467_n 0.0129724f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1004_g N_VGND_c_469_n 0.00430908f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A1_M1006_g N_VGND_c_471_n 0.00383152f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A1_M1004_g N_VGND_c_472_n 0.00817122f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A1_M1006_g N_VGND_c_472_n 0.00761264f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A1_M1004_g N_A_225_74#_c_520_n 0.00347348f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A1_M1004_g N_A_225_74#_c_540_n 0.00831216f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_M1004_g N_A_225_74#_c_522_n 0.0116199f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A1_c_202_n N_A_225_74#_c_522_n 0.0166004f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A1_c_203_n N_A_225_74#_c_522_n 6.21754e-19 $X=2.415 $Y=1.515 $X2=0
+ $Y2=0
cc_217 N_A1_M1004_g N_A_225_74#_c_523_n 0.00158144f $X=2.415 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_c_202_n N_A_225_74#_c_523_n 0.010051f $X=2.415 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A1_c_203_n N_A_225_74#_c_523_n 7.04412e-19 $X=2.415 $Y=1.515 $X2=0
+ $Y2=0
cc_220 N_A1_M1006_g N_A_225_74#_c_525_n 0.012998f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_c_204_n N_A_225_74#_c_525_n 0.00425672f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_222 N_A1_c_205_n N_A_225_74#_c_525_n 0.0443322f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_223 N_A1_M1006_g N_A_225_74#_c_526_n 0.00159319f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A2_M1002_g N_VPWR_c_346_n 0.00335119f $X=2.91 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A2_M1003_g N_VPWR_c_346_n 0.00333896f $X=3.36 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A2_M1002_g N_VPWR_c_339_n 0.00421887f $X=2.91 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A2_M1003_g N_VPWR_c_339_n 0.00422843f $X=3.36 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A2_M1002_g N_Y_c_403_n 0.0112423f $X=2.91 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A2_M1002_g N_A_510_368#_c_438_n 0.00904673f $X=2.91 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A2_M1003_g N_A_510_368#_c_438_n 0.0135711f $X=3.36 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A2_M1002_g N_A_510_368#_c_444_n 6.46121e-19 $X=2.91 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A2_M1003_g N_A_510_368#_c_444_n 0.00948577f $X=3.36 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A2_M1002_g N_A_510_368#_c_439_n 0.00730021f $X=2.91 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A2_M1003_g N_A_510_368#_c_439_n 6.05623e-19 $X=3.36 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A2_M1005_g N_VGND_c_466_n 0.00261709f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A2_M1005_g N_VGND_c_467_n 4.66963e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A2_M1010_g N_VGND_c_467_n 0.00999938f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A2_M1005_g N_VGND_c_470_n 0.00461464f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A2_M1010_g N_VGND_c_470_n 0.00383152f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_M1005_g N_VGND_c_472_n 0.00908164f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1010_g N_VGND_c_472_n 0.0075754f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1005_g N_A_225_74#_c_540_n 8.0819e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A2_M1005_g N_A_225_74#_c_522_n 0.0142114f $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_c_286_n N_A_225_74#_c_522_n 0.0189798f $X=3.03 $Y=1.515 $X2=0 $Y2=0
cc_245 N_A2_c_287_n N_A_225_74#_c_522_n 3.40811e-19 $X=3.375 $Y=1.515 $X2=0
+ $Y2=0
cc_246 N_A2_M1005_g N_A_225_74#_c_524_n 4.00651e-19 $X=2.945 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A2_M1010_g N_A_225_74#_c_524_n 3.92313e-19 $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1010_g N_A_225_74#_c_525_n 0.0172653f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1010_g N_A_225_74#_c_527_n 9.49306e-19 $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_c_286_n N_A_225_74#_c_527_n 0.0137234f $X=3.03 $Y=1.515 $X2=0 $Y2=0
cc_251 N_A2_c_287_n N_A_225_74#_c_527_n 7.88639e-19 $X=3.375 $Y=1.515 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_340_n N_Y_c_397_n 0.0174388f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_253 N_VPWR_c_341_n N_Y_c_397_n 0.01174f $X=2.165 $Y=2.815 $X2=0 $Y2=0
cc_254 N_VPWR_c_345_n N_Y_c_397_n 0.0109793f $X=1.98 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_339_n N_Y_c_397_n 0.00901959f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_M1009_s N_Y_c_403_n 0.0103282f $X=2.01 $Y=1.84 $X2=0 $Y2=0
cc_257 N_VPWR_c_341_n N_Y_c_403_n 0.0204006f $X=2.165 $Y=2.815 $X2=0 $Y2=0
cc_258 N_VPWR_c_340_n Y 0.016521f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_259 N_VPWR_c_343_n N_A_510_368#_c_438_n 0.0103534f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_346_n N_A_510_368#_c_438_n 0.0595904f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_339_n N_A_510_368#_c_438_n 0.0328069f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_341_n N_A_510_368#_c_439_n 0.0207727f $X=2.165 $Y=2.815 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_346_n N_A_510_368#_c_439_n 0.0225565f $X=3.955 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_339_n N_A_510_368#_c_439_n 0.0123454f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_343_n N_A_225_74#_c_525_n 0.00464454f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_Y_c_403_n N_A_510_368#_M1001_d 0.00332066f $X=3.05 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_267 N_Y_M1002_d N_A_510_368#_c_438_n 0.00165831f $X=3 $Y=1.84 $X2=0 $Y2=0
cc_268 N_Y_c_403_n N_A_510_368#_c_438_n 0.00464895f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_269 N_Y_c_433_p N_A_510_368#_c_438_n 0.0114967f $X=3.135 $Y=2.46 $X2=0 $Y2=0
cc_270 N_Y_c_403_n N_A_510_368#_c_439_n 0.0164176f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_271 N_Y_M1007_s N_A_225_74#_c_520_n 0.00184993f $X=1.56 $Y=0.37 $X2=0 $Y2=0
cc_272 N_Y_c_395_n N_A_225_74#_c_520_n 0.0129924f $X=1.7 $Y=0.8 $X2=0 $Y2=0
cc_273 N_Y_c_395_n N_A_225_74#_c_523_n 0.00932276f $X=1.7 $Y=0.8 $X2=0 $Y2=0
cc_274 N_VGND_c_465_n N_A_225_74#_c_519_n 0.027945f $X=0.71 $Y=0.675 $X2=0 $Y2=0
cc_275 N_VGND_c_466_n N_A_225_74#_c_520_n 0.011924f $X=2.7 $Y=0.675 $X2=0 $Y2=0
cc_276 N_VGND_c_469_n N_A_225_74#_c_520_n 0.0613638f $X=2.535 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_472_n N_A_225_74#_c_520_n 0.034015f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_465_n N_A_225_74#_c_521_n 0.0121616f $X=0.71 $Y=0.675 $X2=0
+ $Y2=0
cc_279 N_VGND_c_469_n N_A_225_74#_c_521_n 0.0233048f $X=2.535 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_472_n N_A_225_74#_c_521_n 0.0126653f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_281 N_VGND_M1004_s N_A_225_74#_c_522_n 0.00293722f $X=2.49 $Y=0.37 $X2=0
+ $Y2=0
cc_282 N_VGND_c_466_n N_A_225_74#_c_522_n 0.0216414f $X=2.7 $Y=0.675 $X2=0 $Y2=0
cc_283 N_VGND_c_466_n N_A_225_74#_c_524_n 0.00129758f $X=2.7 $Y=0.675 $X2=0
+ $Y2=0
cc_284 N_VGND_c_467_n N_A_225_74#_c_524_n 0.0171736f $X=3.59 $Y=0.645 $X2=0
+ $Y2=0
cc_285 N_VGND_c_470_n N_A_225_74#_c_524_n 0.00749631f $X=3.425 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_472_n N_A_225_74#_c_524_n 0.0062048f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_M1010_s N_A_225_74#_c_525_n 0.00176461f $X=3.45 $Y=0.37 $X2=0
+ $Y2=0
cc_288 N_VGND_c_467_n N_A_225_74#_c_525_n 0.0170777f $X=3.59 $Y=0.645 $X2=0
+ $Y2=0
cc_289 N_VGND_c_467_n N_A_225_74#_c_526_n 0.017215f $X=3.59 $Y=0.645 $X2=0 $Y2=0
cc_290 N_VGND_c_471_n N_A_225_74#_c_526_n 0.011066f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_c_472_n N_A_225_74#_c_526_n 0.00915947f $X=4.08 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__fah_1.spice
* Created: Wed Sep  2 12:09:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fah_1.pex.spice"
.subckt sky130_fd_sc_ms__fah_1  VNB VPB CI B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* CI	CI
* VPB	VPB
* VNB	VNB
MM1026 N_VGND_M1026_d N_A_83_21#_M1026_g N_SUM_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.206342 AS=0.2072 PD=1.51217 PS=2.04 NRD=36.288 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1012 N_A_231_132#_M1012_d N_CI_M1012_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.2016 AS=0.178458 PD=1.91 PS=1.30783 NRD=2.808 NRS=41.964 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_A_410_58#_M1008_g N_COUT_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.313857 AS=0.2072 PD=1.72667 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1025 N_A_644_104#_M1025_d N_A_231_132#_M1025_g N_VGND_M1008_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.23505 AS=0.271443 PD=2.02 PS=1.49333 NRD=14.988 NRS=111.552
+ M=1 R=4.26667 SA=75001.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1001 N_A_410_58#_M1001_d N_A_811_379#_M1001_g N_A_879_55#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.131975 AS=0.28315 PD=1.205 PS=3.17 NRD=0 NRS=72.636 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1016 N_A_231_132#_M1016_d N_A_1023_379#_M1016_g N_A_410_58#_M1001_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.131975 PD=0.92 PS=1.205 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75000.5 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_A_83_21#_M1002_d N_A_811_379#_M1002_g N_A_231_132#_M1016_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.11875 AS=0.0896 PD=1.08 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_644_104#_M1020_d N_A_1023_379#_M1020_g N_A_83_21#_M1002_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.11875 PD=1.85 PS=1.08 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_B_M1023_g N_A_879_55#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3136 AS=0.2109 PD=2.51 PS=2.05 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1006 N_A_1023_379#_M1006_d N_A_879_55#_M1006_g N_A_1660_374#_M1006_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.24825 AS=0.2568 PD=1.49 PS=2.17 NRD=62.412
+ NRS=15.936 M=1 R=4.26667 SA=75000.3 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1027 N_A_1852_374#_M1027_d N_B_M1027_g N_A_1023_379#_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1524 AS=0.24825 PD=1.16 PS=1.49 NRD=15.936 NRS=62.412 M=1
+ R=4.26667 SA=75001 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1004 N_A_811_379#_M1004_d N_A_879_55#_M1004_g N_A_1852_374#_M1027_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.3264 AS=0.1524 PD=1.66 PS=1.16 NRD=61.872 NRS=15.936 M=1
+ R=4.26667 SA=75001.6 SB=75002 A=0.096 P=1.58 MULT=1
MM1024 N_A_1660_374#_M1024_d N_B_M1024_g N_A_811_379#_M1004_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.12007 AS=0.3264 PD=1.02029 PS=1.66 NRD=15.468 NRS=76.872 M=1
+ R=4.26667 SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1022_d N_A_2342_48#_M1022_g N_A_1660_374#_M1024_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2875 AS=0.13883 PD=2.33 PS=1.17971 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75002.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_1852_374#_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.208 PD=1.02 PS=1.93 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1014 N_A_2342_48#_M1014_d N_A_M1014_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1216 PD=1.85 PS=1.02 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VPWR_M1015_d N_A_83_21#_M1015_g N_SUM_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.281426 AS=0.3136 PD=1.7117 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1000 N_A_231_132#_M1000_d N_CI_M1000_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.251274 PD=2.56 PS=1.5283 NRD=0 NRS=44.7978 M=1 R=5.55556
+ SA=90000.9 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_410_58#_M1007_g N_COUT_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.306164 AS=0.45085 PD=1.92302 PS=3.26 NRD=38.3953 NRS=14.9326 M=1
+ R=6.22222 SA=90000.3 SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1003 N_A_644_104#_M1003_d N_A_231_132#_M1003_g N_VPWR_M1007_d VPB PSHORT
+ L=0.18 W=1 AD=0.288655 AS=0.273361 PD=1.74457 PS=1.71698 NRD=15.7403
+ NRS=43.0051 M=1 R=5.55556 SA=90000.9 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1017 N_A_83_21#_M1017_d N_A_811_379#_M1017_g N_A_644_104#_M1003_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.3696 AS=0.24247 PD=1.72 PS=1.46543 NRD=0 NRS=54.7857 M=1
+ R=4.66667 SA=90001.5 SB=90003.1 A=0.1512 P=2.04 MULT=1
MM1028 N_A_231_132#_M1028_d N_A_1023_379#_M1028_g N_A_83_21#_M1017_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.394012 AS=0.3696 PD=1.98 PS=1.72 NRD=0 NRS=141.879 M=1
+ R=4.66667 SA=90002.6 SB=90002 A=0.1512 P=2.04 MULT=1
MM1010 N_A_410_58#_M1010_d N_A_811_379#_M1010_g N_A_231_132#_M1028_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2415 AS=0.394012 PD=1.415 PS=1.98 NRD=0 NRS=97.1013 M=1
+ R=4.66667 SA=90002.7 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1019 N_A_879_55#_M1019_d N_A_1023_379#_M1019_g N_A_410_58#_M1010_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.160371 AS=0.2415 PD=1.26429 PS=1.415 NRD=19.1484
+ NRS=70.3487 M=1 R=4.66667 SA=90003.4 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1021 N_VPWR_M1021_d N_B_M1021_g N_A_879_55#_M1019_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.213829 PD=2.9 PS=1.68571 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90003 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1013 N_A_811_379#_M1013_d N_A_879_55#_M1013_g N_A_1660_374#_M1013_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1344 AS=0.2352 PD=1.16 PS=2.24 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90003.4 A=0.1512 P=2.04 MULT=1
MM1011 N_A_1852_374#_M1011_d N_B_M1011_g N_A_811_379#_M1013_d VPB PSHORT L=0.18
+ W=0.84 AD=0.648075 AS=0.1344 PD=2.365 PS=1.16 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1005 N_A_1023_379#_M1005_d N_A_879_55#_M1005_g N_A_1852_374#_M1011_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.648075 PD=1.11 PS=2.365 NRD=0 NRS=71.511
+ M=1 R=4.66667 SA=90002.3 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1009 N_A_1660_374#_M1009_d N_B_M1009_g N_A_1023_379#_M1005_d VPB PSHORT L=0.18
+ W=0.84 AD=0.147 AS=0.1134 PD=1.23857 PS=1.11 NRD=4.6886 NRS=0 M=1 R=4.66667
+ SA=90002.8 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1029 N_VPWR_M1029_d N_A_2342_48#_M1029_g N_A_1660_374#_M1009_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.4683 AS=0.196 PD=3.28 PS=1.65143 NRD=15.2281 NRS=4.3931 M=1
+ R=6.22222 SA=90002.5 SB=90000.3 A=0.2016 P=2.6 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_1852_374#_M1030_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1031 N_A_2342_48#_M1031_d N_A_M1031_g N_VPWR_M1030_d VPB PSHORT L=0.18 W=1
+ AD=0.285 AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=26.8204 P=33.14
*
.include "sky130_fd_sc_ms__fah_1.pxi.spice"
*
.ends
*
*

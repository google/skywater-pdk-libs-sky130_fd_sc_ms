* File: sky130_fd_sc_ms__fahcon_1.pex.spice
* Created: Wed Sep  2 12:09:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A 3 6 8 11 13
r39 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.515
+ $X2=0.54 $Y2=1.68
r40 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.515
+ $X2=0.54 $Y2=1.35
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.515 $X2=0.54 $Y2=1.515
r42 8 12 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.54 $Y2=1.565
r43 6 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.545 $Y=2.4
+ $X2=0.545 $Y2=1.68
r44 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.87
+ $X2=0.495 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_27_100# 1 2 3 4 15 17 19 22 28 30 34 38
+ 39 40 45 47 48 49 51 52 55 56 60
c124 60 0 2.01518e-20 $X=1.365 $Y=1.515
c125 51 0 1.53129e-19 $X=2.565 $Y=1.97
c126 34 0 7.413e-20 $X=1.08 $Y=1.515
r127 59 60 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.365 $Y2=1.515
r128 55 56 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.81
+ $X2=2.61 $Y2=0.725
r129 51 52 5.26587 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.587 $Y=1.97
+ $X2=2.587 $Y2=1.805
r130 47 48 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=2.115
+ $X2=0.285 $Y2=1.95
r131 43 55 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.61 $Y=0.89 $X2=2.61
+ $Y2=0.81
r132 43 52 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=2.61 $Y=0.89
+ $X2=2.61 $Y2=1.805
r133 41 56 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.53 $Y=0.425
+ $X2=2.53 $Y2=0.725
r134 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=0.34
+ $X2=2.53 $Y2=0.425
r135 39 40 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=2.445 $Y=0.34
+ $X2=1.245 $Y2=0.34
r136 38 49 5.44924 $w=1.87e-07 $l=1.85e-07 $layer=LI1_cond $X=1.16 $Y=0.98
+ $X2=0.975 $Y2=0.98
r137 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.16 $Y=0.425
+ $X2=1.245 $Y2=0.34
r138 37 38 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.16 $Y=0.425
+ $X2=1.16 $Y2=0.98
r139 35 59 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.08 $Y=1.515
+ $X2=1.13 $Y2=1.515
r140 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.515 $X2=1.08 $Y2=1.515
r141 32 49 5.44924 $w=1.87e-07 $l=2.45764e-07 $layer=LI1_cond $X=1.077 $Y=1.18
+ $X2=0.975 $Y2=0.98
r142 32 34 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=1.077 $Y=1.18
+ $X2=1.077 $Y2=1.515
r143 31 45 1.76993 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.08
+ $X2=0.225 $Y2=1.08
r144 30 49 1.11122 $w=2e-07 $l=1e-07 $layer=LI1_cond $X=0.975 $Y=1.08 $X2=0.975
+ $Y2=0.98
r145 30 31 33.8273 $w=1.98e-07 $l=6.1e-07 $layer=LI1_cond $X=0.975 $Y=1.08
+ $X2=0.365 $Y2=1.08
r146 26 47 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=0.285 $Y=2.15
+ $X2=0.285 $Y2=2.115
r147 26 28 19.1594 $w=3.98e-07 $l=6.65e-07 $layer=LI1_cond $X=0.285 $Y=2.15
+ $X2=0.285 $Y2=2.815
r148 24 45 4.67858 $w=2.25e-07 $l=1.24499e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.225 $Y2=1.08
r149 24 48 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.17 $Y2=1.95
r150 20 45 4.67858 $w=2.25e-07 $l=1e-07 $layer=LI1_cond $X=0.225 $Y=0.98
+ $X2=0.225 $Y2=1.08
r151 20 22 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.225 $Y=0.98
+ $X2=0.225 $Y2=0.645
r152 17 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.365 $Y2=1.515
r153 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.365 $Y2=0.92
r154 13 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.68
+ $X2=1.13 $Y2=1.515
r155 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.13 $Y=1.68
+ $X2=1.13 $Y2=2.34
r156 4 51 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.825 $X2=2.565 $Y2=1.97
r157 3 47 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.115
r158 3 28 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r159 2 55 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.665 $X2=2.61 $Y2=0.81
r160 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.5 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_336_263# 1 2 9 14 15 16 19 24 26 28 29 35
+ 41 48 49
c105 49 0 9.91361e-20 $X=4.207 $Y=1.805
c106 41 0 1.41326e-19 $X=3.115 $Y=0.405
c107 26 0 7.413e-20 $X=1.775 $Y=1.465
c108 15 0 3.57245e-21 $X=2.75 $Y=0.22
r109 48 49 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=4.207 $Y=1.97
+ $X2=4.207 $Y2=1.805
r110 46 49 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.125 $Y=1.01
+ $X2=4.125 $Y2=1.805
r111 45 46 16.4522 $w=6.93e-07 $l=4.95e-07 $layer=LI1_cond $X=4.387 $Y=0.515
+ $X2=4.387 $Y2=1.01
r112 39 53 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.932 $Y=0.39
+ $X2=2.932 $Y2=0.555
r113 38 41 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=0.405
+ $X2=3.115 $Y2=0.405
r114 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=0.39 $X2=2.95 $Y2=0.39
r115 33 48 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=4.207 $Y=1.972
+ $X2=4.207 $Y2=1.97
r116 33 35 28.4843 $w=3.33e-07 $l=8.28e-07 $layer=LI1_cond $X=4.207 $Y=1.972
+ $X2=4.207 $Y2=2.8
r117 29 45 3.01171 $w=6.93e-07 $l=1.75e-07 $layer=LI1_cond $X=4.387 $Y=0.34
+ $X2=4.387 $Y2=0.515
r118 29 41 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.04 $Y=0.34
+ $X2=3.115 $Y2=0.34
r119 27 28 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.8 $Y=1.38 $X2=2.8
+ $Y2=1.53
r120 25 26 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.775 $Y=1.315
+ $X2=1.775 $Y2=1.465
r121 24 27 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.825 $Y=0.985
+ $X2=2.825 $Y2=1.38
r122 24 53 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.825 $Y=0.985
+ $X2=2.825 $Y2=0.555
r123 19 28 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=2.79 $Y=2.245
+ $X2=2.79 $Y2=1.53
r124 15 39 26.8759 $w=3.65e-07 $l=1.7e-07 $layer=POLY_cond $X=2.932 $Y=0.22
+ $X2=2.932 $Y2=0.39
r125 15 16 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.75 $Y=0.22
+ $X2=1.87 $Y2=0.22
r126 14 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.795 $Y=0.92
+ $X2=1.795 $Y2=1.315
r127 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.795 $Y=0.295
+ $X2=1.87 $Y2=0.22
r128 11 14 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.795 $Y=0.295
+ $X2=1.795 $Y2=0.92
r129 9 26 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=1.77 $Y=2.245
+ $X2=1.77 $Y2=1.465
r130 2 48 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.825 $X2=4.21 $Y2=1.97
r131 2 35 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=1.825 $X2=4.21 $Y2=2.8
r132 1 45 60.6667 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=3
+ $X=4.105 $Y=0.37 $X2=4.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%B 4 7 9 10 14 17 19 22 23 24 27 29 31 33 36
+ 40 43 45 46 47 48 53 54
c139 53 0 3.00527e-20 $X=4.9 $Y=1.385
c140 43 0 1.08015e-19 $X=2.355 $Y=1.615
c141 27 0 1.73957e-19 $X=4.435 $Y=2.385
c142 17 0 2.22531e-19 $X=3.43 $Y=0.985
c143 7 0 1.79307e-20 $X=2.385 $Y=0.985
r144 52 54 25.6578 $w=2.63e-07 $l=1.4e-07 $layer=POLY_cond $X=4.9 $Y=1.385
+ $X2=5.04 $Y2=1.385
r145 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.385 $X2=4.9 $Y2=1.385
r146 50 52 16.4943 $w=2.63e-07 $l=9e-08 $layer=POLY_cond $X=4.81 $Y=1.385
+ $X2=4.9 $Y2=1.385
r147 48 53 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.56 $Y=1.365 $X2=4.9
+ $Y2=1.365
r148 44 45 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.407 $Y=1.6
+ $X2=3.407 $Y2=1.75
r149 42 43 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.355 $Y=1.465
+ $X2=2.355 $Y2=1.615
r150 38 54 44.9011 $w=2.63e-07 $l=3.16938e-07 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.04 $Y2=1.385
r151 38 40 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.285 $Y2=0.69
r152 34 54 11.6845 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=1.385
r153 34 36 347.895 $w=1.8e-07 $l=8.95e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=2.445
r154 31 50 15.8942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.22
+ $X2=4.81 $Y2=1.385
r155 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.81 $Y=1.22
+ $X2=4.81 $Y2=0.74
r156 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.525 $Y=1.475
+ $X2=4.435 $Y2=1.475
r157 29 50 22.5691 $w=2.63e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.735 $Y=1.475
+ $X2=4.81 $Y2=1.385
r158 29 30 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.735 $Y=1.475
+ $X2=4.525 $Y2=1.475
r159 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.55
+ $X2=4.435 $Y2=1.475
r160 25 27 324.573 $w=1.8e-07 $l=8.35e-07 $layer=POLY_cond $X=4.435 $Y=1.55
+ $X2=4.435 $Y2=2.385
r161 23 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.345 $Y=1.475
+ $X2=4.435 $Y2=1.475
r162 23 24 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.345 $Y=1.475
+ $X2=3.99 $Y2=1.475
r163 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.915 $Y=1.55
+ $X2=3.99 $Y2=1.475
r164 21 22 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=3.915 $Y=1.55
+ $X2=3.915 $Y2=3.035
r165 20 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.49 $Y=3.11 $X2=3.4
+ $Y2=3.11
r166 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=3.11
+ $X2=3.915 $Y2=3.035
r167 19 20 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.84 $Y=3.11
+ $X2=3.49 $Y2=3.11
r168 17 44 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.43 $Y=0.985
+ $X2=3.43 $Y2=1.6
r169 14 45 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.4 $Y=2.245
+ $X2=3.4 $Y2=1.75
r170 12 46 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.4 $Y=3.035 $X2=3.4
+ $Y2=3.11
r171 12 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=3.4 $Y=3.035
+ $X2=3.4 $Y2=2.245
r172 9 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.31 $Y=3.11 $X2=3.4
+ $Y2=3.11
r173 9 10 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.31 $Y=3.11
+ $X2=2.43 $Y2=3.11
r174 7 42 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.385 $Y=0.985
+ $X2=2.385 $Y2=1.465
r175 4 43 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.34 $Y=2.245
+ $X2=2.34 $Y2=1.615
r176 2 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.34 $Y=3.035
+ $X2=2.43 $Y2=3.11
r177 2 4 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.34 $Y=3.035
+ $X2=2.34 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_374_120# 1 2 9 13 16 20 23 25 26 28 31 34
+ 36 37 43 46 48 50 55 56 57 59 60 61 62 63 64 71 74 76 81 87 97
c256 63 0 1.54021e-19 $X=9.215 $Y=0.925
c257 61 0 1.05698e-19 $X=6.815 $Y=0.925
c258 59 0 1.11588e-19 $X=5.855 $Y=0.925
c259 55 0 8.9203e-20 $X=9.58 $Y=1.425
c260 50 0 3.00527e-20 $X=5.702 $Y=1.475
c261 43 0 2.01518e-20 $X=2.01 $Y=1.745
c262 34 0 1.54205e-19 $X=6.977 $Y=1.287
c263 20 0 3.23497e-19 $X=9.5 $Y=2.26
c264 16 0 9.08104e-20 $X=9.455 $Y=0.79
r265 77 97 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=9.36 $Y=0.925
+ $X2=9.56 $Y2=0.925
r266 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0.925
+ $X2=9.36 $Y2=0.925
r267 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0.925
+ $X2=6.96 $Y2=0.925
r268 71 91 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6 $Y=0.925 $X2=5.75
+ $Y2=0.925
r269 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0.925 $X2=6
+ $Y2=0.925
r270 66 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.925
r271 64 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=0.925
+ $X2=6.96 $Y2=0.925
r272 63 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=9.36 $Y2=0.925
r273 63 64 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=7.105 $Y2=0.925
r274 62 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=0.925
+ $X2=6 $Y2=0.925
r275 61 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=0.925
+ $X2=6.96 $Y2=0.925
r276 61 62 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=6.815 $Y=0.925
+ $X2=6.145 $Y2=0.925
r277 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.925
+ $X2=2.16 $Y2=0.925
r278 59 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=6 $Y2=0.925
r279 59 60 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=2.305 $Y2=0.925
r280 56 85 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.562 $Y=1.425
+ $X2=9.562 $Y2=1.59
r281 56 84 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.562 $Y=1.425
+ $X2=9.562 $Y2=1.26
r282 55 57 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=9.582 $Y=1.425
+ $X2=9.582 $Y2=1.26
r283 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.58
+ $Y=1.425 $X2=9.58 $Y2=1.425
r284 53 74 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=6.947 $Y=1.13
+ $X2=6.947 $Y2=0.925
r285 49 81 26.3208 $w=2.93e-07 $l=1.6e-07 $layer=POLY_cond $X=5.735 $Y=1.64
+ $X2=5.575 $Y2=1.64
r286 48 50 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.702 $Y=1.64
+ $X2=5.702 $Y2=1.475
r287 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.735
+ $Y=1.64 $X2=5.735 $Y2=1.64
r288 45 87 12.8415 $w=3.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.1 $Y=1.15 $X2=2.1
+ $Y2=0.76
r289 45 46 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=2.1 $Y=1.15
+ $X2=2.1 $Y2=1.325
r290 41 43 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.775 $Y=1.745
+ $X2=2.01 $Y2=1.745
r291 39 97 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.56 $Y=1.04
+ $X2=9.56 $Y2=0.925
r292 39 57 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.56 $Y=1.04
+ $X2=9.56 $Y2=1.26
r293 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.985
+ $Y=1.295 $X2=6.985 $Y2=1.295
r294 34 53 6.1958 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=6.977 $Y=1.287
+ $X2=6.977 $Y2=1.13
r295 34 36 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=6.977 $Y=1.287
+ $X2=6.977 $Y2=1.295
r296 32 91 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.75 $Y=1.04
+ $X2=5.75 $Y2=0.925
r297 32 50 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.75 $Y=1.04
+ $X2=5.75 $Y2=1.475
r298 31 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=1.66
+ $X2=2.01 $Y2=1.745
r299 31 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.01 $Y=1.66
+ $X2=2.01 $Y2=1.325
r300 26 28 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.86 $Y=2.65
+ $X2=3.095 $Y2=2.65
r301 25 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.775 $Y=2.565
+ $X2=1.86 $Y2=2.65
r302 24 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=1.83
+ $X2=1.775 $Y2=1.745
r303 24 25 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.775 $Y=1.83
+ $X2=1.775 $Y2=2.565
r304 23 37 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.985 $Y=1.13
+ $X2=6.985 $Y2=1.295
r305 20 85 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=9.5 $Y=2.26 $X2=9.5
+ $Y2=1.59
r306 16 84 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=9.455 $Y=0.79 $X2=9.455
+ $Y2=1.26
r307 13 23 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.925 $Y=0.69
+ $X2=6.925 $Y2=1.13
r308 7 81 14.174 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.805
+ $X2=5.575 $Y2=1.64
r309 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.575 $Y=1.805
+ $X2=5.575 $Y2=2.525
r310 2 28 600 $w=1.7e-07 $l=9.26283e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.825 $X2=3.095 $Y2=2.65
r311 1 87 91 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.6 $X2=2.09 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_372_365# 1 2 9 13 17 19 23 25 28 33 34 35
+ 36 43 45 52 56 57 62
c168 57 0 6.54889e-20 $X=8.64 $Y=1.465
c169 56 0 1.54021e-19 $X=8.64 $Y=1.465
c170 23 0 1.11511e-19 $X=9.05 $Y=2.26
c171 19 0 8.9203e-20 $X=8.96 $Y=1.555
c172 9 0 1.54205e-19 $X=6.215 $Y=0.69
r173 56 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.64 $Y=1.465
+ $X2=8.64 $Y2=1.555
r174 56 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.64 $Y=1.465
+ $X2=8.64 $Y2=1.3
r175 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.64
+ $Y=1.465 $X2=8.64 $Y2=1.465
r176 50 52 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.23 $Y=1.715
+ $X2=6.445 $Y2=1.715
r177 48 50 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.215 $Y=1.715
+ $X2=6.23 $Y2=1.715
r178 46 57 7.95652 $w=3.68e-07 $l=2.95973e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.64 $Y2=1.54
r179 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.665
r180 43 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.445
+ $Y=1.715 $X2=6.445 $Y2=1.715
r181 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r182 39 62 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=0.81
r183 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r184 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.665
+ $X2=6.48 $Y2=1.665
r185 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=8.88 $Y2=1.665
r186 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=6.625 $Y2=1.665
r187 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r188 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r189 33 34 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=3.265 $Y2=1.665
r190 32 39 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.11 $Y=2.225
+ $X2=3.11 $Y2=1.665
r191 28 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.115 $Y=2.195
+ $X2=2.115 $Y2=2.31
r192 26 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.31
+ $X2=2.115 $Y2=2.31
r193 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.945 $Y=2.31
+ $X2=3.11 $Y2=2.225
r194 25 26 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.945 $Y=2.31
+ $X2=2.2 $Y2=2.31
r195 21 23 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=9.05 $Y=1.63
+ $X2=9.05 $Y2=2.26
r196 20 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.805 $Y=1.555
+ $X2=8.64 $Y2=1.555
r197 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.96 $Y=1.555
+ $X2=9.05 $Y2=1.63
r198 19 20 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=8.96 $Y=1.555
+ $X2=8.805 $Y2=1.555
r199 17 58 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=8.645 $Y=0.79
+ $X2=8.645 $Y2=1.3
r200 11 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.88
+ $X2=6.23 $Y2=1.715
r201 11 13 250.718 $w=1.8e-07 $l=6.45e-07 $layer=POLY_cond $X=6.23 $Y=1.88
+ $X2=6.23 $Y2=2.525
r202 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.215 $Y=1.55
+ $X2=6.215 $Y2=1.715
r203 7 9 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.215 $Y=1.55
+ $X2=6.215 $Y2=0.69
r204 2 28 600 $w=1.7e-07 $l=4.80885e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.825 $X2=2.115 $Y2=2.195
r205 1 62 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.9
+ $Y=0.665 $X2=3.11 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%CI 3 5 8 12 14 16 17 18 25
c63 25 0 6.54889e-20 $X=7.955 $Y=1.46
c64 8 0 2.79202e-20 $X=7.625 $Y=0.69
r65 23 25 19.9388 $w=2.78e-07 $l=1.15e-07 $layer=POLY_cond $X=7.84 $Y=1.46
+ $X2=7.955 $Y2=1.46
r66 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.84
+ $Y=1.385 $X2=7.84 $Y2=1.385
r67 21 23 37.277 $w=2.78e-07 $l=2.15e-07 $layer=POLY_cond $X=7.625 $Y=1.46
+ $X2=7.84 $Y2=1.46
r68 18 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.84 $Y=1.295 $X2=7.84
+ $Y2=1.385
r69 14 25 31.2086 $w=2.78e-07 $l=3.1749e-07 $layer=POLY_cond $X=8.135 $Y=1.22
+ $X2=7.955 $Y2=1.46
r70 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.135 $Y=1.22
+ $X2=8.135 $Y2=0.74
r71 10 25 12.9618 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=7.955 $Y=1.7
+ $X2=7.955 $Y2=1.46
r72 10 12 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=7.955 $Y=1.7 $X2=7.955
+ $Y2=2.4
r73 6 21 17.1848 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.625 $Y=1.22
+ $X2=7.625 $Y2=1.46
r74 6 8 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.625 $Y=1.22
+ $X2=7.625 $Y2=0.69
r75 3 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.45 $Y=1.88 $X2=7.45
+ $Y2=1.79
r76 3 5 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.45 $Y=1.88 $X2=7.45
+ $Y2=2.46
r77 1 21 32.9424 $w=2.78e-07 $l=1.9e-07 $layer=POLY_cond $X=7.435 $Y=1.46
+ $X2=7.625 $Y2=1.46
r78 1 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.435 $Y=1.55
+ $X2=7.435 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_1609_368# 1 2 3 12 16 19 21 24 28 32 35
+ 38 39 41 44 45 49 50
c115 44 0 1.11511e-19 $X=9.725 $Y=1.985
c116 39 0 1.25754e-19 $X=8.18 $Y=2.405
c117 38 0 2.79202e-20 $X=8.18 $Y=1.82
r118 50 52 0.995868 $w=2.42e-07 $l=5e-09 $layer=POLY_cond $X=10.12 $Y=1.425
+ $X2=10.115 $Y2=1.425
r119 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.12
+ $Y=1.425 $X2=10.12 $Y2=1.425
r120 46 49 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=9.945 $Y=1.425
+ $X2=10.12 $Y2=1.425
r121 44 45 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.795 $Y=1.985
+ $X2=9.795 $Y2=1.82
r122 41 42 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=0.965
+ $X2=8.345 $Y2=1.13
r123 38 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.26 $Y=1.82
+ $X2=8.26 $Y2=1.13
r124 36 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.945 $Y=1.59
+ $X2=9.945 $Y2=1.425
r125 36 45 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.945 $Y=1.59
+ $X2=9.945 $Y2=1.82
r126 34 44 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=9.795 $Y=2.055
+ $X2=9.795 $Y2=1.985
r127 34 35 6.74385 $w=4.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.795 $Y=2.055
+ $X2=9.795 $Y2=2.32
r128 33 39 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=2.405
+ $X2=8.18 $Y2=2.405
r129 32 35 8.97637 $w=1.7e-07 $l=2.74226e-07 $layer=LI1_cond $X=9.56 $Y=2.405
+ $X2=9.795 $Y2=2.32
r130 32 33 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=9.56 $Y=2.405
+ $X2=8.345 $Y2=2.405
r131 26 41 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=8.345 $Y=0.96
+ $X2=8.345 $Y2=0.965
r132 26 28 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=8.345 $Y=0.96
+ $X2=8.345 $Y2=0.515
r133 22 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.18 $Y=2.49
+ $X2=8.18 $Y2=2.405
r134 22 24 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.18 $Y=2.49
+ $X2=8.18 $Y2=2.815
r135 21 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.18 $Y=1.985
+ $X2=8.18 $Y2=1.82
r136 19 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.18 $Y=2.32
+ $X2=8.18 $Y2=2.405
r137 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.18 $Y=2.32
+ $X2=8.18 $Y2=1.985
r138 14 50 77.6777 $w=2.42e-07 $l=4.65242e-07 $layer=POLY_cond $X=10.51 $Y=1.59
+ $X2=10.12 $Y2=1.425
r139 14 16 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=10.51 $Y=1.59
+ $X2=10.51 $Y2=2.46
r140 10 52 13.9682 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.115 $Y=1.26
+ $X2=10.115 $Y2=1.425
r141 10 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=10.115 $Y=1.26
+ $X2=10.115 $Y2=0.79
r142 3 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.59
+ $Y=1.84 $X2=9.725 $Y2=1.985
r143 2 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.045
+ $Y=1.84 $X2=8.18 $Y2=2.815
r144 2 21 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.045
+ $Y=1.84 $X2=8.18 $Y2=1.985
r145 1 41 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.21
+ $Y=0.37 $X2=8.35 $Y2=0.965
r146 1 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.21
+ $Y=0.37 $X2=8.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_1744_94# 1 2 9 13 16 18 19 20 24 25 26 32
+ 33 36 37 38
c109 32 0 1.51844e-19 $X=9.275 $Y=1.985
c110 26 0 9.08104e-20 $X=10.325 $Y=0.665
r111 37 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.975 $Y=1.465
+ $X2=10.975 $Y2=1.63
r112 37 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.975 $Y=1.465
+ $X2=10.975 $Y2=1.3
r113 36 38 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=10.952 $Y=1.465
+ $X2=10.952 $Y2=1.3
r114 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.975
+ $Y=1.465 $X2=10.975 $Y2=1.465
r115 32 33 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=9.247 $Y=1.985
+ $X2=9.247 $Y2=1.82
r116 27 38 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=10.895 $Y=0.75
+ $X2=10.895 $Y2=1.3
r117 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.81 $Y=0.665
+ $X2=10.895 $Y2=0.75
r118 25 26 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.81 $Y=0.665
+ $X2=10.325 $Y2=0.665
r119 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.24 $Y=0.58
+ $X2=10.325 $Y2=0.665
r120 23 24 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.24 $Y=0.425
+ $X2=10.24 $Y2=0.58
r121 21 33 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=9.22 $Y=1.38
+ $X2=9.22 $Y2=1.82
r122 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.155 $Y=0.34
+ $X2=10.24 $Y2=0.425
r123 19 20 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=10.155 $Y=0.34
+ $X2=9.105 $Y2=0.34
r124 16 21 13.83 $w=2.47e-07 $l=3.69648e-07 $layer=LI1_cond $X=8.94 $Y=1.172
+ $X2=9.22 $Y2=1.38
r125 16 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.94 $Y=0.965
+ $X2=8.94 $Y2=0.615
r126 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.94 $Y=0.425
+ $X2=9.105 $Y2=0.34
r127 15 18 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=8.94 $Y=0.425
+ $X2=8.94 $Y2=0.615
r128 13 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.025 $Y=0.74
+ $X2=11.025 $Y2=1.3
r129 9 42 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.015 $Y=2.4
+ $X2=11.015 $Y2=1.63
r130 2 32 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.84 $X2=9.275 $Y2=1.985
r131 1 18 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.47 $X2=8.94 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%VPWR 1 2 3 4 17 23 29 35 38 39 40 42 54 63
+ 64 67 70 73
r94 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r95 70 71 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 64 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r98 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r99 61 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.9 $Y=3.33
+ $X2=10.775 $Y2=3.33
r100 61 63 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.9 $Y=3.33
+ $X2=11.28 $Y2=3.33
r101 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r102 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r103 57 60 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r104 56 59 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r105 56 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 54 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.775 $Y2=3.33
r107 54 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.32 $Y2=3.33
r108 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 49 52 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=4.71 $Y2=3.33
r114 47 49 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=5.04 $Y2=3.33
r115 46 71 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 46 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 45 46 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r119 43 45 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 42 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.71 $Y2=3.33
r121 42 45 218.23 $w=1.68e-07 $l=3.345e-06 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 40 53 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 40 50 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.04 $Y2=3.33
r124 38 52 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.645 $Y=3.33
+ $X2=7.44 $Y2=3.33
r125 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.645 $Y=3.33
+ $X2=7.73 $Y2=3.33
r126 37 56 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.815 $Y=3.33
+ $X2=7.92 $Y2=3.33
r127 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=3.33
+ $X2=7.73 $Y2=3.33
r128 33 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.775 $Y=3.245
+ $X2=10.775 $Y2=3.33
r129 33 35 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=10.775 $Y=3.245
+ $X2=10.775 $Y2=2.265
r130 29 32 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.73 $Y=2.105
+ $X2=7.73 $Y2=2.815
r131 27 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.73 $Y=3.245
+ $X2=7.73 $Y2=3.33
r132 27 32 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.73 $Y=3.245
+ $X2=7.73 $Y2=2.815
r133 23 26 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.71 $Y=1.97
+ $X2=4.71 $Y2=2.385
r134 21 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=3.245
+ $X2=4.71 $Y2=3.33
r135 21 26 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.71 $Y=3.245
+ $X2=4.71 $Y2=2.385
r136 17 20 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.82 $Y=2.115
+ $X2=0.82 $Y2=2.815
r137 15 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r138 15 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.815
r139 4 35 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=10.6
+ $Y=1.96 $X2=10.735 $Y2=2.265
r140 3 32 400 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.96 $X2=7.73 $Y2=2.815
r141 3 29 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.96 $X2=7.73 $Y2=2.105
r142 2 26 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=4.525
+ $Y=1.825 $X2=4.71 $Y2=2.385
r143 2 23 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.825 $X2=4.71 $Y2=1.97
r144 1 20 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.82 $Y2=2.815
r145 1 17 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=0.635
+ $Y=1.84 $X2=0.82 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_244_368# 1 2 3 4 16 18 23 25 26 29 33 35
c68 25 0 1.73957e-19 $X=3.46 $Y=2.99
r69 34 35 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.547 $Y=1.32
+ $X2=1.547 $Y2=1.49
r70 33 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.435 $Y=1.85
+ $X2=1.435 $Y2=1.49
r71 29 32 38.1953 $w=3.48e-07 $l=1.16e-06 $layer=LI1_cond $X=3.635 $Y=0.81
+ $X2=3.635 $Y2=1.97
r72 27 32 30.7867 $w=3.48e-07 $l=9.35e-07 $layer=LI1_cond $X=3.635 $Y=2.905
+ $X2=3.635 $Y2=1.97
r73 25 27 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=3.46 $Y=2.99
+ $X2=3.635 $Y2=2.905
r74 25 26 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=3.46 $Y=2.99
+ $X2=1.52 $Y2=2.99
r75 23 34 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.58 $Y=0.76
+ $X2=1.58 $Y2=1.32
r76 16 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=2.015
+ $X2=1.355 $Y2=1.85
r77 16 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.355 $Y=2.015
+ $X2=1.355 $Y2=2.695
r78 14 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=2.905
+ $X2=1.52 $Y2=2.99
r79 14 18 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.355 $Y=2.905
+ $X2=1.355 $Y2=2.695
r80 4 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=1.825 $X2=3.625 $Y2=1.97
r81 3 18 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.355 $Y2=2.695
r82 3 16 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.84 $X2=1.355 $Y2=2.015
r83 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.665 $X2=3.645 $Y2=0.81
r84 1 23 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=1.44
+ $Y=0.6 $X2=1.58 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_1026_389# 1 2 9 14 15 17 20 21 24
c55 17 0 1.05698e-19 $X=5.985 $Y=0.555
r56 22 24 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.315 $Y=1.22
+ $X2=5.41 $Y2=1.22
r57 20 21 7.76373 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.265 $Y=2.12
+ $X2=5.265 $Y2=1.975
r58 15 17 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=5.495 $Y=0.515
+ $X2=5.985 $Y2=0.515
r59 14 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=1.135
+ $X2=5.41 $Y2=1.22
r60 13 15 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.41 $Y=0.64
+ $X2=5.495 $Y2=0.515
r61 13 14 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.41 $Y=0.64
+ $X2=5.41 $Y2=1.135
r62 11 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=1.305
+ $X2=5.315 $Y2=1.22
r63 11 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.315 $Y=1.305
+ $X2=5.315 $Y2=1.975
r64 7 20 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=5.265 $Y=2.14 $X2=5.265
+ $Y2=2.12
r65 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.265 $Y=2.14
+ $X2=5.265 $Y2=2.46
r66 2 20 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.13
+ $Y=1.945 $X2=5.265 $Y2=2.12
r67 2 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.13
+ $Y=1.945 $X2=5.265 $Y2=2.46
r68 1 17 91 $w=1.7e-07 $l=7.11512e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.37 $X2=5.985 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%COUT_N 1 2 12 13 18 20
r55 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.485 $Y=1.21
+ $X2=6.485 $Y2=0.515
r56 15 18 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.09 $Y=1.295
+ $X2=6.485 $Y2=1.295
r57 12 13 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.982 $Y=2.25
+ $X2=5.982 $Y2=2.085
r58 9 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=1.38 $X2=6.09
+ $Y2=1.295
r59 9 13 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.09 $Y=1.38
+ $X2=6.09 $Y2=2.085
r60 2 12 300 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=2 $X=5.665
+ $Y=2.105 $X2=5.955 $Y2=2.25
r61 1 20 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=6.29
+ $Y=0.37 $X2=6.485 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_1264_421# 1 2 7 15 18 19
r47 18 19 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=7.39 $Y=2.085
+ $X2=7.39 $Y2=0.96
r48 13 19 7.30505 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=0.795
+ $X2=7.41 $Y2=0.96
r49 13 15 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.41 $Y=0.795
+ $X2=7.41 $Y2=0.515
r50 9 12 10.6147 $w=8.83e-07 $l=7.7e-07 $layer=LI1_cond $X=6.455 $Y=2.527
+ $X2=7.225 $Y2=2.527
r51 7 18 12.0616 $w=8.85e-07 $l=4.82632e-07 $layer=LI1_cond $X=7.305 $Y=2.527
+ $X2=7.39 $Y2=2.085
r52 7 12 1.10282 $w=8.83e-07 $l=8e-08 $layer=LI1_cond $X=7.305 $Y=2.527
+ $X2=7.225 $Y2=2.527
r53 2 12 200 $w=1.7e-07 $l=9.74808e-07 $layer=licon1_PDIFF $count=3 $X=6.32
+ $Y=2.105 $X2=7.225 $Y2=2.25
r54 2 9 200 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=3 $X=6.32
+ $Y=2.105 $X2=6.455 $Y2=2.25
r55 1 15 91 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_NDIFF $count=2 $X=7 $Y=0.37
+ $X2=7.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%A_1719_368# 1 2 3 10 14 16 17 21 25 27 33
c65 33 0 1.71654e-19 $X=10.54 $Y=1.845
r66 27 29 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.74 $Y=2.825
+ $X2=8.74 $Y2=2.955
r67 25 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.54 $Y=1.76
+ $X2=10.54 $Y2=1.845
r68 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.54 $Y=1.09
+ $X2=10.54 $Y2=1.76
r69 21 23 32.0876 $w=2.53e-07 $l=7.1e-07 $layer=LI1_cond $X=10.327 $Y=2.105
+ $X2=10.327 $Y2=2.815
r70 19 23 2.48566 $w=2.53e-07 $l=5.5e-08 $layer=LI1_cond $X=10.327 $Y=2.87
+ $X2=10.327 $Y2=2.815
r71 18 33 13.8963 $w=1.68e-07 $l=2.13e-07 $layer=LI1_cond $X=10.327 $Y=1.845
+ $X2=10.54 $Y2=1.845
r72 18 21 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=10.327 $Y=1.93
+ $X2=10.327 $Y2=2.105
r73 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.455 $Y=1.005
+ $X2=10.54 $Y2=1.09
r74 16 17 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=10.455 $Y=1.005
+ $X2=9.985 $Y2=1.005
r75 12 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.9 $Y=0.92
+ $X2=9.985 $Y2=1.005
r76 12 14 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=9.9 $Y=0.92 $X2=9.9
+ $Y2=0.84
r77 11 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.905 $Y=2.955
+ $X2=8.74 $Y2=2.955
r78 10 19 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=10.2 $Y=2.955
+ $X2=10.327 $Y2=2.87
r79 10 11 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=10.2 $Y=2.955
+ $X2=8.905 $Y2=2.955
r80 3 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.96 $X2=10.285 $Y2=2.815
r81 3 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.96 $X2=10.285 $Y2=2.105
r82 2 27 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=8.595
+ $Y=1.84 $X2=8.74 $Y2=2.825
r83 1 14 182 $w=1.7e-07 $l=5.23259e-07 $layer=licon1_NDIFF $count=1 $X=9.53
+ $Y=0.47 $X2=9.9 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%SUM 1 2 9 13 14 15 16 23 32
r28 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=11.255 $Y=2
+ $X2=11.255 $Y2=2.035
r29 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=11.255 $Y=2.405
+ $X2=11.255 $Y2=2.775
r30 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=2
r31 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=1.82
r32 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.405
r33 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.035
r34 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.35 $Y=1.13
+ $X2=11.35 $Y2=1.82
r35 7 13 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=11.295 $Y=0.99
+ $X2=11.295 $Y2=1.13
r36 7 9 19.5504 $w=2.78e-07 $l=4.75e-07 $layer=LI1_cond $X=11.295 $Y=0.99
+ $X2=11.295 $Y2=0.515
r37 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=1.985
r38 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=2.815
r39 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.1
+ $Y=0.37 $X2=11.24 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCON_1%VGND 1 2 3 4 14 17 21 24 25 29 31 37 44 52
+ 59 60 63 66 70
r108 70 73 9.3636 $w=3.98e-07 $l=3.25e-07 $layer=LI1_cond $X=10.695 $Y=0
+ $X2=10.695 $Y2=0.325
r109 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r110 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r111 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r112 60 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r113 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r114 57 70 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.895 $Y=0 $X2=10.695
+ $Y2=0
r115 57 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r116 56 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r117 56 67 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=7.92 $Y2=0
r118 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r119 53 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.87
+ $Y2=0
r120 53 55 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=7.995 $Y=0
+ $X2=10.32 $Y2=0
r121 52 70 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.495 $Y=0 $X2=10.695
+ $Y2=0
r122 52 55 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.32 $Y2=0
r123 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r124 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r125 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r126 47 50 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r127 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r128 45 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.03
+ $Y2=0
r129 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.52 $Y2=0
r130 44 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.87
+ $Y2=0
r131 44 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r132 43 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r133 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r134 40 43 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.72 $Y=0 $X2=4.56
+ $Y2=0
r135 39 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=4.56
+ $Y2=0
r136 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r137 37 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=5.03
+ $Y2=0
r138 37 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=4.56
+ $Y2=0
r139 35 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r140 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r141 31 51 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r142 31 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r143 26 29 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.63 $Y=0.645
+ $X2=0.725 $Y2=0.645
r144 24 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r145 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.63
+ $Y2=0
r146 23 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.72
+ $Y2=0
r147 23 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.63
+ $Y2=0
r148 19 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0
r149 19 21 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.495
r150 15 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r151 15 17 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.655
r152 14 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0.48
+ $X2=0.63 $Y2=0.645
r153 13 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0
r154 13 14 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0.48
r155 4 73 182 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=1 $X=10.19
+ $Y=0.47 $X2=10.695 $Y2=0.325
r156 3 21 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=7.7
+ $Y=0.37 $X2=7.91 $Y2=0.495
r157 2 17 182 $w=1.7e-07 $l=3.65992e-07 $layer=licon1_NDIFF $count=1 $X=4.885
+ $Y=0.37 $X2=5.07 $Y2=0.655
r158 1 29 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.5 $X2=0.725 $Y2=0.645
.ends


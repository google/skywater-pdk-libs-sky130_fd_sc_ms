* File: sky130_fd_sc_ms__nor2_2.pex.spice
* Created: Wed Sep  2 12:15:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR2_2%B 3 6 7 9 11 13 14 16 17
c38 17 0 6.90346e-20 $X=0.24 $Y=1.295
c39 9 0 1.87992e-19 $X=0.995 $Y=1.765
r40 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.385 $X2=0.28 $Y2=1.385
r41 17 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=1.295 $X2=0.28
+ $Y2=1.385
r42 15 16 27.7067 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=0.547 $Y=1.69
+ $X2=0.547 $Y2=1.765
r43 13 20 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.455 $Y=1.385
+ $X2=0.28 $Y2=1.385
r44 13 15 112.674 $w=1.85e-07 $l=3.05e-07 $layer=POLY_cond $X=0.547 $Y=1.385
+ $X2=0.547 $Y2=1.69
r45 13 14 63.6015 $w=1.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.547 $Y=1.385
+ $X2=0.547 $Y2=1.22
r46 9 11 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=2.4
r47 8 15 7.77431 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=0.64 $Y=1.69
+ $X2=0.547 $Y2=1.69
r48 7 9 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.905 $Y=1.69
+ $X2=0.995 $Y2=1.765
r49 7 8 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.905 $Y=1.69
+ $X2=0.64 $Y2=1.69
r50 6 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=0.74
+ $X2=0.565 $Y2=1.22
r51 3 16 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=0.545 $Y=2.4
+ $X2=0.545 $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_2%A 1 3 4 5 8 12 14 15 16 22 28 30
c46 5 0 6.90346e-20 $X=1.07 $Y=1.26
r47 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.44 $X2=1.97 $Y2=1.44
r48 26 28 8.79562 $w=4.11e-07 $l=7.5e-08 $layer=POLY_cond $X=1.895 $Y=1.395
+ $X2=1.97 $Y2=1.395
r49 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=0.42 $X2=1.97 $Y2=0.42
r50 20 28 8.00104 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.97 $Y=1.185
+ $X2=1.97 $Y2=1.395
r51 20 22 133.769 $w=3.3e-07 $l=7.65e-07 $layer=POLY_cond $X=1.97 $Y=1.185
+ $X2=1.97 $Y2=0.42
r52 16 29 4.35714 $w=4.06e-07 $l=1.45e-07 $layer=LI1_cond $X=2.04 $Y=1.295
+ $X2=2.04 $Y2=1.44
r53 16 31 3.37457 $w=4.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=1.295
+ $X2=2.04 $Y2=1.175
r54 15 31 6.36212 $w=4.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.04 $Y=0.925
+ $X2=2.04 $Y2=1.175
r55 15 30 6.36212 $w=4.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.04 $Y=0.925
+ $X2=2.04 $Y2=0.675
r56 14 30 3.36005 $w=4.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=0.555
+ $X2=2.04 $Y2=0.675
r57 14 23 4.03676 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.04 $Y=0.555
+ $X2=2.04 $Y2=0.42
r58 10 26 22.1098 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.895 $Y=1.605
+ $X2=1.895 $Y2=1.395
r59 10 12 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=1.895 $Y=1.605
+ $X2=1.895 $Y2=2.4
r60 6 26 52.7737 $w=4.11e-07 $l=4.5e-07 $layer=POLY_cond $X=1.445 $Y=1.395
+ $X2=1.895 $Y2=1.395
r61 6 8 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=1.445 $Y=1.59
+ $X2=1.445 $Y2=2.4
r62 4 6 31.0118 $w=4.11e-07 $l=1.74284e-07 $layer=POLY_cond $X=1.355 $Y=1.26
+ $X2=1.445 $Y2=1.395
r63 4 5 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.355 $Y=1.26
+ $X2=1.07 $Y2=1.26
r64 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=1.07 $Y2=1.26
r65 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_2%A_35_368# 1 2 3 12 16 17 24 25 28
r37 28 30 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.12 $Y=1.985
+ $X2=2.12 $Y2=2.815
r38 26 28 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.12 $Y=1.945 $X2=2.12
+ $Y2=1.985
r39 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.955 $Y=1.86
+ $X2=2.12 $Y2=1.945
r40 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.955 $Y=1.86
+ $X2=1.305 $Y2=1.86
r41 21 23 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.22 $Y=1.985
+ $X2=1.22 $Y2=2.815
r42 19 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.22 $Y=2.905 $X2=1.22
+ $Y2=2.815
r43 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=1.945
+ $X2=1.305 $Y2=1.86
r44 18 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.22 $Y=1.945 $X2=1.22
+ $Y2=1.985
r45 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=2.99
+ $X2=1.22 $Y2=2.905
r46 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.135 $Y=2.99
+ $X2=0.405 $Y2=2.99
r47 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r48 10 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.405 $Y2=2.99
r49 10 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r50 3 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=2.815
r51 3 28 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=1.985
r52 2 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.84 $X2=1.22 $Y2=2.815
r53 2 21 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.84 $X2=1.22 $Y2=1.985
r54 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r55 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_2%Y 1 2 9 11 12 18
r23 16 18 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.775 $Y=1.99
+ $X2=0.775 $Y2=2.035
r24 11 16 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.775 $Y=1.97
+ $X2=0.775 $Y2=1.99
r25 11 24 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.775 $Y=1.97
+ $X2=0.775 $Y2=1.82
r26 11 12 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=0.775 $Y=2.055
+ $X2=0.775 $Y2=2.405
r27 11 18 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.775 $Y=2.055
+ $X2=0.775 $Y2=2.035
r28 9 24 45.5739 $w=3.28e-07 $l=1.305e-06 $layer=LI1_cond $X=0.78 $Y=0.515
+ $X2=0.78 $Y2=1.82
r29 2 11 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=1.985
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_2%VPWR 1 6 9 10 11 21 22
c26 6 0 1.87992e-19 $X=1.67 $Y=2.28
r27 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 14 18 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 11 15 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 9 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 9 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.63 $Y2=3.33
r35 8 21 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 8 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.63 $Y2=3.33
r37 4 10 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r38 4 6 44.4843 $w=2.48e-07 $l=9.65e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.28
r39 1 6 300 $w=1.7e-07 $l=5.02991e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.84 $X2=1.67 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_2%VGND 1 2 7 9 13 15 17 24 25 31
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r30 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r31 22 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=2.16
+ $Y2=0
r32 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r33 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 18 28 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r35 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r36 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r37 17 20 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r38 15 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r39 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r40 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r42 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.515
r43 7 28 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r44 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r45 2 13 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r46 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends


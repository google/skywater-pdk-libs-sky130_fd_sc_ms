* File: sky130_fd_sc_ms__ha_2.pxi.spice
* Created: Fri Aug 28 17:37:22 2020
* 
x_PM_SKY130_FD_SC_MS__HA_2%B N_B_c_113_n N_B_M1014_g N_B_M1016_g N_B_c_106_n
+ N_B_M1007_g N_B_c_107_n N_B_M1010_g N_B_c_108_n N_B_c_109_n N_B_c_110_n
+ N_B_c_111_n N_B_c_123_p B B B B PM_SKY130_FD_SC_MS__HA_2%B
x_PM_SKY130_FD_SC_MS__HA_2%A N_A_M1009_g N_A_M1015_g N_A_M1001_g N_A_M1005_g A
+ N_A_c_194_n PM_SKY130_FD_SC_MS__HA_2%A
x_PM_SKY130_FD_SC_MS__HA_2%A_27_74# N_A_27_74#_M1016_s N_A_27_74#_M1014_d
+ N_A_27_74#_M1017_g N_A_27_74#_c_264_n N_A_27_74#_M1013_g N_A_27_74#_M1006_g
+ N_A_27_74#_M1000_g N_A_27_74#_M1011_g N_A_27_74#_M1008_g N_A_27_74#_c_251_n
+ N_A_27_74#_c_252_n N_A_27_74#_c_253_n N_A_27_74#_c_254_n N_A_27_74#_c_255_n
+ N_A_27_74#_c_256_n N_A_27_74#_c_257_n N_A_27_74#_c_324_p N_A_27_74#_c_258_n
+ N_A_27_74#_c_315_p N_A_27_74#_c_291_n N_A_27_74#_c_259_n N_A_27_74#_c_293_n
+ N_A_27_74#_c_260_n N_A_27_74#_c_261_n N_A_27_74#_c_262_n N_A_27_74#_c_263_n
+ PM_SKY130_FD_SC_MS__HA_2%A_27_74#
x_PM_SKY130_FD_SC_MS__HA_2%A_394_388# N_A_394_388#_M1017_s N_A_394_388#_M1010_d
+ N_A_394_388#_M1002_g N_A_394_388#_c_412_n N_A_394_388#_M1004_g
+ N_A_394_388#_M1003_g N_A_394_388#_c_414_n N_A_394_388#_M1012_g
+ N_A_394_388#_c_423_n N_A_394_388#_c_491_p N_A_394_388#_c_415_n
+ N_A_394_388#_c_416_n N_A_394_388#_c_417_n N_A_394_388#_c_466_p
+ N_A_394_388#_c_418_n N_A_394_388#_c_419_n N_A_394_388#_c_420_n
+ PM_SKY130_FD_SC_MS__HA_2%A_394_388#
x_PM_SKY130_FD_SC_MS__HA_2%VPWR N_VPWR_M1014_s N_VPWR_M1015_d N_VPWR_M1013_d
+ N_VPWR_M1003_s N_VPWR_M1011_s N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n VPWR N_VPWR_c_506_n
+ N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n
+ N_VPWR_c_512_n N_VPWR_c_499_n PM_SKY130_FD_SC_MS__HA_2%VPWR
x_PM_SKY130_FD_SC_MS__HA_2%SUM N_SUM_M1004_d N_SUM_M1002_d N_SUM_c_571_n
+ N_SUM_c_567_n SUM SUM N_SUM_c_569_n PM_SKY130_FD_SC_MS__HA_2%SUM
x_PM_SKY130_FD_SC_MS__HA_2%COUT N_COUT_M1000_d N_COUT_M1006_d N_COUT_c_601_n
+ N_COUT_c_598_n COUT COUT COUT PM_SKY130_FD_SC_MS__HA_2%COUT
x_PM_SKY130_FD_SC_MS__HA_2%VGND N_VGND_M1009_d N_VGND_M1007_d N_VGND_M1004_s
+ N_VGND_M1012_s N_VGND_M1008_s N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n
+ N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ N_VGND_c_640_n N_VGND_c_641_n VGND N_VGND_c_642_n N_VGND_c_643_n
+ N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n
+ PM_SKY130_FD_SC_MS__HA_2%VGND
x_PM_SKY130_FD_SC_MS__HA_2%A_278_74# N_A_278_74#_M1001_d N_A_278_74#_M1017_d
+ N_A_278_74#_c_705_n N_A_278_74#_c_706_n N_A_278_74#_c_707_n
+ N_A_278_74#_c_708_n N_A_278_74#_c_709_n PM_SKY130_FD_SC_MS__HA_2%A_278_74#
cc_1 VNB N_B_M1016_g 0.0297382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B_c_106_n 0.0173977f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.185
cc_3 VNB N_B_c_107_n 0.04926f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.78
cc_4 VNB N_B_c_108_n 0.00167339f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_5 VNB N_B_c_109_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.615
cc_6 VNB N_B_c_110_n 0.0137652f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_7 VNB N_B_c_111_n 0.0387783f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_8 VNB B 0.00154267f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_9 VNB N_A_M1009_g 0.0232343f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.88
cc_10 VNB N_A_M1001_g 0.0249069f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_11 VNB N_A_c_194_n 0.034228f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.63
cc_12 VNB N_A_27_74#_M1017_g 0.0257234f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_13 VNB N_A_27_74#_M1006_g 0.001465f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.615
cc_14 VNB N_A_27_74#_M1000_g 0.0207917f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.63
cc_15 VNB N_A_27_74#_M1011_g 0.00166756f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_16 VNB N_A_27_74#_M1008_g 0.026707f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_17 VNB N_A_27_74#_c_251_n 0.00327664f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.32
cc_18 VNB N_A_27_74#_c_252_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_253_n 0.00469558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_254_n 0.00942532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_255_n 0.0023864f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.3
cc_22 VNB N_A_27_74#_c_256_n 0.0286895f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.63
cc_23 VNB N_A_27_74#_c_257_n 9.06092e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.42
cc_24 VNB N_A_27_74#_c_258_n 0.0748099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_259_n 0.00120577f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.42
cc_26 VNB N_A_27_74#_c_260_n 0.00146718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_261_n 0.00717931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_262_n 0.00509894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_263_n 0.0730235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_394_388#_M1002_g 0.00669167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_394_388#_c_412_n 0.0198259f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_32 VNB N_A_394_388#_M1003_g 0.00602725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_394_388#_c_414_n 0.017136f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.32
cc_34 VNB N_A_394_388#_c_415_n 0.003372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_394_388#_c_416_n 0.00102048f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.42
cc_36 VNB N_A_394_388#_c_417_n 0.00213328f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_37 VNB N_A_394_388#_c_418_n 0.0119963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_394_388#_c_419_n 0.0608476f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.63
cc_39 VNB N_A_394_388#_c_420_n 0.037587f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.42
cc_40 VNB N_VPWR_c_499_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_SUM_c_567_n 0.00990022f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_42 VNB N_COUT_c_598_n 0.00134727f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_43 VNB COUT 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.78
cc_44 VNB COUT 0.00417716f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.44
cc_45 VNB N_VGND_c_632_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.32
cc_46 VNB N_VGND_c_633_n 0.00851745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_634_n 0.00938716f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_48 VNB N_VGND_c_635_n 0.00493915f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.42
cc_49 VNB N_VGND_c_636_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_50 VNB N_VGND_c_637_n 0.0450391f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.32
cc_51 VNB N_VGND_c_638_n 0.0291765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_639_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_640_n 0.016486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_641_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_55 VNB N_VGND_c_642_n 0.0353722f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=2.42
cc_56 VNB N_VGND_c_643_n 0.0180771f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.42
cc_57 VNB N_VGND_c_644_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_645_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_646_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_647_n 0.34251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_278_74#_c_705_n 0.0101103f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_62 VNB N_A_278_74#_c_706_n 0.00817638f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_63 VNB N_A_278_74#_c_707_n 0.013117f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.78
cc_64 VNB N_A_278_74#_c_708_n 0.00353599f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.44
cc_65 VNB N_A_278_74#_c_709_n 0.00359387f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_66 VPB N_B_c_113_n 0.0220706f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.88
cc_67 VPB N_B_c_107_n 0.0135149f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.78
cc_68 VPB N_B_M1010_g 0.0260723f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=2.44
cc_69 VPB N_B_c_108_n 0.00744368f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_70 VPB N_B_c_109_n 0.00148678f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.615
cc_71 VPB B 0.0338726f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=2.32
cc_72 VPB N_A_M1015_g 0.0198464f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_73 VPB N_A_M1005_g 0.0216783f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=2.44
cc_74 VPB A 0.00483519f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_75 VPB N_A_c_194_n 0.0146214f $X=-0.19 $Y=1.66 $X2=0.21 $Y2=1.63
cc_76 VPB N_A_27_74#_c_264_n 0.0290231f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=2.44
cc_77 VPB N_A_27_74#_M1006_g 0.0213324f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.615
cc_78 VPB N_A_27_74#_M1011_g 0.0245596f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.465
cc_79 VPB N_A_27_74#_c_251_n 0.00862625f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=2.32
cc_80 VPB N_A_27_74#_c_255_n 0.0021267f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.3
cc_81 VPB N_A_27_74#_c_257_n 0.0060413f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.42
cc_82 VPB N_A_27_74#_c_259_n 0.00773025f $X=-0.19 $Y=1.66 $X2=0.21 $Y2=2.42
cc_83 VPB N_A_394_388#_M1002_g 0.0250091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_394_388#_M1003_g 0.0218669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_394_388#_c_423_n 0.0105005f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.615
cc_86 VPB N_A_394_388#_c_417_n 0.00644789f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=2.32
cc_87 VPB N_VPWR_c_500_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_501_n 0.0207459f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.32
cc_89 VPB N_VPWR_c_502_n 0.00454028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_503_n 0.00261656f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.465
cc_91 VPB N_VPWR_c_504_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.465
cc_92 VPB N_VPWR_c_505_n 0.02067f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=2.42
cc_93 VPB N_VPWR_c_506_n 0.0180749f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=2.32
cc_94 VPB N_VPWR_c_507_n 0.017758f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.615
cc_95 VPB N_VPWR_c_508_n 0.0177589f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=2.42
cc_96 VPB N_VPWR_c_509_n 0.00734065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_510_n 0.0533445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_511_n 0.0220885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_512_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_499_n 0.0880503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_SUM_c_567_n 0.00286068f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_102 VPB N_SUM_c_569_n 0.00403418f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.32
cc_103 VPB N_COUT_c_601_n 0.00359349f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=1.185
cc_104 VPB N_COUT_c_598_n 8.08081e-19 $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_105 N_B_M1016_g N_A_M1009_g 0.0340417f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B_c_110_n N_A_M1009_g 2.56105e-19 $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_107 N_B_c_113_n N_A_M1015_g 0.0429944f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_108 N_B_c_108_n N_A_M1015_g 0.00462911f $X=0.505 $Y=1.79 $X2=0 $Y2=0
cc_109 N_B_c_123_p N_A_M1015_g 0.0192692f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_110 N_B_c_106_n N_A_M1001_g 0.0312814f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_111 N_B_c_107_n N_A_M1001_g 0.00903936f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_112 N_B_M1010_g N_A_M1005_g 0.0402713f $X=1.88 $Y=2.44 $X2=0 $Y2=0
cc_113 N_B_c_123_p N_A_M1005_g 0.0196319f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_114 N_B_c_107_n A 0.00116491f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_115 N_B_c_109_n A 0.0124081f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_116 N_B_c_123_p A 0.00965235f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_117 N_B_c_107_n N_A_c_194_n 0.0402713f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_118 N_B_c_109_n N_A_c_194_n 0.00505747f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_119 N_B_c_111_n N_A_c_194_n 0.0386708f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_120 N_B_c_123_p N_A_c_194_n 7.54049e-19 $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_121 N_B_c_123_p N_A_27_74#_M1014_d 0.00478714f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_122 N_B_M1016_g N_A_27_74#_c_252_n 0.0123382f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B_c_113_n N_A_27_74#_c_253_n 6.25944e-19 $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_124 N_B_M1016_g N_A_27_74#_c_253_n 0.0108371f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_125 N_B_c_110_n N_A_27_74#_c_253_n 0.00746443f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_126 N_B_M1016_g N_A_27_74#_c_254_n 0.00113234f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B_c_110_n N_A_27_74#_c_254_n 0.0272661f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_128 N_B_c_111_n N_A_27_74#_c_254_n 0.00467885f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_129 N_B_c_113_n N_A_27_74#_c_255_n 0.0014999f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_130 N_B_c_110_n N_A_27_74#_c_255_n 0.025258f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_131 N_B_c_111_n N_A_27_74#_c_255_n 0.00348918f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_132 B N_A_27_74#_c_255_n 0.0137441f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_133 N_B_c_106_n N_A_27_74#_c_256_n 0.00565175f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_134 N_B_c_107_n N_A_27_74#_c_256_n 0.0152606f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_135 N_B_c_109_n N_A_27_74#_c_256_n 0.0256551f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_136 N_B_c_107_n N_A_27_74#_c_257_n 0.0038093f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_137 N_B_M1010_g N_A_27_74#_c_257_n 0.00277051f $X=1.88 $Y=2.44 $X2=0 $Y2=0
cc_138 N_B_c_109_n N_A_27_74#_c_257_n 0.054424f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_139 N_B_c_123_p N_A_27_74#_c_257_n 0.00159069f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_140 N_B_c_107_n N_A_27_74#_c_258_n 0.0123225f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_141 N_B_M1010_g N_A_27_74#_c_291_n 9.46803e-19 $X=1.88 $Y=2.44 $X2=0 $Y2=0
cc_142 N_B_c_123_p N_A_27_74#_c_291_n 0.0153274f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_143 N_B_c_113_n N_A_27_74#_c_293_n 0.00396863f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_144 N_B_c_123_p N_A_27_74#_c_293_n 0.0155211f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_145 B N_A_27_74#_c_293_n 0.00872339f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_146 N_B_M1016_g N_A_27_74#_c_260_n 0.0036485f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_147 N_B_c_107_n N_A_27_74#_c_261_n 0.00506711f $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_148 N_B_c_109_n N_A_27_74#_c_261_n 0.0134933f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_149 N_B_c_109_n N_A_394_388#_M1010_d 0.00412198f $X=1.955 $Y=1.615 $X2=0
+ $Y2=0
cc_150 N_B_c_123_p N_A_394_388#_M1010_d 0.00468291f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_151 N_B_c_123_p N_VPWR_M1014_s 0.001789f $X=1.79 $Y=2.42 $X2=-0.19 $Y2=-0.245
cc_152 B N_VPWR_M1014_s 0.0100702f $X=0.155 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_153 N_B_c_123_p N_VPWR_M1015_d 0.0058179f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_154 N_B_c_113_n N_VPWR_c_501_n 0.0105188f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_155 N_B_c_123_p N_VPWR_c_501_n 0.0071545f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_156 B N_VPWR_c_501_n 0.0148608f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_157 N_B_c_113_n N_VPWR_c_502_n 0.00105093f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_158 N_B_M1010_g N_VPWR_c_502_n 0.0018217f $X=1.88 $Y=2.44 $X2=0 $Y2=0
cc_159 N_B_c_123_p N_VPWR_c_502_n 0.0211976f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_160 N_B_c_113_n N_VPWR_c_506_n 0.00547402f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_161 N_B_M1010_g N_VPWR_c_510_n 0.00676105f $X=1.88 $Y=2.44 $X2=0 $Y2=0
cc_162 N_B_c_113_n N_VPWR_c_499_n 0.00536634f $X=0.505 $Y=1.88 $X2=0 $Y2=0
cc_163 N_B_M1010_g N_VPWR_c_499_n 0.00647345f $X=1.88 $Y=2.44 $X2=0 $Y2=0
cc_164 N_B_c_123_p N_VPWR_c_499_n 0.0474698f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_165 B N_VPWR_c_499_n 6.43314e-19 $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_166 N_B_c_123_p A_310_388# 0.00742025f $X=1.79 $Y=2.42 $X2=-0.19 $Y2=-0.245
cc_167 N_B_M1016_g N_VGND_c_632_n 0.00126873f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B_c_106_n N_VGND_c_632_n 0.00106137f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_169 N_B_c_106_n N_VGND_c_633_n 0.00970106f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_170 N_B_M1016_g N_VGND_c_638_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B_c_106_n N_VGND_c_640_n 0.00383152f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_172 N_B_M1016_g N_VGND_c_647_n 0.00824638f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B_c_106_n N_VGND_c_647_n 0.00369368f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_174 N_B_c_106_n N_A_278_74#_c_705_n 0.0113476f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_175 N_B_c_107_n N_A_278_74#_c_705_n 5.76956e-19 $X=1.88 $Y=1.78 $X2=0 $Y2=0
cc_176 N_B_c_106_n N_A_278_74#_c_706_n 0.0028624f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_177 N_B_c_106_n N_A_278_74#_c_708_n 5.73857e-19 $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_178 N_A_M1009_g N_A_27_74#_c_252_n 0.00248918f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_M1009_g N_A_27_74#_c_253_n 2.23249e-19 $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_M1009_g N_A_27_74#_c_255_n 0.00308843f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_M1015_g N_A_27_74#_c_255_n 0.00507269f $X=0.955 $Y=2.42 $X2=0 $Y2=0
cc_182 N_A_M1005_g N_A_27_74#_c_255_n 9.45948e-19 $X=1.46 $Y=2.44 $X2=0 $Y2=0
cc_183 A N_A_27_74#_c_255_n 0.0236139f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A_c_194_n N_A_27_74#_c_255_n 0.0114373f $X=1.315 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A_M1009_g N_A_27_74#_c_256_n 0.00934412f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_M1001_g N_A_27_74#_c_256_n 0.0137825f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_187 A N_A_27_74#_c_256_n 0.0242166f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A_c_194_n N_A_27_74#_c_256_n 0.00851165f $X=1.315 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A_M1015_g N_A_27_74#_c_293_n 0.0040933f $X=0.955 $Y=2.42 $X2=0 $Y2=0
cc_190 N_A_M1005_g N_A_27_74#_c_293_n 7.85429e-19 $X=1.46 $Y=2.44 $X2=0 $Y2=0
cc_191 N_A_M1009_g N_A_27_74#_c_260_n 0.0106214f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_M1001_g N_A_27_74#_c_260_n 0.00156882f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_M1015_g N_VPWR_c_501_n 0.00105204f $X=0.955 $Y=2.42 $X2=0 $Y2=0
cc_194 N_A_M1015_g N_VPWR_c_502_n 0.00966588f $X=0.955 $Y=2.42 $X2=0 $Y2=0
cc_195 N_A_M1005_g N_VPWR_c_502_n 0.0101071f $X=1.46 $Y=2.44 $X2=0 $Y2=0
cc_196 N_A_M1015_g N_VPWR_c_506_n 0.00547402f $X=0.955 $Y=2.42 $X2=0 $Y2=0
cc_197 N_A_M1005_g N_VPWR_c_510_n 0.00562069f $X=1.46 $Y=2.44 $X2=0 $Y2=0
cc_198 N_A_M1015_g N_VPWR_c_499_n 0.00536634f $X=0.955 $Y=2.42 $X2=0 $Y2=0
cc_199 N_A_M1005_g N_VPWR_c_499_n 0.0054305f $X=1.46 $Y=2.44 $X2=0 $Y2=0
cc_200 N_A_M1009_g N_VGND_c_632_n 0.00876864f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_M1001_g N_VGND_c_632_n 0.00891708f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_M1001_g N_VGND_c_633_n 0.00106137f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_M1009_g N_VGND_c_638_n 0.00383152f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_M1001_g N_VGND_c_640_n 0.00383152f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_M1009_g N_VGND_c_647_n 0.0075725f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_M1001_g N_VGND_c_647_n 0.006806f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_M1009_g N_A_278_74#_c_705_n 8.11834e-19 $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_M1001_g N_A_278_74#_c_705_n 0.00416578f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_27_74#_c_257_n N_A_394_388#_M1010_d 0.0119319f $X=2.375 $Y=2.34 $X2=0
+ $Y2=0
cc_210 N_A_27_74#_c_315_p N_A_394_388#_M1010_d 0.0198666f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_211 N_A_27_74#_c_291_n N_A_394_388#_M1010_d 0.00708664f $X=2.46 $Y=2.425
+ $X2=0 $Y2=0
cc_212 N_A_27_74#_c_264_n N_A_394_388#_M1002_g 0.0125885f $X=3.02 $Y=1.88 $X2=0
+ $Y2=0
cc_213 N_A_27_74#_c_315_p N_A_394_388#_M1002_g 0.0191336f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_214 N_A_27_74#_c_315_p N_A_394_388#_M1003_g 0.0129745f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_215 N_A_27_74#_c_263_n N_A_394_388#_M1003_g 0.0508297f $X=5.265 $Y=1.465
+ $X2=0 $Y2=0
cc_216 N_A_27_74#_M1000_g N_A_394_388#_c_414_n 0.0282033f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_A_27_74#_c_264_n N_A_394_388#_c_423_n 0.016741f $X=3.02 $Y=1.88 $X2=0
+ $Y2=0
cc_218 N_A_27_74#_c_257_n N_A_394_388#_c_423_n 0.0202358f $X=2.375 $Y=2.34 $X2=0
+ $Y2=0
cc_219 N_A_27_74#_c_324_p N_A_394_388#_c_423_n 0.0196011f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_220 N_A_27_74#_c_258_n N_A_394_388#_c_423_n 0.0063963f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_221 N_A_27_74#_c_315_p N_A_394_388#_c_423_n 0.0559474f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_222 N_A_27_74#_M1017_g N_A_394_388#_c_415_n 0.012478f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_27_74#_c_264_n N_A_394_388#_c_415_n 7.36618e-19 $X=3.02 $Y=1.88 $X2=0
+ $Y2=0
cc_224 N_A_27_74#_c_324_p N_A_394_388#_c_415_n 0.0136762f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_225 N_A_27_74#_c_258_n N_A_394_388#_c_415_n 0.00191708f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_226 N_A_27_74#_c_324_p N_A_394_388#_c_416_n 0.0136463f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_227 N_A_27_74#_c_258_n N_A_394_388#_c_416_n 0.00391672f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_228 N_A_27_74#_c_264_n N_A_394_388#_c_417_n 0.00304252f $X=3.02 $Y=1.88 $X2=0
+ $Y2=0
cc_229 N_A_27_74#_c_258_n N_A_394_388#_c_417_n 0.00722092f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_230 N_A_27_74#_M1017_g N_A_394_388#_c_418_n 0.00421066f $X=2.935 $Y=0.74
+ $X2=0 $Y2=0
cc_231 N_A_27_74#_c_324_p N_A_394_388#_c_418_n 0.0167012f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_232 N_A_27_74#_c_258_n N_A_394_388#_c_418_n 0.00118728f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_233 N_A_27_74#_M1017_g N_A_394_388#_c_419_n 0.00275209f $X=2.935 $Y=0.74
+ $X2=0 $Y2=0
cc_234 N_A_27_74#_c_324_p N_A_394_388#_c_419_n 0.00106912f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_235 N_A_27_74#_c_258_n N_A_394_388#_c_419_n 0.0158741f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_236 N_A_27_74#_c_263_n N_A_394_388#_c_420_n 0.012752f $X=5.265 $Y=1.465 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_c_315_p N_VPWR_M1013_d 0.0230736f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_238 N_A_27_74#_c_315_p N_VPWR_M1003_s 0.00325968f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_239 N_A_27_74#_c_315_p N_VPWR_M1011_s 0.00960768f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_240 N_A_27_74#_c_259_n N_VPWR_M1011_s 0.022026f $X=5.47 $Y=2.34 $X2=0 $Y2=0
cc_241 N_A_27_74#_M1006_g N_VPWR_c_503_n 0.0103068f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A_27_74#_M1011_g N_VPWR_c_503_n 0.00119973f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_315_p N_VPWR_c_503_n 0.0166216f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_244 N_A_27_74#_M1006_g N_VPWR_c_505_n 0.00119973f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A_27_74#_M1011_g N_VPWR_c_505_n 0.011438f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_315_p N_VPWR_c_505_n 0.0155081f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_247 N_A_27_74#_M1006_g N_VPWR_c_508_n 0.00460063f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_27_74#_M1011_g N_VPWR_c_508_n 0.00460063f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_27_74#_c_264_n N_VPWR_c_510_n 0.00562069f $X=3.02 $Y=1.88 $X2=0 $Y2=0
cc_250 N_A_27_74#_c_264_n N_VPWR_c_511_n 0.022365f $X=3.02 $Y=1.88 $X2=0 $Y2=0
cc_251 N_A_27_74#_c_315_p N_VPWR_c_511_n 0.0510767f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_c_264_n N_VPWR_c_499_n 0.00539454f $X=3.02 $Y=1.88 $X2=0 $Y2=0
cc_253 N_A_27_74#_M1006_g N_VPWR_c_499_n 0.00455838f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_27_74#_M1011_g N_VPWR_c_499_n 0.00455838f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A_27_74#_c_315_p N_VPWR_c_499_n 0.0615639f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_256 N_A_27_74#_c_291_n N_VPWR_c_499_n 0.00678047f $X=2.46 $Y=2.425 $X2=0
+ $Y2=0
cc_257 N_A_27_74#_c_315_p N_SUM_M1002_d 0.00474508f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_258 N_A_27_74#_M1000_g N_SUM_c_571_n 0.00141692f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_27_74#_M1006_g N_SUM_c_567_n 0.00162105f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_27_74#_M1000_g N_SUM_c_567_n 0.00177272f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_27_74#_c_315_p N_SUM_c_567_n 0.0124479f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_262 N_A_27_74#_c_263_n N_SUM_c_567_n 0.00456353f $X=5.265 $Y=1.465 $X2=0
+ $Y2=0
cc_263 N_A_27_74#_c_315_p N_SUM_c_569_n 0.0270781f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_264 N_A_27_74#_c_315_p N_COUT_M1006_d 0.00474103f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_265 N_A_27_74#_M1006_g N_COUT_c_601_n 0.00556879f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_266 N_A_27_74#_M1011_g N_COUT_c_601_n 0.00630301f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_267 N_A_27_74#_c_315_p N_COUT_c_601_n 0.0166124f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_268 N_A_27_74#_c_259_n N_COUT_c_601_n 0.0126742f $X=5.47 $Y=2.34 $X2=0 $Y2=0
cc_269 N_A_27_74#_c_263_n N_COUT_c_601_n 7.98008e-19 $X=5.265 $Y=1.465 $X2=0
+ $Y2=0
cc_270 N_A_27_74#_M1006_g N_COUT_c_598_n 0.00362606f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A_27_74#_M1000_g N_COUT_c_598_n 0.00331881f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_272 N_A_27_74#_M1011_g N_COUT_c_598_n 0.00115534f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_27_74#_M1008_g N_COUT_c_598_n 0.002587f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_27_74#_c_259_n N_COUT_c_598_n 0.00661557f $X=5.47 $Y=2.34 $X2=0 $Y2=0
cc_275 N_A_27_74#_c_262_n N_COUT_c_598_n 0.0235661f $X=5.39 $Y=1.465 $X2=0 $Y2=0
cc_276 N_A_27_74#_c_263_n N_COUT_c_598_n 0.0157146f $X=5.265 $Y=1.465 $X2=0
+ $Y2=0
cc_277 N_A_27_74#_M1000_g COUT 0.00892916f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A_27_74#_M1008_g COUT 0.00788704f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A_27_74#_M1000_g COUT 0.00203717f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_27_74#_M1008_g COUT 0.00327512f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_27_74#_c_263_n COUT 0.00209846f $X=5.265 $Y=1.465 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_253_n A_114_74# 0.0039014f $X=0.72 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_283 N_A_27_74#_c_260_n A_114_74# 0.0018016f $X=0.805 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_27_74#_c_252_n N_VGND_c_632_n 0.00792017f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_285 N_A_27_74#_c_256_n N_VGND_c_632_n 0.00968283f $X=2.29 $Y=1.195 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_M1017_g N_VGND_c_634_n 0.00144451f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_M1000_g N_VGND_c_635_n 0.00294833f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_M1008_g N_VGND_c_637_n 0.00647412f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_262_n N_VGND_c_637_n 0.0140864f $X=5.39 $Y=1.465 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_263_n N_VGND_c_637_n 0.00125053f $X=5.265 $Y=1.465 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_c_252_n N_VGND_c_638_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_292 N_A_27_74#_M1017_g N_VGND_c_642_n 0.00278247f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_M1000_g N_VGND_c_644_n 0.00434272f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_M1008_g N_VGND_c_644_n 0.00434272f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_M1017_g N_VGND_c_647_n 0.00363424f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_M1000_g N_VGND_c_647_n 0.00820382f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_M1008_g N_VGND_c_647_n 0.00823942f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_252_n N_VGND_c_647_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_256_n N_A_278_74#_c_705_n 0.0613147f $X=2.29 $Y=1.195 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_324_p N_A_278_74#_c_705_n 2.30459e-19 $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_258_n N_A_278_74#_c_705_n 6.05904e-19 $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_261_n N_A_278_74#_c_705_n 0.0158527f $X=2.375 $Y=1.36 $X2=0
+ $Y2=0
cc_303 N_A_27_74#_M1017_g N_A_278_74#_c_706_n 0.00317277f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_M1017_g N_A_278_74#_c_707_n 0.0131176f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_M1017_g N_A_278_74#_c_709_n 0.00549447f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_394_388#_c_423_n N_VPWR_M1013_d 0.00935782f $X=3.32 $Y=2.045 $X2=0
+ $Y2=0
cc_307 N_A_394_388#_M1002_g N_VPWR_c_503_n 0.00120108f $X=3.905 $Y=2.4 $X2=0
+ $Y2=0
cc_308 N_A_394_388#_M1003_g N_VPWR_c_503_n 0.0102839f $X=4.355 $Y=2.4 $X2=0
+ $Y2=0
cc_309 N_A_394_388#_M1002_g N_VPWR_c_507_n 0.00460063f $X=3.905 $Y=2.4 $X2=0
+ $Y2=0
cc_310 N_A_394_388#_M1003_g N_VPWR_c_507_n 0.00460063f $X=4.355 $Y=2.4 $X2=0
+ $Y2=0
cc_311 N_A_394_388#_M1002_g N_VPWR_c_511_n 0.0116314f $X=3.905 $Y=2.4 $X2=0
+ $Y2=0
cc_312 N_A_394_388#_M1003_g N_VPWR_c_511_n 0.00119308f $X=4.355 $Y=2.4 $X2=0
+ $Y2=0
cc_313 N_A_394_388#_M1002_g N_VPWR_c_499_n 0.00454199f $X=3.905 $Y=2.4 $X2=0
+ $Y2=0
cc_314 N_A_394_388#_M1003_g N_VPWR_c_499_n 0.00455838f $X=4.355 $Y=2.4 $X2=0
+ $Y2=0
cc_315 N_A_394_388#_c_412_n N_SUM_c_571_n 0.00614403f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_316 N_A_394_388#_c_414_n N_SUM_c_571_n 0.015895f $X=4.405 $Y=1.22 $X2=0 $Y2=0
cc_317 N_A_394_388#_c_466_p N_SUM_c_571_n 0.021978f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_318 N_A_394_388#_c_418_n N_SUM_c_571_n 0.00394508f $X=3.405 $Y=1.025 $X2=0
+ $Y2=0
cc_319 N_A_394_388#_c_420_n N_SUM_c_571_n 0.00361918f $X=4.355 $Y=1.385 $X2=0
+ $Y2=0
cc_320 N_A_394_388#_c_414_n N_SUM_c_567_n 0.00438312f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_321 N_A_394_388#_c_466_p N_SUM_c_567_n 0.0256364f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_322 N_A_394_388#_c_420_n N_SUM_c_567_n 0.00807539f $X=4.355 $Y=1.385 $X2=0
+ $Y2=0
cc_323 N_A_394_388#_M1002_g N_SUM_c_569_n 0.00789648f $X=3.905 $Y=2.4 $X2=0
+ $Y2=0
cc_324 N_A_394_388#_M1003_g N_SUM_c_569_n 0.0184199f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A_394_388#_c_423_n N_SUM_c_569_n 0.00983061f $X=3.32 $Y=2.045 $X2=0
+ $Y2=0
cc_326 N_A_394_388#_c_417_n N_SUM_c_569_n 0.00362678f $X=3.405 $Y=1.92 $X2=0
+ $Y2=0
cc_327 N_A_394_388#_c_466_p N_SUM_c_569_n 0.02017f $X=4.165 $Y=1.385 $X2=0 $Y2=0
cc_328 N_A_394_388#_c_420_n N_SUM_c_569_n 0.0031095f $X=4.355 $Y=1.385 $X2=0
+ $Y2=0
cc_329 N_A_394_388#_M1003_g N_COUT_c_601_n 2.50611e-19 $X=4.355 $Y=2.4 $X2=0
+ $Y2=0
cc_330 N_A_394_388#_c_414_n COUT 0.00104911f $X=4.405 $Y=1.22 $X2=0 $Y2=0
cc_331 N_A_394_388#_c_412_n N_VGND_c_634_n 0.0123991f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_332 N_A_394_388#_c_414_n N_VGND_c_634_n 0.00143104f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_333 N_A_394_388#_c_466_p N_VGND_c_634_n 0.0104044f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_334 N_A_394_388#_c_419_n N_VGND_c_634_n 0.0054838f $X=3.815 $Y=1.385 $X2=0
+ $Y2=0
cc_335 N_A_394_388#_c_412_n N_VGND_c_635_n 0.00143325f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_336 N_A_394_388#_c_414_n N_VGND_c_635_n 0.0106835f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_337 N_A_394_388#_c_412_n N_VGND_c_643_n 0.00383152f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_338 N_A_394_388#_c_414_n N_VGND_c_643_n 0.00383152f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_339 N_A_394_388#_c_412_n N_VGND_c_647_n 0.00758019f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_340 N_A_394_388#_c_414_n N_VGND_c_647_n 0.00758019f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_341 N_A_394_388#_c_415_n N_A_278_74#_M1017_d 0.00884481f $X=3.32 $Y=1.025
+ $X2=0 $Y2=0
cc_342 N_A_394_388#_c_491_p N_A_278_74#_c_705_n 0.0140951f $X=2.72 $Y=0.85 $X2=0
+ $Y2=0
cc_343 N_A_394_388#_c_491_p N_A_278_74#_c_706_n 0.0129062f $X=2.72 $Y=0.85 $X2=0
+ $Y2=0
cc_344 N_A_394_388#_M1017_s N_A_278_74#_c_707_n 0.00297651f $X=2.575 $Y=0.615
+ $X2=0 $Y2=0
cc_345 N_A_394_388#_c_412_n N_A_278_74#_c_707_n 6.04331e-19 $X=3.925 $Y=1.22
+ $X2=0 $Y2=0
cc_346 N_A_394_388#_c_491_p N_A_278_74#_c_707_n 0.0124436f $X=2.72 $Y=0.85 $X2=0
+ $Y2=0
cc_347 N_A_394_388#_c_415_n N_A_278_74#_c_707_n 0.00339819f $X=3.32 $Y=1.025
+ $X2=0 $Y2=0
cc_348 N_A_394_388#_c_412_n N_A_278_74#_c_709_n 0.0013469f $X=3.925 $Y=1.22
+ $X2=0 $Y2=0
cc_349 N_A_394_388#_c_415_n N_A_278_74#_c_709_n 0.0214975f $X=3.32 $Y=1.025
+ $X2=0 $Y2=0
cc_350 N_VPWR_M1003_s N_SUM_c_567_n 0.00228363f $X=4.445 $Y=1.84 $X2=0 $Y2=0
cc_351 N_SUM_c_567_n N_COUT_c_601_n 0.0128877f $X=4.59 $Y=1.82 $X2=0 $Y2=0
cc_352 N_SUM_c_571_n COUT 0.0119219f $X=4.505 $Y=0.965 $X2=0 $Y2=0
cc_353 N_SUM_c_567_n COUT 0.0476603f $X=4.59 $Y=1.82 $X2=0 $Y2=0
cc_354 N_SUM_c_571_n N_VGND_M1012_s 0.00322251f $X=4.505 $Y=0.965 $X2=0 $Y2=0
cc_355 N_SUM_c_567_n N_VGND_M1012_s 5.69077e-19 $X=4.59 $Y=1.82 $X2=0 $Y2=0
cc_356 N_SUM_c_571_n N_VGND_c_635_n 0.0142284f $X=4.505 $Y=0.965 $X2=0 $Y2=0
cc_357 COUT N_VGND_c_635_n 0.0136308f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_358 COUT N_VGND_c_637_n 0.0293763f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_359 COUT N_VGND_c_644_n 0.0144922f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_360 COUT N_VGND_c_647_n 0.0118826f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_361 N_VGND_M1007_d N_A_278_74#_c_705_n 0.00443918f $X=1.82 $Y=0.37 $X2=0
+ $Y2=0
cc_362 N_VGND_c_633_n N_A_278_74#_c_705_n 0.0213709f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_363 N_VGND_c_647_n N_A_278_74#_c_705_n 0.0221192f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_633_n N_A_278_74#_c_706_n 0.0138372f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_365 N_VGND_c_634_n N_A_278_74#_c_707_n 0.0121616f $X=3.71 $Y=0.53 $X2=0 $Y2=0
cc_366 N_VGND_c_642_n N_A_278_74#_c_707_n 0.0561641f $X=3.545 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_647_n N_A_278_74#_c_707_n 0.0315987f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_633_n N_A_278_74#_c_708_n 0.0150383f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_VGND_c_642_n N_A_278_74#_c_708_n 0.0121935f $X=3.545 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_647_n N_A_278_74#_c_708_n 0.00661049f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_634_n N_A_278_74#_c_709_n 0.0191805f $X=3.71 $Y=0.53 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dlclkp_1.pex.spice
* Created: Fri Aug 28 17:25:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%A_83_260# 1 2 9 13 15 16 17 19 20 22 24 25
+ 27 29 31 36
c96 36 0 1.96644e-19 $X=0.6 $Y=1.465
c97 24 0 1.41993e-19 $X=1.47 $Y=2.55
c98 19 0 5.23846e-20 $X=1.385 $Y=2.055
r99 36 39 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.465
+ $X2=0.59 $Y2=1.63
r100 36 38 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.465
+ $X2=0.59 $Y2=1.3
r101 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.465 $X2=0.6 $Y2=1.465
r102 29 31 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.555 $Y=2.715
+ $X2=1.99 $Y2=2.715
r103 25 27 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.555 $Y=0.815
+ $X2=1.98 $Y2=0.815
r104 24 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.47 $Y=2.55
+ $X2=1.555 $Y2=2.715
r105 23 24 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.47 $Y=2.14
+ $X2=1.47 $Y2=2.55
r106 21 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.47 $Y=0.98
+ $X2=1.555 $Y2=0.815
r107 21 22 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.47 $Y=0.98
+ $X2=1.47 $Y2=1.13
r108 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.385 $Y=2.055
+ $X2=1.47 $Y2=2.14
r109 19 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.385 $Y=2.055
+ $X2=0.785 $Y2=2.055
r110 18 35 10.5903 $w=2.88e-07 $l=3.2596e-07 $layer=LI1_cond $X=0.785 $Y=1.215
+ $X2=0.61 $Y2=1.465
r111 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.385 $Y=1.215
+ $X2=1.47 $Y2=1.13
r112 17 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.385 $Y=1.215
+ $X2=0.785 $Y2=1.215
r113 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.97
+ $X2=0.785 $Y2=2.055
r114 15 35 9.02084 $w=2.88e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=1.63
+ $X2=0.61 $Y2=1.465
r115 15 16 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.7 $Y=1.63 $X2=0.7
+ $Y2=1.97
r116 13 38 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.3
r117 9 39 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.63
r118 2 31 600 $w=1.7e-07 $l=8.77553e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.96 $X2=1.99 $Y2=2.715
r119 1 27 182 $w=1.7e-07 $l=5.27304e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.4 $X2=1.98 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%GATE 3 7 9 12
c44 9 0 2.38625e-19 $X=1.2 $Y=1.665
c45 3 0 4.2292e-19 $X=1.215 $Y=2.46
r46 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.635
+ $X2=1.17 $Y2=1.8
r47 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.635
+ $X2=1.17 $Y2=1.47
r48 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.635 $X2=1.17 $Y2=1.635
r49 7 14 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.26 $Y=0.72 $X2=1.26
+ $Y2=1.47
r50 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.215 $Y=2.46
+ $X2=1.215 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%A_315_54# 1 2 7 9 12 16 20 24 25 27 28 31
+ 33 34 38 40 43 47 48 50
c120 31 0 1.94378e-19 $X=2.3 $Y=2.215
c121 28 0 3.01509e-19 $X=1.995 $Y=2.215
c122 25 0 4.19812e-20 $X=1.83 $Y=1.315
c123 24 0 1.803e-19 $X=1.83 $Y=1.315
c124 20 0 1.44503e-20 $X=3.335 $Y=0.995
c125 7 0 1.29101e-19 $X=1.65 $Y=1.15
r126 48 61 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.665
+ $X2=3.27 $Y2=1.83
r127 48 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.665
+ $X2=3.27 $Y2=1.5
r128 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.665 $X2=3.27 $Y2=1.665
r129 44 47 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.115 $Y=1.665
+ $X2=3.27 $Y2=1.665
r130 41 43 10.2439 $w=3.13e-07 $l=2.8e-07 $layer=LI1_cond $X=4.102 $Y=2.39
+ $X2=4.102 $Y2=2.11
r131 40 51 6.12936 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=4.102 $Y=2.102
+ $X2=4.102 $Y2=1.945
r132 40 43 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=4.102 $Y=2.102
+ $X2=4.102 $Y2=2.11
r133 38 51 32.1354 $w=2.58e-07 $l=7.25e-07 $layer=LI1_cond $X=4.075 $Y=1.22
+ $X2=4.075 $Y2=1.945
r134 35 50 3.70735 $w=2.5e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.2 $Y=2.475
+ $X2=3.115 $Y2=2.305
r135 34 41 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=3.945 $Y=2.475
+ $X2=4.102 $Y2=2.39
r136 34 35 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.945 $Y=2.475
+ $X2=3.2 $Y2=2.475
r137 33 50 2.76166 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.115 $Y=2.05
+ $X2=3.115 $Y2=2.305
r138 32 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=1.83
+ $X2=3.115 $Y2=1.665
r139 32 33 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.115 $Y=1.83
+ $X2=3.115 $Y2=2.05
r140 31 58 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=2.215
+ $X2=2.3 $Y2=2.38
r141 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=2.215 $X2=2.3 $Y2=2.215
r142 28 30 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.995 $Y=2.215
+ $X2=2.3 $Y2=2.215
r143 27 50 3.70735 $w=2.5e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.03 $Y=2.215
+ $X2=3.115 $Y2=2.305
r144 27 30 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=3.03 $Y=2.215
+ $X2=2.3 $Y2=2.215
r145 25 52 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.83 $Y=1.315
+ $X2=1.65 $Y2=1.315
r146 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.315 $X2=1.83 $Y2=1.315
r147 22 28 6.90553 $w=3.3e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.86 $Y=2.05
+ $X2=1.995 $Y2=2.215
r148 22 24 31.3721 $w=2.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.86 $Y=2.05
+ $X2=1.86 $Y2=1.315
r149 20 60 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.335 $Y=0.995
+ $X2=3.335 $Y2=1.5
r150 16 61 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.31 $Y=2.41
+ $X2=3.31 $Y2=1.83
r151 12 58 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.345 $Y=2.75
+ $X2=2.345 $Y2=2.38
r152 7 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.15
+ $X2=1.65 $Y2=1.315
r153 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.65 $Y=1.15 $X2=1.65
+ $Y2=0.72
r154 2 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.965 $X2=4.095 $Y2=2.11
r155 1 38 182 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.625 $X2=4.115 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%A_309_338# 1 2 7 9 10 11 14 18 19 21 22 25
+ 28 32 34
c82 32 0 1.11191e-19 $X=3.69 $Y=2.135
c83 28 0 1.85557e-19 $X=3.69 $Y=2.05
c84 14 0 1.23395e-19 $X=2.31 $Y=0.83
r85 30 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.535 $Y=2.135
+ $X2=3.69 $Y2=2.135
r86 28 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.05
+ $X2=3.69 $Y2=2.135
r87 27 34 3.84343 $w=2.4e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.69 $Y=1.33
+ $X2=3.62 $Y2=1.245
r88 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.69 $Y=1.33
+ $X2=3.69 $Y2=2.05
r89 23 34 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.16 $X2=3.62
+ $Y2=1.245
r90 23 25 14.4985 $w=3.08e-07 $l=3.9e-07 $layer=LI1_cond $X=3.62 $Y=1.16
+ $X2=3.62 $Y2=0.77
r91 21 34 2.60907 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.465 $Y=1.245
+ $X2=3.62 $Y2=1.245
r92 21 22 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.465 $Y=1.245
+ $X2=2.535 $Y2=1.245
r93 19 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.37 $Y=1.675 $X2=2.37
+ $Y2=1.765
r94 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.675
+ $X2=2.37 $Y2=1.51
r95 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.675 $X2=2.37 $Y2=1.675
r96 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.37 $Y=1.33
+ $X2=2.535 $Y2=1.245
r97 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.37 $Y=1.33
+ $X2=2.37 $Y2=1.675
r98 14 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.31 $Y=0.83
+ $X2=2.31 $Y2=1.51
r99 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=2.37 $Y2=1.765
r100 10 11 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=1.725 $Y2=1.765
r101 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.635 $Y=1.84
+ $X2=1.725 $Y2=1.765
r102 7 9 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=1.635 $Y=1.84
+ $X2=1.635 $Y2=2.46
r103 2 30 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.99 $X2=3.535 $Y2=2.135
r104 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.625 $X2=3.55 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%CLK 1 3 4 6 9 11 13 14 15 23
c44 23 0 1.11691e-19 $X=4.845 $Y=1.677
c45 15 0 1.36678e-19 $X=5.04 $Y=1.665
c46 1 0 1.85557e-19 $X=4.32 $Y=1.88
r47 23 24 1.83503 $w=3.94e-07 $l=1.5e-08 $layer=POLY_cond $X=4.845 $Y=1.677
+ $X2=4.86 $Y2=1.677
r48 21 23 11.0102 $w=3.94e-07 $l=9e-08 $layer=POLY_cond $X=4.755 $Y=1.677
+ $X2=4.845 $Y2=1.677
r49 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.64 $X2=4.755 $Y2=1.64
r50 19 21 51.3807 $w=3.94e-07 $l=4.2e-07 $layer=POLY_cond $X=4.335 $Y=1.677
+ $X2=4.755 $Y2=1.677
r51 18 19 1.83503 $w=3.94e-07 $l=1.5e-08 $layer=POLY_cond $X=4.32 $Y=1.677
+ $X2=4.335 $Y2=1.677
r52 15 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.04 $Y=1.64
+ $X2=4.755 $Y2=1.64
r53 14 22 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.56 $Y=1.64
+ $X2=4.755 $Y2=1.64
r54 11 24 21.1025 $w=1.8e-07 $l=2.03e-07 $layer=POLY_cond $X=4.86 $Y=1.88
+ $X2=4.86 $Y2=1.677
r55 11 13 135.228 $w=1.8e-07 $l=5.05e-07 $layer=POLY_cond $X=4.86 $Y=1.88
+ $X2=4.86 $Y2=2.385
r56 7 23 25.4929 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=4.845 $Y=1.475
+ $X2=4.845 $Y2=1.677
r57 7 9 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.845 $Y=1.475
+ $X2=4.845 $Y2=0.945
r58 4 19 25.4929 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=4.335 $Y=1.475
+ $X2=4.335 $Y2=1.677
r59 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.335 $Y=1.475
+ $X2=4.335 $Y2=0.995
r60 1 18 21.1025 $w=1.8e-07 $l=2.03e-07 $layer=POLY_cond $X=4.32 $Y=1.88
+ $X2=4.32 $Y2=1.677
r61 1 3 135.228 $w=1.8e-07 $l=5.05e-07 $layer=POLY_cond $X=4.32 $Y=1.88 $X2=4.32
+ $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%A_27_74# 1 2 10 13 17 22 25 29 31 32 34 37
+ 43 45 48 50 51 54 55 57 59 61
c134 57 0 1.37846e-19 $X=2.79 $Y=0.345
c135 54 0 1.19531e-19 $X=0.28 $Y=1.985
c136 45 0 1.29101e-19 $X=1.045 $Y=0.875
c137 34 0 1.36678e-19 $X=5.285 $Y=1.49
c138 31 0 1.11191e-19 $X=2.785 $Y=2.08
r139 58 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.345
+ $X2=2.79 $Y2=0.51
r140 58 61 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.345
+ $X2=2.79 $Y2=0.18
r141 57 59 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0.382
+ $X2=2.625 $Y2=0.382
r142 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=0.345 $X2=2.79 $Y2=0.345
r143 54 55 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=1.82
r144 52 55 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.18 $Y=1.13
+ $X2=0.18 $Y2=1.82
r145 51 52 11.4519 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.27 $Y=0.875
+ $X2=0.27 $Y2=1.13
r146 50 59 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=1.215 $Y=0.34
+ $X2=2.625 $Y2=0.34
r147 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.215 $Y2=0.34
r148 47 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.13 $Y2=0.79
r149 46 51 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=0.875
+ $X2=0.27 $Y2=0.875
r150 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.045 $Y=0.875
+ $X2=1.13 $Y2=0.79
r151 45 46 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.045 $Y=0.875
+ $X2=0.445 $Y2=0.875
r152 41 54 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=1.985
r153 41 43 27.0001 $w=3.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=2.815
r154 35 51 2.79879 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=0.79
+ $X2=0.27 $Y2=0.875
r155 35 37 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.27 $Y=0.79
+ $X2=0.27 $Y2=0.515
r156 33 34 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.285 $Y=1.34
+ $X2=5.285 $Y2=1.49
r157 31 32 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.785 $Y=2.08
+ $X2=2.785 $Y2=2.23
r158 27 29 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.7 $Y=1.19
+ $X2=2.82 $Y2=1.19
r159 25 34 347.895 $w=1.8e-07 $l=8.95e-07 $layer=POLY_cond $X=5.32 $Y=2.385
+ $X2=5.32 $Y2=1.49
r160 22 33 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.235 $Y=0.945
+ $X2=5.235 $Y2=1.34
r161 19 22 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.235 $Y=0.255
+ $X2=5.235 $Y2=0.945
r162 18 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=0.18
+ $X2=2.79 $Y2=0.18
r163 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.16 $Y=0.18
+ $X2=5.235 $Y2=0.255
r164 17 18 1130.65 $w=1.5e-07 $l=2.205e-06 $layer=POLY_cond $X=5.16 $Y=0.18
+ $X2=2.955 $Y2=0.18
r165 15 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.82 $Y=1.265
+ $X2=2.82 $Y2=1.19
r166 15 31 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.82 $Y=1.265
+ $X2=2.82 $Y2=2.08
r167 13 32 202.129 $w=1.8e-07 $l=5.2e-07 $layer=POLY_cond $X=2.765 $Y=2.75
+ $X2=2.765 $Y2=2.23
r168 10 64 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.7 $Y=0.83 $X2=2.7
+ $Y2=0.51
r169 8 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.115 $X2=2.7
+ $Y2=1.19
r170 8 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.7 $Y=1.115
+ $X2=2.7 $Y2=0.83
r171 2 54 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r172 2 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r173 1 37 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%A_990_393# 1 2 9 13 15 16 21 24 27 31 33 35
c63 35 0 1.11691e-19 $X=5.285 $Y=1.12
r64 31 33 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.095 $Y=2.06
+ $X2=5.45 $Y2=2.06
r65 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.87
+ $Y=1.465 $X2=5.87 $Y2=1.465
r66 25 35 0.364692 $w=3.3e-07 $l=4.82571e-07 $layer=LI1_cond $X=5.615 $Y=1.465
+ $X2=5.285 $Y2=1.12
r67 25 27 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.615 $Y=1.465
+ $X2=5.87 $Y2=1.465
r68 24 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=1.975
+ $X2=5.45 $Y2=2.06
r69 23 35 6.46576 $w=2.5e-07 $l=5.86728e-07 $layer=LI1_cond $X=5.45 $Y=1.63
+ $X2=5.285 $Y2=1.12
r70 23 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.45 $Y=1.63
+ $X2=5.45 $Y2=1.975
r71 19 35 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.45 $Y=1.12
+ $X2=5.285 $Y2=1.12
r72 19 21 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.45 $Y=1.12
+ $X2=5.45 $Y2=0.77
r73 15 28 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=6.055 $Y=1.465
+ $X2=5.87 $Y2=1.465
r74 15 16 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.055 $Y=1.465
+ $X2=6.055 $Y2=1.3
r75 11 16 34.7346 $w=1.65e-07 $l=1.7e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=6.055 $Y2=1.3
r76 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=6.225 $Y2=0.74
r77 7 16 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=6.145 $Y=1.63
+ $X2=6.055 $Y2=1.3
r78 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.145 $Y=1.63
+ $X2=6.145 $Y2=2.4
r79 2 31 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.965 $X2=5.095 $Y2=2.14
r80 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.31
+ $Y=0.625 $X2=5.45 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%VPWR 1 2 3 4 15 19 23 27 32 33 34 36 41 49
+ 59 60 63 66 69
r84 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r86 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r88 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 57 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 54 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=4.595 $Y2=3.33
r92 54 56 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 50 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33 $X2=3
+ $Y2=3.33
r96 50 52 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.595 $Y2=3.33
r98 49 52 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r99 48 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r104 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r106 42 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33 $X2=3
+ $Y2=3.33
r108 41 47 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r111 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r112 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 34 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 34 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 32 56 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.705 $Y=3.33
+ $X2=5.52 $Y2=3.33
r116 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.705 $Y=3.33
+ $X2=5.87 $Y2=3.33
r117 31 59 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.035 $Y=3.33
+ $X2=6.48 $Y2=3.33
r118 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.035 $Y=3.33
+ $X2=5.87 $Y2=3.33
r119 27 30 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=5.87 $Y=2.11
+ $X2=5.87 $Y2=2.815
r120 25 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=3.245
+ $X2=5.87 $Y2=3.33
r121 25 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.87 $Y=3.245
+ $X2=5.87 $Y2=2.815
r122 21 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=3.33
r123 21 23 38.5894 $w=3.28e-07 $l=1.105e-06 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=2.14
r124 17 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=3.33
r125 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.815
r126 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r127 13 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.475
r128 4 30 600 $w=1.7e-07 $l=1.05523e-06 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.965 $X2=5.87 $Y2=2.815
r129 4 27 300 $w=1.7e-07 $l=5.27541e-07 $layer=licon1_PDIFF $count=2 $X=5.41
+ $Y=1.965 $X2=5.87 $Y2=2.11
r130 3 23 300 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=1.965 $X2=4.595 $Y2=2.14
r131 2 19 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=2.54 $X2=3 $Y2=2.815
r132 1 15 300 $w=1.7e-07 $l=7.21595e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%GCLK 1 2 9 11 12 13 14 22
r19 14 31 1.15244 $w=3.98e-07 $l=4e-08 $layer=LI1_cond $X=6.405 $Y=2.775
+ $X2=6.405 $Y2=2.815
r20 13 14 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=6.405 $Y=2.405
+ $X2=6.405 $Y2=2.775
r21 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=6.405 $Y=2.035
+ $X2=6.405 $Y2=2.405
r22 12 22 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=6.405 $Y=2.035
+ $X2=6.405 $Y2=1.985
r23 11 34 3.70031 $w=3.98e-07 $l=1.15e-07 $layer=LI1_cond $X=6.405 $Y=1.665
+ $X2=6.405 $Y2=1.55
r24 11 22 6.00917 $w=5.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.405 $Y=1.75
+ $X2=6.405 $Y2=1.985
r25 9 34 36.1448 $w=3.28e-07 $l=1.035e-06 $layer=LI1_cond $X=6.44 $Y=0.515
+ $X2=6.44 $Y2=1.55
r26 2 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.235
+ $Y=1.84 $X2=6.37 $Y2=2.815
r27 2 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.235
+ $Y=1.84 $X2=6.37 $Y2=1.985
r28 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3 $Y=0.37
+ $X2=6.44 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLCLKP_1%VGND 1 2 3 4 15 17 22 25 29 32 33 34 36 48
+ 52 59 60 63 66 69
r83 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r84 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r85 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 60 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r87 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r88 57 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.97
+ $Y2=0
r89 57 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=6.48
+ $Y2=0
r90 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r91 56 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r92 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r93 53 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.55
+ $Y2=0
r94 53 55 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=5.52
+ $Y2=0
r95 52 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.845 $Y=0 $X2=5.97
+ $Y2=0
r96 52 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=0 $X2=5.52
+ $Y2=0
r97 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r98 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r99 48 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=0 $X2=4.55
+ $Y2=0
r100 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.385 $Y=0
+ $X2=4.08 $Y2=0
r101 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r102 44 47 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r103 44 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r104 43 46 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r105 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r106 41 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.75
+ $Y2=0
r107 41 43 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r108 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r109 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 36 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.75
+ $Y2=0
r111 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r112 34 51 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r113 34 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r114 32 46 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.12
+ $Y2=0
r115 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.21
+ $Y2=0
r116 31 50 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.295 $Y=0
+ $X2=4.08 $Y2=0
r117 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.21
+ $Y2=0
r118 27 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0
r119 27 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.515
r120 23 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=0.085
+ $X2=4.55 $Y2=0
r121 23 25 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.55 $Y=0.085
+ $X2=4.55 $Y2=0.77
r122 21 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r123 21 22 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.685
r124 17 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.125 $Y=0.81
+ $X2=3.21 $Y2=0.685
r125 17 19 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.125 $Y=0.81
+ $X2=3.015 $Y2=0.81
r126 13 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r127 13 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.455
r128 4 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.37 $X2=6.01 $Y2=0.515
r129 3 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.625 $X2=4.55 $Y2=0.77
r130 2 19 182 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.62 $X2=3.015 $Y2=0.77
r131 1 15 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.79 $Y2=0.455
.ends


* File: sky130_fd_sc_ms__a31oi_2.spice
* Created: Fri Aug 28 17:07:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a31oi_2.pex.spice"
.subckt sky130_fd_sc_ms__a31oi_2  VNB VPB A3 A2 B1 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* B1	B1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A3_M1006_g N_A_114_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1007 N_A_114_74#_M1006_s N_A2_M1007_g N_A_200_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75003.1 A=0.111 P=1.78 MULT=1
MM1012 N_A_114_74#_M1012_d N_A2_M1012_g N_A_200_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A3_M1011_g N_A_114_74#_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1295 PD=1.16 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.24605 AS=0.1554 PD=1.405 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1000 N_A_200_74#_M1000_d N_A1_M1000_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.24605 PD=1.035 PS=1.405 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1005 N_A_200_74#_M1000_d N_A1_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.2627 PD=1.035 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_368#_M1002_d N_A3_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1568 PD=2.8 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1002_s N_A2_M1003_g N_A_27_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1568 AS=0.1736 PD=1.4 PS=1.43 NRD=0.8668 NRS=6.1464 M=1 R=6.22222
+ SA=90000.6 SB=90003 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_27_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1736 PD=1.44 PS=1.43 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1004 N_A_27_368#_M1004_d N_A3_M1004_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1568 AS=0.1792 PD=1.4 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.6
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g N_A_27_368#_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1013 N_Y_M1009_d N_B1_M1013_g N_A_27_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_27_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1010_d N_A1_M1014_g N_A_27_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX15_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__a31oi_2.pxi.spice"
*
.ends
*
*

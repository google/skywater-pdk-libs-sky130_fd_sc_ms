* File: sky130_fd_sc_ms__o211a_2.pxi.spice
* Created: Wed Sep  2 12:20:08 2020
* 
x_PM_SKY130_FD_SC_MS__O211A_2%C1 N_C1_M1007_g N_C1_c_69_n N_C1_M1011_g C1
+ N_C1_c_71_n PM_SKY130_FD_SC_MS__O211A_2%C1
x_PM_SKY130_FD_SC_MS__O211A_2%B1 N_B1_M1004_g N_B1_M1006_g B1 N_B1_c_94_n
+ N_B1_c_95_n PM_SKY130_FD_SC_MS__O211A_2%B1
x_PM_SKY130_FD_SC_MS__O211A_2%A2 N_A2_M1010_g N_A2_M1005_g A2 N_A2_c_133_n
+ PM_SKY130_FD_SC_MS__O211A_2%A2
x_PM_SKY130_FD_SC_MS__O211A_2%A1 N_A1_M1008_g N_A1_M1000_g A1 N_A1_c_170_n
+ N_A1_c_171_n PM_SKY130_FD_SC_MS__O211A_2%A1
x_PM_SKY130_FD_SC_MS__O211A_2%A_27_368# N_A_27_368#_M1011_s N_A_27_368#_M1007_s
+ N_A_27_368#_M1006_d N_A_27_368#_c_215_n N_A_27_368#_M1001_g
+ N_A_27_368#_c_208_n N_A_27_368#_M1003_g N_A_27_368#_c_209_n
+ N_A_27_368#_M1002_g N_A_27_368#_c_211_n N_A_27_368#_M1009_g
+ N_A_27_368#_c_218_n N_A_27_368#_c_219_n N_A_27_368#_c_226_n
+ N_A_27_368#_c_212_n N_A_27_368#_c_220_n N_A_27_368#_c_248_n
+ N_A_27_368#_c_213_n N_A_27_368#_c_221_n N_A_27_368#_c_214_n
+ N_A_27_368#_c_242_n PM_SKY130_FD_SC_MS__O211A_2%A_27_368#
x_PM_SKY130_FD_SC_MS__O211A_2%VPWR N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_M1002_s
+ N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n VPWR
+ N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n
+ N_VPWR_c_328_n PM_SKY130_FD_SC_MS__O211A_2%VPWR
x_PM_SKY130_FD_SC_MS__O211A_2%X N_X_M1003_d N_X_M1001_d N_X_c_380_n N_X_c_381_n
+ N_X_c_377_n X X X X X PM_SKY130_FD_SC_MS__O211A_2%X
x_PM_SKY130_FD_SC_MS__O211A_2%A_195_74# N_A_195_74#_M1004_d N_A_195_74#_M1000_d
+ N_A_195_74#_c_411_n N_A_195_74#_c_408_n N_A_195_74#_c_409_n
+ PM_SKY130_FD_SC_MS__O211A_2%A_195_74#
x_PM_SKY130_FD_SC_MS__O211A_2%VGND N_VGND_M1010_d N_VGND_M1003_s N_VGND_M1009_s
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND
+ N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n
+ N_VGND_c_444_n PM_SKY130_FD_SC_MS__O211A_2%VGND
cc_1 VNB N_C1_M1007_g 0.00908106f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_2 VNB N_C1_c_69_n 0.0226984f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_3 VNB C1 0.00891253f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_C1_c_71_n 0.0579203f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.385
cc_5 VNB N_B1_M1004_g 0.0246592f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_6 VNB N_B1_c_94_n 0.0217959f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_7 VNB N_B1_c_95_n 0.00613118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_M1010_g 0.0267529f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_9 VNB A2 0.00508898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_133_n 0.0216956f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_11 VNB N_A1_M1000_g 0.0290764f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_12 VNB N_A1_c_170_n 0.0317836f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.385
cc_13 VNB N_A1_c_171_n 0.00231998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_208_n 0.0161558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_368#_c_209_n 0.089659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_368#_M1002_g 0.00671474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_368#_c_211_n 0.0184695f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_18 VNB N_A_27_368#_c_212_n 0.0284016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_368#_c_213_n 0.00677368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_368#_c_214_n 0.0341051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_328_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_377_n 5.40438e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.385
cc_23 VNB X 0.00210995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 8.99291e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_195_74#_c_408_n 0.0028557f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_26 VNB N_A_195_74#_c_409_n 0.00734199f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.385
cc_27 VNB N_VGND_c_435_n 0.00560579f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_28 VNB N_VGND_c_436_n 0.0129885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_437_n 0.0115487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_438_n 0.0510963f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_31 VNB N_VGND_c_439_n 0.0423577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_440_n 0.0210122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_441_n 0.0172134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_442_n 0.00477896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_443_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_444_n 0.236934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_C1_M1007_g 0.031632f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.34
cc_38 VPB N_B1_M1006_g 0.0211858f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_39 VPB N_B1_c_94_n 0.00538978f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_40 VPB N_B1_c_95_n 0.00520645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A2_M1005_g 0.0205116f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_42 VPB A2 0.00410495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A2_c_133_n 0.00539227f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_44 VPB N_A1_M1008_g 0.0232335f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.34
cc_45 VPB N_A1_c_170_n 0.00839136f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.385
cc_46 VPB N_A1_c_171_n 0.00294054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_368#_c_215_n 0.0209853f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_48 VPB N_A_27_368#_c_209_n 0.0130583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_368#_M1002_g 0.0273944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_368#_c_218_n 0.0144246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_27_368#_c_219_n 0.0315273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_368#_c_220_n 0.00292787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_368#_c_221_n 0.00196231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_329_n 0.0198204f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_55 VPB N_VPWR_c_330_n 0.0162037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_331_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_332_n 0.0685527f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_58 VPB N_VPWR_c_333_n 0.0193716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_334_n 0.0325983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_335_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_336_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_337_n 0.0134384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_328_n 0.0785034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_X_c_380_n 0.0032582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_X_c_381_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_66 VPB N_X_c_377_n 0.00116354f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.385
cc_67 N_C1_c_69_n N_B1_M1004_g 0.0568681f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_68 C1 N_B1_M1004_g 6.12064e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_C1_M1007_g N_B1_M1006_g 0.0198491f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_70 N_C1_c_71_n N_B1_c_94_n 0.0203372f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_71 C1 N_B1_c_95_n 0.0164128f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_C1_c_71_n N_B1_c_95_n 0.00879395f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_73 N_C1_M1007_g N_A_27_368#_c_218_n 0.0040552f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_74 C1 N_A_27_368#_c_218_n 0.0196739f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_C1_c_71_n N_A_27_368#_c_218_n 0.00223706f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_76 N_C1_M1007_g N_A_27_368#_c_219_n 0.0107867f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_77 N_C1_M1007_g N_A_27_368#_c_226_n 0.0179323f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_78 N_C1_M1007_g N_A_27_368#_c_220_n 3.80819e-19 $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_79 N_C1_c_69_n N_A_27_368#_c_214_n 0.0264367f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_80 C1 N_A_27_368#_c_214_n 0.0241619f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_C1_c_71_n N_A_27_368#_c_214_n 0.00198571f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_82 N_C1_M1007_g N_VPWR_c_329_n 0.00344602f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_83 N_C1_M1007_g N_VPWR_c_333_n 0.00567889f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_84 N_C1_M1007_g N_VPWR_c_328_n 0.00610055f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_85 N_C1_c_69_n N_VGND_c_439_n 0.00291513f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_86 N_C1_c_69_n N_VGND_c_444_n 0.00362434f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_87 N_B1_M1004_g N_A2_M1010_g 0.0298942f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_88 N_B1_M1006_g N_A2_M1005_g 0.0137343f $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_89 N_B1_M1006_g A2 3.86431e-19 $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_90 N_B1_c_94_n A2 4.14478e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_91 N_B1_c_95_n A2 0.029447f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B1_c_94_n N_A2_c_133_n 0.0214219f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B1_c_95_n N_A2_c_133_n 4.13845e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B1_M1006_g N_A_27_368#_c_218_n 5.99214e-19 $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_95 N_B1_M1006_g N_A_27_368#_c_219_n 3.88951e-19 $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_96 N_B1_M1006_g N_A_27_368#_c_226_n 0.0141191f $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_97 N_B1_c_94_n N_A_27_368#_c_226_n 7.06531e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_98 N_B1_c_95_n N_A_27_368#_c_226_n 0.0353078f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_99 N_B1_M1004_g N_A_27_368#_c_212_n 0.0147907f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B1_c_94_n N_A_27_368#_c_212_n 0.00462669f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B1_c_95_n N_A_27_368#_c_212_n 0.0263338f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_102 N_B1_M1006_g N_A_27_368#_c_220_n 0.00998372f $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_103 N_B1_M1004_g N_A_27_368#_c_214_n 0.00255489f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_104 N_B1_c_95_n N_A_27_368#_c_214_n 0.0153286f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B1_M1006_g N_A_27_368#_c_242_n 5.79575e-19 $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_106 N_B1_c_95_n N_A_27_368#_c_242_n 0.00158553f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B1_M1006_g N_VPWR_c_329_n 0.00349261f $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_108 N_B1_M1006_g N_VPWR_c_334_n 0.005765f $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_109 N_B1_M1006_g N_VPWR_c_328_n 0.00610055f $X=1.035 $Y=2.34 $X2=0 $Y2=0
cc_110 N_B1_M1004_g N_A_195_74#_c_408_n 0.00267731f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_111 N_B1_M1004_g N_VGND_c_439_n 0.00461464f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B1_M1004_g N_VGND_c_444_n 0.00909821f $X=0.9 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A2_M1005_g N_A1_M1008_g 0.055528f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_114 N_A2_M1010_g N_A1_M1000_g 0.0308987f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_115 A2 N_A1_c_170_n 0.00312425f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A2_c_133_n N_A1_c_170_n 0.02078f $X=1.5 $Y=1.515 $X2=0 $Y2=0
cc_117 A2 N_A1_c_171_n 0.0349136f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A2_c_133_n N_A1_c_171_n 2.77744e-19 $X=1.5 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A2_M1010_g N_A_27_368#_c_212_n 0.0114661f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_120 A2 N_A_27_368#_c_212_n 0.0352799f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A2_c_133_n N_A_27_368#_c_212_n 0.00442969f $X=1.5 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A2_M1005_g N_A_27_368#_c_220_n 0.0150264f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_123 N_A2_M1005_g N_A_27_368#_c_248_n 0.0130112f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_124 A2 N_A_27_368#_c_248_n 0.0255673f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_c_133_n N_A_27_368#_c_248_n 3.33288e-19 $X=1.5 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A2_M1005_g N_A_27_368#_c_242_n 8.84614e-19 $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_127 A2 N_A_27_368#_c_242_n 0.00602891f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A2_c_133_n N_A_27_368#_c_242_n 2.83572e-19 $X=1.5 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A2_M1005_g N_VPWR_c_330_n 0.00219965f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_130 N_A2_M1005_g N_VPWR_c_334_n 0.00567889f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_131 N_A2_M1005_g N_VPWR_c_328_n 0.00610055f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_132 N_A2_M1010_g N_A_195_74#_c_411_n 0.00989989f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_M1010_g N_A_195_74#_c_408_n 0.00739554f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A2_M1010_g N_A_195_74#_c_409_n 6.56032e-19 $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A2_M1010_g N_VGND_c_435_n 0.00400267f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A2_M1010_g N_VGND_c_439_n 0.00325937f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A2_M1010_g N_VGND_c_444_n 0.00413498f $X=1.41 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A1_M1008_g N_A_27_368#_c_215_n 0.00602916f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_139 N_A1_M1008_g N_A_27_368#_c_209_n 9.85093e-19 $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_140 N_A1_M1000_g N_A_27_368#_c_209_n 0.00356504f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A1_c_170_n N_A_27_368#_c_209_n 0.021153f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A1_c_171_n N_A_27_368#_c_209_n 9.27871e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A1_M1000_g N_A_27_368#_c_212_n 0.0151825f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_c_170_n N_A_27_368#_c_212_n 0.0025845f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_171_n N_A_27_368#_c_212_n 0.0249861f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A1_M1008_g N_A_27_368#_c_220_n 0.00249437f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_147 N_A1_M1008_g N_A_27_368#_c_248_n 0.020527f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_148 N_A1_c_170_n N_A_27_368#_c_248_n 0.00119851f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A1_c_171_n N_A_27_368#_c_248_n 0.0235732f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A1_M1000_g N_A_27_368#_c_213_n 0.00103826f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A1_c_170_n N_A_27_368#_c_213_n 0.00102181f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A1_c_171_n N_A_27_368#_c_213_n 0.0178205f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A1_M1008_g N_A_27_368#_c_221_n 0.00313163f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_154 N_A1_c_171_n N_A_27_368#_c_221_n 0.00964975f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A1_M1008_g N_VPWR_c_330_n 0.0171459f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_156 N_A1_M1008_g N_VPWR_c_334_n 0.00492916f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_157 N_A1_M1008_g N_VPWR_c_328_n 0.00511769f $X=1.965 $Y=2.34 $X2=0 $Y2=0
cc_158 N_A1_M1000_g N_A_195_74#_c_411_n 0.00966375f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A1_M1000_g N_A_195_74#_c_408_n 6.37625e-19 $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_M1000_g N_A_195_74#_c_409_n 0.00876423f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A1_M1000_g N_VGND_c_435_n 0.0040624f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A1_M1000_g N_VGND_c_436_n 0.00369425f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A1_M1000_g N_VGND_c_440_n 0.00324657f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_M1000_g N_VGND_c_444_n 0.00416919f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_27_368#_c_226_n N_VPWR_M1007_d 0.00505363f $X=1.105 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_166 N_A_27_368#_c_248_n N_VPWR_M1008_d 0.0213148f $X=2.505 $Y=2.035 $X2=0
+ $Y2=0
cc_167 N_A_27_368#_c_221_n N_VPWR_M1008_d 0.00299745f $X=2.59 $Y=1.95 $X2=0
+ $Y2=0
cc_168 N_A_27_368#_c_219_n N_VPWR_c_329_n 0.0221782f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_169 N_A_27_368#_c_226_n N_VPWR_c_329_n 0.0200142f $X=1.105 $Y=2.035 $X2=0
+ $Y2=0
cc_170 N_A_27_368#_c_220_n N_VPWR_c_329_n 0.0221782f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_171 N_A_27_368#_c_215_n N_VPWR_c_330_n 0.00456059f $X=2.835 $Y=1.725 $X2=0
+ $Y2=0
cc_172 N_A_27_368#_c_209_n N_VPWR_c_330_n 0.00140425f $X=3.285 $Y=1.575 $X2=0
+ $Y2=0
cc_173 N_A_27_368#_c_220_n N_VPWR_c_330_n 0.0162312f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_174 N_A_27_368#_c_248_n N_VPWR_c_330_n 0.0493417f $X=2.505 $Y=2.035 $X2=0
+ $Y2=0
cc_175 N_A_27_368#_c_213_n N_VPWR_c_330_n 8.04659e-19 $X=2.59 $Y=1.63 $X2=0
+ $Y2=0
cc_176 N_A_27_368#_c_209_n N_VPWR_c_332_n 0.00135549f $X=3.285 $Y=1.575 $X2=0
+ $Y2=0
cc_177 N_A_27_368#_M1002_g N_VPWR_c_332_n 0.00546761f $X=3.285 $Y=2.4 $X2=0
+ $Y2=0
cc_178 N_A_27_368#_c_219_n N_VPWR_c_333_n 0.00975961f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_179 N_A_27_368#_c_220_n N_VPWR_c_334_n 0.00971074f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_180 N_A_27_368#_c_215_n N_VPWR_c_335_n 0.005209f $X=2.835 $Y=1.725 $X2=0
+ $Y2=0
cc_181 N_A_27_368#_M1002_g N_VPWR_c_335_n 0.005209f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_27_368#_c_215_n N_VPWR_c_328_n 0.00986727f $X=2.835 $Y=1.725 $X2=0
+ $Y2=0
cc_183 N_A_27_368#_M1002_g N_VPWR_c_328_n 0.00985497f $X=3.285 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A_27_368#_c_219_n N_VPWR_c_328_n 0.0111753f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_185 N_A_27_368#_c_220_n N_VPWR_c_328_n 0.0111559f $X=1.27 $Y=2.715 $X2=0
+ $Y2=0
cc_186 N_A_27_368#_c_248_n A_317_368# 0.00917813f $X=2.505 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_27_368#_c_215_n N_X_c_380_n 0.00387883f $X=2.835 $Y=1.725 $X2=0 $Y2=0
cc_188 N_A_27_368#_M1002_g N_X_c_380_n 0.00215936f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_27_368#_c_248_n N_X_c_380_n 0.011477f $X=2.505 $Y=2.035 $X2=0 $Y2=0
cc_190 N_A_27_368#_c_221_n N_X_c_380_n 0.00786825f $X=2.59 $Y=1.95 $X2=0 $Y2=0
cc_191 N_A_27_368#_c_215_n N_X_c_381_n 0.0184403f $X=2.835 $Y=1.725 $X2=0 $Y2=0
cc_192 N_A_27_368#_M1002_g N_X_c_381_n 0.0127634f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_27_368#_c_209_n N_X_c_377_n 0.0166008f $X=3.285 $Y=1.575 $X2=0 $Y2=0
cc_194 N_A_27_368#_M1002_g N_X_c_377_n 0.0122469f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_27_368#_c_221_n N_X_c_377_n 0.00878562f $X=2.59 $Y=1.95 $X2=0 $Y2=0
cc_196 N_A_27_368#_c_208_n X 0.0131366f $X=2.93 $Y=1.185 $X2=0 $Y2=0
cc_197 N_A_27_368#_c_211_n X 0.00191951f $X=3.36 $Y=1.185 $X2=0 $Y2=0
cc_198 N_A_27_368#_c_208_n X 0.00341227f $X=2.93 $Y=1.185 $X2=0 $Y2=0
cc_199 N_A_27_368#_c_213_n X 0.00625242f $X=2.59 $Y=1.63 $X2=0 $Y2=0
cc_200 N_A_27_368#_c_208_n X 5.79411e-19 $X=2.93 $Y=1.185 $X2=0 $Y2=0
cc_201 N_A_27_368#_c_209_n X 0.0205638f $X=3.285 $Y=1.575 $X2=0 $Y2=0
cc_202 N_A_27_368#_c_213_n X 0.0319634f $X=2.59 $Y=1.63 $X2=0 $Y2=0
cc_203 N_A_27_368#_c_212_n N_A_195_74#_M1004_d 0.00261503f $X=2.505 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_204 N_A_27_368#_c_212_n N_A_195_74#_M1000_d 0.0027574f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_205 N_A_27_368#_c_212_n N_A_195_74#_c_411_n 0.0387834f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_206 N_A_27_368#_c_212_n N_A_195_74#_c_408_n 0.0208988f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_207 N_A_27_368#_c_214_n N_A_195_74#_c_408_n 0.0012754f $X=0.295 $Y=0.515
+ $X2=0 $Y2=0
cc_208 N_A_27_368#_c_212_n N_A_195_74#_c_409_n 0.0214503f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_209 N_A_27_368#_c_212_n N_VGND_M1010_d 0.00342819f $X=2.505 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_210 N_A_27_368#_c_213_n N_VGND_M1003_s 0.00210817f $X=2.59 $Y=1.63 $X2=0
+ $Y2=0
cc_211 N_A_27_368#_c_208_n N_VGND_c_436_n 0.00505083f $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_212 N_A_27_368#_c_209_n N_VGND_c_436_n 0.00370338f $X=3.285 $Y=1.575 $X2=0
+ $Y2=0
cc_213 N_A_27_368#_c_213_n N_VGND_c_436_n 0.016027f $X=2.59 $Y=1.63 $X2=0 $Y2=0
cc_214 N_A_27_368#_c_208_n N_VGND_c_438_n 6.08778e-19 $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_215 N_A_27_368#_c_211_n N_VGND_c_438_n 0.015817f $X=3.36 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A_27_368#_c_214_n N_VGND_c_439_n 0.0282878f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_217 N_A_27_368#_c_208_n N_VGND_c_441_n 0.00434272f $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_218 N_A_27_368#_c_211_n N_VGND_c_441_n 0.00383152f $X=3.36 $Y=1.185 $X2=0
+ $Y2=0
cc_219 N_A_27_368#_c_208_n N_VGND_c_444_n 0.00825283f $X=2.93 $Y=1.185 $X2=0
+ $Y2=0
cc_220 N_A_27_368#_c_211_n N_VGND_c_444_n 0.0075754f $X=3.36 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_27_368#_c_214_n N_VGND_c_444_n 0.0230808f $X=0.295 $Y=0.515 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_332_n N_X_c_380_n 0.0450694f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_223 N_VPWR_c_330_n N_X_c_381_n 0.026776f $X=2.56 $Y=2.375 $X2=0 $Y2=0
cc_224 N_VPWR_c_335_n N_X_c_381_n 0.0144623f $X=3.395 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_328_n N_X_c_381_n 0.0118344f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_226 X N_VGND_c_436_n 0.0176099f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_227 X N_VGND_c_438_n 0.0300842f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_228 X N_VGND_c_441_n 0.0112174f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_229 X N_VGND_c_444_n 0.00922837f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_230 N_A_195_74#_c_411_n N_VGND_M1010_d 0.0070032f $X=2.02 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_195_74#_c_411_n N_VGND_c_435_n 0.017876f $X=2.02 $Y=0.755 $X2=0 $Y2=0
cc_232 N_A_195_74#_c_408_n N_VGND_c_435_n 0.00638631f $X=1.19 $Y=0.595 $X2=0
+ $Y2=0
cc_233 N_A_195_74#_c_409_n N_VGND_c_435_n 0.00861021f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
cc_234 N_A_195_74#_c_409_n N_VGND_c_436_n 0.035653f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
cc_235 N_A_195_74#_c_411_n N_VGND_c_439_n 0.00230811f $X=2.02 $Y=0.755 $X2=0
+ $Y2=0
cc_236 N_A_195_74#_c_408_n N_VGND_c_439_n 0.0142392f $X=1.19 $Y=0.595 $X2=0
+ $Y2=0
cc_237 N_A_195_74#_c_411_n N_VGND_c_440_n 0.00340448f $X=2.02 $Y=0.755 $X2=0
+ $Y2=0
cc_238 N_A_195_74#_c_409_n N_VGND_c_440_n 0.0142249f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0
cc_239 N_A_195_74#_c_411_n N_VGND_c_444_n 0.0113875f $X=2.02 $Y=0.755 $X2=0
+ $Y2=0
cc_240 N_A_195_74#_c_408_n N_VGND_c_444_n 0.0118911f $X=1.19 $Y=0.595 $X2=0
+ $Y2=0
cc_241 N_A_195_74#_c_409_n N_VGND_c_444_n 0.011867f $X=2.185 $Y=0.595 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o221a_4.spice
* Created: Fri Aug 28 17:57:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o221a_4.pex.spice"
.subckt sky130_fd_sc_ms__o221a_4  VNB VPB C1 B2 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1012 N_A_27_125#_M1012_d N_C1_M1012_g N_A_114_125#_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1014 N_A_27_125#_M1014_d N_C1_M1014_g N_A_114_125#_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_27_125#_M1014_d N_B1_M1001_g N_A_300_125#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.1008 PD=0.99 PS=0.955 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1004 N_A_300_125#_M1001_s N_B2_M1004_g N_A_27_125#_M1004_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1008 AS=0.1008 PD=0.955 PS=0.955 NRD=6.552 NRS=6.552 M=1 R=4.26667
+ SA=75001.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1025 N_A_300_125#_M1025_d N_B2_M1025_g N_A_27_125#_M1004_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0912 AS=0.1008 PD=0.925 PS=0.955 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_27_125#_M1011_d N_B1_M1011_g N_A_300_125#_M1025_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0.936 M=1 R=4.26667
+ SA=75002.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_300_125#_M1006_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_300_125#_M1006_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75000.6
+ SB=75003.1 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1009_d N_A2_M1010_g N_A_300_125#_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_A1_M1018_g N_A_300_125#_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.142377 AS=0.0896 PD=1.08058 PS=0.92 NRD=15.468 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1018_d N_A_114_125#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.164623 AS=0.10545 PD=1.24942 PS=1.025 NRD=10.536 NRS=0.804 M=1 R=4.93333
+ SA=75001.8 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_114_125#_M1005_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.10545 PD=1.16 PS=1.025 NRD=5.664 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1005_d N_A_114_125#_M1022_g N_X_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_114_125#_M1027_g N_X_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1015 N_A_114_125#_M1015_d N_C1_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90006.9 A=0.18 P=2.36 MULT=1
MM1016 N_A_114_125#_M1015_d N_C1_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.1375 PD=1.27 PS=1.275 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90006.4 A=0.18 P=2.36 MULT=1
MM1008 N_A_300_387#_M1008_d N_B1_M1008_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.1575 AS=0.1375 PD=1.315 PS=1.275 NRD=7.8603 NRS=0 M=1 R=5.55556
+ SA=90001.1 SB=90006 A=0.18 P=2.36 MULT=1
MM1019 N_A_114_125#_M1019_d N_B2_M1019_g N_A_300_387#_M1008_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.1575 PD=1.27 PS=1.315 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90005.5 A=0.18 P=2.36 MULT=1
MM1021 N_A_114_125#_M1019_d N_B2_M1021_g N_A_300_387#_M1021_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1023 N_A_300_387#_M1021_s N_B1_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.3775 PD=1.27 PS=1.755 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.5
+ SB=90004.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_766_387#_M1013_d N_A1_M1013_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1
+ AD=0.1475 AS=0.3775 PD=1.295 PS=1.755 NRD=0 NRS=0 M=1 R=5.55556 SA=90003.4
+ SB=90003.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_114_125#_M1007_d N_A2_M1007_g N_A_766_387#_M1013_d VPB PSHORT L=0.18
+ W=1 AD=0.1475 AS=0.1475 PD=1.295 PS=1.295 NRD=3.9203 NRS=3.9203 M=1 R=5.55556
+ SA=90003.9 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1017 N_A_114_125#_M1007_d N_A2_M1017_g N_A_766_387#_M1017_s VPB PSHORT L=0.18
+ W=1 AD=0.1475 AS=0.16 PD=1.295 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90004.4 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1024 N_A_766_387#_M1017_s N_A1_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.167453 PD=1.32 PS=1.36321 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90004.9 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_114_125#_M1000_g N_VPWR_M1024_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1932 AS=0.187547 PD=1.465 PS=1.52679 NRD=12.2928 NRS=0 M=1 R=6.22222
+ SA=90004.8 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1003 N_X_M1000_d N_A_114_125#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1932 AS=0.1512 PD=1.465 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.3
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1020 N_X_M1020_d N_A_114_125#_M1020_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.182 AS=0.1512 PD=1.445 PS=1.39 NRD=8.7862 NRS=0 M=1 R=6.22222 SA=90005.8
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1026 N_X_M1020_d N_A_114_125#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.182 AS=0.3136 PD=1.445 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_140 VPB 0 1.22796e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__o221a_4.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__dlygate4sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlygate4sd1_1 A VGND VNB VPB VPWR X
M1000 VPWR a_288_74# a_405_138# VPB pshort w=1e+06u l=180000u
+  ad=9.874e+11p pd=6.28e+06u as=5.8e+11p ps=3.16e+06u
M1001 X a_405_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1002 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1003 VGND a_288_74# a_405_138# VNB nlowvt w=420000u l=150000u
+  ad=5.384e+11p pd=4.48e+06u as=2.562e+11p ps=2.06e+06u
M1004 VPWR A a_28_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 X a_405_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1007 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


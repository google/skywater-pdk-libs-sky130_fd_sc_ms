* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2_8 A B VGND VNB VPB VPWR Y
X0 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* NGSPICE file created from sky130_fd_sc_ms__xor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__xor2_1 A B VGND VNB VPB VPWR X
M1000 a_161_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=7.168e+11p ps=5.58e+06u
M1001 a_194_125# B a_161_392# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1002 VGND B a_194_125# VNB nlowvt w=550000u l=150000u
+  ad=8.846e+11p pd=6.8e+06u as=3.5475e+11p ps=2.39e+06u
M1003 VPWR A a_355_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.168e+11p ps=5.76e+06u
M1004 a_455_87# A VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1005 X B a_455_87# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1006 a_355_368# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_194_125# a_355_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.696e+11p pd=2.9e+06u as=0p ps=0u
M1008 a_194_125# A VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_194_125# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


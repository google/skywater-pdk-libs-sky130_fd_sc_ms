* File: sky130_fd_sc_ms__a222o_1.pxi.spice
* Created: Fri Aug 28 17:01:54 2020
* 
x_PM_SKY130_FD_SC_MS__A222O_1%C1 N_C1_M1001_g N_C1_M1005_g C1 C1 N_C1_c_82_n
+ N_C1_c_83_n N_C1_c_84_n PM_SKY130_FD_SC_MS__A222O_1%C1
x_PM_SKY130_FD_SC_MS__A222O_1%C2 N_C2_c_110_n N_C2_M1000_g N_C2_M1009_g C2
+ N_C2_c_113_n PM_SKY130_FD_SC_MS__A222O_1%C2
x_PM_SKY130_FD_SC_MS__A222O_1%B2 N_B2_M1008_g N_B2_M1006_g N_B2_c_149_n
+ N_B2_c_153_n B2 N_B2_c_151_n PM_SKY130_FD_SC_MS__A222O_1%B2
x_PM_SKY130_FD_SC_MS__A222O_1%B1 N_B1_c_197_n N_B1_M1010_g N_B1_M1007_g
+ N_B1_c_193_n B1 B1 N_B1_c_194_n N_B1_c_195_n N_B1_c_196_n
+ PM_SKY130_FD_SC_MS__A222O_1%B1
x_PM_SKY130_FD_SC_MS__A222O_1%A1 N_A1_M1004_g N_A1_M1011_g N_A1_c_234_n
+ N_A1_c_239_n A1 N_A1_c_236_n N_A1_c_237_n PM_SKY130_FD_SC_MS__A222O_1%A1
x_PM_SKY130_FD_SC_MS__A222O_1%A2 N_A2_M1003_g N_A2_M1012_g A2 N_A2_c_270_n
+ N_A2_c_271_n PM_SKY130_FD_SC_MS__A222O_1%A2
x_PM_SKY130_FD_SC_MS__A222O_1%A_32_74# N_A_32_74#_M1005_s N_A_32_74#_M1007_d
+ N_A_32_74#_M1001_d N_A_32_74#_M1013_g N_A_32_74#_M1002_g N_A_32_74#_c_309_n
+ N_A_32_74#_c_320_n N_A_32_74#_c_310_n N_A_32_74#_c_317_n N_A_32_74#_c_348_n
+ N_A_32_74#_c_311_n N_A_32_74#_c_332_n N_A_32_74#_c_312_n N_A_32_74#_c_336_n
+ N_A_32_74#_c_313_n N_A_32_74#_c_314_n N_A_32_74#_c_315_n
+ PM_SKY130_FD_SC_MS__A222O_1%A_32_74#
x_PM_SKY130_FD_SC_MS__A222O_1%A_27_390# N_A_27_390#_M1001_s N_A_27_390#_M1009_d
+ N_A_27_390#_M1010_d N_A_27_390#_c_413_n N_A_27_390#_c_414_n
+ N_A_27_390#_c_415_n N_A_27_390#_c_416_n N_A_27_390#_c_417_n
+ N_A_27_390#_c_418_n N_A_27_390#_c_419_n PM_SKY130_FD_SC_MS__A222O_1%A_27_390#
x_PM_SKY130_FD_SC_MS__A222O_1%A_340_390# N_A_340_390#_M1008_d
+ N_A_340_390#_M1011_d N_A_340_390#_c_456_n N_A_340_390#_c_457_n
+ N_A_340_390#_c_458_n N_A_340_390#_c_459_n
+ PM_SKY130_FD_SC_MS__A222O_1%A_340_390#
x_PM_SKY130_FD_SC_MS__A222O_1%VPWR N_VPWR_M1011_s N_VPWR_M1012_d N_VPWR_c_490_n
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n VPWR N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_489_n N_VPWR_c_497_n PM_SKY130_FD_SC_MS__A222O_1%VPWR
x_PM_SKY130_FD_SC_MS__A222O_1%X N_X_M1002_d N_X_M1013_d N_X_c_538_n N_X_c_539_n
+ X X X X N_X_c_540_n PM_SKY130_FD_SC_MS__A222O_1%X
x_PM_SKY130_FD_SC_MS__A222O_1%VGND N_VGND_M1000_d N_VGND_M1003_d VGND
+ N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n
+ PM_SKY130_FD_SC_MS__A222O_1%VGND
cc_1 VNB N_C1_M1001_g 0.014917f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.45
cc_2 VNB N_C1_c_82_n 0.0415775f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_3 VNB N_C1_c_83_n 0.0243057f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_4 VNB N_C1_c_84_n 0.0238394f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.12
cc_5 VNB N_C2_c_110_n 0.0211034f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.45
cc_6 VNB N_C2_M1009_g 0.0126102f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_7 VNB C2 0.00372322f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_C2_c_113_n 0.0473823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B2_M1006_g 0.0250785f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_B2_c_149_n 0.00756866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B2 0.00699165f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.285
cc_12 VNB N_B2_c_151_n 0.0286514f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.12
cc_13 VNB N_B1_c_193_n 0.0136647f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_B1_c_194_n 0.0401895f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.12
cc_15 VNB N_B1_c_195_n 0.00896147f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.45
cc_16 VNB N_B1_c_196_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.285
cc_17 VNB N_A1_c_234_n 0.0130874f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB A1 0.00802928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_236_n 0.0303908f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_20 VNB N_A1_c_237_n 0.0235136f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.45
cc_21 VNB N_A2_M1012_g 0.0114015f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_22 VNB A2 0.00857517f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_A2_c_270_n 0.0290381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_271_n 0.0188217f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_25 VNB N_A_32_74#_M1013_g 0.00189489f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.285
cc_26 VNB N_A_32_74#_M1002_g 0.0292321f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.45
cc_27 VNB N_A_32_74#_c_309_n 0.0189692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_32_74#_c_310_n 0.00721971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_32_74#_c_311_n 0.00282281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_32_74#_c_312_n 0.00768644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_32_74#_c_313_n 0.00712101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_32_74#_c_314_n 0.00281093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_32_74#_c_315_n 0.0351299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_489_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_538_n 0.0265168f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_X_c_539_n 0.0133911f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_37 VNB N_X_c_540_n 0.0246923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_566_n 0.0703162f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_39 VNB N_VGND_c_567_n 0.0189863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_568_n 0.271043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_569_n 0.0299712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_570_n 0.0244424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_C1_M1001_g 0.0371429f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.45
cc_44 VPB N_C1_c_83_n 0.00822918f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_45 VPB N_C2_M1009_g 0.0293033f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_46 VPB C2 0.00305182f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_47 VPB N_B2_c_149_n 0.0014731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_B2_c_153_n 0.0333842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB B2 0.00262299f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.285
cc_50 VPB N_B1_c_197_n 0.029221f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.45
cc_51 VPB N_B1_c_193_n 0.0086808f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_52 VPB N_B1_c_195_n 0.00739206f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.45
cc_53 VPB N_A1_c_234_n 0.0018398f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_54 VPB N_A1_c_239_n 0.037424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A2_M1012_g 0.0282634f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_56 VPB N_A_32_74#_M1013_g 0.0304608f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.285
cc_57 VPB N_A_32_74#_c_317_n 0.00254837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_32_74#_c_312_n 0.00547856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_27_390#_c_413_n 0.0363365f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.285
cc_60 VPB N_A_27_390#_c_414_n 0.00345944f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.45
cc_61 VPB N_A_27_390#_c_415_n 0.00969566f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.285
cc_62 VPB N_A_27_390#_c_416_n 0.00667471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_390#_c_417_n 0.0074121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_390#_c_418_n 0.00562516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_390#_c_419_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_340_390#_c_456_n 0.0146376f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_67 VPB N_A_340_390#_c_457_n 0.00677663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_340_390#_c_458_n 0.00249873f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_69 VPB N_A_340_390#_c_459_n 0.0067196f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.45
cc_70 VPB N_VPWR_c_490_n 0.0178662f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_71 VPB N_VPWR_c_491_n 0.0155643f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_72 VPB N_VPWR_c_492_n 0.0679541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_493_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_74 VPB N_VPWR_c_494_n 0.0200251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_495_n 0.0189562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_489_n 0.0897449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_497_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB X 0.0133306f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_79 VPB X 0.0413779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_X_c_540_n 0.00766684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 N_C1_c_84_n N_C2_c_110_n 0.0266007f $X=0.407 $Y=1.12 $X2=-0.19 $Y2=-0.245
cc_82 N_C1_M1001_g N_C2_M1009_g 0.0155401f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_83 N_C1_c_82_n N_C2_c_113_n 0.0421408f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_84 N_C1_c_84_n N_A_32_74#_c_309_n 0.00793201f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_85 N_C1_c_83_n N_A_32_74#_c_320_n 0.0059763f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_86 N_C1_c_84_n N_A_32_74#_c_320_n 0.00946381f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_87 N_C1_c_82_n N_A_32_74#_c_310_n 0.00158451f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_88 N_C1_c_83_n N_A_32_74#_c_310_n 0.026304f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_89 N_C1_c_84_n N_A_32_74#_c_310_n 7.14797e-19 $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_90 N_C1_M1001_g N_A_32_74#_c_317_n 0.0068306f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_91 N_C1_c_82_n N_A_32_74#_c_317_n 0.0068306f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_92 N_C1_c_83_n N_A_32_74#_c_312_n 0.0513051f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_93 N_C1_c_84_n N_A_32_74#_c_312_n 0.0068306f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_94 N_C1_M1001_g N_A_27_390#_c_413_n 0.0148218f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_95 N_C1_c_82_n N_A_27_390#_c_413_n 6.60882e-19 $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_96 N_C1_c_83_n N_A_27_390#_c_413_n 0.0263936f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_97 N_C1_M1001_g N_A_27_390#_c_414_n 0.0123263f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_98 N_C1_M1001_g N_A_27_390#_c_415_n 0.00311011f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_99 N_C1_M1001_g N_VPWR_c_492_n 0.00468821f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_100 N_C1_M1001_g N_VPWR_c_489_n 0.00651205f $X=0.505 $Y=2.45 $X2=0 $Y2=0
cc_101 N_C1_c_84_n N_VGND_c_568_n 0.00437003f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_102 N_C1_c_84_n N_VGND_c_569_n 0.00434272f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_103 N_C1_c_84_n N_VGND_c_570_n 0.00126064f $X=0.407 $Y=1.12 $X2=0 $Y2=0
cc_104 C2 N_B2_M1006_g 3.3883e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_C2_c_113_n N_B2_M1006_g 0.0016358f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_106 N_C2_M1009_g N_B2_c_153_n 0.0153398f $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_107 C2 N_B2_c_153_n 5.04794e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_C2_M1009_g B2 6.69477e-19 $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_109 C2 B2 0.0465362f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C2_c_113_n B2 9.0494e-19 $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_111 N_C2_M1009_g N_B2_c_151_n 0.0066094f $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_112 C2 N_B2_c_151_n 0.00116331f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_C2_c_113_n N_B2_c_151_n 0.0175466f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_114 N_C2_c_110_n N_A_32_74#_c_309_n 0.00159871f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_115 N_C2_M1009_g N_A_32_74#_c_317_n 0.0123612f $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_116 N_C2_c_113_n N_A_32_74#_c_317_n 0.00364036f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_117 N_C2_c_110_n N_A_32_74#_c_332_n 0.0040045f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_118 N_C2_c_110_n N_A_32_74#_c_312_n 0.00811889f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_119 C2 N_A_32_74#_c_312_n 0.0475893f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_120 N_C2_c_113_n N_A_32_74#_c_312_n 0.0129514f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_121 N_C2_c_110_n N_A_32_74#_c_336_n 0.0111662f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_122 C2 N_A_32_74#_c_336_n 0.0256857f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_123 N_C2_c_113_n N_A_32_74#_c_336_n 0.00982054f $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_124 N_C2_M1009_g N_A_27_390#_c_413_n 9.45651e-19 $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_125 N_C2_M1009_g N_A_27_390#_c_414_n 0.0150018f $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_126 C2 N_A_27_390#_c_416_n 0.0156932f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_C2_c_113_n N_A_27_390#_c_416_n 6.89403e-19 $X=1.11 $Y=1.285 $X2=0 $Y2=0
cc_128 N_C2_M1009_g N_VPWR_c_492_n 0.0046885f $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_129 N_C2_M1009_g N_VPWR_c_489_n 0.00651205f $X=1.11 $Y=2.45 $X2=0 $Y2=0
cc_130 N_C2_c_110_n N_VGND_c_568_n 0.00369441f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_131 N_C2_c_110_n N_VGND_c_569_n 0.00383152f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_132 N_C2_c_110_n N_VGND_c_570_n 0.0102512f $X=0.91 $Y=1.12 $X2=0 $Y2=0
cc_133 N_B2_c_153_n N_B1_c_197_n 0.0240899f $X=1.635 $Y=1.84 $X2=-0.19
+ $Y2=-0.245
cc_134 N_B2_c_149_n N_B1_c_193_n 0.00738059f $X=1.635 $Y=1.69 $X2=0 $Y2=0
cc_135 B2 N_B1_c_193_n 0.00200975f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B2_c_151_n N_B1_c_193_n 0.012376f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_137 N_B2_M1006_g N_B1_c_194_n 0.012376f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_138 B2 N_B1_c_194_n 0.00122615f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_139 N_B2_M1006_g N_B1_c_195_n 3.3231e-19 $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_140 N_B2_c_149_n N_B1_c_195_n 2.23407e-19 $X=1.635 $Y=1.69 $X2=0 $Y2=0
cc_141 B2 N_B1_c_195_n 0.0307418f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B2_c_151_n N_B1_c_195_n 3.65571e-19 $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_143 N_B2_M1006_g N_B1_c_196_n 0.0467273f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_144 N_B2_c_153_n N_A_32_74#_c_317_n 2.00604e-19 $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_145 N_B2_M1006_g N_A_32_74#_c_336_n 0.0136055f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_146 B2 N_A_32_74#_c_336_n 0.0204678f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B2_c_151_n N_A_32_74#_c_336_n 0.00426176f $X=1.765 $Y=1.345 $X2=0 $Y2=0
cc_148 N_B2_M1006_g N_A_32_74#_c_313_n 0.0016437f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_149 N_B2_c_153_n N_A_27_390#_c_416_n 0.0143035f $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_150 N_B2_c_153_n N_A_27_390#_c_417_n 0.0122641f $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_151 N_B2_c_153_n N_A_27_390#_c_418_n 7.916e-19 $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_152 N_B2_c_153_n N_A_27_390#_c_419_n 0.00223192f $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_153 N_B2_c_153_n N_A_340_390#_c_459_n 8.838e-19 $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_154 B2 N_A_340_390#_c_459_n 0.0192235f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B2_c_151_n N_A_340_390#_c_459_n 8.10809e-19 $X=1.765 $Y=1.345 $X2=0
+ $Y2=0
cc_156 N_B2_c_153_n N_VPWR_c_492_n 0.00468821f $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_157 N_B2_c_153_n N_VPWR_c_489_n 0.00651205f $X=1.635 $Y=1.84 $X2=0 $Y2=0
cc_158 N_B2_M1006_g N_VGND_c_566_n 0.00383152f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_159 N_B2_M1006_g N_VGND_c_568_n 0.00369533f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_160 N_B2_M1006_g N_VGND_c_570_n 0.0101986f $X=1.855 $Y=0.69 $X2=0 $Y2=0
cc_161 N_B1_c_195_n N_A1_c_234_n 0.00933156f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_162 N_B1_c_193_n A1 2.03024e-19 $X=2.2 $Y=1.79 $X2=0 $Y2=0
cc_163 N_B1_c_194_n A1 3.06869e-19 $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_164 N_B1_c_195_n A1 0.0331959f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_165 N_B1_c_194_n N_A1_c_236_n 0.0101376f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_166 N_B1_c_195_n N_A1_c_236_n 0.00134319f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_167 N_B1_c_195_n N_A_32_74#_c_336_n 0.0434877f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_168 N_B1_c_196_n N_A_32_74#_c_336_n 0.00961672f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_169 N_B1_c_194_n N_A_32_74#_c_313_n 0.00162761f $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_170 N_B1_c_196_n N_A_32_74#_c_313_n 0.00978938f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_171 N_B1_c_197_n N_A_27_390#_c_416_n 9.95405e-19 $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_172 N_B1_c_197_n N_A_27_390#_c_417_n 0.0153742f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_173 N_B1_c_197_n N_A_27_390#_c_418_n 0.00936514f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_174 N_B1_c_197_n N_A_340_390#_c_456_n 0.0220843f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_175 N_B1_c_194_n N_A_340_390#_c_456_n 8.177e-19 $X=2.385 $Y=1.285 $X2=0 $Y2=0
cc_176 N_B1_c_195_n N_A_340_390#_c_456_n 0.0419391f $X=2.385 $Y=1.285 $X2=0
+ $Y2=0
cc_177 N_B1_c_197_n N_A_340_390#_c_459_n 0.0100455f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_178 N_B1_c_197_n N_VPWR_c_490_n 0.00175982f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_179 N_B1_c_197_n N_VPWR_c_492_n 0.00468821f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_180 N_B1_c_197_n N_VPWR_c_489_n 0.00651205f $X=2.2 $Y=1.88 $X2=0 $Y2=0
cc_181 N_B1_c_196_n N_VGND_c_566_n 0.00432706f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_182 N_B1_c_196_n N_VGND_c_568_n 0.00438903f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_183 N_B1_c_196_n N_VGND_c_570_n 0.00122056f $X=2.345 $Y=1.12 $X2=0 $Y2=0
cc_184 N_A1_c_234_n N_A2_M1012_g 0.00876246f $X=3.227 $Y=1.69 $X2=0 $Y2=0
cc_185 N_A1_c_239_n N_A2_M1012_g 0.0180859f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_186 N_A1_c_234_n A2 5.72071e-19 $X=3.227 $Y=1.69 $X2=0 $Y2=0
cc_187 A1 A2 0.0253547f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A1_c_236_n A2 0.00148118f $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_189 A1 N_A2_c_270_n 4.13361e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_236_n N_A2_c_270_n 0.0324045f $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_191 N_A1_c_237_n N_A2_c_271_n 0.0324045f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_192 N_A1_c_237_n N_A_32_74#_c_348_n 0.00806212f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_193 A1 N_A_32_74#_c_313_n 0.023365f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A1_c_236_n N_A_32_74#_c_313_n 0.00400401f $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_195 N_A1_c_237_n N_A_32_74#_c_313_n 0.00976723f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_196 N_A1_c_239_n N_A_340_390#_c_456_n 0.0192234f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_197 A1 N_A_340_390#_c_456_n 0.0114042f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A1_c_236_n N_A_340_390#_c_456_n 9.0515e-19 $X=3.09 $Y=1.285 $X2=0 $Y2=0
cc_199 N_A1_c_239_n N_A_340_390#_c_457_n 0.0049331f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_200 N_A1_c_239_n N_A_340_390#_c_458_n 0.0154495f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_201 N_A1_c_239_n N_VPWR_c_490_n 0.00538235f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_202 N_A1_c_239_n N_VPWR_c_494_n 0.00624523f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_203 N_A1_c_239_n N_VPWR_c_489_n 0.006378f $X=3.227 $Y=1.84 $X2=0 $Y2=0
cc_204 N_A1_c_237_n N_VGND_c_566_n 0.00557855f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_205 N_A1_c_237_n N_VGND_c_568_n 0.00438903f $X=3.09 $Y=1.12 $X2=0 $Y2=0
cc_206 N_A2_M1012_g N_A_32_74#_M1013_g 0.021709f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_207 N_A2_c_270_n N_A_32_74#_M1002_g 0.00426644f $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_208 N_A2_c_271_n N_A_32_74#_M1002_g 0.0133207f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_209 A2 N_A_32_74#_c_348_n 0.0228539f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A2_c_270_n N_A_32_74#_c_348_n 0.00452134f $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_211 N_A2_c_271_n N_A_32_74#_c_348_n 0.012296f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_212 A2 N_A_32_74#_c_311_n 0.0124561f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A2_c_270_n N_A_32_74#_c_311_n 6.3503e-19 $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_214 N_A2_c_271_n N_A_32_74#_c_311_n 0.00310754f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_215 N_A2_c_271_n N_A_32_74#_c_313_n 0.00162108f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_216 N_A2_M1012_g N_A_32_74#_c_314_n 0.00221602f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_217 A2 N_A_32_74#_c_314_n 0.0183844f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A2_c_270_n N_A_32_74#_c_314_n 5.13863e-19 $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_219 N_A2_M1012_g N_A_32_74#_c_315_n 0.00951623f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_220 A2 N_A_32_74#_c_315_n 4.88188e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A2_c_270_n N_A_32_74#_c_315_n 0.00945972f $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_222 N_A2_M1012_g N_A_340_390#_c_457_n 0.00374986f $X=3.71 $Y=2.415 $X2=0
+ $Y2=0
cc_223 A2 N_A_340_390#_c_457_n 0.00872764f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_224 N_A2_c_270_n N_A_340_390#_c_457_n 7.51809e-19 $X=3.66 $Y=1.285 $X2=0
+ $Y2=0
cc_225 N_A2_M1012_g N_A_340_390#_c_458_n 0.0103697f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_226 N_A2_M1012_g N_VPWR_c_491_n 0.00958834f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_227 N_A2_M1012_g N_VPWR_c_494_n 0.00624523f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_228 N_A2_M1012_g N_VPWR_c_489_n 0.006378f $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_229 N_A2_M1012_g X 5.48264e-19 $X=3.71 $Y=2.415 $X2=0 $Y2=0
cc_230 N_A2_c_271_n N_VGND_c_566_n 0.0178758f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_231 N_A2_c_271_n N_VGND_c_568_n 0.00371083f $X=3.66 $Y=1.12 $X2=0 $Y2=0
cc_232 N_A_32_74#_c_317_n N_A_27_390#_c_413_n 0.0415807f $X=0.885 $Y=2.095 $X2=0
+ $Y2=0
cc_233 N_A_32_74#_M1001_d N_A_27_390#_c_414_n 0.00536354f $X=0.595 $Y=1.95 $X2=0
+ $Y2=0
cc_234 N_A_32_74#_c_317_n N_A_27_390#_c_414_n 0.0204485f $X=0.885 $Y=2.095 $X2=0
+ $Y2=0
cc_235 N_A_32_74#_c_317_n N_A_27_390#_c_416_n 0.0309585f $X=0.885 $Y=2.095 $X2=0
+ $Y2=0
cc_236 N_A_32_74#_M1013_g N_VPWR_c_491_n 0.00413104f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_32_74#_c_314_n N_VPWR_c_491_n 0.00886523f $X=4.205 $Y=1.465 $X2=0
+ $Y2=0
cc_238 N_A_32_74#_c_315_n N_VPWR_c_491_n 0.00304496f $X=4.205 $Y=1.465 $X2=0
+ $Y2=0
cc_239 N_A_32_74#_M1013_g N_VPWR_c_495_n 0.005209f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A_32_74#_M1013_g N_VPWR_c_489_n 0.00990469f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_32_74#_M1002_g N_X_c_538_n 0.0138767f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_32_74#_c_311_n N_X_c_538_n 0.00750685f $X=4.1 $Y=1.3 $X2=0 $Y2=0
cc_243 N_A_32_74#_M1002_g N_X_c_539_n 0.00299691f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_32_74#_c_314_n N_X_c_539_n 0.00111755f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_245 N_A_32_74#_c_315_n N_X_c_539_n 2.41927e-19 $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_246 N_A_32_74#_M1013_g X 0.00412821f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_32_74#_c_314_n X 0.00102175f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_248 N_A_32_74#_M1013_g X 0.0128933f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_32_74#_M1002_g N_X_c_540_n 0.00255192f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_32_74#_c_311_n N_X_c_540_n 0.00541114f $X=4.1 $Y=1.3 $X2=0 $Y2=0
cc_251 N_A_32_74#_c_314_n N_X_c_540_n 0.0249107f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_252 N_A_32_74#_c_315_n N_X_c_540_n 0.0125816f $X=4.205 $Y=1.465 $X2=0 $Y2=0
cc_253 N_A_32_74#_c_320_n A_119_74# 0.00383368f $X=0.72 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_254 N_A_32_74#_c_332_n A_119_74# 0.00130602f $X=0.805 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_255 N_A_32_74#_c_312_n A_119_74# 6.66187e-19 $X=0.885 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_256 N_A_32_74#_c_336_n N_VGND_M1000_d 0.0224135f $X=2.295 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_257 N_A_32_74#_c_348_n N_VGND_M1003_d 0.0163508f $X=4.015 $Y=0.865 $X2=0
+ $Y2=0
cc_258 N_A_32_74#_c_311_n N_VGND_M1003_d 0.00355979f $X=4.1 $Y=1.3 $X2=0 $Y2=0
cc_259 N_A_32_74#_M1002_g N_VGND_c_566_n 0.00583725f $X=4.305 $Y=0.74 $X2=0
+ $Y2=0
cc_260 N_A_32_74#_c_348_n N_VGND_c_566_n 0.0401368f $X=4.015 $Y=0.865 $X2=0
+ $Y2=0
cc_261 N_A_32_74#_c_313_n N_VGND_c_566_n 0.0496465f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_262 N_A_32_74#_c_315_n N_VGND_c_566_n 4.00439e-19 $X=4.205 $Y=1.465 $X2=0
+ $Y2=0
cc_263 N_A_32_74#_M1002_g N_VGND_c_567_n 0.00434272f $X=4.305 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_32_74#_M1002_g N_VGND_c_568_n 0.00826002f $X=4.305 $Y=0.74 $X2=0
+ $Y2=0
cc_265 N_A_32_74#_c_309_n N_VGND_c_568_n 0.0119472f $X=0.305 $Y=0.515 $X2=0
+ $Y2=0
cc_266 N_A_32_74#_c_320_n N_VGND_c_568_n 0.0081717f $X=0.72 $Y=0.865 $X2=0 $Y2=0
cc_267 N_A_32_74#_c_348_n N_VGND_c_568_n 0.0180838f $X=4.015 $Y=0.865 $X2=0
+ $Y2=0
cc_268 N_A_32_74#_c_332_n N_VGND_c_568_n 0.00663982f $X=0.805 $Y=0.865 $X2=0
+ $Y2=0
cc_269 N_A_32_74#_c_336_n N_VGND_c_568_n 0.0210815f $X=2.295 $Y=0.64 $X2=0 $Y2=0
cc_270 N_A_32_74#_c_313_n N_VGND_c_568_n 0.0308511f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_271 N_A_32_74#_c_309_n N_VGND_c_569_n 0.0144324f $X=0.305 $Y=0.515 $X2=0
+ $Y2=0
cc_272 N_A_32_74#_c_309_n N_VGND_c_570_n 0.00836615f $X=0.305 $Y=0.515 $X2=0
+ $Y2=0
cc_273 N_A_32_74#_c_336_n N_VGND_c_570_n 0.0545917f $X=2.295 $Y=0.64 $X2=0 $Y2=0
cc_274 N_A_32_74#_c_313_n N_VGND_c_570_n 0.00952048f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_275 N_A_32_74#_c_336_n A_386_74# 0.0072096f $X=2.295 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_32_74#_c_348_n A_651_74# 0.0072096f $X=4.015 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_27_390#_c_417_n N_A_340_390#_M1008_d 0.00322579f $X=2.26 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_278 N_A_27_390#_M1010_d N_A_340_390#_c_456_n 0.00543715f $X=2.29 $Y=1.95
+ $X2=0 $Y2=0
cc_279 N_A_27_390#_c_418_n N_A_340_390#_c_456_n 0.0219147f $X=2.425 $Y=2.465
+ $X2=0 $Y2=0
cc_280 N_A_27_390#_c_416_n N_A_340_390#_c_459_n 0.00833462f $X=1.385 $Y=2.095
+ $X2=0 $Y2=0
cc_281 N_A_27_390#_c_417_n N_A_340_390#_c_459_n 0.022225f $X=2.26 $Y=2.99 $X2=0
+ $Y2=0
cc_282 N_A_27_390#_c_418_n N_A_340_390#_c_459_n 0.0287016f $X=2.425 $Y=2.465
+ $X2=0 $Y2=0
cc_283 N_A_27_390#_c_417_n N_VPWR_c_490_n 0.0121617f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_284 N_A_27_390#_c_418_n N_VPWR_c_490_n 0.0407547f $X=2.425 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_27_390#_c_414_n N_VPWR_c_492_n 0.0489082f $X=1.22 $Y=2.99 $X2=0 $Y2=0
cc_286 N_A_27_390#_c_415_n N_VPWR_c_492_n 0.0235512f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_287 N_A_27_390#_c_417_n N_VPWR_c_492_n 0.0683624f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_288 N_A_27_390#_c_419_n N_VPWR_c_492_n 0.0235512f $X=1.385 $Y=2.99 $X2=0
+ $Y2=0
cc_289 N_A_27_390#_c_414_n N_VPWR_c_489_n 0.0289441f $X=1.22 $Y=2.99 $X2=0 $Y2=0
cc_290 N_A_27_390#_c_415_n N_VPWR_c_489_n 0.0128119f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_27_390#_c_417_n N_VPWR_c_489_n 0.0393297f $X=2.26 $Y=2.99 $X2=0 $Y2=0
cc_292 N_A_27_390#_c_419_n N_VPWR_c_489_n 0.0128119f $X=1.385 $Y=2.99 $X2=0
+ $Y2=0
cc_293 N_A_340_390#_c_456_n N_VPWR_M1011_s 0.0102346f $X=3.32 $Y=2.045 $X2=-0.19
+ $Y2=1.66
cc_294 N_A_340_390#_c_456_n N_VPWR_c_490_n 0.0238156f $X=3.32 $Y=2.045 $X2=0
+ $Y2=0
cc_295 N_A_340_390#_c_458_n N_VPWR_c_490_n 0.0246172f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_296 N_A_340_390#_c_457_n N_VPWR_c_491_n 0.00896489f $X=3.485 $Y=2.13 $X2=0
+ $Y2=0
cc_297 N_A_340_390#_c_458_n N_VPWR_c_491_n 0.026664f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_298 N_A_340_390#_c_458_n N_VPWR_c_494_n 0.0122272f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_299 N_A_340_390#_c_458_n N_VPWR_c_489_n 0.0117276f $X=3.485 $Y=2.77 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_491_n X 0.0419219f $X=4.02 $Y=2.06 $X2=0 $Y2=0
cc_301 N_VPWR_c_495_n X 0.0156645f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_c_489_n X 0.0128976f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_303 N_X_c_538_n N_VGND_c_566_n 0.0107229f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_304 N_X_c_538_n N_VGND_c_567_n 0.0156794f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_305 N_X_c_538_n N_VGND_c_568_n 0.0129217f $X=4.52 $Y=0.515 $X2=0 $Y2=0

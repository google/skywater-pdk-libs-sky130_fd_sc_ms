* NGSPICE file created from sky130_fd_sc_ms__sdfxtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sdfxtp_2 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_1707_496# a_846_74# a_1595_424# VPB pshort w=420000u l=180000u
+  ad=2.562e+11p pd=2.06e+06u as=2.754e+11p ps=2.44e+06u
M1001 a_1044_100# a_634_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=3.045e+11p pd=2.29e+06u as=3.528e+11p ps=3.36e+06u
M1002 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=2.72693e+12p pd=2.061e+07u as=1.792e+11p ps=1.84e+06u
M1003 a_1595_424# a_634_74# a_1287_320# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.2e+11p ps=2.68e+06u
M1004 VGND SCD a_442_74# VNB nlowvt w=420000u l=150000u
+  ad=1.84785e+12p pd=1.542e+07u as=1.008e+11p ps=1.32e+06u
M1005 VGND a_1829_398# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.13e+06u
M1006 a_301_74# D a_219_453# VPB pshort w=640000u l=180000u
+  ad=4.472e+11p pd=3.71e+06u as=1.536e+11p ps=1.76e+06u
M1007 a_1219_100# a_846_74# a_1044_100# VNB nlowvt w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=0p ps=0u
M1008 a_1287_320# a_1044_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=3.795e+11p pd=2.48e+06u as=0p ps=0u
M1009 a_1829_398# a_1595_424# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1010 VGND a_1287_320# a_1219_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1595_424# a_846_74# a_1287_320# VNB nlowvt w=550000u l=150000u
+  ad=1.8825e+11p pd=1.82e+06u as=0p ps=0u
M1012 a_634_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1013 a_442_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_1829_398# a_1707_496# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_223_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1016 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1829_398# a_1595_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 VPWR SCD a_442_453# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1019 a_846_74# a_634_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 VPWR a_1287_320# a_1213_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.554e+11p ps=1.58e+06u
M1021 a_1787_74# a_634_74# a_1595_424# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1022 VGND a_1829_398# a_1787_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1044_100# a_846_74# a_301_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1024 Q a_1829_398# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1213_508# a_634_74# a_1044_100# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_1829_398# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 a_1287_320# a_1044_100# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_1829_398# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_442_453# a_27_74# a_301_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_846_74# a_634_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1031 a_634_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1032 a_219_453# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
.ends


* File: sky130_fd_sc_ms__or2b_2.pex.spice
* Created: Fri Aug 28 18:06:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR2B_2%B_N 3 7 9 12 13
c29 7 0 1.58544e-19 $X=0.5 $Y=0.835
c30 3 0 8.6078e-20 $X=0.505 $Y=2.26
r31 12 15 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.515
+ $X2=0.407 $Y2=1.68
r32 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.515
+ $X2=0.407 $Y2=1.35
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r34 9 13 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r35 7 14 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.5 $Y=0.835 $X2=0.5
+ $Y2=1.35
r36 3 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.505 $Y=2.26
+ $X2=0.505 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_2%A_187_48# 1 2 9 13 17 21 25 26 29 31 35 40 41
+ 42 44 46 47
r107 49 50 59.8804 $w=3.26e-07 $l=4.05e-07 $layer=POLY_cond $X=1.04 $Y=1.465
+ $X2=1.445 $Y2=1.465
r108 48 49 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=1.01 $Y=1.465
+ $X2=1.04 $Y2=1.465
r109 46 47 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=1.985
+ $X2=3.075 $Y2=1.82
r110 41 52 11.089 $w=3.26e-07 $l=7.5e-08 $layer=POLY_cond $X=1.63 $Y=1.465
+ $X2=1.705 $Y2=1.465
r111 41 50 27.3528 $w=3.26e-07 $l=1.85e-07 $layer=POLY_cond $X=1.63 $Y=1.465
+ $X2=1.445 $Y2=1.465
r112 40 42 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=1.465
+ $X2=1.63 $Y2=1.3
r113 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.465 $X2=1.63 $Y2=1.465
r114 37 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=1.15
+ $X2=3.19 $Y2=1.82
r115 33 46 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.075 $Y2=1.985
r116 33 35 19.4475 $w=3.98e-07 $l=6.75e-07 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.075 $Y2=2.695
r117 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=1.065
+ $X2=2.57 $Y2=1.065
r118 31 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=1.065
+ $X2=3.19 $Y2=1.15
r119 31 32 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.065
+ $X2=2.735 $Y2=1.065
r120 27 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0.98
+ $X2=2.57 $Y2=1.065
r121 27 29 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.57 $Y=0.98
+ $X2=2.57 $Y2=0.515
r122 25 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=1.065
+ $X2=2.57 $Y2=1.065
r123 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.405 $Y=1.065
+ $X2=1.795 $Y2=1.065
r124 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.71 $Y=1.15
+ $X2=1.795 $Y2=1.065
r125 23 42 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.15
+ $X2=1.71 $Y2=1.3
r126 19 52 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.63
+ $X2=1.705 $Y2=1.465
r127 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.705 $Y=1.63
+ $X2=1.705 $Y2=2.4
r128 15 50 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.3
+ $X2=1.445 $Y2=1.465
r129 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.445 $Y=1.3
+ $X2=1.445 $Y2=0.74
r130 11 49 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.63
+ $X2=1.04 $Y2=1.465
r131 11 13 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.04 $Y=1.63
+ $X2=1.04 $Y2=2.4
r132 7 48 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.3 $X2=1.01
+ $Y2=1.465
r133 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.01 $Y=1.3 $X2=1.01
+ $Y2=0.74
r134 2 46 400 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=3.04 $Y2=1.985
r135 2 35 400 $w=1.7e-07 $l=9.74192e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=3.04 $Y2=2.695
r136 1 29 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.37 $X2=2.57 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_2%A 3 7 9 12 13
c38 13 0 1.44053e-19 $X=2.2 $Y=1.515
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.515
+ $X2=2.2 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.515
+ $X2=2.2 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.2
+ $Y=1.515 $X2=2.2 $Y2=1.515
r42 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=1.515
r43 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.29 $Y=0.69 $X2=2.29
+ $Y2=1.35
r44 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.275 $Y=2.34
+ $X2=2.275 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_2%A_27_368# 1 2 9 13 17 19 20 22 23 24 26 33 34
c92 9 0 1.44053e-19 $X=2.695 $Y=2.34
r93 34 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.485
+ $X2=2.77 $Y2=1.65
r94 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.485
+ $X2=2.77 $Y2=1.32
r95 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.485 $X2=2.77 $Y2=1.485
r96 30 33 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.62 $Y=1.485
+ $X2=2.77 $Y2=1.485
r97 28 29 10.9863 $w=5.83e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=2.325
+ $X2=0.805 $Y2=2.325
r98 25 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=1.65
+ $X2=2.62 $Y2=1.485
r99 25 26 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.62 $Y=1.65 $X2=2.62
+ $Y2=2.24
r100 24 29 8.57219 $w=5.83e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=2.325
+ $X2=0.805 $Y2=2.325
r101 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.535 $Y=2.325
+ $X2=2.62 $Y2=2.24
r102 23 24 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=2.535 $Y=2.325
+ $X2=0.89 $Y2=2.325
r103 22 29 8.13184 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=2.325
r104 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.805 $Y2=1.95
r105 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.805 $Y2=1.18
r106 19 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.45 $Y2=1.095
r107 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.45 $Y2=1.095
r108 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.285 $Y2=0.835
r109 13 37 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.785 $Y=0.69
+ $X2=2.785 $Y2=1.32
r110 9 38 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=2.695 $Y=2.34
+ $X2=2.695 $Y2=1.65
r111 2 28 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r112 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.56 $X2=0.285 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_2%VPWR 1 2 11 15 18 19 20 30 31 34
r34 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r38 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r40 22 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r41 20 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 20 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 20 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 18 24 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r46 17 27 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r48 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r49 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.78
r50 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r51 9 11 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.78
r52 2 15 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.84 $X2=1.93 $Y2=2.78
r53 1 11 600 $w=1.7e-07 $l=1.04422e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_2%X 1 2 8 9 11 13 14 25
c37 14 0 1.16427e-19 $X=1.115 $Y=0.84
c38 9 0 8.6078e-20 $X=1.23 $Y=1.945
c39 8 0 4.21169e-20 $X=1.145 $Y=1.82
r40 18 25 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.225 $Y=0.965
+ $X2=1.225 $Y2=0.925
r41 14 27 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=1.225 $Y=0.987
+ $X2=1.225 $Y2=1.13
r42 14 18 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=1.225 $Y=0.987
+ $X2=1.225 $Y2=0.965
r43 14 25 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=1.225 $Y=0.902
+ $X2=1.225 $Y2=0.925
r44 13 14 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=1.225 $Y=0.515
+ $X2=1.225 $Y2=0.902
r45 9 11 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.23 $Y=1.945
+ $X2=1.37 $Y2=1.945
r46 8 9 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.145 $Y=1.82
+ $X2=1.23 $Y2=1.945
r47 8 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.145 $Y=1.82
+ $X2=1.145 $Y2=1.13
r48 2 11 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.37 $Y2=1.985
r49 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.37 $X2=1.225 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r47 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r50 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 35 43 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=1.897
+ $Y2=0
r52 35 37 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.64
+ $Y2=0
r53 34 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r54 34 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r55 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r56 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 30 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.755
+ $Y2=0
r58 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r59 29 43 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.897
+ $Y2=0
r60 29 32 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.2
+ $Y2=0
r61 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 24 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.755
+ $Y2=0
r64 24 26 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r65 22 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r66 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r67 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 18 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r69 18 20 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.645
r70 14 43 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.897 $Y=0.085
+ $X2=1.897 $Y2=0
r71 14 16 9.92302 $w=6.73e-07 $l=5.6e-07 $layer=LI1_cond $X=1.897 $Y=0.085
+ $X2=1.897 $Y2=0.645
r72 10 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r73 10 12 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.675
r74 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.37 $X2=3 $Y2=0.645
r75 2 16 91 $w=1.7e-07 $l=6.7361e-07 $layer=licon1_NDIFF $count=2 $X=1.52
+ $Y=0.37 $X2=2.07 $Y2=0.645
r76 1 12 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.675
.ends


* File: sky130_fd_sc_ms__o31ai_2.pxi.spice
* Created: Fri Aug 28 18:03:00 2020
* 
x_PM_SKY130_FD_SC_MS__O31AI_2%A1 N_A1_M1013_g N_A1_M1000_g N_A1_M1001_g
+ N_A1_c_82_n N_A1_M1015_g A1 A1 A1 N_A1_c_84_n PM_SKY130_FD_SC_MS__O31AI_2%A1
x_PM_SKY130_FD_SC_MS__O31AI_2%A2 N_A2_c_134_n N_A2_M1002_g N_A2_M1006_g
+ N_A2_c_135_n N_A2_M1004_g N_A2_M1010_g A2 A2 N_A2_c_133_n
+ PM_SKY130_FD_SC_MS__O31AI_2%A2
x_PM_SKY130_FD_SC_MS__O31AI_2%A3 N_A3_M1003_g N_A3_c_186_n N_A3_M1009_g
+ N_A3_M1011_g N_A3_M1005_g A3 N_A3_c_188_n N_A3_c_189_n N_A3_c_190_n
+ PM_SKY130_FD_SC_MS__O31AI_2%A3
x_PM_SKY130_FD_SC_MS__O31AI_2%B1 N_B1_M1007_g N_B1_M1012_g N_B1_M1008_g
+ N_B1_M1014_g N_B1_c_250_n B1 N_B1_c_252_n PM_SKY130_FD_SC_MS__O31AI_2%B1
x_PM_SKY130_FD_SC_MS__O31AI_2%A_28_368# N_A_28_368#_M1000_s N_A_28_368#_M1001_s
+ N_A_28_368#_M1004_s N_A_28_368#_c_303_n N_A_28_368#_c_304_n
+ N_A_28_368#_c_309_n N_A_28_368#_c_305_n N_A_28_368#_c_319_n
+ N_A_28_368#_c_315_n N_A_28_368#_c_306_n PM_SKY130_FD_SC_MS__O31AI_2%A_28_368#
x_PM_SKY130_FD_SC_MS__O31AI_2%VPWR N_VPWR_M1000_d N_VPWR_M1012_d N_VPWR_c_344_n
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n VPWR N_VPWR_c_348_n
+ N_VPWR_c_349_n N_VPWR_c_343_n N_VPWR_c_351_n PM_SKY130_FD_SC_MS__O31AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O31AI_2%A_300_368# N_A_300_368#_M1002_d
+ N_A_300_368#_M1009_d N_A_300_368#_c_402_n N_A_300_368#_c_392_n
+ N_A_300_368#_c_393_n N_A_300_368#_c_398_n
+ PM_SKY130_FD_SC_MS__O31AI_2%A_300_368#
x_PM_SKY130_FD_SC_MS__O31AI_2%Y N_Y_M1007_d N_Y_M1009_s N_Y_M1011_s N_Y_M1014_s
+ N_Y_c_418_n N_Y_c_415_n N_Y_c_416_n N_Y_c_430_n N_Y_c_449_n N_Y_c_434_n
+ N_Y_c_419_n N_Y_c_420_n N_Y_c_421_n N_Y_c_417_n N_Y_c_444_n Y Y
+ PM_SKY130_FD_SC_MS__O31AI_2%Y
x_PM_SKY130_FD_SC_MS__O31AI_2%A_27_74# N_A_27_74#_M1013_s N_A_27_74#_M1015_s
+ N_A_27_74#_M1010_s N_A_27_74#_M1005_s N_A_27_74#_M1008_s N_A_27_74#_c_490_n
+ N_A_27_74#_c_491_n N_A_27_74#_c_492_n N_A_27_74#_c_493_n N_A_27_74#_c_494_n
+ N_A_27_74#_c_518_n N_A_27_74#_c_525_n N_A_27_74#_c_529_n N_A_27_74#_c_495_n
+ N_A_27_74#_c_496_n N_A_27_74#_c_497_n N_A_27_74#_c_498_n N_A_27_74#_c_499_n
+ PM_SKY130_FD_SC_MS__O31AI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O31AI_2%VGND N_VGND_M1013_d N_VGND_M1006_d N_VGND_M1003_d
+ N_VGND_c_571_n N_VGND_c_572_n N_VGND_c_573_n VGND N_VGND_c_574_n
+ N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n
+ N_VGND_c_580_n PM_SKY130_FD_SC_MS__O31AI_2%VGND
cc_1 VNB N_A1_M1013_g 0.0339584f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_c_82_n 0.0157773f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.185
cc_3 VNB A1 0.0218337f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_A1_c_84_n 0.0578087f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.432
cc_5 VNB N_A2_M1006_g 0.0254433f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_6 VNB N_A2_M1010_g 0.0253921f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.185
cc_7 VNB A2 0.00408815f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A2_c_133_n 0.0493981f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.432
cc_9 VNB N_A3_M1003_g 0.0254342f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A3_c_186_n 0.0119391f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_11 VNB N_A3_M1005_g 0.0262448f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_A3_c_188_n 0.0144872f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.432
cc_13 VNB N_A3_c_189_n 0.00217772f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_14 VNB N_A3_c_190_n 0.0395308f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.432
cc_15 VNB N_B1_M1007_g 0.0205226f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_B1_M1008_g 0.0255449f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_17 VNB N_B1_c_250_n 0.00219487f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB B1 0.0102709f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.432
cc_19 VNB N_B1_c_252_n 0.0843705f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.185
cc_20 VNB N_VPWR_c_343_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_415_n 0.0147535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_416_n 8.30186e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_417_n 0.00570061f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_24 VNB N_A_27_74#_c_490_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_25 VNB N_A_27_74#_c_491_n 0.00263637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_492_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_493_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.432
cc_28 VNB N_A_27_74#_c_494_n 0.010404f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_29 VNB N_A_27_74#_c_495_n 0.0126811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_496_n 0.00163372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_497_n 0.0222992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_498_n 0.00322614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_499_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_571_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_572_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_36 VNB N_VGND_c_573_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_37 VNB N_VGND_c_574_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.432
cc_38 VNB N_VGND_c_575_n 0.0387921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_576_n 0.271117f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_40 VNB N_VGND_c_577_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_578_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_579_n 0.0182584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_580_n 0.0206062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_A1_M1000_g 0.0267788f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_45 VPB N_A1_M1001_g 0.0208126f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_46 VPB A1 0.0142305f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_47 VPB N_A1_c_84_n 0.00473899f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.432
cc_48 VPB N_A2_c_134_n 0.0192985f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_49 VPB N_A2_c_135_n 0.0222065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB A2 0.00776607f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_51 VPB N_A2_c_133_n 0.0100204f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.432
cc_52 VPB N_A3_M1009_g 0.0244315f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.68
cc_53 VPB N_A3_M1011_g 0.0210273f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.185
cc_54 VPB N_A3_c_189_n 0.00433668f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_55 VPB N_A3_c_190_n 0.00500772f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.432
cc_56 VPB N_B1_M1012_g 0.022329f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_57 VPB N_B1_M1014_g 0.0298893f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_58 VPB B1 0.00389529f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.432
cc_59 VPB N_B1_c_252_n 0.00624797f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.185
cc_60 VPB N_A_28_368#_c_303_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_61 VPB N_A_28_368#_c_304_n 0.0339247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_28_368#_c_305_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_63 VPB N_A_28_368#_c_306_n 0.00759181f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_64 VPB N_VPWR_c_344_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.68
cc_65 VPB N_VPWR_c_345_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.185
cc_66 VPB N_VPWR_c_346_n 0.0787949f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_67 VPB N_VPWR_c_347_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_68 VPB N_VPWR_c_348_n 0.0181665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_349_n 0.0201062f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_70 VPB N_VPWR_c_343_n 0.0755913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_351_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_300_368#_c_392_n 0.0202557f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_73 VPB N_A_300_368#_c_393_n 0.00254693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_Y_c_418_n 0.00580164f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_75 VPB N_Y_c_419_n 0.007175f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_76 VPB N_Y_c_420_n 0.0390534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_Y_c_421_n 0.00567808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_Y_c_417_n 0.00290204f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_79 VPB Y 0.00275585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 N_A1_M1001_g N_A2_c_134_n 0.0114319f $X=0.96 $Y=2.4 $X2=-0.19 $Y2=-0.245
cc_81 N_A1_c_82_n N_A2_M1006_g 0.0195161f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_82 N_A1_c_84_n N_A2_M1006_g 0.00742259f $X=0.96 $Y=1.432 $X2=0 $Y2=0
cc_83 A1 A2 0.0288692f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A1_c_84_n A2 2.5596e-19 $X=0.96 $Y=1.432 $X2=0 $Y2=0
cc_85 A1 N_A2_c_133_n 0.00505372f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A1_c_84_n N_A2_c_133_n 0.0114319f $X=0.96 $Y=1.432 $X2=0 $Y2=0
cc_87 A1 N_A_28_368#_c_303_n 0.0213698f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A1_M1000_g N_A_28_368#_c_304_n 4.69176e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A1_M1000_g N_A_28_368#_c_309_n 0.0142562f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A1_M1001_g N_A_28_368#_c_309_n 0.012931f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_91 A1 N_A_28_368#_c_309_n 0.0435425f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A1_c_84_n N_A_28_368#_c_309_n 4.90767e-19 $X=0.96 $Y=1.432 $X2=0 $Y2=0
cc_93 N_A1_M1000_g N_A_28_368#_c_305_n 6.74232e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A1_M1001_g N_A_28_368#_c_305_n 0.0121322f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A1_M1001_g N_A_28_368#_c_315_n 8.84614e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_96 A1 N_A_28_368#_c_315_n 0.0209326f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A1_M1000_g N_VPWR_c_344_n 0.0153844f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A1_M1001_g N_VPWR_c_344_n 0.002979f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A1_M1001_g N_VPWR_c_346_n 0.005209f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A1_M1000_g N_VPWR_c_348_n 0.00460063f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A1_M1000_g N_VPWR_c_343_n 0.00912313f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A1_M1001_g N_VPWR_c_343_n 0.00982376f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A1_M1013_g N_A_27_74#_c_490_n 0.0104846f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A1_c_82_n N_A_27_74#_c_490_n 6.72835e-19 $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_105 N_A1_M1013_g N_A_27_74#_c_491_n 0.0118691f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A1_c_82_n N_A_27_74#_c_491_n 0.0115835f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_107 A1 N_A_27_74#_c_491_n 0.0506639f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A1_c_84_n N_A_27_74#_c_491_n 0.0112285f $X=0.96 $Y=1.432 $X2=0 $Y2=0
cc_109 N_A1_M1013_g N_A_27_74#_c_492_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_110 A1 N_A_27_74#_c_492_n 0.0286342f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A1_M1013_g N_A_27_74#_c_493_n 6.72835e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A1_c_82_n N_A_27_74#_c_493_n 0.00981147f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_113 N_A1_c_82_n N_A_27_74#_c_498_n 0.0014252f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_114 A1 N_A_27_74#_c_498_n 0.0179197f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A1_M1013_g N_VGND_c_571_n 0.00613492f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A1_c_82_n N_VGND_c_571_n 0.00475299f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_117 N_A1_c_82_n N_VGND_c_572_n 0.00434272f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_118 N_A1_M1013_g N_VGND_c_574_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A1_M1013_g N_VGND_c_576_n 0.00824951f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_c_82_n N_VGND_c_576_n 0.00821391f $X=1.065 $Y=1.185 $X2=0 $Y2=0
cc_121 N_A2_M1010_g N_A3_M1003_g 0.0130706f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_122 A2 N_A3_c_186_n 0.00174805f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A2_c_133_n N_A3_c_186_n 0.0130706f $X=1.86 $Y=1.537 $X2=0 $Y2=0
cc_124 A2 N_A3_c_190_n 0.00153959f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_c_134_n N_A_28_368#_c_305_n 0.0119229f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_126 N_A2_c_135_n N_A_28_368#_c_305_n 6.58809e-19 $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_127 N_A2_c_134_n N_A_28_368#_c_319_n 0.0172416f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_128 N_A2_c_135_n N_A_28_368#_c_319_n 0.012931f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_129 A2 N_A_28_368#_c_319_n 0.025169f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A2_c_133_n N_A_28_368#_c_319_n 5.40988e-19 $X=1.86 $Y=1.537 $X2=0 $Y2=0
cc_131 N_A2_c_134_n N_A_28_368#_c_315_n 0.00184802f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_132 N_A2_c_134_n N_A_28_368#_c_306_n 5.73047e-19 $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_133 N_A2_c_135_n N_A_28_368#_c_306_n 0.011119f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_134 A2 N_A_28_368#_c_306_n 0.0263958f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A2_c_133_n N_A_28_368#_c_306_n 7.05594e-19 $X=1.86 $Y=1.537 $X2=0 $Y2=0
cc_136 N_A2_c_134_n N_VPWR_c_346_n 0.005209f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_137 N_A2_c_135_n N_VPWR_c_346_n 0.00333926f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_138 N_A2_c_134_n N_VPWR_c_343_n 0.00983474f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_139 N_A2_c_135_n N_VPWR_c_343_n 0.0042782f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_140 N_A2_c_135_n N_A_300_368#_c_392_n 0.0158247f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_141 N_A2_c_134_n N_A_300_368#_c_393_n 0.0032006f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_142 N_A2_c_135_n N_Y_c_421_n 0.00445005f $X=1.86 $Y=1.725 $X2=0 $Y2=0
cc_143 A2 N_Y_c_417_n 0.0198017f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A2_M1006_g N_A_27_74#_c_493_n 0.00981147f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_M1010_g N_A_27_74#_c_493_n 6.72835e-19 $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1006_g N_A_27_74#_c_494_n 0.0155035f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_M1010_g N_A_27_74#_c_494_n 0.0134273f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_148 A2 N_A_27_74#_c_494_n 0.0558786f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A2_c_133_n N_A_27_74#_c_494_n 0.00625968f $X=1.86 $Y=1.537 $X2=0 $Y2=0
cc_150 N_A2_M1010_g N_A_27_74#_c_518_n 0.00342095f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1006_g N_A_27_74#_c_498_n 0.00249368f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_c_133_n N_A_27_74#_c_498_n 0.00381239f $X=1.86 $Y=1.537 $X2=0 $Y2=0
cc_153 N_A2_M1006_g N_A_27_74#_c_499_n 6.72158e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1010_g N_A_27_74#_c_499_n 0.00637016f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1006_g N_VGND_c_572_n 0.00434272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1006_g N_VGND_c_573_n 0.00475299f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_M1010_g N_VGND_c_573_n 0.00613492f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1006_g N_VGND_c_576_n 0.00821391f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1010_g N_VGND_c_576_n 0.00821391f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1010_g N_VGND_c_579_n 0.00434272f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A3_M1005_g N_B1_M1007_g 0.0307304f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A3_M1011_g N_B1_M1012_g 0.0139583f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A3_c_189_n N_B1_M1012_g 0.00213915f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A3_c_189_n N_B1_c_250_n 0.0203452f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A3_c_190_n N_B1_c_250_n 4.12636e-19 $X=3.37 $Y=1.515 $X2=0 $Y2=0
cc_166 N_A3_M1005_g N_B1_c_252_n 0.021601f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A3_c_189_n N_B1_c_252_n 4.14586e-19 $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A3_M1009_g N_VPWR_c_346_n 0.00333896f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A3_M1011_g N_VPWR_c_346_n 0.00517089f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A3_M1009_g N_VPWR_c_343_n 0.00427818f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A3_M1011_g N_VPWR_c_343_n 0.00979141f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A3_M1009_g N_A_300_368#_c_392_n 0.0156999f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A3_M1011_g N_A_300_368#_c_392_n 0.00436192f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A3_M1009_g N_A_300_368#_c_398_n 0.0134366f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A3_M1011_g N_A_300_368#_c_398_n 0.00732498f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A3_M1005_g N_Y_c_415_n 0.0123777f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A3_c_189_n N_Y_c_415_n 0.0331911f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A3_c_190_n N_Y_c_415_n 0.0119562f $X=3.37 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A3_M1003_g N_Y_c_416_n 0.00388066f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A3_M1009_g N_Y_c_430_n 0.0169639f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A3_M1011_g N_Y_c_430_n 0.0142562f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A3_c_189_n N_Y_c_430_n 0.0300318f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A3_c_190_n N_Y_c_430_n 4.90767e-19 $X=3.37 $Y=1.515 $X2=0 $Y2=0
cc_184 N_A3_M1005_g N_Y_c_434_n 9.17327e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A3_c_186_n N_Y_c_421_n 0.00650414f $X=2.57 $Y=1.425 $X2=0 $Y2=0
cc_186 N_A3_M1009_g N_Y_c_421_n 0.00529166f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A3_M1003_g N_Y_c_417_n 0.00627755f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A3_M1009_g N_Y_c_417_n 0.00418434f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A3_M1011_g N_Y_c_417_n 8.85973e-19 $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A3_M1005_g N_Y_c_417_n 0.00426386f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A3_c_188_n N_Y_c_417_n 0.0104157f $X=2.805 $Y=1.515 $X2=0 $Y2=0
cc_192 N_A3_c_189_n N_Y_c_417_n 0.0318332f $X=3.28 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A3_c_190_n N_Y_c_417_n 0.00907424f $X=3.37 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A3_M1011_g N_Y_c_444_n 0.0026629f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A3_M1003_g N_A_27_74#_c_494_n 0.0040258f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A3_M1003_g N_A_27_74#_c_518_n 0.00728117f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A3_M1003_g N_A_27_74#_c_525_n 0.0147088f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A3_M1005_g N_A_27_74#_c_525_n 0.0117184f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A3_c_188_n N_A_27_74#_c_525_n 7.07703e-19 $X=2.805 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A3_c_190_n N_A_27_74#_c_525_n 4.51931e-19 $X=3.37 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A3_M1005_g N_A_27_74#_c_529_n 0.00793893f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A3_M1005_g N_A_27_74#_c_496_n 0.00368639f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A3_M1003_g N_A_27_74#_c_499_n 0.0111378f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_M1005_g N_VGND_c_575_n 0.00321293f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A3_M1003_g N_VGND_c_576_n 0.00414829f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1005_g N_VGND_c_576_n 0.00414843f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_M1003_g N_VGND_c_579_n 0.00324657f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_M1003_g N_VGND_c_580_n 0.00790404f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_M1005_g N_VGND_c_580_n 0.00576111f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B1_M1012_g N_VPWR_c_345_n 0.00307681f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B1_M1014_g N_VPWR_c_345_n 0.00307681f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_212 N_B1_M1012_g N_VPWR_c_346_n 0.005209f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_213 N_B1_M1014_g N_VPWR_c_349_n 0.005209f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B1_M1012_g N_VPWR_c_343_n 0.00982832f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_215 N_B1_M1014_g N_VPWR_c_343_n 0.00986008f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_216 N_B1_M1012_g N_A_300_368#_c_392_n 4.66732e-19 $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_217 N_B1_M1007_g N_Y_c_415_n 0.0116769f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_218 N_B1_M1008_g N_Y_c_415_n 0.00283624f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B1_c_250_n N_Y_c_415_n 0.0392202f $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_220 N_B1_c_252_n N_Y_c_415_n 0.004978f $X=4.295 $Y=1.49 $X2=0 $Y2=0
cc_221 N_B1_M1012_g N_Y_c_449_n 0.012931f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B1_M1014_g N_Y_c_449_n 0.0129082f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_223 N_B1_c_250_n N_Y_c_449_n 0.0371523f $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_224 N_B1_c_252_n N_Y_c_449_n 0.00207739f $X=4.295 $Y=1.49 $X2=0 $Y2=0
cc_225 N_B1_M1007_g N_Y_c_434_n 0.00625675f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B1_M1014_g N_Y_c_419_n 8.69327e-19 $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_227 N_B1_c_250_n N_Y_c_419_n 7.98247e-19 $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_228 B1 N_Y_c_419_n 0.0259384f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_229 N_B1_c_252_n N_Y_c_419_n 0.00192045f $X=4.295 $Y=1.49 $X2=0 $Y2=0
cc_230 N_B1_M1012_g N_Y_c_420_n 6.82021e-19 $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_231 N_B1_M1014_g N_Y_c_420_n 0.0136905f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_232 N_B1_M1012_g N_Y_c_444_n 0.00339139f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_233 N_B1_M1014_g N_Y_c_444_n 2.91133e-19 $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_234 N_B1_c_250_n N_Y_c_444_n 0.00561722f $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_235 N_B1_c_252_n N_Y_c_444_n 0.00160183f $X=4.295 $Y=1.49 $X2=0 $Y2=0
cc_236 N_B1_M1012_g Y 0.0112049f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_237 N_B1_M1014_g Y 3.89903e-19 $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B1_M1007_g N_A_27_74#_c_495_n 0.0107757f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_M1008_g N_A_27_74#_c_495_n 0.0140969f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1007_g N_A_27_74#_c_497_n 8.96536e-19 $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B1_M1008_g N_A_27_74#_c_497_n 0.00715938f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B1_c_250_n N_A_27_74#_c_497_n 3.7446e-19 $X=4.365 $Y=1.515 $X2=0 $Y2=0
cc_243 B1 N_A_27_74#_c_497_n 0.0260711f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_244 N_B1_c_252_n N_A_27_74#_c_497_n 0.00172989f $X=4.295 $Y=1.49 $X2=0 $Y2=0
cc_245 N_B1_M1007_g N_VGND_c_575_n 0.00278271f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B1_M1008_g N_VGND_c_575_n 0.00278266f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B1_M1007_g N_VGND_c_576_n 0.00354005f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B1_M1008_g N_VGND_c_576_n 0.00357648f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_28_368#_c_309_n N_VPWR_M1000_d 0.00314376f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_250 N_A_28_368#_c_304_n N_VPWR_c_344_n 0.0224614f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_28_368#_c_309_n N_VPWR_c_344_n 0.0148589f $X=1.02 $Y=2.035 $X2=0
+ $Y2=0
cc_252 N_A_28_368#_c_305_n N_VPWR_c_344_n 0.0234083f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_253 N_A_28_368#_c_305_n N_VPWR_c_346_n 0.0144623f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_A_28_368#_c_304_n N_VPWR_c_348_n 0.011066f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_255 N_A_28_368#_c_304_n N_VPWR_c_343_n 0.00915947f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_256 N_A_28_368#_c_305_n N_VPWR_c_343_n 0.0118344f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_257 N_A_28_368#_c_319_n N_A_300_368#_M1002_d 0.00335f $X=1.92 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_258 N_A_28_368#_c_319_n N_A_300_368#_c_402_n 0.0126919f $X=1.92 $Y=2.035
+ $X2=0 $Y2=0
cc_259 N_A_28_368#_M1004_s N_A_300_368#_c_392_n 0.00266942f $X=1.95 $Y=1.84
+ $X2=0 $Y2=0
cc_260 N_A_28_368#_c_306_n N_A_300_368#_c_392_n 0.0205035f $X=2.085 $Y=2.115
+ $X2=0 $Y2=0
cc_261 N_A_28_368#_c_305_n N_A_300_368#_c_393_n 0.00327031f $X=1.185 $Y=2.815
+ $X2=0 $Y2=0
cc_262 N_A_28_368#_c_306_n N_Y_c_418_n 0.0377581f $X=2.085 $Y=2.115 $X2=0 $Y2=0
cc_263 N_A_28_368#_c_306_n N_Y_c_421_n 0.0113228f $X=2.085 $Y=2.115 $X2=0 $Y2=0
cc_264 N_VPWR_c_346_n N_A_300_368#_c_392_n 0.101986f $X=3.985 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_343_n N_A_300_368#_c_392_n 0.0574792f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_346_n N_A_300_368#_c_393_n 0.0121867f $X=3.985 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_343_n N_A_300_368#_c_393_n 0.00660921f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_268 N_VPWR_M1012_d N_Y_c_449_n 0.00311483f $X=3.935 $Y=1.84 $X2=0 $Y2=0
cc_269 N_VPWR_c_345_n N_Y_c_449_n 0.0126919f $X=4.07 $Y=2.355 $X2=0 $Y2=0
cc_270 N_VPWR_c_345_n N_Y_c_420_n 0.0266644f $X=4.07 $Y=2.355 $X2=0 $Y2=0
cc_271 N_VPWR_c_349_n N_Y_c_420_n 0.014549f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_343_n N_Y_c_420_n 0.0119743f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_c_345_n Y 0.0266644f $X=4.07 $Y=2.355 $X2=0 $Y2=0
cc_274 N_VPWR_c_346_n Y 0.014549f $X=3.985 $Y=3.33 $X2=0 $Y2=0
cc_275 N_VPWR_c_343_n Y 0.0119743f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_276 N_A_300_368#_c_392_n N_Y_M1009_s 0.00266942f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_277 N_A_300_368#_c_392_n N_Y_c_418_n 0.0184743f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_278 N_A_300_368#_M1009_d N_Y_c_430_n 0.00314376f $X=2.985 $Y=1.84 $X2=0 $Y2=0
cc_279 N_A_300_368#_c_398_n N_Y_c_430_n 0.0170259f $X=3.12 $Y=2.455 $X2=0 $Y2=0
cc_280 N_A_300_368#_c_392_n Y 0.0039531f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_281 N_Y_c_415_n N_A_27_74#_M1005_s 0.00176461f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_282 N_Y_c_416_n N_A_27_74#_c_494_n 0.012289f $X=2.835 $Y=1.095 $X2=0 $Y2=0
cc_283 N_Y_c_415_n N_A_27_74#_c_525_n 0.0528952f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_284 N_Y_c_416_n N_A_27_74#_c_525_n 0.013831f $X=2.835 $Y=1.095 $X2=0 $Y2=0
cc_285 N_Y_M1007_d N_A_27_74#_c_495_n 0.00237956f $X=3.875 $Y=0.37 $X2=0 $Y2=0
cc_286 N_Y_c_415_n N_A_27_74#_c_495_n 0.0030313f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_287 N_Y_c_434_n N_A_27_74#_c_495_n 0.0166105f $X=4.015 $Y=0.775 $X2=0 $Y2=0
cc_288 N_Y_c_415_n N_VGND_M1003_d 0.00581259f $X=3.85 $Y=1.095 $X2=0 $Y2=0
cc_289 N_Y_c_416_n N_VGND_M1003_d 0.00372663f $X=2.835 $Y=1.095 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_491_n N_VGND_M1013_d 0.00369983f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_27_74#_c_494_n N_VGND_M1006_d 0.00369983f $X=2.115 $Y=1.095 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_c_525_n N_VGND_M1003_d 0.0164865f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_490_n N_VGND_c_571_n 0.0186136f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_491_n N_VGND_c_571_n 0.0233713f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_493_n N_VGND_c_571_n 0.0186136f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_493_n N_VGND_c_572_n 0.0144922f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_493_n N_VGND_c_573_n 0.0186136f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_494_n N_VGND_c_573_n 0.0233713f $X=2.115 $Y=1.095 $X2=0
+ $Y2=0
cc_299 N_A_27_74#_c_499_n N_VGND_c_573_n 0.0186136f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_490_n N_VGND_c_574_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_525_n N_VGND_c_575_n 0.00236055f $X=3.42 $Y=0.755 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_495_n N_VGND_c_575_n 0.0665294f $X=4.35 $Y=0.34 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_496_n N_VGND_c_575_n 0.0176331f $X=3.67 $Y=0.34 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_490_n N_VGND_c_576_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_493_n N_VGND_c_576_n 0.0118826f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_525_n N_VGND_c_576_n 0.0113479f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_495_n N_VGND_c_576_n 0.0370234f $X=4.35 $Y=0.34 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_496_n N_VGND_c_576_n 0.00956698f $X=3.67 $Y=0.34 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_499_n N_VGND_c_576_n 0.0118826f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_525_n N_VGND_c_579_n 0.0023667f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_499_n N_VGND_c_579_n 0.0144922f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_525_n N_VGND_c_580_n 0.0468302f $X=3.42 $Y=0.755 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_496_n N_VGND_c_580_n 0.0119157f $X=3.67 $Y=0.34 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_499_n N_VGND_c_580_n 0.00620201f $X=2.28 $Y=0.515 $X2=0
+ $Y2=0

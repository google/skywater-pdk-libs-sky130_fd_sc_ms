* File: sky130_fd_sc_ms__a41oi_4.pxi.spice
* Created: Fri Aug 28 17:10:08 2020
* 
x_PM_SKY130_FD_SC_MS__A41OI_4%B1 N_B1_M1015_g N_B1_c_157_n N_B1_M1002_g
+ N_B1_c_158_n N_B1_M1007_g N_B1_M1032_g N_B1_c_159_n N_B1_M1009_g N_B1_c_154_n
+ N_B1_c_161_n N_B1_M1012_g B1 B1 B1 N_B1_c_155_n N_B1_c_156_n
+ PM_SKY130_FD_SC_MS__A41OI_4%B1
x_PM_SKY130_FD_SC_MS__A41OI_4%A1 N_A1_c_227_n N_A1_M1020_g N_A1_c_228_n
+ N_A1_c_229_n N_A1_c_235_n N_A1_M1000_g N_A1_c_230_n N_A1_M1022_g N_A1_c_236_n
+ N_A1_M1010_g N_A1_c_231_n N_A1_M1026_g N_A1_c_237_n N_A1_M1013_g N_A1_c_232_n
+ N_A1_M1036_g N_A1_c_238_n N_A1_M1014_g A1 A1 N_A1_c_233_n N_A1_c_234_n
+ PM_SKY130_FD_SC_MS__A41OI_4%A1
x_PM_SKY130_FD_SC_MS__A41OI_4%A2 N_A2_c_335_n N_A2_M1005_g N_A2_M1003_g
+ N_A2_c_337_n N_A2_M1006_g N_A2_M1019_g N_A2_c_339_n N_A2_M1023_g N_A2_M1024_g
+ N_A2_c_341_n N_A2_M1027_g N_A2_M1025_g N_A2_c_343_n A2 A2 N_A2_c_344_n
+ N_A2_c_345_n N_A2_c_351_n PM_SKY130_FD_SC_MS__A41OI_4%A2
x_PM_SKY130_FD_SC_MS__A41OI_4%A3 N_A3_M1029_g N_A3_M1008_g N_A3_M1030_g
+ N_A3_M1018_g N_A3_M1034_g N_A3_M1021_g N_A3_M1035_g N_A3_M1033_g A3 A3 A3 A3
+ A3 N_A3_c_435_n PM_SKY130_FD_SC_MS__A41OI_4%A3
x_PM_SKY130_FD_SC_MS__A41OI_4%A4 N_A4_M1001_g N_A4_M1004_g N_A4_M1011_g
+ N_A4_M1016_g N_A4_M1031_g N_A4_M1017_g N_A4_M1037_g N_A4_M1028_g A4 A4 A4 A4
+ N_A4_c_523_n PM_SKY130_FD_SC_MS__A41OI_4%A4
x_PM_SKY130_FD_SC_MS__A41OI_4%A_27_368# N_A_27_368#_M1002_s N_A_27_368#_M1007_s
+ N_A_27_368#_M1012_s N_A_27_368#_M1010_d N_A_27_368#_M1014_d
+ N_A_27_368#_M1019_s N_A_27_368#_M1025_s N_A_27_368#_M1030_s
+ N_A_27_368#_M1035_s N_A_27_368#_M1011_s N_A_27_368#_M1037_s
+ N_A_27_368#_c_595_n N_A_27_368#_c_596_n N_A_27_368#_c_597_n
+ N_A_27_368#_c_616_n N_A_27_368#_c_598_n N_A_27_368#_c_620_n
+ N_A_27_368#_c_621_n N_A_27_368#_c_628_n N_A_27_368#_c_630_n
+ N_A_27_368#_c_633_n N_A_27_368#_c_634_n N_A_27_368#_c_599_n
+ N_A_27_368#_c_649_n N_A_27_368#_c_600_n N_A_27_368#_c_658_n
+ N_A_27_368#_c_601_n N_A_27_368#_c_674_n N_A_27_368#_c_602_n
+ N_A_27_368#_c_682_n N_A_27_368#_c_603_n N_A_27_368#_c_697_n
+ N_A_27_368#_c_604_n N_A_27_368#_c_705_n N_A_27_368#_c_605_n
+ N_A_27_368#_c_606_n N_A_27_368#_c_607_n N_A_27_368#_c_608_n
+ N_A_27_368#_c_642_n N_A_27_368#_c_609_n N_A_27_368#_c_671_n
+ N_A_27_368#_c_690_n N_A_27_368#_c_694_n N_A_27_368#_c_713_n
+ PM_SKY130_FD_SC_MS__A41OI_4%A_27_368#
x_PM_SKY130_FD_SC_MS__A41OI_4%Y N_Y_M1015_s N_Y_M1020_d N_Y_M1026_d N_Y_M1002_d
+ N_Y_M1009_d N_Y_c_787_n N_Y_c_788_n N_Y_c_789_n N_Y_c_858_n N_Y_c_790_n
+ N_Y_c_791_n N_Y_c_833_n N_Y_c_834_n N_Y_c_811_n N_Y_c_815_n N_Y_c_794_n
+ N_Y_c_842_n Y N_Y_c_792_n Y PM_SKY130_FD_SC_MS__A41OI_4%Y
x_PM_SKY130_FD_SC_MS__A41OI_4%VPWR N_VPWR_M1000_s N_VPWR_M1013_s N_VPWR_M1003_d
+ N_VPWR_M1024_d N_VPWR_M1029_d N_VPWR_M1034_d N_VPWR_M1001_d N_VPWR_M1031_d
+ N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n
+ N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_901_n
+ N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n N_VPWR_c_906_n
+ VPWR N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n N_VPWR_c_891_n
+ N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n N_VPWR_c_914_n N_VPWR_c_915_n
+ N_VPWR_c_916_n N_VPWR_c_917_n PM_SKY130_FD_SC_MS__A41OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A41OI_4%VGND N_VGND_M1015_d N_VGND_M1032_d N_VGND_M1004_s
+ N_VGND_M1017_s N_VGND_c_1034_n N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n
+ N_VGND_c_1038_n VGND N_VGND_c_1039_n N_VGND_c_1040_n N_VGND_c_1041_n
+ N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n PM_SKY130_FD_SC_MS__A41OI_4%VGND
x_PM_SKY130_FD_SC_MS__A41OI_4%A_325_74# N_A_325_74#_M1020_s N_A_325_74#_M1022_s
+ N_A_325_74#_M1036_s N_A_325_74#_M1006_s N_A_325_74#_M1027_s
+ N_A_325_74#_c_1133_n N_A_325_74#_c_1134_n N_A_325_74#_c_1135_n
+ N_A_325_74#_c_1136_n N_A_325_74#_c_1137_n N_A_325_74#_c_1138_n
+ N_A_325_74#_c_1139_n N_A_325_74#_c_1140_n
+ PM_SKY130_FD_SC_MS__A41OI_4%A_325_74#
x_PM_SKY130_FD_SC_MS__A41OI_4%A_852_74# N_A_852_74#_M1005_d N_A_852_74#_M1023_d
+ N_A_852_74#_M1008_s N_A_852_74#_M1021_s N_A_852_74#_c_1196_n
+ N_A_852_74#_c_1197_n PM_SKY130_FD_SC_MS__A41OI_4%A_852_74#
x_PM_SKY130_FD_SC_MS__A41OI_4%A_1235_74# N_A_1235_74#_M1008_d
+ N_A_1235_74#_M1018_d N_A_1235_74#_M1033_d N_A_1235_74#_M1016_d
+ N_A_1235_74#_M1028_d N_A_1235_74#_c_1227_n N_A_1235_74#_c_1228_n
+ N_A_1235_74#_c_1229_n N_A_1235_74#_c_1230_n N_A_1235_74#_c_1231_n
+ N_A_1235_74#_c_1232_n N_A_1235_74#_c_1233_n N_A_1235_74#_c_1234_n
+ N_A_1235_74#_c_1235_n PM_SKY130_FD_SC_MS__A41OI_4%A_1235_74#
cc_1 VNB N_B1_M1015_g 0.0315575f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_M1032_g 0.0315591f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_B1_c_154_n 0.015937f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.64
cc_4 VNB N_B1_c_155_n 0.0184974f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_5 VNB N_B1_c_156_n 0.0718552f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.532
cc_6 VNB N_A1_c_227_n 0.01857f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_7 VNB N_A1_c_228_n 0.0132358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_229_n 0.00839791f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.715
cc_9 VNB N_A1_c_230_n 0.0179822f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_10 VNB N_A1_c_231_n 0.0176901f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.715
cc_11 VNB N_A1_c_232_n 0.0157849f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_12 VNB N_A1_c_233_n 0.00231182f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_13 VNB N_A1_c_234_n 0.112919f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_14 VNB N_A2_c_335_n 0.0166764f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_15 VNB N_A2_M1003_g 4.25593e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_16 VNB N_A2_c_337_n 0.0158586f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.715
cc_17 VNB N_A2_M1019_g 4.96947e-19 $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_18 VNB N_A2_c_339_n 0.015257f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.715
cc_19 VNB N_A2_M1024_g 4.96305e-19 $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.715
cc_20 VNB N_A2_c_341_n 0.0199171f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_21 VNB N_A2_M1025_g 4.6008e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_343_n 0.00252762f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.532
cc_23 VNB N_A2_c_344_n 0.125066f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_24 VNB N_A2_c_345_n 0.00352257f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_25 VNB N_A3_M1008_g 0.0320084f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_26 VNB N_A3_M1018_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.715
cc_27 VNB N_A3_M1021_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_A3_M1033_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.532
cc_29 VNB A3 0.00908404f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.532
cc_30 VNB N_A3_c_435_n 0.0809135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A4_M1004_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_32 VNB N_A4_M1016_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.715
cc_33 VNB N_A4_M1017_g 0.0230771f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_A4_M1028_g 0.0331137f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.532
cc_35 VNB A4 0.0166485f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.532
cc_36 VNB N_A4_c_523_n 0.074341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_787_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.64
cc_38 VNB N_Y_c_788_n 0.0168364f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_39 VNB N_Y_c_789_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_40 VNB N_Y_c_790_n 0.0105726f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.532
cc_41 VNB N_Y_c_791_n 0.00412271f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.532
cc_42 VNB N_Y_c_792_n 8.52578e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VPWR_c_891_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_1034_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_45 VNB N_VGND_c_1035_n 0.043326f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.715
cc_46 VNB N_VGND_c_1036_n 0.0107076f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.64
cc_47 VNB N_VGND_c_1037_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_48 VNB N_VGND_c_1038_n 0.00574819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1039_n 0.018855f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.532
cc_50 VNB N_VGND_c_1040_n 0.163203f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.532
cc_51 VNB N_VGND_c_1041_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1042_n 0.0188218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1043_n 0.533259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1044_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1045_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1046_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_325_74#_c_1133_n 0.00384069f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.64
cc_58 VNB N_A_325_74#_c_1134_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=1.955
+ $Y2=1.715
cc_59 VNB N_A_325_74#_c_1135_n 0.00417961f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_60 VNB N_A_325_74#_c_1136_n 0.00437333f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_61 VNB N_A_325_74#_c_1137_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_325_74#_c_1138_n 0.0133561f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_63 VNB N_A_325_74#_c_1139_n 0.00496413f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.532
cc_64 VNB N_A_325_74#_c_1140_n 0.00609172f $X=-0.19 $Y=-0.245 $X2=1.265
+ $Y2=1.515
cc_65 VNB N_A_852_74#_c_1196_n 0.00251362f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_66 VNB N_A_852_74#_c_1197_n 0.0283516f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_67 VNB N_A_1235_74#_c_1227_n 0.00754101f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_68 VNB N_A_1235_74#_c_1228_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.955
+ $Y2=1.715
cc_69 VNB N_A_1235_74#_c_1229_n 0.00323033f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_70 VNB N_A_1235_74#_c_1230_n 0.00517531f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.58
cc_71 VNB N_A_1235_74#_c_1231_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1235_74#_c_1232_n 0.0134691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1235_74#_c_1233_n 0.0266181f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.515
cc_74 VNB N_A_1235_74#_c_1234_n 0.00523512f $X=-0.19 $Y=-0.245 $X2=1.265
+ $Y2=1.515
cc_75 VNB N_A_1235_74#_c_1235_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.565
cc_76 VPB N_B1_c_157_n 0.0236174f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.715
cc_77 VPB N_B1_c_158_n 0.0190417f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.715
cc_78 VPB N_B1_c_159_n 0.0187981f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.715
cc_79 VPB N_B1_c_154_n 0.00519579f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.64
cc_80 VPB N_B1_c_161_n 0.0174829f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.715
cc_81 VPB N_B1_c_155_n 0.0144606f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_82 VPB N_B1_c_156_n 0.0162884f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.532
cc_83 VPB N_A1_c_235_n 0.01814f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_84 VPB N_A1_c_236_n 0.0184193f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_85 VPB N_A1_c_237_n 0.0179167f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.64
cc_86 VPB N_A1_c_238_n 0.0184747f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_87 VPB N_A1_c_233_n 0.0070377f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_88 VPB N_A1_c_234_n 0.0306284f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_89 VPB N_A2_M1003_g 0.0224783f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_90 VPB N_A2_M1019_g 0.0230178f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_91 VPB N_A2_M1024_g 0.0229387f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.715
cc_92 VPB N_A2_M1025_g 0.0228646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A2_c_345_n 0.00251835f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.565
cc_94 VPB N_A2_c_351_n 0.00341355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A3_M1029_g 0.0213808f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_96 VPB N_A3_M1030_g 0.0210664f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_97 VPB N_A3_M1034_g 0.0210667f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.64
cc_98 VPB N_A3_M1035_g 0.0219312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB A3 0.013906f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.532
cc_100 VPB N_A3_c_435_n 0.0172592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A4_M1001_g 0.0213266f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_102 VPB N_A4_M1011_g 0.020498f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_103 VPB N_A4_M1031_g 0.020498f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.64
cc_104 VPB N_A4_M1037_g 0.027583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB A4 0.0156573f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.532
cc_106 VPB N_A4_c_523_n 0.0118911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_368#_c_595_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.532
cc_108 VPB N_A_27_368#_c_596_n 0.00237811f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.532
cc_109 VPB N_A_27_368#_c_597_n 0.00971634f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.532
cc_110 VPB N_A_27_368#_c_598_n 0.00388794f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_111 VPB N_A_27_368#_c_599_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_368#_c_600_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_368#_c_601_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_368#_c_602_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_368#_c_603_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_368#_c_604_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_368#_c_605_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_368#_c_606_n 0.0352219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_368#_c_607_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_368#_c_608_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_368#_c_609_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_Y_c_790_n 0.00244544f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.532
cc_123 VPB N_Y_c_794_n 0.00263228f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_124 VPB Y 8.18243e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_892_n 0.00928334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_893_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.532
cc_127 VPB N_VPWR_c_894_n 0.00888637f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_128 VPB N_VPWR_c_895_n 0.0198086f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.532
cc_129 VPB N_VPWR_c_896_n 0.00891028f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_130 VPB N_VPWR_c_897_n 0.0199677f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.532
cc_131 VPB N_VPWR_c_898_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_132 VPB N_VPWR_c_899_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_900_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_901_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_902_n 0.0081889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_903_n 0.00499798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_904_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_905_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_906_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_907_n 0.0604926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_908_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_909_n 0.0202453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_891_n 0.0971579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_911_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_912_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_913_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_914_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_915_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_916_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_917_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 N_B1_c_154_n N_A1_c_229_n 0.00883023f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_152 N_B1_c_161_n N_A1_c_235_n 0.0285934f $X=1.955 $Y=1.715 $X2=0 $Y2=0
cc_153 N_B1_c_154_n N_A1_c_233_n 2.0015e-19 $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_154 N_B1_c_154_n N_A1_c_234_n 0.00994134f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_155 N_B1_c_156_n N_A1_c_234_n 0.00226331f $X=1.595 $Y=1.532 $X2=0 $Y2=0
cc_156 N_B1_c_157_n N_A_27_368#_c_595_n 0.0124591f $X=0.51 $Y=1.715 $X2=0 $Y2=0
cc_157 N_B1_c_158_n N_A_27_368#_c_595_n 6.09213e-19 $X=1.005 $Y=1.715 $X2=0
+ $Y2=0
cc_158 N_B1_c_155_n N_A_27_368#_c_595_n 0.0254478f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_159 N_B1_c_157_n N_A_27_368#_c_596_n 0.012228f $X=0.51 $Y=1.715 $X2=0 $Y2=0
cc_160 N_B1_c_158_n N_A_27_368#_c_596_n 0.0144896f $X=1.005 $Y=1.715 $X2=0 $Y2=0
cc_161 N_B1_c_157_n N_A_27_368#_c_597_n 0.00282152f $X=0.51 $Y=1.715 $X2=0 $Y2=0
cc_162 N_B1_c_159_n N_A_27_368#_c_616_n 0.00915505f $X=1.505 $Y=1.715 $X2=0
+ $Y2=0
cc_163 N_B1_c_161_n N_A_27_368#_c_616_n 5.73047e-19 $X=1.955 $Y=1.715 $X2=0
+ $Y2=0
cc_164 N_B1_c_159_n N_A_27_368#_c_598_n 0.0116345f $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_165 N_B1_c_161_n N_A_27_368#_c_598_n 0.0135505f $X=1.955 $Y=1.715 $X2=0 $Y2=0
cc_166 N_B1_c_161_n N_A_27_368#_c_620_n 0.00244698f $X=1.955 $Y=1.715 $X2=0
+ $Y2=0
cc_167 N_B1_c_159_n N_A_27_368#_c_621_n 5.18977e-19 $X=1.505 $Y=1.715 $X2=0
+ $Y2=0
cc_168 N_B1_c_161_n N_A_27_368#_c_621_n 0.00706265f $X=1.955 $Y=1.715 $X2=0
+ $Y2=0
cc_169 N_B1_c_159_n N_A_27_368#_c_607_n 0.00214324f $X=1.505 $Y=1.715 $X2=0
+ $Y2=0
cc_170 N_B1_M1015_g N_Y_c_787_n 0.00838277f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B1_M1032_g N_Y_c_787_n 0.00350341f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B1_M1032_g N_Y_c_788_n 0.0167736f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B1_c_154_n N_Y_c_788_n 0.00520299f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_174 N_B1_c_155_n N_Y_c_788_n 0.041974f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_175 N_B1_c_156_n N_Y_c_788_n 0.0158526f $X=1.595 $Y=1.532 $X2=0 $Y2=0
cc_176 N_B1_M1015_g N_Y_c_789_n 0.00502286f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B1_c_155_n N_Y_c_789_n 0.0282341f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_178 N_B1_c_156_n N_Y_c_789_n 0.0041619f $X=1.595 $Y=1.532 $X2=0 $Y2=0
cc_179 N_B1_c_159_n N_Y_c_790_n 0.00137886f $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_180 N_B1_c_154_n N_Y_c_790_n 0.0103123f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_181 N_B1_c_161_n N_Y_c_790_n 0.00323799f $X=1.955 $Y=1.715 $X2=0 $Y2=0
cc_182 N_B1_c_155_n N_Y_c_790_n 0.0186051f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_183 N_B1_c_156_n N_Y_c_790_n 0.00298455f $X=1.595 $Y=1.532 $X2=0 $Y2=0
cc_184 N_B1_c_154_n N_Y_c_791_n 3.06452e-19 $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_185 N_B1_c_158_n N_Y_c_811_n 0.0112855f $X=1.005 $Y=1.715 $X2=0 $Y2=0
cc_186 N_B1_c_159_n N_Y_c_811_n 7.25672e-19 $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_187 N_B1_c_155_n N_Y_c_811_n 0.0244752f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_188 N_B1_c_156_n N_Y_c_811_n 9.01473e-19 $X=1.595 $Y=1.532 $X2=0 $Y2=0
cc_189 N_B1_c_158_n N_Y_c_815_n 0.0132272f $X=1.005 $Y=1.715 $X2=0 $Y2=0
cc_190 N_B1_c_159_n N_Y_c_815_n 0.0192717f $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_191 N_B1_c_155_n N_Y_c_815_n 0.0333532f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_192 N_B1_c_156_n N_Y_c_815_n 8.28211e-19 $X=1.595 $Y=1.532 $X2=0 $Y2=0
cc_193 N_B1_c_159_n N_Y_c_794_n 5.29908e-19 $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_194 N_B1_c_154_n N_Y_c_794_n 0.00242746f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_195 N_B1_c_161_n N_Y_c_794_n 0.0157103f $X=1.955 $Y=1.715 $X2=0 $Y2=0
cc_196 N_B1_c_157_n N_VPWR_c_907_n 0.00333901f $X=0.51 $Y=1.715 $X2=0 $Y2=0
cc_197 N_B1_c_158_n N_VPWR_c_907_n 0.00333926f $X=1.005 $Y=1.715 $X2=0 $Y2=0
cc_198 N_B1_c_159_n N_VPWR_c_907_n 0.00333896f $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_199 N_B1_c_161_n N_VPWR_c_907_n 0.00333896f $X=1.955 $Y=1.715 $X2=0 $Y2=0
cc_200 N_B1_c_157_n N_VPWR_c_891_n 0.00426886f $X=0.51 $Y=1.715 $X2=0 $Y2=0
cc_201 N_B1_c_158_n N_VPWR_c_891_n 0.00423617f $X=1.005 $Y=1.715 $X2=0 $Y2=0
cc_202 N_B1_c_159_n N_VPWR_c_891_n 0.00423173f $X=1.505 $Y=1.715 $X2=0 $Y2=0
cc_203 N_B1_c_161_n N_VPWR_c_891_n 0.00422796f $X=1.955 $Y=1.715 $X2=0 $Y2=0
cc_204 N_B1_M1015_g N_VGND_c_1035_n 0.00647381f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B1_c_155_n N_VGND_c_1035_n 0.0179756f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_206 N_B1_M1015_g N_VGND_c_1036_n 6.83978e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B1_M1032_g N_VGND_c_1036_n 0.012834f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B1_M1015_g N_VGND_c_1039_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B1_M1032_g N_VGND_c_1039_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B1_M1015_g N_VGND_c_1043_n 0.008246f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B1_M1032_g N_VGND_c_1043_n 0.00758198f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B1_M1032_g N_A_325_74#_c_1133_n 8.38994e-19 $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_B1_M1032_g N_A_325_74#_c_1135_n 7.24903e-19 $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A1_c_232_n N_A2_c_335_n 0.0123861f $X=3.685 $Y=1.205 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A1_c_238_n N_A2_M1003_g 0.00909593f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_216 N_A1_c_234_n N_A2_c_344_n 0.0260014f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_217 N_A1_c_238_n N_A2_c_345_n 0.00138267f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_218 N_A1_c_234_n N_A2_c_345_n 0.00895648f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_219 N_A1_c_235_n N_A_27_368#_c_598_n 0.00338824f $X=2.405 $Y=1.745 $X2=0
+ $Y2=0
cc_220 N_A1_c_235_n N_A_27_368#_c_620_n 8.84614e-19 $X=2.405 $Y=1.745 $X2=0
+ $Y2=0
cc_221 N_A1_c_235_n N_A_27_368#_c_621_n 0.00726463f $X=2.405 $Y=1.745 $X2=0
+ $Y2=0
cc_222 N_A1_c_236_n N_A_27_368#_c_621_n 3.69413e-19 $X=2.955 $Y=1.745 $X2=0
+ $Y2=0
cc_223 N_A1_c_235_n N_A_27_368#_c_628_n 0.0132511f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_224 N_A1_c_236_n N_A_27_368#_c_628_n 0.0132511f $X=2.955 $Y=1.745 $X2=0 $Y2=0
cc_225 N_A1_c_237_n N_A_27_368#_c_630_n 0.0130047f $X=3.405 $Y=1.745 $X2=0 $Y2=0
cc_226 N_A1_c_238_n N_A_27_368#_c_630_n 0.0172228f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_227 N_A1_c_234_n N_A_27_368#_c_630_n 8.47014e-19 $X=3.685 $Y=1.475 $X2=0
+ $Y2=0
cc_228 N_A1_c_238_n N_A_27_368#_c_633_n 0.00267871f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_229 N_A1_c_237_n N_A_27_368#_c_634_n 7.88686e-19 $X=3.405 $Y=1.745 $X2=0
+ $Y2=0
cc_230 N_A1_c_238_n N_A_27_368#_c_634_n 0.00345837f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_231 N_A1_c_237_n N_A_27_368#_c_599_n 5.31941e-19 $X=3.405 $Y=1.745 $X2=0
+ $Y2=0
cc_232 N_A1_c_238_n N_A_27_368#_c_599_n 0.00792151f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_233 N_A1_c_235_n N_A_27_368#_c_608_n 3.85457e-19 $X=2.405 $Y=1.745 $X2=0
+ $Y2=0
cc_234 N_A1_c_236_n N_A_27_368#_c_608_n 0.00951626f $X=2.955 $Y=1.745 $X2=0
+ $Y2=0
cc_235 N_A1_c_237_n N_A_27_368#_c_608_n 0.00958507f $X=3.405 $Y=1.745 $X2=0
+ $Y2=0
cc_236 N_A1_c_238_n N_A_27_368#_c_608_n 5.43202e-19 $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_237 N_A1_c_238_n N_A_27_368#_c_642_n 4.64231e-19 $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_238 N_A1_c_227_n N_Y_c_790_n 0.00133985f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_239 N_A1_c_228_n N_Y_c_790_n 0.00843072f $X=2.285 $Y=1.28 $X2=0 $Y2=0
cc_240 N_A1_c_229_n N_Y_c_790_n 0.00605915f $X=2.06 $Y=1.28 $X2=0 $Y2=0
cc_241 N_A1_c_235_n N_Y_c_790_n 0.00100621f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_242 N_A1_c_230_n N_Y_c_790_n 5.00179e-19 $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_243 N_A1_c_233_n N_Y_c_790_n 0.0341985f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A1_c_234_n N_Y_c_790_n 0.00153936f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_245 N_A1_c_227_n N_Y_c_791_n 0.0129676f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_246 N_A1_c_228_n N_Y_c_791_n 0.00643692f $X=2.285 $Y=1.28 $X2=0 $Y2=0
cc_247 N_A1_c_230_n N_Y_c_791_n 0.00641298f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_248 N_A1_c_233_n N_Y_c_791_n 0.0114135f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A1_c_230_n N_Y_c_833_n 0.0054833f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_250 N_A1_c_228_n N_Y_c_834_n 0.00385069f $X=2.285 $Y=1.28 $X2=0 $Y2=0
cc_251 N_A1_c_235_n N_Y_c_834_n 0.0121787f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_252 N_A1_c_236_n N_Y_c_834_n 0.0121787f $X=2.955 $Y=1.745 $X2=0 $Y2=0
cc_253 N_A1_c_237_n N_Y_c_834_n 0.0155276f $X=3.405 $Y=1.745 $X2=0 $Y2=0
cc_254 N_A1_c_238_n N_Y_c_834_n 0.0016208f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_255 N_A1_c_233_n N_Y_c_834_n 0.0693964f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A1_c_234_n N_Y_c_834_n 0.00177205f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_257 N_A1_c_235_n N_Y_c_794_n 0.0031019f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_258 N_A1_c_231_n N_Y_c_842_n 0.00605027f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_259 N_A1_c_232_n N_Y_c_842_n 0.0047069f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_260 N_A1_c_234_n N_Y_c_842_n 0.00196781f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_261 N_A1_c_236_n Y 8.3732e-19 $X=2.955 $Y=1.745 $X2=0 $Y2=0
cc_262 N_A1_c_237_n Y 0.00556536f $X=3.405 $Y=1.745 $X2=0 $Y2=0
cc_263 N_A1_c_238_n Y 0.00450986f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_264 N_A1_c_234_n Y 0.0167559f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_265 N_A1_c_231_n N_Y_c_792_n 0.00263107f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_266 N_A1_c_232_n N_Y_c_792_n 0.00413936f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_267 N_A1_c_233_n N_Y_c_792_n 0.0331256f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A1_c_234_n N_Y_c_792_n 0.0204398f $X=3.685 $Y=1.475 $X2=0 $Y2=0
cc_269 N_A1_c_235_n N_VPWR_c_892_n 0.00168541f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_270 N_A1_c_236_n N_VPWR_c_892_n 0.00361707f $X=2.955 $Y=1.745 $X2=0 $Y2=0
cc_271 N_A1_c_236_n N_VPWR_c_893_n 0.005209f $X=2.955 $Y=1.745 $X2=0 $Y2=0
cc_272 N_A1_c_237_n N_VPWR_c_893_n 0.005209f $X=3.405 $Y=1.745 $X2=0 $Y2=0
cc_273 N_A1_c_237_n N_VPWR_c_894_n 0.00307655f $X=3.405 $Y=1.745 $X2=0 $Y2=0
cc_274 N_A1_c_238_n N_VPWR_c_894_n 0.00317456f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_275 N_A1_c_238_n N_VPWR_c_895_n 0.005209f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_276 N_A1_c_235_n N_VPWR_c_907_n 0.00517089f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_277 N_A1_c_235_n N_VPWR_c_891_n 0.00977848f $X=2.405 $Y=1.745 $X2=0 $Y2=0
cc_278 N_A1_c_236_n N_VPWR_c_891_n 0.00982526f $X=2.955 $Y=1.745 $X2=0 $Y2=0
cc_279 N_A1_c_237_n N_VPWR_c_891_n 0.009828f $X=3.405 $Y=1.745 $X2=0 $Y2=0
cc_280 N_A1_c_238_n N_VPWR_c_891_n 0.00982351f $X=3.91 $Y=1.745 $X2=0 $Y2=0
cc_281 N_A1_c_227_n N_VGND_c_1036_n 0.00179989f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_282 N_A1_c_227_n N_VGND_c_1040_n 0.00278247f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_283 N_A1_c_230_n N_VGND_c_1040_n 0.00278271f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_284 N_A1_c_231_n N_VGND_c_1040_n 0.00278271f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_285 N_A1_c_232_n N_VGND_c_1040_n 0.00278271f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_286 N_A1_c_227_n N_VGND_c_1043_n 0.00359084f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_287 N_A1_c_230_n N_VGND_c_1043_n 0.00356595f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_288 N_A1_c_231_n N_VGND_c_1043_n 0.00355937f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_289 N_A1_c_232_n N_VGND_c_1043_n 0.0035414f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_290 N_A1_c_227_n N_A_325_74#_c_1133_n 0.00690005f $X=1.985 $Y=1.205 $X2=0
+ $Y2=0
cc_291 N_A1_c_230_n N_A_325_74#_c_1133_n 4.62714e-19 $X=2.485 $Y=1.205 $X2=0
+ $Y2=0
cc_292 N_A1_c_227_n N_A_325_74#_c_1134_n 0.00831967f $X=1.985 $Y=1.205 $X2=0
+ $Y2=0
cc_293 N_A1_c_230_n N_A_325_74#_c_1134_n 0.0136015f $X=2.485 $Y=1.205 $X2=0
+ $Y2=0
cc_294 N_A1_c_227_n N_A_325_74#_c_1135_n 0.00395315f $X=1.985 $Y=1.205 $X2=0
+ $Y2=0
cc_295 N_A1_c_230_n N_A_325_74#_c_1136_n 7.29988e-19 $X=2.485 $Y=1.205 $X2=0
+ $Y2=0
cc_296 N_A1_c_231_n N_A_325_74#_c_1136_n 7.86496e-19 $X=3.255 $Y=1.205 $X2=0
+ $Y2=0
cc_297 N_A1_c_233_n N_A_325_74#_c_1136_n 0.0373748f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_298 N_A1_c_234_n N_A_325_74#_c_1136_n 0.0136525f $X=3.685 $Y=1.475 $X2=0
+ $Y2=0
cc_299 N_A1_c_231_n N_A_325_74#_c_1137_n 0.0132525f $X=3.255 $Y=1.205 $X2=0
+ $Y2=0
cc_300 N_A1_c_232_n N_A_325_74#_c_1137_n 0.0133672f $X=3.685 $Y=1.205 $X2=0
+ $Y2=0
cc_301 N_A1_c_232_n N_A_325_74#_c_1140_n 0.00272146f $X=3.685 $Y=1.205 $X2=0
+ $Y2=0
cc_302 N_A1_c_234_n N_A_325_74#_c_1140_n 0.00579192f $X=3.685 $Y=1.475 $X2=0
+ $Y2=0
cc_303 N_A2_M1025_g N_A3_M1029_g 0.0112375f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A2_M1024_g A3 5.8843e-19 $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A2_M1025_g A3 0.00451503f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A2_c_343_n A3 0.018331f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_307 N_A2_c_344_n A3 0.00601056f $X=5.545 $Y=1.427 $X2=0 $Y2=0
cc_308 N_A2_c_343_n N_A3_c_435_n 2.09661e-19 $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_309 N_A2_c_344_n N_A3_c_435_n 0.0136196f $X=5.545 $Y=1.427 $X2=0 $Y2=0
cc_310 N_A2_M1003_g N_A_27_368#_c_633_n 8.84614e-19 $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A2_c_344_n N_A_27_368#_c_633_n 4.50786e-19 $X=5.545 $Y=1.427 $X2=0
+ $Y2=0
cc_312 N_A2_c_345_n N_A_27_368#_c_633_n 0.0236942f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_313 N_A2_M1003_g N_A_27_368#_c_634_n 0.00354169f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_314 N_A2_M1019_g N_A_27_368#_c_634_n 4.47398e-19 $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_315 N_A2_M1003_g N_A_27_368#_c_599_n 0.00672608f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A2_M1003_g N_A_27_368#_c_649_n 0.0132818f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_317 N_A2_M1019_g N_A_27_368#_c_649_n 0.0140162f $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_318 N_A2_c_343_n N_A_27_368#_c_649_n 0.0104059f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_319 N_A2_c_344_n N_A_27_368#_c_649_n 0.00103811f $X=5.545 $Y=1.427 $X2=0
+ $Y2=0
cc_320 N_A2_c_345_n N_A_27_368#_c_649_n 0.0268831f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_321 N_A2_M1003_g N_A_27_368#_c_600_n 6.17654e-19 $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_322 N_A2_M1019_g N_A_27_368#_c_600_n 0.0124872f $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_323 N_A2_M1024_g N_A_27_368#_c_600_n 0.0127647f $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_324 N_A2_M1025_g N_A_27_368#_c_600_n 6.3785e-19 $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A2_M1024_g N_A_27_368#_c_658_n 0.0139615f $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_326 N_A2_M1025_g N_A_27_368#_c_658_n 0.017354f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_327 N_A2_c_343_n N_A_27_368#_c_658_n 0.0154424f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_328 N_A2_c_344_n N_A_27_368#_c_658_n 0.00346396f $X=5.545 $Y=1.427 $X2=0
+ $Y2=0
cc_329 N_A2_M1024_g N_A_27_368#_c_601_n 6.10838e-19 $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_330 N_A2_M1025_g N_A_27_368#_c_601_n 0.0116523f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_331 N_A2_M1003_g N_A_27_368#_c_642_n 0.00204617f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_332 N_A2_M1003_g N_A_27_368#_c_609_n 6.06588e-19 $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_333 N_A2_M1019_g N_A_27_368#_c_609_n 0.00372949f $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_334 N_A2_M1024_g N_A_27_368#_c_609_n 0.00370988f $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A2_M1025_g N_A_27_368#_c_609_n 6.08944e-19 $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A2_c_343_n N_A_27_368#_c_609_n 0.0275631f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_337 N_A2_c_344_n N_A_27_368#_c_609_n 0.00245159f $X=5.545 $Y=1.427 $X2=0
+ $Y2=0
cc_338 N_A2_M1025_g N_A_27_368#_c_671_n 0.00105412f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_339 N_A2_c_345_n Y 0.0134646f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_340 N_A2_c_335_n N_Y_c_792_n 0.00102246f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_341 N_A2_c_345_n N_Y_c_792_n 0.0112767f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_342 N_A2_M1003_g N_VPWR_c_895_n 0.005209f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A2_M1003_g N_VPWR_c_896_n 0.00308519f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_344 N_A2_M1019_g N_VPWR_c_896_n 0.00316363f $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_345 N_A2_M1019_g N_VPWR_c_897_n 0.005209f $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_346 N_A2_M1024_g N_VPWR_c_897_n 0.005209f $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_347 N_A2_M1024_g N_VPWR_c_898_n 0.00306788f $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A2_M1025_g N_VPWR_c_898_n 0.00318542f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_349 N_A2_M1025_g N_VPWR_c_899_n 0.005209f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_350 N_A2_M1003_g N_VPWR_c_891_n 0.00982957f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A2_M1019_g N_VPWR_c_891_n 0.00982398f $X=4.87 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A2_M1024_g N_VPWR_c_891_n 0.00982754f $X=5.32 $Y=2.4 $X2=0 $Y2=0
cc_353 N_A2_M1025_g N_VPWR_c_891_n 0.00982193f $X=5.82 $Y=2.4 $X2=0 $Y2=0
cc_354 N_A2_c_335_n N_VGND_c_1040_n 0.00278247f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_355 N_A2_c_337_n N_VGND_c_1040_n 0.00278271f $X=4.685 $Y=1.205 $X2=0 $Y2=0
cc_356 N_A2_c_339_n N_VGND_c_1040_n 0.00278271f $X=5.115 $Y=1.205 $X2=0 $Y2=0
cc_357 N_A2_c_341_n N_VGND_c_1040_n 0.00278271f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_358 N_A2_c_335_n N_VGND_c_1043_n 0.00354796f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_359 N_A2_c_337_n N_VGND_c_1043_n 0.00354087f $X=4.685 $Y=1.205 $X2=0 $Y2=0
cc_360 N_A2_c_339_n N_VGND_c_1043_n 0.00353428f $X=5.115 $Y=1.205 $X2=0 $Y2=0
cc_361 N_A2_c_341_n N_VGND_c_1043_n 0.00358427f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_362 N_A2_c_335_n N_A_325_74#_c_1138_n 0.016033f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_363 N_A2_c_337_n N_A_325_74#_c_1138_n 0.0144954f $X=4.685 $Y=1.205 $X2=0
+ $Y2=0
cc_364 N_A2_c_339_n N_A_325_74#_c_1138_n 0.0136457f $X=5.115 $Y=1.205 $X2=0
+ $Y2=0
cc_365 N_A2_c_341_n N_A_325_74#_c_1138_n 0.014579f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_366 N_A2_c_335_n N_A_325_74#_c_1140_n 0.0106f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_367 N_A2_c_337_n N_A_325_74#_c_1140_n 8.0943e-19 $X=4.685 $Y=1.205 $X2=0
+ $Y2=0
cc_368 N_A2_c_345_n N_A_325_74#_c_1140_n 0.0139392f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_369 N_A2_c_335_n N_A_852_74#_c_1197_n 0.00183659f $X=4.185 $Y=1.205 $X2=0
+ $Y2=0
cc_370 N_A2_c_337_n N_A_852_74#_c_1197_n 0.013333f $X=4.685 $Y=1.205 $X2=0 $Y2=0
cc_371 N_A2_c_339_n N_A_852_74#_c_1197_n 0.0133316f $X=5.115 $Y=1.205 $X2=0
+ $Y2=0
cc_372 N_A2_c_341_n N_A_852_74#_c_1197_n 0.017437f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_373 N_A2_c_344_n N_A_852_74#_c_1197_n 0.020743f $X=5.545 $Y=1.427 $X2=0 $Y2=0
cc_374 N_A2_c_345_n N_A_852_74#_c_1197_n 0.0946862f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_375 N_A2_c_341_n N_A_1235_74#_c_1234_n 5.88287e-19 $X=5.545 $Y=1.205 $X2=0
+ $Y2=0
cc_376 N_A3_M1035_g N_A4_M1001_g 0.0108583f $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_377 N_A3_M1033_g N_A4_M1004_g 0.019323f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_378 A3 A4 0.0284998f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_379 N_A3_c_435_n A4 2.63965e-19 $X=7.825 $Y=1.515 $X2=0 $Y2=0
cc_380 A3 N_A4_c_523_n 0.00412885f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_381 N_A3_c_435_n N_A4_c_523_n 0.0193511f $X=7.825 $Y=1.515 $X2=0 $Y2=0
cc_382 N_A3_M1029_g N_A_27_368#_c_601_n 0.012177f $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_383 N_A3_M1030_g N_A_27_368#_c_601_n 6.3785e-19 $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_384 N_A3_M1029_g N_A_27_368#_c_674_n 0.0132272f $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_385 N_A3_M1030_g N_A_27_368#_c_674_n 0.0132272f $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_386 A3 N_A_27_368#_c_674_n 0.0431694f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_387 N_A3_c_435_n N_A_27_368#_c_674_n 7.54246e-19 $X=7.825 $Y=1.515 $X2=0
+ $Y2=0
cc_388 N_A3_M1029_g N_A_27_368#_c_602_n 6.10838e-19 $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_389 N_A3_M1030_g N_A_27_368#_c_602_n 0.0116961f $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_390 N_A3_M1034_g N_A_27_368#_c_602_n 0.0121813f $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_391 N_A3_M1035_g N_A_27_368#_c_602_n 6.3785e-19 $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_392 N_A3_M1034_g N_A_27_368#_c_682_n 0.0132272f $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A3_M1035_g N_A_27_368#_c_682_n 0.0132272f $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_394 A3 N_A_27_368#_c_682_n 0.0431694f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_395 N_A3_c_435_n N_A_27_368#_c_682_n 7.5354e-19 $X=7.825 $Y=1.515 $X2=0 $Y2=0
cc_396 N_A3_M1034_g N_A_27_368#_c_603_n 6.10838e-19 $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A3_M1035_g N_A_27_368#_c_603_n 0.0116908f $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A3_M1029_g N_A_27_368#_c_671_n 8.84614e-19 $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_399 A3 N_A_27_368#_c_671_n 0.0231426f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_400 N_A3_M1030_g N_A_27_368#_c_690_n 8.84614e-19 $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_401 N_A3_M1034_g N_A_27_368#_c_690_n 8.84614e-19 $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_402 A3 N_A_27_368#_c_690_n 0.0235495f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_403 N_A3_c_435_n N_A_27_368#_c_690_n 5.48413e-19 $X=7.825 $Y=1.515 $X2=0
+ $Y2=0
cc_404 N_A3_M1035_g N_A_27_368#_c_694_n 8.84614e-19 $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_405 A3 N_A_27_368#_c_694_n 0.0197305f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_406 N_A3_c_435_n N_A_27_368#_c_694_n 4.05442e-19 $X=7.825 $Y=1.515 $X2=0
+ $Y2=0
cc_407 N_A3_M1029_g N_VPWR_c_899_n 0.005209f $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_408 N_A3_M1029_g N_VPWR_c_900_n 0.00306788f $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_409 N_A3_M1030_g N_VPWR_c_900_n 0.00318542f $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_410 N_A3_M1030_g N_VPWR_c_901_n 0.005209f $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A3_M1034_g N_VPWR_c_901_n 0.005209f $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_412 N_A3_M1034_g N_VPWR_c_902_n 0.00306788f $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_413 N_A3_M1035_g N_VPWR_c_902_n 0.00187311f $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A3_M1035_g N_VPWR_c_903_n 5.1469e-19 $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_415 N_A3_M1035_g N_VPWR_c_908_n 0.005209f $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_416 N_A3_M1029_g N_VPWR_c_891_n 0.00982865f $X=6.27 $Y=2.4 $X2=0 $Y2=0
cc_417 N_A3_M1030_g N_VPWR_c_891_n 0.00982082f $X=6.77 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A3_M1034_g N_VPWR_c_891_n 0.00982754f $X=7.22 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A3_M1035_g N_VPWR_c_891_n 0.00982648f $X=7.72 $Y=2.4 $X2=0 $Y2=0
cc_420 N_A3_M1033_g N_VGND_c_1037_n 6.35276e-19 $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_421 N_A3_M1008_g N_VGND_c_1040_n 0.00291649f $X=6.535 $Y=0.74 $X2=0 $Y2=0
cc_422 N_A3_M1018_g N_VGND_c_1040_n 0.00291649f $X=6.965 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A3_M1021_g N_VGND_c_1040_n 0.00291649f $X=7.395 $Y=0.74 $X2=0 $Y2=0
cc_424 N_A3_M1033_g N_VGND_c_1040_n 0.00291649f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A3_M1008_g N_VGND_c_1043_n 0.0036412f $X=6.535 $Y=0.74 $X2=0 $Y2=0
cc_426 N_A3_M1018_g N_VGND_c_1043_n 0.00359121f $X=6.965 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A3_M1021_g N_VGND_c_1043_n 0.00359121f $X=7.395 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A3_M1033_g N_VGND_c_1043_n 0.00359219f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A3_M1008_g N_A_325_74#_c_1138_n 0.00326143f $X=6.535 $Y=0.74 $X2=0
+ $Y2=0
cc_430 N_A3_M1021_g N_A_852_74#_c_1196_n 0.00207464f $X=7.395 $Y=0.74 $X2=0
+ $Y2=0
cc_431 N_A3_M1033_g N_A_852_74#_c_1196_n 0.00466497f $X=7.825 $Y=0.74 $X2=0
+ $Y2=0
cc_432 N_A3_c_435_n N_A_852_74#_c_1196_n 0.00258952f $X=7.825 $Y=1.515 $X2=0
+ $Y2=0
cc_433 N_A3_M1008_g N_A_852_74#_c_1197_n 0.0177225f $X=6.535 $Y=0.74 $X2=0 $Y2=0
cc_434 N_A3_M1018_g N_A_852_74#_c_1197_n 0.0136379f $X=6.965 $Y=0.74 $X2=0 $Y2=0
cc_435 N_A3_M1021_g N_A_852_74#_c_1197_n 0.0118331f $X=7.395 $Y=0.74 $X2=0 $Y2=0
cc_436 A3 N_A_852_74#_c_1197_n 0.125425f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_437 N_A3_c_435_n N_A_852_74#_c_1197_n 0.0123736f $X=7.825 $Y=1.515 $X2=0
+ $Y2=0
cc_438 N_A3_M1008_g N_A_1235_74#_c_1227_n 0.00891446f $X=6.535 $Y=0.74 $X2=0
+ $Y2=0
cc_439 N_A3_M1018_g N_A_1235_74#_c_1227_n 0.0103412f $X=6.965 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A3_M1021_g N_A_1235_74#_c_1227_n 0.0102518f $X=7.395 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A3_M1033_g N_A_1235_74#_c_1227_n 0.014175f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_442 N_A3_M1033_g N_A_1235_74#_c_1230_n 0.0017668f $X=7.825 $Y=0.74 $X2=0
+ $Y2=0
cc_443 A3 N_A_1235_74#_c_1230_n 0.00721346f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_444 N_A3_M1008_g N_A_1235_74#_c_1234_n 0.0018597f $X=6.535 $Y=0.74 $X2=0
+ $Y2=0
cc_445 N_A4_M1001_g N_A_27_368#_c_697_n 0.0188185f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_446 N_A4_M1011_g N_A_27_368#_c_697_n 0.012931f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_447 A4 N_A_27_368#_c_697_n 0.0301004f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_448 N_A4_c_523_n N_A_27_368#_c_697_n 4.89356e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_449 N_A4_M1001_g N_A_27_368#_c_604_n 6.6858e-19 $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_450 N_A4_M1011_g N_A_27_368#_c_604_n 0.0120649f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_451 N_A4_M1031_g N_A_27_368#_c_604_n 0.0119382f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_452 N_A4_M1037_g N_A_27_368#_c_604_n 6.50516e-19 $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_453 N_A4_M1031_g N_A_27_368#_c_705_n 0.012931f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_454 N_A4_M1037_g N_A_27_368#_c_705_n 0.012931f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_455 A4 N_A_27_368#_c_705_n 0.0391869f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_456 N_A4_c_523_n N_A_27_368#_c_705_n 4.90767e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_457 N_A4_M1037_g N_A_27_368#_c_605_n 8.84614e-19 $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_458 A4 N_A_27_368#_c_605_n 0.0259449f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_459 N_A4_M1031_g N_A_27_368#_c_606_n 6.50516e-19 $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_460 N_A4_M1037_g N_A_27_368#_c_606_n 0.0121004f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_461 N_A4_M1011_g N_A_27_368#_c_713_n 8.84614e-19 $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_462 N_A4_M1031_g N_A_27_368#_c_713_n 8.84614e-19 $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_463 A4 N_A_27_368#_c_713_n 0.0235495f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_464 N_A4_c_523_n N_A_27_368#_c_713_n 5.54777e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_465 N_A4_M1001_g N_VPWR_c_903_n 0.0121308f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A4_M1011_g N_VPWR_c_903_n 0.002979f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_467 N_A4_M1031_g N_VPWR_c_904_n 0.0027763f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_468 N_A4_M1037_g N_VPWR_c_904_n 0.0027763f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_469 N_A4_M1011_g N_VPWR_c_905_n 0.005209f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_470 N_A4_M1031_g N_VPWR_c_905_n 0.005209f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A4_M1001_g N_VPWR_c_908_n 0.00460063f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_472 N_A4_M1037_g N_VPWR_c_909_n 0.005209f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_473 N_A4_M1001_g N_VPWR_c_891_n 0.00909121f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_474 N_A4_M1011_g N_VPWR_c_891_n 0.00982266f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_475 N_A4_M1031_g N_VPWR_c_891_n 0.00982266f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_476 N_A4_M1037_g N_VPWR_c_891_n 0.00986025f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A4_M1004_g N_VGND_c_1037_n 0.010782f $X=8.255 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A4_M1016_g N_VGND_c_1037_n 0.0106755f $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_479 N_A4_M1017_g N_VGND_c_1037_n 4.71636e-19 $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_480 N_A4_M1016_g N_VGND_c_1038_n 4.71636e-19 $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_481 N_A4_M1017_g N_VGND_c_1038_n 0.0105384f $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_482 N_A4_M1028_g N_VGND_c_1038_n 0.00392488f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_483 N_A4_M1004_g N_VGND_c_1040_n 0.00383152f $X=8.255 $Y=0.74 $X2=0 $Y2=0
cc_484 N_A4_M1016_g N_VGND_c_1041_n 0.00383152f $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_485 N_A4_M1017_g N_VGND_c_1041_n 0.00383152f $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_486 N_A4_M1028_g N_VGND_c_1042_n 0.00461464f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_487 N_A4_M1004_g N_VGND_c_1043_n 0.00757637f $X=8.255 $Y=0.74 $X2=0 $Y2=0
cc_488 N_A4_M1016_g N_VGND_c_1043_n 0.0075754f $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_489 N_A4_M1017_g N_VGND_c_1043_n 0.0075754f $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_490 N_A4_M1028_g N_VGND_c_1043_n 0.00911481f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_491 N_A4_M1004_g N_A_1235_74#_c_1229_n 0.0161035f $X=8.255 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_A4_M1016_g N_A_1235_74#_c_1229_n 0.0130453f $X=8.685 $Y=0.74 $X2=0
+ $Y2=0
cc_493 A4 N_A_1235_74#_c_1229_n 0.0398909f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_494 N_A4_c_523_n N_A_1235_74#_c_1229_n 0.00443556f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_495 N_A4_M1016_g N_A_1235_74#_c_1231_n 3.92313e-19 $X=8.685 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A4_M1017_g N_A_1235_74#_c_1231_n 3.92313e-19 $X=9.115 $Y=0.74 $X2=0
+ $Y2=0
cc_497 N_A4_M1017_g N_A_1235_74#_c_1232_n 0.0133256f $X=9.115 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A4_M1028_g N_A_1235_74#_c_1232_n 0.0146212f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_499 A4 N_A_1235_74#_c_1232_n 0.0766773f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_500 N_A4_c_523_n N_A_1235_74#_c_1232_n 0.00333587f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_501 N_A4_M1028_g N_A_1235_74#_c_1233_n 0.00160529f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_502 A4 N_A_1235_74#_c_1235_n 0.0146029f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_503 N_A4_c_523_n N_A_1235_74#_c_1235_n 0.00236901f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_504 N_A_27_368#_c_596_n N_Y_M1002_d 0.00213667f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_505 N_A_27_368#_c_598_n N_Y_M1009_d 0.00165831f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_506 N_A_27_368#_c_598_n N_Y_c_858_n 0.0117822f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_507 N_A_27_368#_M1012_s N_Y_c_834_n 0.00415381f $X=2.045 $Y=1.84 $X2=0 $Y2=0
cc_508 N_A_27_368#_M1010_d N_Y_c_834_n 0.00312423f $X=3.045 $Y=1.84 $X2=0 $Y2=0
cc_509 N_A_27_368#_c_628_n N_Y_c_834_n 0.0388605f $X=3.015 $Y=2.375 $X2=0 $Y2=0
cc_510 N_A_27_368#_c_630_n N_Y_c_834_n 0.023434f $X=3.97 $Y=2.375 $X2=0 $Y2=0
cc_511 N_A_27_368#_c_633_n N_Y_c_834_n 0.0108532f $X=4.135 $Y=2.12 $X2=0 $Y2=0
cc_512 N_A_27_368#_c_608_n N_Y_c_834_n 0.0171986f $X=3.18 $Y=2.375 $X2=0 $Y2=0
cc_513 N_A_27_368#_c_596_n N_Y_c_811_n 0.0173278f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_514 N_A_27_368#_M1007_s N_Y_c_815_n 0.00409304f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_515 N_A_27_368#_c_616_n N_Y_c_815_n 0.0189268f $X=1.28 $Y=2.405 $X2=0 $Y2=0
cc_516 N_A_27_368#_M1012_s N_Y_c_794_n 0.0014799f $X=2.045 $Y=1.84 $X2=0 $Y2=0
cc_517 N_A_27_368#_c_620_n N_Y_c_794_n 0.0172445f $X=2.18 $Y=2.46 $X2=0 $Y2=0
cc_518 N_A_27_368#_c_628_n N_VPWR_M1000_s 0.00534161f $X=3.015 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_519 N_A_27_368#_c_630_n N_VPWR_M1013_s 0.00532869f $X=3.97 $Y=2.375 $X2=0
+ $Y2=0
cc_520 N_A_27_368#_c_649_n N_VPWR_M1003_d 0.00445863f $X=4.93 $Y=2.035 $X2=0
+ $Y2=0
cc_521 N_A_27_368#_c_658_n N_VPWR_M1024_d 0.00549703f $X=5.88 $Y=2.035 $X2=0
+ $Y2=0
cc_522 N_A_27_368#_c_674_n N_VPWR_M1029_d 0.00410979f $X=6.83 $Y=2.035 $X2=0
+ $Y2=0
cc_523 N_A_27_368#_c_682_n N_VPWR_M1034_d 0.00410979f $X=7.78 $Y=2.035 $X2=0
+ $Y2=0
cc_524 N_A_27_368#_c_697_n N_VPWR_M1001_d 0.00314376f $X=8.73 $Y=2.035 $X2=0
+ $Y2=0
cc_525 N_A_27_368#_c_705_n N_VPWR_M1031_d 0.00314376f $X=9.63 $Y=2.035 $X2=0
+ $Y2=0
cc_526 N_A_27_368#_c_598_n N_VPWR_c_892_n 0.0119238f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_527 N_A_27_368#_c_628_n N_VPWR_c_892_n 0.0208278f $X=3.015 $Y=2.375 $X2=0
+ $Y2=0
cc_528 N_A_27_368#_c_608_n N_VPWR_c_892_n 0.0139233f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_529 N_A_27_368#_c_608_n N_VPWR_c_893_n 0.0144776f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_530 N_A_27_368#_c_630_n N_VPWR_c_894_n 0.0171667f $X=3.97 $Y=2.375 $X2=0
+ $Y2=0
cc_531 N_A_27_368#_c_599_n N_VPWR_c_894_n 0.0135735f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_532 N_A_27_368#_c_608_n N_VPWR_c_894_n 0.0122069f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_533 N_A_27_368#_c_599_n N_VPWR_c_895_n 0.0144623f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_534 N_A_27_368#_c_599_n N_VPWR_c_896_n 0.0177747f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_535 N_A_27_368#_c_649_n N_VPWR_c_896_n 0.0175734f $X=4.93 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_A_27_368#_c_600_n N_VPWR_c_896_n 0.0254585f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_537 N_A_27_368#_c_600_n N_VPWR_c_897_n 0.0144623f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_538 N_A_27_368#_c_600_n N_VPWR_c_898_n 0.0234083f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_539 N_A_27_368#_c_658_n N_VPWR_c_898_n 0.0167599f $X=5.88 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_A_27_368#_c_601_n N_VPWR_c_898_n 0.0266484f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_541 N_A_27_368#_c_601_n N_VPWR_c_899_n 0.0144623f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_542 N_A_27_368#_c_601_n N_VPWR_c_900_n 0.0234083f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_543 N_A_27_368#_c_674_n N_VPWR_c_900_n 0.0167599f $X=6.83 $Y=2.035 $X2=0
+ $Y2=0
cc_544 N_A_27_368#_c_602_n N_VPWR_c_900_n 0.0266484f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_545 N_A_27_368#_c_602_n N_VPWR_c_901_n 0.0144623f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_546 N_A_27_368#_c_602_n N_VPWR_c_902_n 0.0234083f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_547 N_A_27_368#_c_682_n N_VPWR_c_902_n 0.0167599f $X=7.78 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_A_27_368#_c_603_n N_VPWR_c_902_n 0.0266484f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_549 N_A_27_368#_c_603_n N_VPWR_c_903_n 0.0256025f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_550 N_A_27_368#_c_697_n N_VPWR_c_903_n 0.0148589f $X=8.73 $Y=2.035 $X2=0
+ $Y2=0
cc_551 N_A_27_368#_c_604_n N_VPWR_c_903_n 0.0234083f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_552 N_A_27_368#_c_604_n N_VPWR_c_904_n 0.0233699f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_553 N_A_27_368#_c_705_n N_VPWR_c_904_n 0.0126919f $X=9.63 $Y=2.035 $X2=0
+ $Y2=0
cc_554 N_A_27_368#_c_606_n N_VPWR_c_904_n 0.0233699f $X=9.795 $Y=2.815 $X2=0
+ $Y2=0
cc_555 N_A_27_368#_c_604_n N_VPWR_c_905_n 0.0144623f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_556 N_A_27_368#_c_596_n N_VPWR_c_907_n 0.0421297f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_557 N_A_27_368#_c_597_n N_VPWR_c_907_n 0.0235688f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_558 N_A_27_368#_c_598_n N_VPWR_c_907_n 0.0592384f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_559 N_A_27_368#_c_607_n N_VPWR_c_907_n 0.0235512f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_560 N_A_27_368#_c_603_n N_VPWR_c_908_n 0.014549f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_561 N_A_27_368#_c_606_n N_VPWR_c_909_n 0.014549f $X=9.795 $Y=2.815 $X2=0
+ $Y2=0
cc_562 N_A_27_368#_c_596_n N_VPWR_c_891_n 0.0236586f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_563 N_A_27_368#_c_597_n N_VPWR_c_891_n 0.0127152f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_564 N_A_27_368#_c_598_n N_VPWR_c_891_n 0.0326137f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_565 N_A_27_368#_c_599_n N_VPWR_c_891_n 0.0118344f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_566 N_A_27_368#_c_600_n N_VPWR_c_891_n 0.0118344f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_567 N_A_27_368#_c_601_n N_VPWR_c_891_n 0.0118344f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_568 N_A_27_368#_c_602_n N_VPWR_c_891_n 0.0118344f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_569 N_A_27_368#_c_603_n N_VPWR_c_891_n 0.0119743f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_570 N_A_27_368#_c_604_n N_VPWR_c_891_n 0.0118344f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_571 N_A_27_368#_c_606_n N_VPWR_c_891_n 0.0119743f $X=9.795 $Y=2.815 $X2=0
+ $Y2=0
cc_572 N_A_27_368#_c_607_n N_VPWR_c_891_n 0.0126924f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_573 N_A_27_368#_c_608_n N_VPWR_c_891_n 0.0118404f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_574 N_Y_c_834_n N_VPWR_M1000_s 0.00513422f $X=3.465 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_575 N_Y_c_834_n N_VPWR_M1013_s 0.00385614f $X=3.465 $Y=2.035 $X2=0 $Y2=0
cc_576 Y N_VPWR_M1013_s 0.00132878f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_577 N_Y_c_788_n N_VGND_M1032_d 0.00299905f $X=1.815 $Y=1.095 $X2=0 $Y2=0
cc_578 N_Y_c_787_n N_VGND_c_1035_n 0.0243474f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_579 N_Y_c_789_n N_VGND_c_1035_n 0.00555794f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_580 N_Y_c_787_n N_VGND_c_1036_n 0.0191765f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_581 N_Y_c_788_n N_VGND_c_1036_n 0.0219406f $X=1.815 $Y=1.095 $X2=0 $Y2=0
cc_582 N_Y_c_787_n N_VGND_c_1039_n 0.0145639f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_583 N_Y_c_787_n N_VGND_c_1043_n 0.0119984f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_584 N_Y_c_788_n N_A_325_74#_M1020_s 0.00258447f $X=1.815 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_585 N_Y_c_791_n N_A_325_74#_M1020_s 4.03947e-19 $X=2.27 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_586 N_Y_c_788_n N_A_325_74#_c_1133_n 0.0216365f $X=1.815 $Y=1.095 $X2=0 $Y2=0
cc_587 N_Y_M1020_d N_A_325_74#_c_1134_n 0.00250873f $X=2.06 $Y=0.37 $X2=0 $Y2=0
cc_588 N_Y_c_791_n N_A_325_74#_c_1134_n 0.00306797f $X=2.27 $Y=1.01 $X2=0 $Y2=0
cc_589 N_Y_c_833_n N_A_325_74#_c_1134_n 0.018913f $X=2.27 $Y=0.76 $X2=0 $Y2=0
cc_590 N_Y_c_791_n N_A_325_74#_c_1136_n 0.00586549f $X=2.27 $Y=1.01 $X2=0 $Y2=0
cc_591 N_Y_c_792_n N_A_325_74#_c_1136_n 0.00343886f $X=3.59 $Y=1.55 $X2=0 $Y2=0
cc_592 N_Y_M1026_d N_A_325_74#_c_1137_n 0.00176461f $X=3.33 $Y=0.37 $X2=0 $Y2=0
cc_593 N_Y_c_842_n N_A_325_74#_c_1137_n 0.0156869f $X=3.47 $Y=0.785 $X2=0 $Y2=0
cc_594 N_Y_c_842_n N_A_325_74#_c_1140_n 0.0194208f $X=3.47 $Y=0.785 $X2=0 $Y2=0
cc_595 N_VGND_c_1036_n N_A_325_74#_c_1133_n 0.027945f $X=1.21 $Y=0.675 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1040_n N_A_325_74#_c_1134_n 0.0423044f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_1043_n N_A_325_74#_c_1134_n 0.0239316f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_1036_n N_A_325_74#_c_1135_n 0.0121616f $X=1.21 $Y=0.675 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1040_n N_A_325_74#_c_1135_n 0.0233048f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_c_1043_n N_A_325_74#_c_1135_n 0.0126653f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1040_n N_A_325_74#_c_1137_n 0.0422287f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1043_n N_A_325_74#_c_1137_n 0.0238173f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_1040_n N_A_325_74#_c_1138_n 0.119831f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1043_n N_A_325_74#_c_1138_n 0.0658365f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_1040_n N_A_325_74#_c_1139_n 0.037994f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_c_1043_n N_A_325_74#_c_1139_n 0.0206052f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_607 N_VGND_c_1040_n N_A_325_74#_c_1140_n 0.0235688f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1043_n N_A_325_74#_c_1140_n 0.0127152f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_c_1043_n N_A_852_74#_c_1197_n 0.0137814f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_610 N_VGND_c_1037_n N_A_1235_74#_c_1228_n 0.00985092f $X=8.47 $Y=0.675 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1040_n N_A_1235_74#_c_1228_n 0.00758556f $X=8.305 $Y=0 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1043_n N_A_1235_74#_c_1228_n 0.00627867f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_613 N_VGND_M1004_s N_A_1235_74#_c_1229_n 0.00176461f $X=8.33 $Y=0.37 $X2=0
+ $Y2=0
cc_614 N_VGND_c_1037_n N_A_1235_74#_c_1229_n 0.0170777f $X=8.47 $Y=0.675 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1037_n N_A_1235_74#_c_1231_n 0.0182488f $X=8.47 $Y=0.675 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1038_n N_A_1235_74#_c_1231_n 0.0182488f $X=9.33 $Y=0.675 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1041_n N_A_1235_74#_c_1231_n 0.00749631f $X=9.165 $Y=0 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1043_n N_A_1235_74#_c_1231_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_M1017_s N_A_1235_74#_c_1232_n 0.00218982f $X=9.19 $Y=0.37 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1038_n N_A_1235_74#_c_1232_n 0.0185459f $X=9.33 $Y=0.675 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1038_n N_A_1235_74#_c_1233_n 0.00129215f $X=9.33 $Y=0.675 $X2=0
+ $Y2=0
cc_622 N_VGND_c_1042_n N_A_1235_74#_c_1233_n 0.011066f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_c_1043_n N_A_1235_74#_c_1233_n 0.00915947f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1040_n N_A_1235_74#_c_1234_n 0.0730035f $X=8.305 $Y=0 $X2=0
+ $Y2=0
cc_625 N_VGND_c_1043_n N_A_1235_74#_c_1234_n 0.0614975f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_626 N_A_325_74#_c_1138_n N_A_852_74#_M1005_d 0.00240933f $X=5.76 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_627 N_A_325_74#_c_1138_n N_A_852_74#_M1023_d 0.00171374f $X=5.76 $Y=0.515
+ $X2=0 $Y2=0
cc_628 N_A_325_74#_M1006_s N_A_852_74#_c_1197_n 0.0017749f $X=4.76 $Y=0.37 $X2=0
+ $Y2=0
cc_629 N_A_325_74#_M1027_s N_A_852_74#_c_1197_n 0.00429177f $X=5.62 $Y=0.37
+ $X2=0 $Y2=0
cc_630 N_A_325_74#_c_1138_n N_A_852_74#_c_1197_n 0.0970525f $X=5.76 $Y=0.515
+ $X2=0 $Y2=0
cc_631 N_A_325_74#_c_1140_n N_A_852_74#_c_1197_n 0.0135819f $X=3.97 $Y=0.515
+ $X2=0 $Y2=0
cc_632 N_A_325_74#_c_1138_n N_A_1235_74#_c_1234_n 0.0202095f $X=5.76 $Y=0.515
+ $X2=0 $Y2=0
cc_633 N_A_852_74#_c_1197_n N_A_1235_74#_M1008_d 0.00429177f $X=7.445 $Y=0.95
+ $X2=-0.19 $Y2=-0.245
cc_634 N_A_852_74#_c_1197_n N_A_1235_74#_M1018_d 0.00185845f $X=7.445 $Y=0.95
+ $X2=0 $Y2=0
cc_635 N_A_852_74#_M1008_s N_A_1235_74#_c_1227_n 0.00187648f $X=6.61 $Y=0.37
+ $X2=0 $Y2=0
cc_636 N_A_852_74#_M1021_s N_A_1235_74#_c_1227_n 0.00179007f $X=7.47 $Y=0.37
+ $X2=0 $Y2=0
cc_637 N_A_852_74#_c_1196_n N_A_1235_74#_c_1227_n 0.016201f $X=7.61 $Y=0.95
+ $X2=0 $Y2=0
cc_638 N_A_852_74#_c_1197_n N_A_1235_74#_c_1227_n 0.0487326f $X=7.445 $Y=0.95
+ $X2=0 $Y2=0
cc_639 N_A_852_74#_c_1196_n N_A_1235_74#_c_1230_n 0.00561736f $X=7.61 $Y=0.95
+ $X2=0 $Y2=0
cc_640 N_A_852_74#_c_1197_n N_A_1235_74#_c_1234_n 0.0208608f $X=7.445 $Y=0.95
+ $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o211ai_4.pex.spice
* Created: Fri Aug 28 17:53:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O211AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 55
r88 54 55 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.87 $Y=1.515
+ $X2=1.925 $Y2=1.515
r89 52 54 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.605 $Y=1.515
+ $X2=1.87 $Y2=1.515
r90 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.605
+ $Y=1.515 $X2=1.605 $Y2=1.515
r91 50 52 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.605 $Y2=1.515
r92 49 50 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.42 $Y=1.515
+ $X2=1.425 $Y2=1.515
r93 48 49 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=0.995 $Y=1.515
+ $X2=1.42 $Y2=1.515
r94 47 48 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.97 $Y=1.515
+ $X2=0.995 $Y2=1.515
r95 45 47 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.97 $Y2=1.515
r96 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r97 43 45 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=0.52 $Y=1.515
+ $X2=0.585 $Y2=1.515
r98 41 43 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.52 $Y2=1.515
r99 36 53 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.605 $Y2=1.565
r100 35 53 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.605 $Y2=1.565
r101 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r102 34 46 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r103 33 46 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r104 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.515
r105 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.74
r106 25 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.68
+ $X2=1.87 $Y2=1.515
r107 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.87 $Y=1.68
+ $X2=1.87 $Y2=2.4
r108 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.515
r109 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r110 17 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.68
+ $X2=1.42 $Y2=1.515
r111 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.42 $Y=1.68
+ $X2=1.42 $Y2=2.4
r112 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r113 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r114 9 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.68
+ $X2=0.97 $Y2=1.515
r115 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.97 $Y=1.68
+ $X2=0.97 $Y2=2.4
r116 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.68
+ $X2=0.52 $Y2=1.515
r117 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.52 $Y=1.68 $X2=0.52
+ $Y2=2.4
r118 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r119 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 33 51
r93 49 51 26.8524 $w=3.59e-07 $l=2e-07 $layer=POLY_cond $X=3.465 $Y=1.537
+ $X2=3.665 $Y2=1.537
r94 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.465
+ $Y=1.515 $X2=3.465 $Y2=1.515
r95 47 49 26.1811 $w=3.59e-07 $l=1.95e-07 $layer=POLY_cond $X=3.27 $Y=1.537
+ $X2=3.465 $Y2=1.537
r96 46 47 7.3844 $w=3.59e-07 $l=5.5e-08 $layer=POLY_cond $X=3.215 $Y=1.537
+ $X2=3.27 $Y2=1.537
r97 45 46 53.0334 $w=3.59e-07 $l=3.95e-07 $layer=POLY_cond $X=2.82 $Y=1.537
+ $X2=3.215 $Y2=1.537
r98 44 45 4.69916 $w=3.59e-07 $l=3.5e-08 $layer=POLY_cond $X=2.785 $Y=1.537
+ $X2=2.82 $Y2=1.537
r99 42 44 45.649 $w=3.59e-07 $l=3.4e-07 $layer=POLY_cond $X=2.445 $Y=1.537
+ $X2=2.785 $Y2=1.537
r100 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.445
+ $Y=1.515 $X2=2.445 $Y2=1.515
r101 40 42 10.0696 $w=3.59e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.537
+ $X2=2.445 $Y2=1.537
r102 39 40 2.01393 $w=3.59e-07 $l=1.5e-08 $layer=POLY_cond $X=2.355 $Y=1.537
+ $X2=2.37 $Y2=1.537
r103 32 33 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r104 32 50 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.465 $Y2=1.565
r105 31 50 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.465 $Y2=1.565
r106 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r107 30 43 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.445 $Y2=1.565
r108 29 43 7.63829 $w=4.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.445 $Y2=1.565
r109 26 51 14.0975 $w=3.59e-07 $l=2.347e-07 $layer=POLY_cond $X=3.77 $Y=1.725
+ $X2=3.665 $Y2=1.537
r110 26 28 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.77 $Y=1.725
+ $X2=3.77 $Y2=2.4
r111 22 51 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.665 $Y=1.35
+ $X2=3.665 $Y2=1.537
r112 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.665 $Y=1.35
+ $X2=3.665 $Y2=0.74
r113 19 47 18.9031 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=3.27 $Y=1.725
+ $X2=3.27 $Y2=1.537
r114 19 21 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.27 $Y=1.725
+ $X2=3.27 $Y2=2.4
r115 15 46 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.215 $Y=1.35
+ $X2=3.215 $Y2=1.537
r116 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.215 $Y=1.35
+ $X2=3.215 $Y2=0.74
r117 12 45 18.9031 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=2.82 $Y=1.725
+ $X2=2.82 $Y2=1.537
r118 12 14 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.82 $Y=1.725
+ $X2=2.82 $Y2=2.4
r119 8 44 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.785 $Y=1.35
+ $X2=2.785 $Y2=1.537
r120 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.785 $Y=1.35
+ $X2=2.785 $Y2=0.74
r121 5 40 18.9031 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=2.37 $Y=1.725
+ $X2=2.37 $Y2=1.537
r122 5 7 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.37 $Y=1.725
+ $X2=2.37 $Y2=2.4
r123 1 39 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=1.537
r124 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%B1 1 3 4 5 6 8 11 15 19 23 25 26 27 40
c72 19 0 1.87397e-19 $X=5.37 $Y=2.4
c73 11 0 1.83484e-19 $X=4.83 $Y=2.4
r74 38 40 10.2119 $w=3.54e-07 $l=7.5e-08 $layer=POLY_cond $X=5.295 $Y=1.432
+ $X2=5.37 $Y2=1.432
r75 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.295
+ $Y=1.515 $X2=5.295 $Y2=1.515
r76 33 35 29.274 $w=3.54e-07 $l=2.15e-07 $layer=POLY_cond $X=4.615 $Y=1.432
+ $X2=4.83 $Y2=1.432
r77 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.615
+ $Y=1.515 $X2=4.615 $Y2=1.515
r78 31 33 12.2542 $w=3.54e-07 $l=9e-08 $layer=POLY_cond $X=4.525 $Y=1.432
+ $X2=4.615 $Y2=1.432
r79 27 39 6.03022 $w=4.28e-07 $l=2.25e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.295 $Y2=1.565
r80 26 39 6.83426 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.295 $Y2=1.565
r81 26 34 11.3904 $w=4.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.615 $Y2=1.565
r82 25 34 1.47406 $w=4.28e-07 $l=5.5e-08 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.615 $Y2=1.565
r83 21 40 2.04237 $w=3.54e-07 $l=1.5e-08 $layer=POLY_cond $X=5.385 $Y=1.432
+ $X2=5.37 $Y2=1.432
r84 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.385 $Y=1.35
+ $X2=5.385 $Y2=0.74
r85 17 40 18.5736 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=5.37 $Y=1.68
+ $X2=5.37 $Y2=1.432
r86 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.37 $Y=1.68
+ $X2=5.37 $Y2=2.4
r87 13 38 46.2938 $w=3.54e-07 $l=3.4e-07 $layer=POLY_cond $X=4.955 $Y=1.432
+ $X2=5.295 $Y2=1.432
r88 13 35 17.0198 $w=3.54e-07 $l=1.25e-07 $layer=POLY_cond $X=4.955 $Y=1.432
+ $X2=4.83 $Y2=1.432
r89 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.955 $Y=1.35
+ $X2=4.955 $Y2=0.74
r90 9 35 18.5736 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=4.83 $Y=1.68
+ $X2=4.83 $Y2=1.432
r91 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.83 $Y=1.68 $X2=4.83
+ $Y2=2.4
r92 6 31 22.9014 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=4.525 $Y=1.185
+ $X2=4.525 $Y2=1.432
r93 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.525 $Y=1.185
+ $X2=4.525 $Y2=0.74
r94 4 31 26.5778 $w=3.54e-07 $l=2.06116e-07 $layer=POLY_cond $X=4.45 $Y=1.26
+ $X2=4.525 $Y2=1.432
r95 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.45 $Y=1.26 $X2=4.17
+ $Y2=1.26
r96 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.095 $Y=1.185
+ $X2=4.17 $Y2=1.26
r97 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.095 $Y=1.185
+ $X2=4.095 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%C1 3 7 11 15 17 21 23 27 29 30 31 32 47
r73 46 47 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.805 $Y=1.515
+ $X2=6.88 $Y2=1.515
r74 44 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.715 $Y=1.515
+ $X2=6.805 $Y2=1.515
r75 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.715
+ $Y=1.515 $X2=6.715 $Y2=1.515
r76 42 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.375 $Y=1.515
+ $X2=6.715 $Y2=1.515
r77 41 42 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.33 $Y=1.515
+ $X2=6.375 $Y2=1.515
r78 39 41 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=6.035 $Y=1.515
+ $X2=6.33 $Y2=1.515
r79 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.035
+ $Y=1.515 $X2=6.035 $Y2=1.515
r80 36 39 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.88 $Y=1.515
+ $X2=6.035 $Y2=1.515
r81 32 45 6.56625 $w=4.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.715 $Y2=1.565
r82 31 45 6.29823 $w=4.28e-07 $l=2.35e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.715 $Y2=1.565
r83 31 40 11.9264 $w=4.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.035 $Y2=1.565
r84 30 40 0.938035 $w=4.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=6.035 $Y2=1.565
r85 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.665 $Y=1.35
+ $X2=7.665 $Y2=0.79
r86 24 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.31 $Y=1.425
+ $X2=7.235 $Y2=1.425
r87 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.59 $Y=1.425
+ $X2=7.665 $Y2=1.35
r88 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.59 $Y=1.425
+ $X2=7.31 $Y2=1.425
r89 19 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.235 $Y=1.35
+ $X2=7.235 $Y2=1.425
r90 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.235 $Y=1.35
+ $X2=7.235 $Y2=0.79
r91 17 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.16 $Y=1.425
+ $X2=7.235 $Y2=1.425
r92 17 47 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.16 $Y=1.425
+ $X2=6.88 $Y2=1.425
r93 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.805 $Y=1.35
+ $X2=6.805 $Y2=1.515
r94 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.805 $Y=1.35
+ $X2=6.805 $Y2=0.79
r95 9 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.375 $Y=1.35
+ $X2=6.375 $Y2=1.515
r96 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.375 $Y=1.35
+ $X2=6.375 $Y2=0.79
r97 5 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.33 $Y=1.68
+ $X2=6.33 $Y2=1.515
r98 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.33 $Y=1.68 $X2=6.33
+ $Y2=2.4
r99 1 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.88 $Y=1.68
+ $X2=5.88 $Y2=1.515
r100 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.88 $Y=1.68 $X2=5.88
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%A_30_368# 1 2 3 4 5 16 18 20 24 26 28 31 32
+ 33 36 38 42 47 50
r72 40 42 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.045 $Y=2.905
+ $X2=4.045 $Y2=2.375
r73 39 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.21 $Y=2.99
+ $X2=3.085 $Y2=2.99
r74 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.88 $Y=2.99
+ $X2=4.045 $Y2=2.905
r75 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.88 $Y=2.99
+ $X2=3.21 $Y2=2.99
r76 34 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=2.905
+ $X2=3.085 $Y2=2.99
r77 34 36 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.085 $Y=2.905
+ $X2=3.085 $Y2=2.455
r78 32 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.96 $Y=2.99
+ $X2=3.085 $Y2=2.99
r79 32 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.96 $Y=2.99 $X2=2.26
+ $Y2=2.99
r80 29 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.095 $Y=2.905
+ $X2=2.26 $Y2=2.99
r81 29 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.095 $Y=2.905
+ $X2=2.095 $Y2=2.815
r82 28 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=2.12
+ $X2=2.095 $Y2=2.035
r83 28 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.095 $Y=2.12
+ $X2=2.095 $Y2=2.815
r84 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=2.035
+ $X2=1.195 $Y2=2.035
r85 26 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=2.035
+ $X2=2.095 $Y2=2.035
r86 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.93 $Y=2.035
+ $X2=1.36 $Y2=2.035
r87 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=2.12
+ $X2=1.195 $Y2=2.035
r88 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.195 $Y=2.12
+ $X2=1.195 $Y2=2.815
r89 21 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=2.035
+ $X2=0.295 $Y2=2.035
r90 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=2.035
+ $X2=1.195 $Y2=2.035
r91 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.03 $Y=2.035
+ $X2=0.46 $Y2=2.035
r92 16 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.295 $Y=2.12
+ $X2=0.295 $Y2=2.035
r93 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.295 $Y=2.12
+ $X2=0.295 $Y2=2.815
r94 5 42 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=3.86
+ $Y=1.84 $X2=4.045 $Y2=2.375
r95 4 36 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=1.84 $X2=3.045 $Y2=2.455
r96 3 49 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.84 $X2=2.095 $Y2=2.115
r97 3 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.84 $X2=2.095 $Y2=2.815
r98 2 47 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.84 $X2=1.195 $Y2=2.115
r99 2 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.84 $X2=1.195 $Y2=2.815
r100 1 45 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.115
r101 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%VPWR 1 2 3 4 5 20 24 28 30 34 36 40 42 44
+ 49 56 57 60 63 66 69 72
r91 73 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 72 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r93 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r94 70 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r95 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r96 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 57 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r101 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r102 54 72 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=7.29 $Y=3.33
+ $X2=6.865 $Y2=3.33
r103 54 56 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.29 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 50 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=1.645 $Y2=3.33
r105 50 52 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=4.08 $Y2=3.33
r106 49 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.605 $Y2=3.33
r107 49 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 48 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r111 45 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=3.33
+ $X2=0.745 $Y2=3.33
r112 45 47 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=3.33 $X2=1.2
+ $Y2=3.33
r113 44 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.645 $Y2=3.33
r114 44 47 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 42 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 42 64 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=1.68 $Y2=3.33
r117 42 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r118 38 72 3.24638 $w=8.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=3.245
+ $X2=6.865 $Y2=3.33
r119 38 40 11.3388 $w=8.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.865 $Y=3.245
+ $X2=6.865 $Y2=2.455
r120 37 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.77 $Y=3.33
+ $X2=5.605 $Y2=3.33
r121 36 72 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=6.44 $Y=3.33
+ $X2=6.865 $Y2=3.33
r122 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.44 $Y=3.33
+ $X2=5.77 $Y2=3.33
r123 32 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=3.245
+ $X2=5.605 $Y2=3.33
r124 32 34 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=5.605 $Y=3.245
+ $X2=5.605 $Y2=2.375
r125 31 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=3.33
+ $X2=4.605 $Y2=3.33
r126 30 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.44 $Y=3.33
+ $X2=5.605 $Y2=3.33
r127 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.44 $Y=3.33
+ $X2=4.77 $Y2=3.33
r128 26 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.605 $Y=3.245
+ $X2=4.605 $Y2=3.33
r129 26 28 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=4.605 $Y=3.245
+ $X2=4.605 $Y2=2.375
r130 22 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=3.33
r131 22 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=2.455
r132 18 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=3.33
r133 18 20 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=2.455
r134 5 40 150 $w=1.7e-07 $l=9.64676e-07 $layer=licon1_PDIFF $count=4 $X=6.42
+ $Y=1.84 $X2=7.125 $Y2=2.455
r135 4 34 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=5.46
+ $Y=1.84 $X2=5.605 $Y2=2.375
r136 3 28 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=4.46
+ $Y=1.84 $X2=4.605 $Y2=2.375
r137 2 24 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=1.84 $X2=1.645 $Y2=2.455
r138 1 20 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.84 $X2=0.745 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%Y 1 2 3 4 5 6 21 25 29 31 35 37 41 43 44 47
+ 52 54 56 58 59 60 61 62 63 77
c95 59 0 1.29151e-19 $X=7.455 $Y=1.095
c96 29 0 3.70881e-19 $X=5.105 $Y=2.815
r97 62 63 9.03161 $w=4.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.79 $Y=2.405
+ $X2=7.79 $Y2=2.775
r98 61 62 5.98354 $w=6.58e-07 $l=2.85e-07 $layer=LI1_cond $X=7.79 $Y=2.12
+ $X2=7.79 $Y2=2.405
r99 60 61 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.7 $Y=1.665 $X2=7.7
+ $Y2=2.035
r100 60 77 9.30395 $w=6.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.7 $Y=1.665
+ $X2=7.7 $Y2=1.55
r101 49 59 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.455 $Y=1.18
+ $X2=7.455 $Y2=1.095
r102 49 77 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=7.455 $Y=1.18
+ $X2=7.455 $Y2=1.55
r103 45 59 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.455 $Y=1.01
+ $X2=7.455 $Y2=1.095
r104 45 47 7.70202 $w=1.78e-07 $l=1.25e-07 $layer=LI1_cond $X=7.455 $Y=1.01
+ $X2=7.455 $Y2=0.885
r105 43 59 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.365 $Y=1.095
+ $X2=7.455 $Y2=1.095
r106 43 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.365 $Y=1.095
+ $X2=6.675 $Y2=1.095
r107 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.59 $Y=1.01
+ $X2=6.675 $Y2=1.095
r108 39 41 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.59 $Y=1.01
+ $X2=6.59 $Y2=0.885
r109 38 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=2.035
+ $X2=6.105 $Y2=2.035
r110 37 61 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.365 $Y=2.035
+ $X2=7.7 $Y2=2.035
r111 37 38 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=7.365 $Y=2.035
+ $X2=6.27 $Y2=2.035
r112 33 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.105 $Y=2.12
+ $X2=6.105 $Y2=2.035
r113 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.105 $Y=2.12
+ $X2=6.105 $Y2=2.815
r114 32 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=2.035
+ $X2=5.105 $Y2=2.035
r115 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.94 $Y=2.035
+ $X2=6.105 $Y2=2.035
r116 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.94 $Y=2.035
+ $X2=5.27 $Y2=2.035
r117 27 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=2.12
+ $X2=5.105 $Y2=2.035
r118 27 29 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.105 $Y=2.12
+ $X2=5.105 $Y2=2.815
r119 26 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=2.035
+ $X2=3.545 $Y2=2.035
r120 25 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.94 $Y=2.035
+ $X2=5.105 $Y2=2.035
r121 25 26 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.94 $Y=2.035
+ $X2=3.71 $Y2=2.035
r122 22 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=2.035
+ $X2=2.595 $Y2=2.035
r123 21 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=2.035
+ $X2=3.545 $Y2=2.035
r124 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.38 $Y=2.035
+ $X2=2.76 $Y2=2.035
r125 6 58 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.84 $X2=6.105 $Y2=2.115
r126 6 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.84 $X2=6.105 $Y2=2.815
r127 5 56 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.84 $X2=5.105 $Y2=2.115
r128 5 29 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.84 $X2=5.105 $Y2=2.815
r129 4 54 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.84 $X2=3.545 $Y2=2.115
r130 3 52 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=2.46
+ $Y=1.84 $X2=2.595 $Y2=2.115
r131 2 47 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=7.31
+ $Y=0.42 $X2=7.45 $Y2=0.885
r132 1 41 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=6.45
+ $Y=0.42 $X2=6.59 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%A_27_74# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 42 44 48 50 52 56 58 59 60 62 65
r111 64 65 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=1
+ $X2=4.905 $Y2=1
r112 54 56 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.6 $Y=1.01 $X2=5.6
+ $Y2=0.86
r113 52 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.435 $Y=1.095
+ $X2=5.6 $Y2=1.01
r114 52 65 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.435 $Y=1.095
+ $X2=4.905 $Y2=1.095
r115 51 62 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=1 $X2=3.88
+ $Y2=1
r116 50 64 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=4.725 $Y=1
+ $X2=4.74 $Y2=1
r117 50 51 24.3294 $w=3.58e-07 $l=7.6e-07 $layer=LI1_cond $X=4.725 $Y=1
+ $X2=3.965 $Y2=1
r118 46 62 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.88 $Y=0.82
+ $X2=3.88 $Y2=1
r119 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.88 $Y=0.82
+ $X2=3.88 $Y2=0.515
r120 45 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=1.095 $X2=3
+ $Y2=1.095
r121 44 62 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.795 $Y=1.095
+ $X2=3.88 $Y2=1
r122 44 45 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.795 $Y=1.095
+ $X2=3.085 $Y2=1.095
r123 40 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=1.01 $X2=3
+ $Y2=1.095
r124 40 42 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3 $Y=1.01 $X2=3
+ $Y2=0.515
r125 39 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.095
+ $X2=2.14 $Y2=1.095
r126 38 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=1.095 $X2=3
+ $Y2=1.095
r127 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.915 $Y=1.095
+ $X2=2.225 $Y2=1.095
r128 34 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.01
+ $X2=2.14 $Y2=1.095
r129 34 36 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.14 $Y=1.01
+ $X2=2.14 $Y2=0.515
r130 33 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.095
+ $X2=1.25 $Y2=1.095
r131 32 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.14 $Y2=1.095
r132 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=1.375 $Y2=1.095
r133 28 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.01
+ $X2=1.25 $Y2=1.095
r134 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.25 $Y=1.01
+ $X2=1.25 $Y2=0.515
r135 26 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=1.25 $Y2=1.095
r136 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=0.445 $Y2=1.095
r137 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r138 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r139 7 56 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.37 $X2=5.6 $Y2=0.86
r140 6 64 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.37 $X2=4.74 $Y2=0.95
r141 5 62 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.74
+ $Y=0.37 $X2=3.88 $Y2=0.965
r142 5 48 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.74
+ $Y=0.37 $X2=3.88 $Y2=0.515
r143 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.86
+ $Y=0.37 $X2=3 $Y2=0.515
r144 3 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r145 2 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r146 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 44
+ 57 58 61 64 67
r94 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r95 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r96 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 57 58 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r98 54 57 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=7.92
+ $Y2=0
r99 54 55 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r100 52 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r101 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r102 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r103 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.57
+ $Y2=0
r104 49 51 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=0
+ $X2=3.12 $Y2=0
r105 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r106 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r107 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r108 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r109 45 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.16 $Y2=0
r110 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.57
+ $Y2=0
r111 44 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.16
+ $Y2=0
r112 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r113 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r114 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r115 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r116 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r117 39 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r118 39 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r119 37 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r120 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r121 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r122 34 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r123 32 58 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r124 32 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r125 30 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=0
+ $X2=3.12 $Y2=0
r126 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.43
+ $Y2=0
r127 29 54 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.6
+ $Y2=0
r128 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.43
+ $Y2=0
r129 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.43 $Y2=0
r130 25 27 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.43 $Y2=0.635
r131 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0
r132 21 23 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0.635
r133 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r134 17 19 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.635
r135 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r136 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.595
r137 4 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.37 $X2=3.43 $Y2=0.635
r138 3 23 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.37 $X2=2.57 $Y2=0.635
r139 2 19 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.635
r140 1 15 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_4%A_834_74# 1 2 3 4 5 20 24 26 30 32 36 40 41
+ 42 43
r66 39 41 8.42273 $w=5.83e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.547
+ $X2=5.255 $Y2=0.547
r67 39 40 3.0054 $w=5.83e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.547
+ $X2=5.085 $Y2=0.547
r68 34 36 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.88 $Y=0.425
+ $X2=7.88 $Y2=0.565
r69 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.185 $Y=0.34
+ $X2=7.02 $Y2=0.34
r70 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=0.34
+ $X2=7.88 $Y2=0.425
r71 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.715 $Y=0.34
+ $X2=7.185 $Y2=0.34
r72 28 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.02 $Y=0.425
+ $X2=7.02 $Y2=0.34
r73 28 30 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.02 $Y=0.425
+ $X2=7.02 $Y2=0.66
r74 27 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.325 $Y=0.34
+ $X2=6.16 $Y2=0.34
r75 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=0.34
+ $X2=7.02 $Y2=0.34
r76 26 27 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.855 $Y=0.34
+ $X2=6.325 $Y2=0.34
r77 22 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=0.425
+ $X2=6.16 $Y2=0.34
r78 22 24 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.16 $Y=0.425
+ $X2=6.16 $Y2=0.565
r79 20 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.995 $Y=0.34
+ $X2=6.16 $Y2=0.34
r80 20 41 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.995 $Y=0.34
+ $X2=5.255 $Y2=0.34
r81 18 40 22.6112 $w=3.93e-07 $l=7.75e-07 $layer=LI1_cond $X=4.31 $Y=0.452
+ $X2=5.085 $Y2=0.452
r82 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.42 $X2=7.88 $Y2=0.565
r83 4 30 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=6.88
+ $Y=0.42 $X2=7.02 $Y2=0.66
r84 3 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.015
+ $Y=0.42 $X2=6.16 $Y2=0.565
r85 2 39 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.37 $X2=5.17 $Y2=0.595
r86 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.17
+ $Y=0.37 $X2=4.31 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__fa_1.pxi.spice
* Created: Fri Aug 28 17:34:44 2020
* 
x_PM_SKY130_FD_SC_MS__FA_1%A_69_260# N_A_69_260#_M1001_d N_A_69_260#_M1004_d
+ N_A_69_260#_M1021_g N_A_69_260#_M1026_g N_A_69_260#_c_160_n
+ N_A_69_260#_c_177_p N_A_69_260#_c_253_p N_A_69_260#_c_165_n
+ N_A_69_260#_c_171_p N_A_69_260#_c_166_n N_A_69_260#_c_161_n
+ N_A_69_260#_c_162_n N_A_69_260#_c_168_n N_A_69_260#_c_163_n
+ N_A_69_260#_c_182_p PM_SKY130_FD_SC_MS__FA_1%A_69_260#
x_PM_SKY130_FD_SC_MS__FA_1%A N_A_M1027_g N_A_M1011_g N_A_M1012_g N_A_M1016_g
+ N_A_M1019_g N_A_M1002_g N_A_M1022_g N_A_c_270_n N_A_c_271_n N_A_M1023_g
+ N_A_c_272_n N_A_c_273_n N_A_c_274_n N_A_c_275_n N_A_c_276_n N_A_c_277_n
+ N_A_c_278_n N_A_c_279_n N_A_c_460_p N_A_c_324_p N_A_c_280_n A N_A_c_282_n
+ N_A_c_283_n N_A_c_284_n N_A_c_285_n PM_SKY130_FD_SC_MS__FA_1%A
x_PM_SKY130_FD_SC_MS__FA_1%CIN N_CIN_M1001_g N_CIN_M1004_g N_CIN_M1008_g
+ N_CIN_M1005_g N_CIN_M1024_g N_CIN_M1020_g N_CIN_c_500_n N_CIN_c_501_n
+ N_CIN_c_502_n N_CIN_c_515_n N_CIN_c_516_n N_CIN_c_517_n N_CIN_c_503_n
+ N_CIN_c_504_n N_CIN_c_505_n CIN N_CIN_c_506_n N_CIN_c_507_n N_CIN_c_508_n
+ PM_SKY130_FD_SC_MS__FA_1%CIN
x_PM_SKY130_FD_SC_MS__FA_1%A_465_249# N_A_465_249#_M1017_d N_A_465_249#_M1013_d
+ N_A_465_249#_M1010_g N_A_465_249#_M1006_g N_A_465_249#_M1007_g
+ N_A_465_249#_c_679_n N_A_465_249#_M1018_g N_A_465_249#_c_680_n
+ N_A_465_249#_c_681_n N_A_465_249#_c_690_n N_A_465_249#_c_699_n
+ N_A_465_249#_c_691_n N_A_465_249#_c_700_n N_A_465_249#_c_714_n
+ N_A_465_249#_c_692_n N_A_465_249#_c_723_n N_A_465_249#_c_682_n
+ N_A_465_249#_c_683_n N_A_465_249#_c_684_n N_A_465_249#_c_685_n
+ N_A_465_249#_c_686_n N_A_465_249#_c_687_n N_A_465_249#_c_742_n
+ PM_SKY130_FD_SC_MS__FA_1%A_465_249#
x_PM_SKY130_FD_SC_MS__FA_1%B N_B_M1000_g N_B_c_875_n N_B_M1003_g N_B_c_877_n
+ N_B_c_878_n N_B_M1014_g N_B_c_865_n N_B_M1025_g N_B_c_880_n N_B_M1017_g
+ N_B_c_867_n N_B_M1013_g N_B_c_882_n N_B_M1009_g N_B_M1015_g N_B_c_870_n
+ N_B_c_884_n N_B_c_871_n N_B_c_885_n B N_B_c_872_n N_B_c_873_n
+ PM_SKY130_FD_SC_MS__FA_1%B
x_PM_SKY130_FD_SC_MS__FA_1%SUM N_SUM_M1026_s N_SUM_M1021_s N_SUM_c_1015_n
+ N_SUM_c_1016_n N_SUM_c_1012_n SUM SUM SUM PM_SKY130_FD_SC_MS__FA_1%SUM
x_PM_SKY130_FD_SC_MS__FA_1%VPWR N_VPWR_M1021_d N_VPWR_M1025_d N_VPWR_M1005_d
+ N_VPWR_M1022_d N_VPWR_M1007_s N_VPWR_c_1035_n N_VPWR_c_1036_n N_VPWR_c_1037_n
+ N_VPWR_c_1038_n N_VPWR_c_1039_n N_VPWR_c_1040_n N_VPWR_c_1041_n VPWR
+ N_VPWR_c_1042_n N_VPWR_c_1043_n N_VPWR_c_1044_n N_VPWR_c_1045_n
+ N_VPWR_c_1046_n N_VPWR_c_1034_n N_VPWR_c_1048_n N_VPWR_c_1049_n
+ N_VPWR_c_1050_n N_VPWR_c_1051_n PM_SKY130_FD_SC_MS__FA_1%VPWR
x_PM_SKY130_FD_SC_MS__FA_1%A_512_347# N_A_512_347#_M1006_d N_A_512_347#_M1012_d
+ N_A_512_347#_c_1152_n N_A_512_347#_c_1144_n N_A_512_347#_c_1147_n
+ N_A_512_347#_c_1145_n PM_SKY130_FD_SC_MS__FA_1%A_512_347#
x_PM_SKY130_FD_SC_MS__FA_1%A_1110_347# N_A_1110_347#_M1020_d
+ N_A_1110_347#_M1009_d N_A_1110_347#_c_1186_n N_A_1110_347#_c_1181_n
+ N_A_1110_347#_c_1185_n N_A_1110_347#_c_1182_n N_A_1110_347#_c_1183_n
+ PM_SKY130_FD_SC_MS__FA_1%A_1110_347#
x_PM_SKY130_FD_SC_MS__FA_1%COUT N_COUT_M1018_d N_COUT_M1007_d COUT COUT COUT
+ COUT COUT COUT COUT COUT PM_SKY130_FD_SC_MS__FA_1%COUT
x_PM_SKY130_FD_SC_MS__FA_1%VGND N_VGND_M1026_d N_VGND_M1014_d N_VGND_M1008_d
+ N_VGND_M1023_d N_VGND_M1018_s N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n
+ N_VGND_c_1229_n VGND N_VGND_c_1230_n N_VGND_c_1231_n N_VGND_c_1232_n
+ N_VGND_c_1233_n N_VGND_c_1234_n N_VGND_c_1235_n N_VGND_c_1236_n
+ N_VGND_c_1237_n N_VGND_c_1238_n N_VGND_c_1239_n PM_SKY130_FD_SC_MS__FA_1%VGND
x_PM_SKY130_FD_SC_MS__FA_1%A_501_75# N_A_501_75#_M1010_d N_A_501_75#_M1016_d
+ N_A_501_75#_c_1341_n N_A_501_75#_c_1338_n N_A_501_75#_c_1346_n
+ PM_SKY130_FD_SC_MS__FA_1%A_501_75#
x_PM_SKY130_FD_SC_MS__FA_1%A_1100_75# N_A_1100_75#_M1024_d N_A_1100_75#_M1015_d
+ N_A_1100_75#_c_1365_n N_A_1100_75#_c_1370_n N_A_1100_75#_c_1380_n
+ N_A_1100_75#_c_1371_n N_A_1100_75#_c_1366_n
+ PM_SKY130_FD_SC_MS__FA_1%A_1100_75#
cc_1 VNB N_A_69_260#_M1021_g 0.00165387f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A_69_260#_M1026_g 0.0264069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_A_69_260#_c_160_n 0.00139797f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_4 VNB N_A_69_260#_c_161_n 0.00272515f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_5 VNB N_A_69_260#_c_162_n 0.0345093f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_6 VNB N_A_69_260#_c_163_n 0.00289452f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.55
cc_7 VNB N_A_M1027_g 0.00638653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_M1011_g 0.0233458f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.63
cc_9 VNB N_A_M1012_g 0.00585096f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_10 VNB N_A_M1019_g 0.00570239f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.665
cc_11 VNB N_A_c_270_n 0.0254757f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.465
cc_12 VNB N_A_c_271_n 0.019979f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_13 VNB N_A_c_272_n 0.0200973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_c_273_n 0.00239261f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.55
cc_15 VNB N_A_c_274_n 0.0327627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_c_275_n 0.00740945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_c_276_n 0.00963516f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_18 VNB N_A_c_277_n 0.00224455f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_19 VNB N_A_c_278_n 0.00811052f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.3
cc_20 VNB N_A_c_279_n 0.0276772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_280_n 0.00338796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A 0.00205822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_282_n 0.0178818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_283_n 0.0324813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_c_284_n 0.0170005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_c_285_n 0.0376182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_CIN_M1001_g 0.0243526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_CIN_M1008_g 0.0252727f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_29 VNB N_CIN_M1024_g 0.025655f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.795
cc_30 VNB N_CIN_c_500_n 0.00103036f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.59
cc_31 VNB N_CIN_c_501_n 0.00370463f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.465
cc_32 VNB N_CIN_c_502_n 0.0223699f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_33 VNB N_CIN_c_503_n 3.94034e-19 $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=2.035
cc_34 VNB N_CIN_c_504_n 0.00392612f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.55
cc_35 VNB N_CIN_c_505_n 3.29665e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_CIN_c_506_n 0.0219645f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.3
cc_37 VNB N_CIN_c_507_n 0.0239451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_CIN_c_508_n 0.00255009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_465_249#_M1010_g 0.0261075f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_40 VNB N_A_465_249#_M1007_g 0.00759298f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.665
cc_41 VNB N_A_465_249#_c_679_n 0.0221372f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.795
cc_42 VNB N_A_465_249#_c_680_n 0.0386285f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.035
cc_43 VNB N_A_465_249#_c_681_n 0.0159332f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.12
cc_44 VNB N_A_465_249#_c_682_n 0.0050609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_465_249#_c_683_n 0.029447f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_46 VNB N_A_465_249#_c_684_n 7.33795e-19 $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_47 VNB N_A_465_249#_c_685_n 0.00629526f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_48 VNB N_A_465_249#_c_686_n 0.00566251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_465_249#_c_687_n 0.0217856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_B_M1000_g 0.0387714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_B_c_865_n 0.00627916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_B_M1025_g 0.020951f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.665
cc_53 VNB N_B_c_867_n 0.00553013f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.12
cc_54 VNB N_B_M1013_g 0.0181796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_B_M1015_g 0.0350093f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.55
cc_56 VNB N_B_c_870_n 0.0168615f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.665
cc_57 VNB N_B_c_871_n 0.014923f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=1.91
cc_58 VNB N_B_c_872_n 0.0426934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_B_c_873_n 0.00483187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_SUM_c_1012_n 0.0246106f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.75
cc_61 VNB SUM 0.0271795f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_62 VNB SUM 0.0094822f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.665
cc_63 VNB N_VPWR_c_1034_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB COUT 0.0263294f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.63
cc_65 VNB COUT 0.00845976f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_66 VNB COUT 0.0269902f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_67 VNB N_VGND_c_1226_n 0.018469f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_68 VNB N_VGND_c_1227_n 0.00826643f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.795
cc_69 VNB N_VGND_c_1228_n 0.00547714f $X=-0.19 $Y=-0.245 $X2=2.245 $Y2=2.59
cc_70 VNB N_VGND_c_1229_n 0.0139843f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_71 VNB N_VGND_c_1230_n 0.0343344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1231_n 0.0555224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1232_n 0.0578707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1233_n 0.019427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1234_n 0.0189924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1235_n 0.467822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1236_n 0.0144116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1237_n 0.00898487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1238_n 0.00477762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1239_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1100_75#_c_1365_n 0.00362777f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.63
cc_82 VNB N_A_1100_75#_c_1366_n 0.00389169f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.3
cc_83 VPB N_A_69_260#_M1021_g 0.0278523f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_84 VPB N_A_69_260#_c_165_n 0.00635828f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.795
cc_85 VPB N_A_69_260#_c_166_n 0.00219645f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_86 VPB N_A_69_260#_c_161_n 4.96285e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_87 VPB N_A_69_260#_c_168_n 0.00188689f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.795
cc_88 VPB N_A_M1027_g 0.0224003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_M1012_g 0.0209766f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_90 VPB N_A_M1019_g 0.0189437f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.665
cc_91 VPB N_A_M1022_g 0.0229867f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_92 VPB N_A_c_280_n 9.06676e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_c_285_n 0.00509374f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_CIN_M1004_g 0.0185843f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.63
cc_95 VPB N_CIN_M1005_g 0.0172776f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.75
cc_96 VPB N_CIN_M1020_g 0.0207922f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.12
cc_97 VPB N_CIN_c_500_n 0.0020408f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_98 VPB N_CIN_c_501_n 0.00190949f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.465
cc_99 VPB N_CIN_c_502_n 0.0048346f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_100 VPB N_CIN_c_515_n 0.0102933f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.795
cc_101 VPB N_CIN_c_516_n 8.36869e-19 $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.795
cc_102 VPB N_CIN_c_517_n 0.00462727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_CIN_c_503_n 6.01613e-19 $X=-0.19 $Y=1.66 $X2=1.14 $Y2=2.035
cc_104 VPB N_CIN_c_504_n 0.00366329f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=0.55
cc_105 VPB N_CIN_c_505_n 0.00315971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_CIN_c_506_n 0.00539003f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.3
cc_107 VPB N_CIN_c_507_n 0.00552786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_CIN_c_508_n 0.00392455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_465_249#_M1006_g 0.0182104f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_110 VPB N_A_465_249#_M1007_g 0.0311934f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=0.665
cc_111 VPB N_A_465_249#_c_690_n 0.00322579f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_112 VPB N_A_465_249#_c_691_n 0.00255223f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_113 VPB N_A_465_249#_c_692_n 9.89315e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_465_249#_c_682_n 0.00417624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_465_249#_c_686_n 0.00348732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_465_249#_c_687_n 0.00539452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_B_M1000_g 0.00518746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B_c_875_n 0.00593513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_B_M1003_g 0.0206748f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_120 VPB N_B_c_877_n 0.0926436f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_121 VPB N_B_c_878_n 0.0140921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_B_M1025_g 0.0361859f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=0.665
cc_123 VPB N_B_c_880_n 0.134922f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.665
cc_124 VPB N_B_M1013_g 0.0359536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_B_c_882_n 0.134592f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.465
cc_126 VPB N_B_M1009_g 0.0372548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_B_c_884_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_B_c_885_n 0.00898883f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=1.91
cc_129 VPB N_B_c_872_n 0.0264488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_B_c_873_n 0.0111011f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_SUM_c_1015_n 0.00919722f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_132 VPB N_SUM_c_1016_n 0.0416689f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_133 VPB N_SUM_c_1012_n 0.00751517f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.75
cc_134 VPB N_VPWR_c_1035_n 0.00837554f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.665
cc_135 VPB N_VPWR_c_1036_n 0.013201f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=2.59
cc_136 VPB N_VPWR_c_1037_n 0.0111988f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_137 VPB N_VPWR_c_1038_n 0.010007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_1039_n 0.0349078f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=0.55
cc_139 VPB N_VPWR_c_1040_n 0.0183142f $X=-0.19 $Y=1.66 $X2=2.245 $Y2=1.91
cc_140 VPB N_VPWR_c_1041_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_1042_n 0.0175529f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.3
cc_142 VPB N_VPWR_c_1043_n 0.0658504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_1044_n 0.0479018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_1045_n 0.0266344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_1046_n 0.0176701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1034_n 0.0921513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_1048_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_1049_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_1050_n 0.00936252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_1051_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_512_347#_c_1144_n 0.00277801f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_152 VPB N_A_512_347#_c_1145_n 0.00260929f $X=-0.19 $Y=1.66 $X2=0.705
+ $Y2=0.665
cc_153 VPB N_A_1110_347#_c_1181_n 0.00272685f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_154 VPB N_A_1110_347#_c_1182_n 0.0045747f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_155 VPB N_A_1110_347#_c_1183_n 0.0120917f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=0.75
cc_156 VPB COUT 0.054872f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_157 N_A_69_260#_M1021_g N_A_M1027_g 0.0255255f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_69_260#_c_165_n N_A_M1027_g 0.0127228f $X=1.055 $Y=1.795 $X2=0 $Y2=0
cc_159 N_A_69_260#_c_171_p N_A_M1027_g 2.3624e-19 $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_160 N_A_69_260#_c_161_n N_A_M1027_g 0.00333696f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A_69_260#_c_162_n N_A_M1027_g 0.00394048f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A_69_260#_c_168_n N_A_M1027_g 0.0114358f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_163 N_A_69_260#_M1026_g N_A_M1011_g 0.0205774f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_69_260#_c_160_n N_A_M1011_g 0.00519091f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_165 N_A_69_260#_c_177_p N_A_M1011_g 0.0119954f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_166 N_A_69_260#_M1001_d N_A_c_272_n 0.00388826f $X=1.965 $Y=0.375 $X2=0 $Y2=0
cc_167 N_A_69_260#_c_177_p N_A_c_272_n 0.0369432f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_168 N_A_69_260#_c_168_n N_A_c_272_n 2.80141e-19 $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_169 N_A_69_260#_c_163_n N_A_c_272_n 0.0209854f $X=2.105 $Y=0.55 $X2=0 $Y2=0
cc_170 N_A_69_260#_c_182_p N_A_c_272_n 0.00237094f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_171 N_A_69_260#_M1026_g N_A_c_278_n 3.94697e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_69_260#_c_160_n N_A_c_278_n 0.0190885f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_173 N_A_69_260#_c_177_p N_A_c_278_n 0.0149495f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A_69_260#_c_165_n N_A_c_278_n 0.0123444f $X=1.055 $Y=1.795 $X2=0 $Y2=0
cc_175 N_A_69_260#_c_161_n N_A_c_278_n 0.0181292f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_176 N_A_69_260#_c_162_n N_A_c_278_n 2.83375e-19 $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_177 N_A_69_260#_c_168_n N_A_c_278_n 0.0133509f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_178 N_A_69_260#_M1026_g N_A_c_279_n 0.00308693f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_69_260#_c_160_n N_A_c_279_n 2.60105e-19 $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_180 N_A_69_260#_c_177_p N_A_c_279_n 6.48184e-19 $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_181 N_A_69_260#_c_165_n N_A_c_279_n 7.93541e-19 $X=1.055 $Y=1.795 $X2=0 $Y2=0
cc_182 N_A_69_260#_c_161_n N_A_c_279_n 0.00100064f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_183 N_A_69_260#_c_162_n N_A_c_279_n 0.0161987f $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_184 N_A_69_260#_c_168_n N_A_c_279_n 0.00300549f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_185 N_A_69_260#_c_177_p N_CIN_M1001_g 0.00835085f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_186 N_A_69_260#_c_163_n N_CIN_M1001_g 0.00569455f $X=2.105 $Y=0.55 $X2=0
+ $Y2=0
cc_187 N_A_69_260#_c_171_p N_CIN_M1004_g 0.0146943f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_188 N_A_69_260#_c_166_n N_CIN_M1004_g 0.0132179f $X=2.245 $Y=2.59 $X2=0 $Y2=0
cc_189 N_A_69_260#_c_182_p N_CIN_M1004_g 0.00521617f $X=2.245 $Y=1.91 $X2=0
+ $Y2=0
cc_190 N_A_69_260#_M1004_d N_CIN_c_515_n 0.00191392f $X=2.11 $Y=1.735 $X2=0
+ $Y2=0
cc_191 N_A_69_260#_c_171_p N_CIN_c_515_n 0.0061202f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_192 N_A_69_260#_c_182_p N_CIN_c_515_n 0.0123284f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_193 N_A_69_260#_c_171_p N_CIN_c_516_n 0.0038604f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_194 N_A_69_260#_c_168_n N_CIN_c_516_n 0.00166828f $X=1.14 $Y=1.795 $X2=0
+ $Y2=0
cc_195 N_A_69_260#_c_182_p N_CIN_c_516_n 9.59784e-19 $X=2.245 $Y=1.91 $X2=0
+ $Y2=0
cc_196 N_A_69_260#_c_171_p N_CIN_c_504_n 0.0184192f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_197 N_A_69_260#_c_168_n N_CIN_c_504_n 0.0020521f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_198 N_A_69_260#_c_182_p N_CIN_c_504_n 0.0032161f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_199 N_A_69_260#_c_171_p N_CIN_c_506_n 6.63963e-19 $X=2.08 $Y=2.035 $X2=0
+ $Y2=0
cc_200 N_A_69_260#_c_163_n N_A_465_249#_M1010_g 0.00476897f $X=2.105 $Y=0.55
+ $X2=0 $Y2=0
cc_201 N_A_69_260#_c_166_n N_A_465_249#_M1006_g 0.00814816f $X=2.245 $Y=2.59
+ $X2=0 $Y2=0
cc_202 N_A_69_260#_c_182_p N_A_465_249#_M1006_g 0.00620517f $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_203 N_A_69_260#_c_182_p N_A_465_249#_c_699_n 0.00375855f $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_204 N_A_69_260#_c_182_p N_A_465_249#_c_700_n 4.07764e-19 $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_205 N_A_69_260#_c_182_p N_A_465_249#_c_686_n 0.0033839f $X=2.245 $Y=1.91
+ $X2=0 $Y2=0
cc_206 N_A_69_260#_c_177_p N_B_M1000_g 0.0107797f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_69_260#_c_168_n N_B_M1000_g 0.00403595f $X=1.14 $Y=1.795 $X2=0 $Y2=0
cc_208 N_A_69_260#_c_163_n N_B_M1000_g 0.00119451f $X=2.105 $Y=0.55 $X2=0 $Y2=0
cc_209 N_A_69_260#_c_182_p N_B_c_875_n 8.24231e-19 $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_210 N_A_69_260#_c_171_p N_B_M1003_g 0.0204934f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_211 N_A_69_260#_c_182_p N_B_M1003_g 0.00303893f $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_212 N_A_69_260#_c_166_n N_B_c_877_n 0.00564972f $X=2.245 $Y=2.59 $X2=0 $Y2=0
cc_213 N_A_69_260#_c_182_p N_B_M1025_g 5.75407e-19 $X=2.245 $Y=1.91 $X2=0 $Y2=0
cc_214 N_A_69_260#_M1021_g N_SUM_c_1015_n 0.00193811f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_215 N_A_69_260#_c_161_n N_SUM_c_1015_n 0.00305802f $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_216 N_A_69_260#_c_162_n N_SUM_c_1015_n 3.91434e-19 $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_217 N_A_69_260#_M1021_g N_SUM_c_1012_n 0.00407785f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_218 N_A_69_260#_M1026_g N_SUM_c_1012_n 0.0034597f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_69_260#_c_160_n N_SUM_c_1012_n 0.00833638f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_220 N_A_69_260#_c_161_n N_SUM_c_1012_n 0.0344362f $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_221 N_A_69_260#_c_162_n N_SUM_c_1012_n 0.00812898f $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_222 N_A_69_260#_M1026_g SUM 0.00206152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_69_260#_c_160_n SUM 0.0136155f $X=0.62 $Y=1.3 $X2=0 $Y2=0
cc_224 N_A_69_260#_c_162_n SUM 8.44384e-19 $X=0.51 $Y=1.465 $X2=0 $Y2=0
cc_225 N_A_69_260#_c_165_n N_VPWR_M1021_d 0.00166894f $X=1.055 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_226 N_A_69_260#_c_161_n N_VPWR_M1021_d 6.97173e-19 $X=0.51 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_69_260#_M1021_g N_VPWR_c_1035_n 0.0199208f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_228 N_A_69_260#_c_165_n N_VPWR_c_1035_n 0.0128182f $X=1.055 $Y=1.795 $X2=0
+ $Y2=0
cc_229 N_A_69_260#_c_161_n N_VPWR_c_1035_n 0.00809274f $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_230 N_A_69_260#_c_162_n N_VPWR_c_1035_n 3.0034e-19 $X=0.51 $Y=1.465 $X2=0
+ $Y2=0
cc_231 N_A_69_260#_M1021_g N_VPWR_c_1042_n 0.00460063f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_232 N_A_69_260#_c_166_n N_VPWR_c_1043_n 0.00741439f $X=2.245 $Y=2.59 $X2=0
+ $Y2=0
cc_233 N_A_69_260#_M1021_g N_VPWR_c_1034_n 0.00912261f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_234 N_A_69_260#_c_166_n N_VPWR_c_1034_n 0.00903331f $X=2.245 $Y=2.59 $X2=0
+ $Y2=0
cc_235 N_A_69_260#_c_171_p A_220_368# 0.0113135f $X=2.08 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_69_260#_c_168_n A_220_368# 0.00456947f $X=1.14 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_237 N_A_69_260#_c_171_p A_321_389# 0.0101896f $X=2.08 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_238 N_A_69_260#_c_166_n N_A_512_347#_c_1144_n 0.0103949f $X=2.245 $Y=2.59
+ $X2=0 $Y2=0
cc_239 N_A_69_260#_c_160_n N_VGND_M1026_d 0.00449182f $X=0.62 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_69_260#_c_177_p N_VGND_M1026_d 0.011913f $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_241 N_A_69_260#_c_253_p N_VGND_M1026_d 8.19949e-19 $X=0.705 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_242 N_A_69_260#_M1026_g N_VGND_c_1230_n 0.00806235f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_69_260#_c_177_p N_VGND_c_1230_n 0.0203993f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_244 N_A_69_260#_c_253_p N_VGND_c_1230_n 0.00778467f $X=0.705 $Y=0.665 $X2=0
+ $Y2=0
cc_245 N_A_69_260#_c_177_p N_VGND_c_1231_n 0.0161153f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_246 N_A_69_260#_c_163_n N_VGND_c_1231_n 0.0137352f $X=2.105 $Y=0.55 $X2=0
+ $Y2=0
cc_247 N_A_69_260#_M1026_g N_VGND_c_1235_n 0.00798259f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_69_260#_c_177_p N_VGND_c_1235_n 0.0279046f $X=1.94 $Y=0.665 $X2=0
+ $Y2=0
cc_249 N_A_69_260#_c_253_p N_VGND_c_1235_n 0.00315983f $X=0.705 $Y=0.665 $X2=0
+ $Y2=0
cc_250 N_A_69_260#_c_163_n N_VGND_c_1235_n 0.0117469f $X=2.105 $Y=0.55 $X2=0
+ $Y2=0
cc_251 N_A_69_260#_c_177_p A_237_75# 0.00339426f $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_69_260#_c_177_p A_315_75# 0.00339426f $X=1.94 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_253 N_A_69_260#_c_163_n N_A_501_75#_c_1338_n 0.0225265f $X=2.105 $Y=0.55
+ $X2=0 $Y2=0
cc_254 N_A_c_272_n N_CIN_M1001_g 0.010684f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_255 N_A_c_273_n N_CIN_M1008_g 0.00149115f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_256 N_A_c_274_n N_CIN_M1008_g 0.00627512f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_257 N_A_c_275_n N_CIN_M1008_g 0.0150364f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_258 N_A_c_324_p N_CIN_M1008_g 3.60835e-19 $X=4.545 $Y=1.012 $X2=0 $Y2=0
cc_259 A N_CIN_M1008_g 0.00111147f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_260 N_A_c_282_n N_CIN_M1008_g 0.0222612f $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_261 N_A_c_283_n N_CIN_M1008_g 0.0045952f $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_262 N_A_c_284_n N_CIN_M1008_g 0.0180648f $X=4.545 $Y=1.125 $X2=0 $Y2=0
cc_263 N_A_M1012_g N_CIN_M1005_g 0.0356843f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_264 N_A_M1019_g N_CIN_M1005_g 0.0430512f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_265 N_A_c_276_n N_CIN_M1024_g 0.01214f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_266 N_A_c_277_n N_CIN_M1024_g 0.00259916f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_267 N_A_c_285_n N_CIN_M1024_g 0.00372458f $X=6.045 $Y=1.185 $X2=0 $Y2=0
cc_268 N_A_M1022_g N_CIN_M1020_g 0.0252605f $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_269 N_A_M1019_g N_CIN_c_500_n 0.00273115f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_270 N_A_c_276_n N_CIN_c_500_n 0.0167049f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_271 A N_CIN_c_500_n 0.0108937f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_272 N_A_c_283_n N_CIN_c_500_n 6.2332e-19 $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_273 N_A_c_276_n N_CIN_c_501_n 0.0361598f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_274 N_A_c_277_n N_CIN_c_501_n 0.00342339f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_275 N_A_c_280_n N_CIN_c_501_n 0.0211108f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A_c_285_n N_CIN_c_501_n 3.27165e-19 $X=6.045 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A_c_276_n N_CIN_c_502_n 0.00438398f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_278 N_A_c_277_n N_CIN_c_502_n 7.67886e-19 $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_279 N_A_c_280_n N_CIN_c_502_n 8.83241e-19 $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_c_285_n N_CIN_c_502_n 0.0180988f $X=6.045 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A_M1012_g N_CIN_c_515_n 0.00651827f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_282 N_A_c_272_n N_CIN_c_515_n 0.0178463f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_283 N_A_c_273_n N_CIN_c_515_n 0.00969257f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_284 N_A_c_275_n N_CIN_c_515_n 0.00728431f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_285 N_A_M1027_g N_CIN_c_516_n 7.69397e-19 $X=1.01 $Y=2.34 $X2=0 $Y2=0
cc_286 N_A_c_272_n N_CIN_c_516_n 0.00192258f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_287 N_A_M1019_g N_CIN_c_517_n 0.00617249f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_288 N_A_c_275_n N_CIN_c_517_n 0.00507703f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_289 N_A_c_276_n N_CIN_c_517_n 0.00614904f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_290 A N_CIN_c_517_n 0.00968886f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_291 N_A_M1019_g N_CIN_c_503_n 0.00135683f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_292 N_A_c_275_n N_CIN_c_503_n 0.0021404f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_293 N_A_M1027_g N_CIN_c_504_n 0.00135687f $X=1.01 $Y=2.34 $X2=0 $Y2=0
cc_294 N_A_c_272_n N_CIN_c_504_n 0.0408998f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_295 N_A_c_278_n N_CIN_c_504_n 0.0123173f $X=1.05 $Y=1.005 $X2=0 $Y2=0
cc_296 N_A_c_279_n N_CIN_c_504_n 3.39404e-19 $X=1.05 $Y=1.385 $X2=0 $Y2=0
cc_297 N_A_M1019_g N_CIN_c_505_n 0.00128569f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_298 N_A_c_276_n N_CIN_c_505_n 0.00210963f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_299 N_A_c_272_n N_CIN_c_506_n 0.00468572f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_300 N_A_M1019_g N_CIN_c_507_n 0.00592873f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_301 N_A_c_273_n N_CIN_c_507_n 7.86199e-19 $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_302 N_A_c_274_n N_CIN_c_507_n 0.0206645f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_303 N_A_c_275_n N_CIN_c_507_n 0.0045209f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_304 A N_CIN_c_507_n 3.40268e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_305 N_A_c_283_n N_CIN_c_507_n 0.0132326f $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_306 N_A_M1012_g N_CIN_c_508_n 0.0023715f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_307 N_A_M1019_g N_CIN_c_508_n 0.00587022f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_308 N_A_c_273_n N_CIN_c_508_n 0.0124273f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_309 N_A_c_274_n N_CIN_c_508_n 0.00148765f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_310 N_A_c_275_n N_CIN_c_508_n 0.0261716f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_311 A N_CIN_c_508_n 0.0145682f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_312 N_A_c_283_n N_CIN_c_508_n 0.00111474f $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_313 N_A_c_276_n N_A_465_249#_M1017_d 0.00176461f $X=5.81 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_c_272_n N_A_465_249#_M1010_g 0.0150305f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_315 N_A_M1012_g N_A_465_249#_c_690_n 0.00184147f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_316 N_A_c_272_n N_A_465_249#_c_690_n 0.00808653f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_317 N_A_M1012_g N_A_465_249#_c_699_n 0.00307561f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_318 N_A_M1012_g N_A_465_249#_c_691_n 0.0141689f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_319 N_A_M1019_g N_A_465_249#_c_691_n 0.020728f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_320 N_A_M1022_g N_A_465_249#_c_691_n 5.7697e-19 $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_321 N_A_c_273_n N_A_465_249#_c_691_n 0.0042328f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_322 N_A_c_274_n N_A_465_249#_c_691_n 6.33241e-19 $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_323 A N_A_465_249#_c_691_n 0.00397556f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_324 N_A_c_283_n N_A_465_249#_c_691_n 4.38407e-19 $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_325 N_A_c_271_n N_A_465_249#_c_714_n 0.0037443f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_326 N_A_c_276_n N_A_465_249#_c_714_n 0.0400333f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_327 N_A_c_280_n N_A_465_249#_c_714_n 0.00489085f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A_c_285_n N_A_465_249#_c_714_n 0.00463693f $X=6.045 $Y=1.185 $X2=0
+ $Y2=0
cc_329 N_A_M1022_g N_A_465_249#_c_692_n 0.0134188f $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_330 N_A_c_270_n N_A_465_249#_c_692_n 0.00268633f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_331 N_A_c_276_n N_A_465_249#_c_692_n 0.00480772f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_332 N_A_c_280_n N_A_465_249#_c_692_n 0.0246553f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_333 N_A_c_285_n N_A_465_249#_c_692_n 0.00335987f $X=6.045 $Y=1.185 $X2=0
+ $Y2=0
cc_334 N_A_c_271_n N_A_465_249#_c_723_n 0.00729181f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_335 N_A_c_276_n N_A_465_249#_c_723_n 0.00366113f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_336 N_A_c_285_n N_A_465_249#_c_723_n 9.62124e-19 $X=6.045 $Y=1.185 $X2=0
+ $Y2=0
cc_337 N_A_M1022_g N_A_465_249#_c_682_n 0.00379848f $X=6.055 $Y=2.235 $X2=0
+ $Y2=0
cc_338 N_A_c_270_n N_A_465_249#_c_682_n 0.0104389f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_339 N_A_c_277_n N_A_465_249#_c_682_n 0.00600815f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_340 N_A_c_280_n N_A_465_249#_c_682_n 0.019392f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A_c_285_n N_A_465_249#_c_682_n 0.00252968f $X=6.045 $Y=1.185 $X2=0
+ $Y2=0
cc_342 N_A_c_270_n N_A_465_249#_c_683_n 0.00113076f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_343 N_A_c_271_n N_A_465_249#_c_683_n 0.00265319f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_344 N_A_c_270_n N_A_465_249#_c_684_n 0.00821163f $X=6.41 $Y=1.185 $X2=0 $Y2=0
cc_345 N_A_c_271_n N_A_465_249#_c_684_n 0.0070169f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_346 N_A_c_276_n N_A_465_249#_c_684_n 0.0114981f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_347 N_A_c_277_n N_A_465_249#_c_684_n 0.00335532f $X=5.895 $Y=1.32 $X2=0 $Y2=0
cc_348 N_A_c_280_n N_A_465_249#_c_684_n 0.00419754f $X=6.045 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A_c_285_n N_A_465_249#_c_684_n 0.00258911f $X=6.045 $Y=1.185 $X2=0
+ $Y2=0
cc_350 N_A_c_272_n N_A_465_249#_c_686_n 0.0313166f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_351 N_A_c_273_n N_A_465_249#_c_686_n 0.00649172f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_352 N_A_c_272_n N_A_465_249#_c_687_n 0.00432533f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_353 N_A_c_276_n N_A_465_249#_c_742_n 0.0161182f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_354 N_A_c_284_n N_A_465_249#_c_742_n 0.00105103f $X=4.545 $Y=1.125 $X2=0
+ $Y2=0
cc_355 N_A_M1027_g N_B_M1000_g 0.0556152f $X=1.01 $Y=2.34 $X2=0 $Y2=0
cc_356 N_A_M1011_g N_B_M1000_g 0.0538361f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_357 N_A_c_272_n N_B_M1000_g 0.0134851f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_358 N_A_c_278_n N_B_M1000_g 0.00373251f $X=1.05 $Y=1.005 $X2=0 $Y2=0
cc_359 N_A_c_279_n N_B_M1000_g 0.0196838f $X=1.05 $Y=1.385 $X2=0 $Y2=0
cc_360 N_A_c_272_n N_B_c_865_n 0.00112223f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_361 N_A_c_273_n N_B_c_865_n 0.00242117f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_362 N_A_c_274_n N_B_c_865_n 0.0167155f $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_363 N_A_c_282_n N_B_c_865_n 8.46159e-19 $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_364 N_A_M1012_g N_B_M1025_g 0.0386479f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_365 N_A_M1012_g N_B_c_880_n 0.0120239f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_366 N_A_M1019_g N_B_c_880_n 0.0124167f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_367 N_A_c_276_n N_B_c_867_n 0.00353286f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_368 A N_B_c_867_n 0.00199957f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_369 N_A_c_283_n N_B_c_867_n 0.0202139f $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_370 N_A_M1019_g N_B_M1013_g 0.0550732f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_371 N_A_M1022_g N_B_c_882_n 0.0123939f $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_372 N_A_c_271_n N_B_M1015_g 0.0176832f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_373 N_A_c_272_n N_B_c_870_n 0.0133079f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_374 N_A_c_282_n N_B_c_870_n 0.0208927f $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_375 N_A_c_276_n N_B_c_871_n 0.011404f $X=5.81 $Y=1.02 $X2=0 $Y2=0
cc_376 N_A_c_284_n N_B_c_871_n 0.0464607f $X=4.545 $Y=1.125 $X2=0 $Y2=0
cc_377 N_A_M1022_g N_B_c_872_n 0.0143519f $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_378 N_A_c_285_n N_B_c_872_n 0.0037349f $X=6.045 $Y=1.185 $X2=0 $Y2=0
cc_379 N_A_M1027_g N_VPWR_c_1035_n 0.00793598f $X=1.01 $Y=2.34 $X2=0 $Y2=0
cc_380 N_A_M1012_g N_VPWR_c_1036_n 0.00408951f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_381 N_A_M1012_g N_VPWR_c_1037_n 6.67826e-19 $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_382 N_A_M1019_g N_VPWR_c_1037_n 0.0138039f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_383 N_A_M1022_g N_VPWR_c_1038_n 0.00854888f $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_384 N_A_M1027_g N_VPWR_c_1043_n 0.0059286f $X=1.01 $Y=2.34 $X2=0 $Y2=0
cc_385 N_A_M1027_g N_VPWR_c_1034_n 0.00610055f $X=1.01 $Y=2.34 $X2=0 $Y2=0
cc_386 N_A_M1012_g N_VPWR_c_1034_n 0.00112709f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_387 N_A_M1019_g N_VPWR_c_1034_n 0.00100812f $X=4.505 $Y=2.235 $X2=0 $Y2=0
cc_388 N_A_M1022_g N_VPWR_c_1034_n 9.76808e-19 $X=6.055 $Y=2.235 $X2=0 $Y2=0
cc_389 N_A_M1012_g N_A_512_347#_c_1147_n 0.010397f $X=3.54 $Y=2.235 $X2=0 $Y2=0
cc_390 N_A_M1012_g N_A_512_347#_c_1145_n 0.00803122f $X=3.54 $Y=2.235 $X2=0
+ $Y2=0
cc_391 N_A_M1022_g N_A_1110_347#_c_1181_n 3.9799e-19 $X=6.055 $Y=2.235 $X2=0
+ $Y2=0
cc_392 N_A_M1022_g N_A_1110_347#_c_1185_n 0.0156586f $X=6.055 $Y=2.235 $X2=0
+ $Y2=0
cc_393 N_A_c_272_n N_VGND_M1014_d 0.00252521f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_394 N_A_c_460_p N_VGND_M1014_d 0.00106822f $X=3.465 $Y=1.005 $X2=0 $Y2=0
cc_395 N_A_c_275_n N_VGND_M1008_d 0.0035226f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_396 N_A_c_324_p N_VGND_M1008_d 0.0011084f $X=4.545 $Y=1.012 $X2=0 $Y2=0
cc_397 N_A_c_282_n N_VGND_c_1226_n 0.00314919f $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_398 N_A_c_275_n N_VGND_c_1227_n 0.0199906f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_399 N_A_c_324_p N_VGND_c_1227_n 0.00871655f $X=4.545 $Y=1.012 $X2=0 $Y2=0
cc_400 N_A_c_283_n N_VGND_c_1227_n 6.06098e-19 $X=4.545 $Y=1.29 $X2=0 $Y2=0
cc_401 N_A_c_284_n N_VGND_c_1227_n 0.016605f $X=4.545 $Y=1.125 $X2=0 $Y2=0
cc_402 N_A_c_271_n N_VGND_c_1228_n 9.17969e-19 $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_403 N_A_M1011_g N_VGND_c_1230_n 0.00407101f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_404 N_A_M1011_g N_VGND_c_1231_n 0.00317047f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_405 N_A_c_271_n N_VGND_c_1232_n 0.0027564f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_406 N_A_c_284_n N_VGND_c_1232_n 0.00379792f $X=4.545 $Y=1.125 $X2=0 $Y2=0
cc_407 N_A_M1011_g N_VGND_c_1235_n 0.00544287f $X=1.11 $Y=0.695 $X2=0 $Y2=0
cc_408 N_A_c_271_n N_VGND_c_1235_n 0.00544287f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_409 N_A_c_282_n N_VGND_c_1235_n 0.00544287f $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_410 N_A_c_284_n N_VGND_c_1235_n 0.00457201f $X=4.545 $Y=1.125 $X2=0 $Y2=0
cc_411 N_A_c_282_n N_VGND_c_1236_n 0.00397421f $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_412 N_A_c_272_n A_237_75# 0.00134267f $X=3.3 $Y=1.005 $X2=-0.19 $Y2=-0.245
cc_413 N_A_c_272_n A_315_75# 0.00134267f $X=3.3 $Y=1.005 $X2=-0.19 $Y2=-0.245
cc_414 N_A_c_272_n N_A_501_75#_M1010_d 0.0026214f $X=3.3 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_415 N_A_c_275_n N_A_501_75#_M1016_d 0.00176461f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_416 N_A_c_274_n N_A_501_75#_c_1341_n 5.87085e-19 $X=3.465 $Y=1.29 $X2=0 $Y2=0
cc_417 N_A_c_460_p N_A_501_75#_c_1341_n 0.0171542f $X=3.465 $Y=1.005 $X2=0 $Y2=0
cc_418 N_A_c_282_n N_A_501_75#_c_1341_n 0.00936066f $X=3.465 $Y=1.125 $X2=0
+ $Y2=0
cc_419 N_A_c_272_n N_A_501_75#_c_1338_n 0.0472581f $X=3.3 $Y=1.005 $X2=0 $Y2=0
cc_420 N_A_c_282_n N_A_501_75#_c_1338_n 7.1726e-19 $X=3.465 $Y=1.125 $X2=0 $Y2=0
cc_421 N_A_c_275_n N_A_501_75#_c_1346_n 0.0144331f $X=4.38 $Y=1.005 $X2=0 $Y2=0
cc_422 N_A_c_460_p N_A_501_75#_c_1346_n 0.00185147f $X=3.465 $Y=1.005 $X2=0
+ $Y2=0
cc_423 N_A_c_282_n N_A_501_75#_c_1346_n 0.00483163f $X=3.465 $Y=1.125 $X2=0
+ $Y2=0
cc_424 N_A_c_284_n N_A_501_75#_c_1346_n 3.54619e-19 $X=4.545 $Y=1.125 $X2=0
+ $Y2=0
cc_425 N_A_c_276_n A_936_75# 0.0048076f $X=5.81 $Y=1.02 $X2=-0.19 $Y2=-0.245
cc_426 N_A_c_276_n N_A_1100_75#_M1024_d 0.00536422f $X=5.81 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_427 N_A_c_271_n N_A_1100_75#_c_1365_n 0.0111244f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_428 N_A_c_285_n N_A_1100_75#_c_1365_n 3.90359e-19 $X=6.045 $Y=1.185 $X2=0
+ $Y2=0
cc_429 N_A_c_271_n N_A_1100_75#_c_1370_n 0.0104474f $X=6.485 $Y=1.11 $X2=0 $Y2=0
cc_430 N_A_c_271_n N_A_1100_75#_c_1371_n 0.00656693f $X=6.485 $Y=1.11 $X2=0
+ $Y2=0
cc_431 N_CIN_c_505_n N_A_465_249#_M1013_d 6.97845e-19 $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_432 N_CIN_M1001_g N_A_465_249#_M1010_g 0.0258374f $X=1.89 $Y=0.695 $X2=0
+ $Y2=0
cc_433 N_CIN_M1004_g N_A_465_249#_M1006_g 0.0151252f $X=2.02 $Y=2.235 $X2=0
+ $Y2=0
cc_434 N_CIN_c_515_n N_A_465_249#_M1006_g 0.0102784f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_435 N_CIN_c_515_n N_A_465_249#_c_690_n 0.0201297f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_436 N_CIN_c_508_n N_A_465_249#_c_690_n 0.00316685f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_437 N_CIN_M1005_g N_A_465_249#_c_691_n 0.0164857f $X=4.045 $Y=2.235 $X2=0
+ $Y2=0
cc_438 N_CIN_M1020_g N_A_465_249#_c_691_n 0.0247886f $X=5.46 $Y=2.235 $X2=0
+ $Y2=0
cc_439 N_CIN_c_500_n N_A_465_249#_c_691_n 0.0116945f $X=5.155 $Y=1.425 $X2=0
+ $Y2=0
cc_440 N_CIN_c_501_n N_A_465_249#_c_691_n 0.0189143f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_441 N_CIN_c_502_n N_A_465_249#_c_691_n 2.57098e-19 $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_442 N_CIN_c_515_n N_A_465_249#_c_691_n 0.0225933f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_443 N_CIN_c_517_n N_A_465_249#_c_691_n 0.0231918f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_444 N_CIN_c_503_n N_A_465_249#_c_691_n 0.00337097f $X=4.225 $Y=1.665 $X2=0
+ $Y2=0
cc_445 N_CIN_c_505_n N_A_465_249#_c_691_n 0.00520956f $X=5.04 $Y=1.665 $X2=0
+ $Y2=0
cc_446 N_CIN_c_507_n N_A_465_249#_c_691_n 4.09008e-19 $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_447 N_CIN_c_508_n N_A_465_249#_c_691_n 0.0165871f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_448 N_CIN_M1024_g N_A_465_249#_c_714_n 0.0107451f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_449 N_CIN_M1020_g N_A_465_249#_c_692_n 0.00656903f $X=5.46 $Y=2.235 $X2=0
+ $Y2=0
cc_450 N_CIN_c_501_n N_A_465_249#_c_692_n 0.00839037f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_451 N_CIN_c_502_n N_A_465_249#_c_692_n 0.0018928f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_452 N_CIN_M1024_g N_A_465_249#_c_723_n 0.00366676f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_453 N_CIN_M1024_g N_A_465_249#_c_684_n 3.99689e-19 $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_454 N_CIN_c_515_n N_A_465_249#_c_686_n 0.0252619f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_455 N_CIN_c_504_n N_A_465_249#_c_686_n 0.021248f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_456 N_CIN_c_506_n N_A_465_249#_c_686_n 3.97232e-19 $X=1.95 $Y=1.41 $X2=0
+ $Y2=0
cc_457 N_CIN_c_504_n N_A_465_249#_c_687_n 3.95958e-19 $X=1.68 $Y=1.665 $X2=0
+ $Y2=0
cc_458 N_CIN_c_506_n N_A_465_249#_c_687_n 0.0215538f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_459 N_CIN_M1024_g N_A_465_249#_c_742_n 0.00851142f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_460 N_CIN_M1001_g N_B_M1000_g 0.0555179f $X=1.89 $Y=0.695 $X2=0 $Y2=0
cc_461 N_CIN_M1004_g N_B_M1000_g 0.00485805f $X=2.02 $Y=2.235 $X2=0 $Y2=0
cc_462 N_CIN_c_516_n N_B_M1000_g 0.00332777f $X=1.825 $Y=1.665 $X2=0 $Y2=0
cc_463 N_CIN_c_504_n N_B_M1000_g 0.011517f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_464 N_CIN_c_506_n N_B_M1000_g 0.0213654f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_465 N_CIN_M1004_g N_B_c_875_n 0.0462101f $X=2.02 $Y=2.235 $X2=0 $Y2=0
cc_466 N_CIN_c_516_n N_B_c_875_n 0.0012981f $X=1.825 $Y=1.665 $X2=0 $Y2=0
cc_467 N_CIN_c_504_n N_B_c_875_n 0.00233633f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_468 N_CIN_M1004_g N_B_c_877_n 0.0123594f $X=2.02 $Y=2.235 $X2=0 $Y2=0
cc_469 N_CIN_c_515_n N_B_M1025_g 0.00282348f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_470 N_CIN_M1005_g N_B_c_880_n 0.0123711f $X=4.045 $Y=2.235 $X2=0 $Y2=0
cc_471 N_CIN_M1024_g N_B_c_867_n 0.00833387f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_472 N_CIN_M1020_g N_B_M1013_g 0.0263212f $X=5.46 $Y=2.235 $X2=0 $Y2=0
cc_473 N_CIN_c_500_n N_B_M1013_g 0.0199831f $X=5.155 $Y=1.425 $X2=0 $Y2=0
cc_474 N_CIN_c_501_n N_B_M1013_g 4.61068e-19 $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_475 N_CIN_c_502_n N_B_M1013_g 0.0214632f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_476 N_CIN_c_505_n N_B_M1013_g 0.00283871f $X=5.04 $Y=1.665 $X2=0 $Y2=0
cc_477 N_CIN_M1020_g N_B_c_882_n 0.0119f $X=5.46 $Y=2.235 $X2=0 $Y2=0
cc_478 N_CIN_M1024_g N_B_c_871_n 0.0214903f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_479 N_CIN_c_515_n N_VPWR_M1025_d 0.00207567f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_480 N_CIN_c_517_n N_VPWR_M1005_d 0.00156921f $X=4.895 $Y=1.665 $X2=0 $Y2=0
cc_481 N_CIN_c_503_n N_VPWR_M1005_d 0.00102642f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_482 N_CIN_c_508_n N_VPWR_M1005_d 7.68641e-19 $X=4.005 $Y=1.41 $X2=0 $Y2=0
cc_483 N_CIN_M1005_g N_VPWR_c_1037_n 0.0103639f $X=4.045 $Y=2.235 $X2=0 $Y2=0
cc_484 N_CIN_M1020_g N_VPWR_c_1038_n 5.32633e-19 $X=5.46 $Y=2.235 $X2=0 $Y2=0
cc_485 N_CIN_M1004_g N_VPWR_c_1034_n 0.00112709f $X=2.02 $Y=2.235 $X2=0 $Y2=0
cc_486 N_CIN_M1005_g N_VPWR_c_1034_n 9.455e-19 $X=4.045 $Y=2.235 $X2=0 $Y2=0
cc_487 N_CIN_M1020_g N_VPWR_c_1034_n 0.00112709f $X=5.46 $Y=2.235 $X2=0 $Y2=0
cc_488 N_CIN_c_515_n A_321_389# 8.6348e-19 $X=3.935 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_489 N_CIN_c_516_n A_321_389# 0.00169585f $X=1.825 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_490 N_CIN_c_504_n A_321_389# 9.79382e-19 $X=1.68 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_491 N_CIN_c_515_n N_A_512_347#_M1006_d 7.22664e-19 $X=3.935 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_492 N_CIN_c_515_n N_A_512_347#_M1012_d 0.00175187f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_493 N_CIN_c_508_n N_A_512_347#_M1012_d 0.00130917f $X=4.005 $Y=1.41 $X2=0
+ $Y2=0
cc_494 N_CIN_c_515_n N_A_512_347#_c_1152_n 0.00184039f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_495 N_CIN_c_515_n N_A_512_347#_c_1147_n 0.00148039f $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_496 N_CIN_M1005_g N_A_512_347#_c_1145_n 6.25506e-19 $X=4.045 $Y=2.235 $X2=0
+ $Y2=0
cc_497 N_CIN_c_517_n A_919_347# 0.00248251f $X=4.895 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_498 N_CIN_c_505_n A_919_347# 9.9595e-19 $X=5.04 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_499 N_CIN_M1020_g N_A_1110_347#_c_1186_n 0.00150746f $X=5.46 $Y=2.235 $X2=0
+ $Y2=0
cc_500 N_CIN_M1020_g N_A_1110_347#_c_1181_n 0.00410545f $X=5.46 $Y=2.235 $X2=0
+ $Y2=0
cc_501 N_CIN_M1008_g N_VGND_c_1226_n 0.00431894f $X=3.96 $Y=0.695 $X2=0 $Y2=0
cc_502 N_CIN_M1008_g N_VGND_c_1227_n 0.0064725f $X=3.96 $Y=0.695 $X2=0 $Y2=0
cc_503 N_CIN_M1001_g N_VGND_c_1231_n 0.00313567f $X=1.89 $Y=0.695 $X2=0 $Y2=0
cc_504 N_CIN_M1024_g N_VGND_c_1232_n 0.00316607f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_505 N_CIN_M1001_g N_VGND_c_1235_n 0.00544287f $X=1.89 $Y=0.695 $X2=0 $Y2=0
cc_506 N_CIN_M1008_g N_VGND_c_1235_n 0.00544287f $X=3.96 $Y=0.695 $X2=0 $Y2=0
cc_507 N_CIN_M1024_g N_VGND_c_1235_n 0.00544287f $X=5.425 $Y=0.695 $X2=0 $Y2=0
cc_508 N_CIN_M1008_g N_A_501_75#_c_1346_n 0.00449722f $X=3.96 $Y=0.695 $X2=0
+ $Y2=0
cc_509 N_CIN_M1024_g N_A_1100_75#_c_1365_n 0.00645788f $X=5.425 $Y=0.695 $X2=0
+ $Y2=0
cc_510 N_A_465_249#_M1006_g N_B_c_877_n 0.0123594f $X=2.47 $Y=2.235 $X2=0 $Y2=0
cc_511 N_A_465_249#_M1006_g N_B_M1025_g 0.0222381f $X=2.47 $Y=2.235 $X2=0 $Y2=0
cc_512 N_A_465_249#_c_690_n N_B_M1025_g 0.0136771f $X=3.03 $Y=1.71 $X2=0 $Y2=0
cc_513 N_A_465_249#_c_699_n N_B_M1025_g 0.0044772f $X=3.115 $Y=1.95 $X2=0 $Y2=0
cc_514 N_A_465_249#_c_700_n N_B_M1025_g 0.00473507f $X=3.2 $Y=2.035 $X2=0 $Y2=0
cc_515 N_A_465_249#_c_686_n N_B_M1025_g 0.00631868f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_516 N_A_465_249#_c_687_n N_B_M1025_g 0.0197606f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_517 N_A_465_249#_c_691_n N_B_M1013_g 0.0296746f $X=5.07 $Y=2.035 $X2=0 $Y2=0
cc_518 N_A_465_249#_c_691_n N_B_c_882_n 0.00400942f $X=5.07 $Y=2.035 $X2=0 $Y2=0
cc_519 N_A_465_249#_c_692_n N_B_M1009_g 0.00417312f $X=6.38 $Y=1.83 $X2=0 $Y2=0
cc_520 N_A_465_249#_c_680_n N_B_M1015_g 0.00323528f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_521 N_A_465_249#_c_682_n N_B_M1015_g 0.00187649f $X=6.465 $Y=1.745 $X2=0
+ $Y2=0
cc_522 N_A_465_249#_c_683_n N_B_M1015_g 0.0136844f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_523 N_A_465_249#_c_685_n N_B_M1015_g 0.00252947f $X=7.875 $Y=1.385 $X2=0
+ $Y2=0
cc_524 N_A_465_249#_M1010_g N_B_c_870_n 0.0225165f $X=2.43 $Y=0.695 $X2=0 $Y2=0
cc_525 N_A_465_249#_c_742_n N_B_c_871_n 0.00617071f $X=5.21 $Y=0.6 $X2=0 $Y2=0
cc_526 N_A_465_249#_M1007_g N_B_c_872_n 0.00241765f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_527 N_A_465_249#_c_680_n N_B_c_872_n 0.0130122f $X=8.055 $Y=1.385 $X2=0 $Y2=0
cc_528 N_A_465_249#_c_682_n N_B_c_872_n 0.00427741f $X=6.465 $Y=1.745 $X2=0
+ $Y2=0
cc_529 N_A_465_249#_c_683_n N_B_c_872_n 0.00363478f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_530 N_A_465_249#_c_685_n N_B_c_872_n 9.69264e-19 $X=7.875 $Y=1.385 $X2=0
+ $Y2=0
cc_531 N_A_465_249#_M1007_g N_B_c_873_n 0.00400384f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_532 N_A_465_249#_c_680_n N_B_c_873_n 9.22207e-19 $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_533 N_A_465_249#_c_692_n N_B_c_873_n 0.00232435f $X=6.38 $Y=1.83 $X2=0 $Y2=0
cc_534 N_A_465_249#_c_682_n N_B_c_873_n 0.0252217f $X=6.465 $Y=1.745 $X2=0 $Y2=0
cc_535 N_A_465_249#_c_683_n N_B_c_873_n 0.0511978f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_536 N_A_465_249#_c_685_n N_B_c_873_n 0.0138522f $X=7.875 $Y=1.385 $X2=0 $Y2=0
cc_537 N_A_465_249#_c_690_n N_VPWR_M1025_d 9.24637e-19 $X=3.03 $Y=1.71 $X2=0
+ $Y2=0
cc_538 N_A_465_249#_c_699_n N_VPWR_M1025_d 0.00188488f $X=3.115 $Y=1.95 $X2=0
+ $Y2=0
cc_539 N_A_465_249#_c_691_n N_VPWR_M1025_d 0.0050235f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_A_465_249#_c_700_n N_VPWR_M1025_d 0.00107668f $X=3.2 $Y=2.035 $X2=0
+ $Y2=0
cc_541 N_A_465_249#_c_691_n N_VPWR_M1005_d 0.00401302f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_542 N_A_465_249#_c_692_n N_VPWR_M1022_d 0.00946701f $X=6.38 $Y=1.83 $X2=0
+ $Y2=0
cc_543 N_A_465_249#_c_691_n N_VPWR_c_1037_n 0.0267454f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_544 N_A_465_249#_M1007_g N_VPWR_c_1039_n 0.0253037f $X=8.145 $Y=2.4 $X2=0
+ $Y2=0
cc_545 N_A_465_249#_c_680_n N_VPWR_c_1039_n 0.00273797f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_546 N_A_465_249#_c_685_n N_VPWR_c_1039_n 0.017603f $X=7.875 $Y=1.385 $X2=0
+ $Y2=0
cc_547 N_A_465_249#_c_691_n N_VPWR_c_1044_n 0.0093693f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_A_465_249#_M1007_g N_VPWR_c_1046_n 0.00460063f $X=8.145 $Y=2.4 $X2=0
+ $Y2=0
cc_549 N_A_465_249#_M1006_g N_VPWR_c_1034_n 0.00112709f $X=2.47 $Y=2.235 $X2=0
+ $Y2=0
cc_550 N_A_465_249#_M1007_g N_VPWR_c_1034_n 0.00912261f $X=8.145 $Y=2.4 $X2=0
+ $Y2=0
cc_551 N_A_465_249#_c_691_n N_VPWR_c_1034_n 0.0115317f $X=5.07 $Y=2.035 $X2=0
+ $Y2=0
cc_552 N_A_465_249#_c_690_n N_A_512_347#_M1006_d 6.05921e-19 $X=3.03 $Y=1.71
+ $X2=-0.19 $Y2=-0.245
cc_553 N_A_465_249#_c_686_n N_A_512_347#_M1006_d 0.00161164f $X=2.49 $Y=1.41
+ $X2=-0.19 $Y2=-0.245
cc_554 N_A_465_249#_c_691_n N_A_512_347#_M1012_d 0.00480643f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_A_465_249#_c_690_n N_A_512_347#_c_1152_n 0.00425453f $X=3.03 $Y=1.71
+ $X2=0 $Y2=0
cc_556 N_A_465_249#_c_686_n N_A_512_347#_c_1152_n 0.0108071f $X=2.49 $Y=1.41
+ $X2=0 $Y2=0
cc_557 N_A_465_249#_c_690_n N_A_512_347#_c_1147_n 0.00378555f $X=3.03 $Y=1.71
+ $X2=0 $Y2=0
cc_558 N_A_465_249#_c_691_n N_A_512_347#_c_1147_n 0.0234498f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_A_465_249#_c_700_n N_A_512_347#_c_1147_n 0.0086513f $X=3.2 $Y=2.035
+ $X2=0 $Y2=0
cc_560 N_A_465_249#_c_691_n N_A_512_347#_c_1145_n 0.0181738f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_561 N_A_465_249#_c_691_n A_919_347# 0.0108851f $X=5.07 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_562 N_A_465_249#_c_692_n N_A_1110_347#_M1020_d 0.0100312f $X=6.38 $Y=1.83
+ $X2=-0.19 $Y2=-0.245
cc_563 N_A_465_249#_c_691_n N_A_1110_347#_c_1186_n 0.0143691f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_564 N_A_465_249#_c_692_n N_A_1110_347#_c_1186_n 0.0197463f $X=6.38 $Y=1.83
+ $X2=0 $Y2=0
cc_565 N_A_465_249#_c_691_n N_A_1110_347#_c_1181_n 0.0391089f $X=5.07 $Y=2.035
+ $X2=0 $Y2=0
cc_566 N_A_465_249#_c_692_n N_A_1110_347#_c_1185_n 0.0388451f $X=6.38 $Y=1.83
+ $X2=0 $Y2=0
cc_567 N_A_465_249#_c_679_n COUT 0.0139505f $X=8.16 $Y=1.22 $X2=0 $Y2=0
cc_568 N_A_465_249#_c_679_n COUT 0.00387556f $X=8.16 $Y=1.22 $X2=0 $Y2=0
cc_569 N_A_465_249#_c_683_n COUT 0.00654086f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_570 N_A_465_249#_c_679_n COUT 0.0251717f $X=8.16 $Y=1.22 $X2=0 $Y2=0
cc_571 N_A_465_249#_c_683_n COUT 0.00131142f $X=7.71 $Y=1.065 $X2=0 $Y2=0
cc_572 N_A_465_249#_c_685_n COUT 0.0238637f $X=7.875 $Y=1.385 $X2=0 $Y2=0
cc_573 N_A_465_249#_c_683_n N_VGND_M1023_d 0.00531596f $X=7.71 $Y=1.065 $X2=0
+ $Y2=0
cc_574 N_A_465_249#_c_683_n N_VGND_M1018_s 0.00320163f $X=7.71 $Y=1.065 $X2=0
+ $Y2=0
cc_575 N_A_465_249#_c_742_n N_VGND_c_1227_n 0.00896174f $X=5.21 $Y=0.6 $X2=0
+ $Y2=0
cc_576 N_A_465_249#_c_679_n N_VGND_c_1229_n 0.00564712f $X=8.16 $Y=1.22 $X2=0
+ $Y2=0
cc_577 N_A_465_249#_c_680_n N_VGND_c_1229_n 0.00116085f $X=8.055 $Y=1.385 $X2=0
+ $Y2=0
cc_578 N_A_465_249#_c_683_n N_VGND_c_1229_n 0.0189083f $X=7.71 $Y=1.065 $X2=0
+ $Y2=0
cc_579 N_A_465_249#_M1010_g N_VGND_c_1231_n 0.00430851f $X=2.43 $Y=0.695 $X2=0
+ $Y2=0
cc_580 N_A_465_249#_c_714_n N_VGND_c_1232_n 0.00284331f $X=6.15 $Y=0.68 $X2=0
+ $Y2=0
cc_581 N_A_465_249#_c_742_n N_VGND_c_1232_n 0.00841586f $X=5.21 $Y=0.6 $X2=0
+ $Y2=0
cc_582 N_A_465_249#_c_679_n N_VGND_c_1234_n 0.00434272f $X=8.16 $Y=1.22 $X2=0
+ $Y2=0
cc_583 N_A_465_249#_M1010_g N_VGND_c_1235_n 0.00544287f $X=2.43 $Y=0.695 $X2=0
+ $Y2=0
cc_584 N_A_465_249#_c_679_n N_VGND_c_1235_n 0.00828888f $X=8.16 $Y=1.22 $X2=0
+ $Y2=0
cc_585 N_A_465_249#_c_714_n N_VGND_c_1235_n 0.00593054f $X=6.15 $Y=0.68 $X2=0
+ $Y2=0
cc_586 N_A_465_249#_c_742_n N_VGND_c_1235_n 0.0109111f $X=5.21 $Y=0.6 $X2=0
+ $Y2=0
cc_587 N_A_465_249#_M1010_g N_A_501_75#_c_1338_n 0.00433986f $X=2.43 $Y=0.695
+ $X2=0 $Y2=0
cc_588 N_A_465_249#_c_714_n N_A_1100_75#_M1024_d 0.0217685f $X=6.15 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_589 N_A_465_249#_c_723_n N_A_1100_75#_M1024_d 0.00690281f $X=6.235 $Y=0.98
+ $X2=-0.19 $Y2=-0.245
cc_590 N_A_465_249#_c_684_n N_A_1100_75#_M1024_d 0.00149425f $X=6.55 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_591 N_A_465_249#_c_683_n N_A_1100_75#_M1015_d 0.00237104f $X=7.71 $Y=1.065
+ $X2=0 $Y2=0
cc_592 N_A_465_249#_c_714_n N_A_1100_75#_c_1365_n 0.0528994f $X=6.15 $Y=0.68
+ $X2=0 $Y2=0
cc_593 N_A_465_249#_c_684_n N_A_1100_75#_c_1365_n 0.00306218f $X=6.55 $Y=1.065
+ $X2=0 $Y2=0
cc_594 N_A_465_249#_c_714_n N_A_1100_75#_c_1370_n 0.0035178f $X=6.15 $Y=0.68
+ $X2=0 $Y2=0
cc_595 N_A_465_249#_c_683_n N_A_1100_75#_c_1380_n 0.0387969f $X=7.71 $Y=1.065
+ $X2=0 $Y2=0
cc_596 N_A_465_249#_c_714_n N_A_1100_75#_c_1371_n 0.0109254f $X=6.15 $Y=0.68
+ $X2=0 $Y2=0
cc_597 N_A_465_249#_c_723_n N_A_1100_75#_c_1371_n 0.00350045f $X=6.235 $Y=0.98
+ $X2=0 $Y2=0
cc_598 N_A_465_249#_c_684_n N_A_1100_75#_c_1371_n 0.00864961f $X=6.55 $Y=1.065
+ $X2=0 $Y2=0
cc_599 N_A_465_249#_c_679_n N_A_1100_75#_c_1366_n 7.49371e-19 $X=8.16 $Y=1.22
+ $X2=0 $Y2=0
cc_600 N_A_465_249#_c_683_n N_A_1100_75#_c_1366_n 0.020765f $X=7.71 $Y=1.065
+ $X2=0 $Y2=0
cc_601 N_B_M1003_g N_VPWR_c_1035_n 0.00700155f $X=1.515 $Y=2.445 $X2=0 $Y2=0
cc_602 N_B_M1025_g N_VPWR_c_1036_n 0.0133115f $X=2.955 $Y=2.235 $X2=0 $Y2=0
cc_603 N_B_c_880_n N_VPWR_c_1036_n 0.0242838f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_604 N_B_c_880_n N_VPWR_c_1037_n 0.0254328f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_605 N_B_M1013_g N_VPWR_c_1037_n 0.0075423f $X=5.01 $Y=2.235 $X2=0 $Y2=0
cc_606 N_B_c_882_n N_VPWR_c_1038_n 0.0430354f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_607 N_B_M1009_g N_VPWR_c_1038_n 0.0222068f $X=6.89 $Y=2.31 $X2=0 $Y2=0
cc_608 N_B_c_880_n N_VPWR_c_1040_n 0.0207894f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_609 N_B_c_878_n N_VPWR_c_1043_n 0.0539698f $X=1.605 $Y=3.15 $X2=0 $Y2=0
cc_610 N_B_c_880_n N_VPWR_c_1044_n 0.0527614f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_611 N_B_c_882_n N_VPWR_c_1045_n 0.0060312f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_612 N_B_c_877_n N_VPWR_c_1034_n 0.0463698f $X=2.865 $Y=3.15 $X2=0 $Y2=0
cc_613 N_B_c_878_n N_VPWR_c_1034_n 0.0134575f $X=1.605 $Y=3.15 $X2=0 $Y2=0
cc_614 N_B_c_880_n N_VPWR_c_1034_n 0.0468212f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_615 N_B_c_882_n N_VPWR_c_1034_n 0.0432123f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_616 N_B_c_884_n N_VPWR_c_1034_n 0.0109459f $X=2.955 $Y=3.15 $X2=0 $Y2=0
cc_617 N_B_c_885_n N_VPWR_c_1034_n 0.0101348f $X=5.01 $Y=3.15 $X2=0 $Y2=0
cc_618 N_B_c_877_n N_A_512_347#_c_1144_n 0.00333139f $X=2.865 $Y=3.15 $X2=0
+ $Y2=0
cc_619 N_B_M1025_g N_A_512_347#_c_1147_n 0.018246f $X=2.955 $Y=2.235 $X2=0 $Y2=0
cc_620 N_B_c_880_n N_A_512_347#_c_1147_n 0.00123931f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_621 N_B_M1025_g N_A_512_347#_c_1145_n 8.71698e-19 $X=2.955 $Y=2.235 $X2=0
+ $Y2=0
cc_622 N_B_c_880_n N_A_512_347#_c_1145_n 0.00598819f $X=4.92 $Y=3.15 $X2=0 $Y2=0
cc_623 N_B_c_882_n N_A_1110_347#_c_1181_n 0.00572149f $X=6.8 $Y=3.15 $X2=0 $Y2=0
cc_624 N_B_M1009_g N_A_1110_347#_c_1185_n 0.0167942f $X=6.89 $Y=2.31 $X2=0 $Y2=0
cc_625 N_B_c_873_n N_A_1110_347#_c_1185_n 0.00852468f $X=7.305 $Y=1.485 $X2=0
+ $Y2=0
cc_626 N_B_c_872_n N_A_1110_347#_c_1182_n 0.00177951f $X=7.305 $Y=1.485 $X2=0
+ $Y2=0
cc_627 N_B_c_873_n N_A_1110_347#_c_1182_n 0.0273707f $X=7.305 $Y=1.485 $X2=0
+ $Y2=0
cc_628 N_B_M1009_g N_A_1110_347#_c_1183_n 0.00380344f $X=6.89 $Y=2.31 $X2=0
+ $Y2=0
cc_629 N_B_c_871_n N_VGND_c_1227_n 0.00171306f $X=5.01 $Y=1.09 $X2=0 $Y2=0
cc_630 N_B_M1015_g N_VGND_c_1228_n 0.00449178f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_631 N_B_M1015_g N_VGND_c_1229_n 0.00562997f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_632 N_B_M1000_g N_VGND_c_1231_n 0.00317047f $X=1.5 $Y=0.695 $X2=0 $Y2=0
cc_633 N_B_c_870_n N_VGND_c_1231_n 0.00313877f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_634 N_B_c_871_n N_VGND_c_1232_n 0.00432196f $X=5.01 $Y=1.09 $X2=0 $Y2=0
cc_635 N_B_M1015_g N_VGND_c_1233_n 0.0032155f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_636 N_B_M1000_g N_VGND_c_1235_n 0.00544287f $X=1.5 $Y=0.695 $X2=0 $Y2=0
cc_637 N_B_M1015_g N_VGND_c_1235_n 0.00544287f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_638 N_B_c_870_n N_VGND_c_1235_n 0.00544287f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_639 N_B_c_871_n N_VGND_c_1235_n 0.00544287f $X=5.01 $Y=1.09 $X2=0 $Y2=0
cc_640 N_B_c_870_n N_VGND_c_1236_n 0.00397421f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_641 N_B_c_870_n N_A_501_75#_c_1341_n 0.0088188f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_642 N_B_c_870_n N_A_501_75#_c_1338_n 0.00440744f $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_643 N_B_c_870_n N_A_501_75#_c_1346_n 8.04385e-19 $X=2.955 $Y=1.09 $X2=0 $Y2=0
cc_644 N_B_M1015_g N_A_1100_75#_c_1370_n 0.00140538f $X=7.21 $Y=0.695 $X2=0
+ $Y2=0
cc_645 N_B_M1015_g N_A_1100_75#_c_1380_n 0.0101012f $X=7.21 $Y=0.695 $X2=0 $Y2=0
cc_646 N_B_M1015_g N_A_1100_75#_c_1366_n 0.00493327f $X=7.21 $Y=0.695 $X2=0
+ $Y2=0
cc_647 N_SUM_c_1016_n N_VPWR_c_1035_n 0.0313231f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_648 N_SUM_c_1016_n N_VPWR_c_1042_n 0.0119584f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_649 N_SUM_c_1016_n N_VPWR_c_1034_n 0.00989813f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_650 SUM N_VGND_c_1230_n 0.0135716f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_651 SUM N_VGND_c_1235_n 0.0102675f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_652 N_VPWR_c_1036_n N_A_512_347#_c_1144_n 0.00129212f $X=3.245 $Y=2.795 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_1043_n N_A_512_347#_c_1144_n 0.00571266f $X=3.08 $Y=3.33 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_1034_n N_A_512_347#_c_1144_n 0.00688066f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_655 N_VPWR_M1025_d N_A_512_347#_c_1147_n 0.00633286f $X=3.045 $Y=1.735 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_1036_n N_A_512_347#_c_1147_n 0.0236753f $X=3.245 $Y=2.795 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_1036_n N_A_512_347#_c_1145_n 0.00502132f $X=3.245 $Y=2.795 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_1037_n N_A_512_347#_c_1145_n 0.0172713f $X=4.27 $Y=2.47 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_1040_n N_A_512_347#_c_1145_n 0.00726814f $X=4.105 $Y=3.33 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_1034_n N_A_512_347#_c_1145_n 0.00888973f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_1038_n N_A_1110_347#_c_1181_n 0.0115183f $X=6.66 $Y=2.6 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_1044_n N_A_1110_347#_c_1181_n 0.00650801f $X=6.12 $Y=3.33 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_1034_n N_A_1110_347#_c_1181_n 0.00784572f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_664 N_VPWR_M1022_d N_A_1110_347#_c_1185_n 0.0205598f $X=6.145 $Y=1.735 $X2=0
+ $Y2=0
cc_665 N_VPWR_c_1038_n N_A_1110_347#_c_1185_n 0.0362096f $X=6.66 $Y=2.6 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_1039_n N_A_1110_347#_c_1182_n 0.0137241f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_1038_n N_A_1110_347#_c_1183_n 0.0143566f $X=6.66 $Y=2.6 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_1039_n N_A_1110_347#_c_1183_n 0.0249394f $X=7.92 $Y=1.985 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_1045_n N_A_1110_347#_c_1183_n 0.0087946f $X=7.755 $Y=3.33 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_1034_n N_A_1110_347#_c_1183_n 0.0106389f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_1039_n COUT 0.0395727f $X=7.92 $Y=1.985 $X2=0 $Y2=0
cc_672 N_VPWR_c_1046_n COUT 0.0112891f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_673 N_VPWR_c_1034_n COUT 0.00934413f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_674 COUT N_VGND_c_1229_n 0.0157813f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_675 COUT N_VGND_c_1234_n 0.0145639f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_676 COUT N_VGND_c_1235_n 0.0119984f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_677 COUT N_A_1100_75#_c_1366_n 0.0011882f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_678 N_VGND_M1014_d N_A_501_75#_c_1341_n 0.00734279f $X=3.015 $Y=0.375 $X2=0
+ $Y2=0
cc_679 N_VGND_c_1226_n N_A_501_75#_c_1341_n 0.0029521f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_680 N_VGND_c_1231_n N_A_501_75#_c_1341_n 0.00294479f $X=3.07 $Y=0 $X2=0 $Y2=0
cc_681 N_VGND_c_1235_n N_A_501_75#_c_1341_n 0.0111994f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_1236_n N_A_501_75#_c_1341_n 0.0243979f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_683 N_VGND_c_1231_n N_A_501_75#_c_1338_n 0.0114153f $X=3.07 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1235_n N_A_501_75#_c_1338_n 0.01383f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_685 N_VGND_c_1226_n N_A_501_75#_c_1346_n 0.00882747f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_686 N_VGND_c_1235_n N_A_501_75#_c_1346_n 0.0110304f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_687 N_VGND_c_1235_n N_A_1100_75#_M1024_d 0.00738975f $X=8.4 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_688 N_VGND_M1023_d N_A_1100_75#_c_1365_n 4.88898e-19 $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_689 N_VGND_c_1228_n N_A_1100_75#_c_1365_n 0.014412f $X=6.915 $Y=0.305 $X2=0
+ $Y2=0
cc_690 N_VGND_c_1232_n N_A_1100_75#_c_1365_n 0.0709494f $X=6.83 $Y=0 $X2=0 $Y2=0
cc_691 N_VGND_c_1235_n N_A_1100_75#_c_1365_n 0.0410407f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_692 N_VGND_M1023_d N_A_1100_75#_c_1370_n 0.00300659f $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_693 N_VGND_c_1228_n N_A_1100_75#_c_1370_n 0.00332933f $X=6.915 $Y=0.305 $X2=0
+ $Y2=0
cc_694 N_VGND_M1023_d N_A_1100_75#_c_1380_n 0.0116084f $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_695 N_VGND_c_1228_n N_A_1100_75#_c_1380_n 0.0188598f $X=6.915 $Y=0.305 $X2=0
+ $Y2=0
cc_696 N_VGND_c_1232_n N_A_1100_75#_c_1380_n 0.00291923f $X=6.83 $Y=0 $X2=0
+ $Y2=0
cc_697 N_VGND_c_1233_n N_A_1100_75#_c_1380_n 0.0025393f $X=7.78 $Y=0 $X2=0 $Y2=0
cc_698 N_VGND_c_1235_n N_A_1100_75#_c_1380_n 0.0105139f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_699 N_VGND_M1023_d N_A_1100_75#_c_1371_n 4.74072e-19 $X=6.56 $Y=0.375 $X2=0
+ $Y2=0
cc_700 N_VGND_c_1229_n N_A_1100_75#_c_1366_n 0.0218711f $X=7.945 $Y=0.605 $X2=0
+ $Y2=0
cc_701 N_VGND_c_1233_n N_A_1100_75#_c_1366_n 0.00810949f $X=7.78 $Y=0 $X2=0
+ $Y2=0
cc_702 N_VGND_c_1235_n N_A_1100_75#_c_1366_n 0.0106855f $X=8.4 $Y=0 $X2=0 $Y2=0

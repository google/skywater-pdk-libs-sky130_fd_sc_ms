* File: sky130_fd_sc_ms__nor2_2.spice
* Created: Fri Aug 28 17:46:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor2_2.pex.spice"
.subckt sky130_fd_sc_ms__nor2_2  VNB VPB B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74 AD=0.2627
+ AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_A_35_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1002_d N_B_M1003_g N_A_35_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_35_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1004_d N_A_M1005_g N_A_35_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__nor2_2.pxi.spice"
*
.ends
*
*

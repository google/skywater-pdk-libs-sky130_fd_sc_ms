* File: sky130_fd_sc_ms__or2_2.pex.spice
* Created: Fri Aug 28 18:06:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR2_2%B 3 5 7 8 15
c26 8 0 1.41453e-19 $X=0.24 $Y=1.295
c27 5 0 1.44963e-19 $X=0.49 $Y=1.22
r28 14 15 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.49 $Y=1.385
+ $X2=0.495 $Y2=1.385
r29 11 14 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.27 $Y=1.385
+ $X2=0.49 $Y2=1.385
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r31 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r32 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.22
+ $X2=0.49 $Y2=1.385
r33 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.49 $Y=1.22 $X2=0.49
+ $Y2=0.79
r34 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=1.385
r35 1 3 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_2%A 3 7 9 10 14 15
c45 14 0 1.41453e-19 $X=0.96 $Y=1.515
r46 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.96 $Y2=1.68
r47 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.96 $Y2=1.35
r48 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.515 $X2=0.96 $Y2=1.515
r49 9 10 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.825 $Y=1.665
+ $X2=0.825 $Y2=2.035
r50 9 15 3.92878 $w=4.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.825 $Y=1.665
+ $X2=0.825 $Y2=1.515
r51 7 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.92 $Y=0.79 $X2=0.92
+ $Y2=1.35
r52 3 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.885 $Y=2.34
+ $X2=0.885 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_2%A_27_368# 1 2 9 13 17 21 25 29 31 35 37 38 40
+ 41 44 45 46 48 49
c100 35 0 1.44963e-19 $X=0.705 $Y=0.615
r101 54 55 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.855 $Y=1.465
+ $X2=1.895 $Y2=1.465
r102 52 54 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.425 $Y=1.465
+ $X2=1.855 $Y2=1.465
r103 49 55 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.13 $Y=1.465
+ $X2=1.895 $Y2=1.465
r104 48 51 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=1.465
+ $X2=2.13 $Y2=1.63
r105 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.465 $X2=2.13 $Y2=1.465
r106 44 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.21 $Y=2.32
+ $X2=2.21 $Y2=1.63
r107 42 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=2.405
+ $X2=1.3 $Y2=2.405
r108 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.125 $Y=2.405
+ $X2=2.21 $Y2=2.32
r109 41 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.125 $Y=2.405
+ $X2=1.385 $Y2=2.405
r110 40 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.32 $X2=1.3
+ $Y2=2.405
r111 39 40 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.3 $Y=1.18
+ $X2=1.3 $Y2=2.32
r112 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.215 $Y=1.095
+ $X2=1.3 $Y2=1.18
r113 37 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.215 $Y=1.095
+ $X2=0.87 $Y2=1.095
r114 33 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.745 $Y=1.01
+ $X2=0.87 $Y2=1.095
r115 33 35 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=0.745 $Y=1.01
+ $X2=0.745 $Y2=0.615
r116 32 45 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.405
+ $X2=0.27 $Y2=2.405
r117 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=1.3 $Y2=2.405
r118 31 32 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=0.435 $Y2=2.405
r119 27 45 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.49
+ $X2=0.27 $Y2=2.405
r120 27 29 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=2.49
+ $X2=0.27 $Y2=2.695
r121 23 45 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.32
+ $X2=0.27 $Y2=2.405
r122 23 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.27 $Y=2.32
+ $X2=0.27 $Y2=1.985
r123 19 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.63
+ $X2=1.895 $Y2=1.465
r124 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.895 $Y=1.63
+ $X2=1.895 $Y2=2.4
r125 15 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.3
+ $X2=1.855 $Y2=1.465
r126 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.855 $Y=1.3
+ $X2=1.855 $Y2=0.74
r127 11 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=1.465
r128 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=0.74
r129 7 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.63
+ $X2=1.425 $Y2=1.465
r130 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.425 $Y=1.63
+ $X2=1.425 $Y2=2.4
r131 2 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.695
r132 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
r133 1 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.47 $X2=0.705 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_2%VPWR 1 2 9 11 13 15 17 22 28 32
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 22 31 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.177 $Y2=3.33
r42 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 15 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 11 31 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.177 $Y2=3.33
r50 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.78
r51 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=3.33
r52 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=2.78
r53 2 13 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=2.78
r54 1 9 600 $w=1.7e-07 $l=1.04647e-06 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.84 $X2=1.2 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_2%X 1 2 7 8 9 10 11
r20 11 30 7.05875 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.985
+ $X2=1.695 $Y2=1.82
r21 10 30 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.675 $Y=1.665
+ $X2=1.675 $Y2=1.82
r22 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.675 $Y=1.295
+ $X2=1.675 $Y2=1.665
r23 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.675 $Y=0.925
+ $X2=1.675 $Y2=1.295
r24 7 8 19.6876 $w=2.38e-07 $l=4.1e-07 $layer=LI1_cond $X=1.675 $Y=0.515
+ $X2=1.675 $Y2=0.925
r25 2 11 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.84 $X2=1.66 $Y2=1.985
r26 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5 $Y=0.37
+ $X2=1.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_2%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r37 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r40 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r42 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r43 29 41 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=2.185
+ $Y2=0
r44 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=1.68
+ $Y2=0
r45 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 25 35 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r48 25 27 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r49 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r50 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r51 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r52 22 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r53 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 18 41 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.185 $Y2=0
r55 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.135 $Y2=0.515
r56 14 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r57 14 16 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.65
r58 10 35 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r59 10 12 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.835
r60 3 20 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.37 $X2=2.135 $Y2=0.515
r61 2 16 182 $w=1.7e-07 $l=2.91419e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.47 $X2=1.21 $Y2=0.65
r62 1 12 182 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.47 $X2=0.275 $Y2=0.835
.ends


* File: sky130_fd_sc_ms__o311ai_1.spice
* Created: Wed Sep  2 12:25:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o311ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o311ai_1  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_A_128_74#_M1003_d N_A1_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.2627 PD=1.045 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_128_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.222 AS=0.11285 PD=1.34 PS=1.045 NRD=27.564 NRS=4.044 M=1 R=4.93333
+ SA=75000.7 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_128_74#_M1009_d N_A3_M1009_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.222 PD=1.09 PS=1.34 NRD=11.34 NRS=24.324 M=1 R=4.93333
+ SA=75001.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1006 A_469_74# N_B1_M1006_g N_A_128_74#_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=16.212 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_C1_M1001_g A_469_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1147 PD=2.05 PS=1.05 NRD=0 NRS=16.212 M=1 R=4.93333 SA=75002.4 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1002 A_141_368# N_A1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90002.3
+ A=0.2016 P=2.6 MULT=1
MM1004 A_225_368# N_A2_M1004_g A_141_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1007_d N_A3_M1007_g A_225_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=20.2122 NRS=24.6053 M=1 R=6.22222 SA=90001.2
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g N_Y_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2184 AS=0.2184 PD=1.51 PS=1.51 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.8
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90002.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__o311ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor4_4.pxi.spice
* Created: Wed Sep  2 12:16:50 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4_4%D N_D_M1001_g N_D_M1002_g N_D_M1003_g N_D_M1004_g
+ N_D_M1022_g N_D_M1006_g D D D N_D_c_111_n N_D_c_106_n
+ PM_SKY130_FD_SC_MS__NOR4_4%D
x_PM_SKY130_FD_SC_MS__NOR4_4%C N_C_M1014_g N_C_M1007_g N_C_M1012_g N_C_M1015_g
+ N_C_M1023_g N_C_M1017_g C C C N_C_c_168_n N_C_c_169_n
+ PM_SKY130_FD_SC_MS__NOR4_4%C
x_PM_SKY130_FD_SC_MS__NOR4_4%B N_B_M1009_g N_B_M1020_g N_B_M1000_g N_B_M1005_g
+ N_B_M1010_g N_B_M1013_g B B B B B B N_B_c_238_n PM_SKY130_FD_SC_MS__NOR4_4%B
x_PM_SKY130_FD_SC_MS__NOR4_4%A N_A_M1008_g N_A_c_311_n N_A_c_312_n N_A_M1016_g
+ N_A_M1011_g N_A_M1018_g N_A_M1021_g N_A_M1019_g A A N_A_c_319_n N_A_c_320_n
+ N_A_c_321_n PM_SKY130_FD_SC_MS__NOR4_4%A
x_PM_SKY130_FD_SC_MS__NOR4_4%A_27_368# N_A_27_368#_M1002_s N_A_27_368#_M1003_s
+ N_A_27_368#_M1006_s N_A_27_368#_M1012_s N_A_27_368#_M1017_s
+ N_A_27_368#_c_386_n N_A_27_368#_c_387_n N_A_27_368#_c_388_n
+ N_A_27_368#_c_395_n N_A_27_368#_c_389_n N_A_27_368#_c_390_n
+ N_A_27_368#_c_403_n N_A_27_368#_c_430_p N_A_27_368#_c_407_n
+ N_A_27_368#_c_391_n N_A_27_368#_c_411_n N_A_27_368#_c_392_n
+ PM_SKY130_FD_SC_MS__NOR4_4%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR4_4%Y N_Y_M1001_s N_Y_M1014_s N_Y_M1009_d N_Y_M1016_d
+ N_Y_M1002_d N_Y_M1004_d N_Y_c_445_n N_Y_c_458_n N_Y_c_456_n N_Y_c_460_n
+ N_Y_c_446_n N_Y_c_447_n N_Y_c_448_n N_Y_c_449_n N_Y_c_450_n N_Y_c_469_n
+ N_Y_c_474_n N_Y_c_451_n N_Y_c_452_n N_Y_c_453_n N_Y_c_454_n Y
+ PM_SKY130_FD_SC_MS__NOR4_4%Y
x_PM_SKY130_FD_SC_MS__NOR4_4%A_499_368# N_A_499_368#_M1007_d
+ N_A_499_368#_M1015_d N_A_499_368#_M1000_d N_A_499_368#_M1010_d
+ N_A_499_368#_c_553_n N_A_499_368#_c_547_n N_A_499_368#_c_548_n
+ N_A_499_368#_c_560_n N_A_499_368#_c_549_n N_A_499_368#_c_567_n
+ N_A_499_368#_c_550_n N_A_499_368#_c_573_n N_A_499_368#_c_551_n
+ N_A_499_368#_c_552_n PM_SKY130_FD_SC_MS__NOR4_4%A_499_368#
x_PM_SKY130_FD_SC_MS__NOR4_4%A_879_368# N_A_879_368#_M1000_s
+ N_A_879_368#_M1005_s N_A_879_368#_M1013_s N_A_879_368#_M1011_d
+ N_A_879_368#_M1019_d N_A_879_368#_c_610_n N_A_879_368#_c_611_n
+ N_A_879_368#_c_618_n N_A_879_368#_c_662_n N_A_879_368#_c_622_n
+ N_A_879_368#_c_612_n N_A_879_368#_c_627_n N_A_879_368#_c_613_n
+ N_A_879_368#_c_641_n N_A_879_368#_c_614_n N_A_879_368#_c_615_n
+ N_A_879_368#_c_628_n N_A_879_368#_c_630_n N_A_879_368#_c_651_n
+ PM_SKY130_FD_SC_MS__NOR4_4%A_879_368#
x_PM_SKY130_FD_SC_MS__NOR4_4%VPWR N_VPWR_M1008_s N_VPWR_M1018_s N_VPWR_c_681_n
+ N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_684_n VPWR N_VPWR_c_685_n
+ N_VPWR_c_686_n N_VPWR_c_680_n N_VPWR_c_688_n PM_SKY130_FD_SC_MS__NOR4_4%VPWR
x_PM_SKY130_FD_SC_MS__NOR4_4%VGND N_VGND_M1001_d N_VGND_M1022_d N_VGND_M1023_d
+ N_VGND_M1020_s N_VGND_M1021_s N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n N_VGND_c_766_n N_VGND_c_767_n
+ N_VGND_c_768_n N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n VGND
+ N_VGND_c_772_n N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n
+ PM_SKY130_FD_SC_MS__NOR4_4%VGND
cc_1 VNB N_D_M1001_g 0.0350087f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_2 VNB N_D_M1022_g 0.033152f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_3 VNB N_D_c_106_n 0.0928911f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.515
cc_4 VNB N_C_M1014_g 0.0340976f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_5 VNB N_C_M1023_g 0.033152f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_6 VNB N_C_c_168_n 0.0012292f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_7 VNB N_C_c_169_n 0.0900674f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.515
cc_8 VNB N_B_M1009_g 0.0244877f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_9 VNB N_B_M1020_g 0.0306733f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_10 VNB B 0.00861277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_238_n 0.121974f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.565
cc_12 VNB N_A_M1008_g 0.00153751f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_13 VNB N_A_c_311_n 0.0206365f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.68
cc_14 VNB N_A_c_312_n 0.0100258f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_15 VNB N_A_M1016_g 0.0318428f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.68
cc_16 VNB N_A_M1011_g 0.00165349f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.68
cc_17 VNB N_A_M1018_g 0.00165685f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.35
cc_18 VNB N_A_M1021_g 0.0293697f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.68
cc_19 VNB N_A_M1019_g 0.00255353f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB A 0.0325254f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_21 VNB N_A_c_319_n 0.0793709f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_22 VNB N_A_c_320_n 0.00425479f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_23 VNB N_A_c_321_n 0.00386031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_445_n 0.00746863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_446_n 0.00675823f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_26 VNB N_Y_c_447_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_27 VNB N_Y_c_448_n 0.0203308f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.515
cc_28 VNB N_Y_c_449_n 0.00374454f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_29 VNB N_Y_c_450_n 0.0197472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_451_n 0.00683417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_452_n 0.0201517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_453_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_454_n 0.00874911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB Y 0.0240186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_680_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_36 VNB N_VGND_c_760_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_761_n 0.0316455f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.74
cc_38 VNB N_VGND_c_762_n 0.00641221f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_39 VNB N_VGND_c_763_n 0.00571437f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_40 VNB N_VGND_c_764_n 0.02962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_765_n 0.028454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_766_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.515
cc_43 VNB N_VGND_c_767_n 0.0389478f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_44 VNB N_VGND_c_768_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.515
cc_45 VNB N_VGND_c_769_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.515
cc_46 VNB N_VGND_c_770_n 0.0252293f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_47 VNB N_VGND_c_771_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_48 VNB N_VGND_c_772_n 0.0376264f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.68
cc_49 VNB N_VGND_c_773_n 0.455329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_774_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_775_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_776_n 0.0126522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_D_M1002_g 0.02307f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_54 VPB N_D_M1003_g 0.0196371f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_55 VPB N_D_M1004_g 0.0202147f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_56 VPB N_D_M1006_g 0.0209373f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_57 VPB N_D_c_111_n 0.00801745f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_58 VPB N_D_c_106_n 0.013373f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.515
cc_59 VPB N_C_M1007_g 0.021023f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_60 VPB N_C_M1012_g 0.0196336f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_61 VPB N_C_M1015_g 0.0196343f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_62 VPB N_C_M1017_g 0.024655f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_63 VPB N_C_c_168_n 0.00755714f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_64 VPB N_C_c_169_n 0.0126363f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.515
cc_65 VPB N_B_M1000_g 0.0252911f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_66 VPB N_B_M1005_g 0.019875f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_67 VPB N_B_M1010_g 0.019875f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_68 VPB N_B_M1013_g 0.0204787f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_69 VPB B 0.0243141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_B_c_238_n 0.0286748f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.565
cc_71 VPB N_A_M1008_g 0.0234328f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=0.74
cc_72 VPB N_A_M1011_g 0.0236033f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.68
cc_73 VPB N_A_M1018_g 0.0236156f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.35
cc_74 VPB N_A_M1019_g 0.0324186f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_75 VPB N_A_27_368#_c_386_n 0.0237653f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_76 VPB N_A_27_368#_c_387_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_368#_c_388_n 0.0100897f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.68
cc_78 VPB N_A_27_368#_c_389_n 0.00474241f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_79 VPB N_A_27_368#_c_390_n 0.00325473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_27_368#_c_391_n 0.00160153f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.68
cc_81 VPB N_A_27_368#_c_392_n 0.00721501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_Y_c_456_n 0.00707089f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_83 VPB Y 0.012933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_499_368#_c_547_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.35
cc_85 VPB N_A_499_368#_c_548_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_86 VPB N_A_499_368#_c_549_n 0.0167491f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_87 VPB N_A_499_368#_c_550_n 0.00403034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_499_368#_c_551_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_89 VPB N_A_499_368#_c_552_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_90 VPB N_A_879_368#_c_610_n 0.00163297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_879_368#_c_611_n 0.00555274f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=0.74
cc_92 VPB N_A_879_368#_c_612_n 0.00220508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_879_368#_c_613_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_94 VPB N_A_879_368#_c_614_n 0.0153056f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_95 VPB N_A_879_368#_c_615_n 0.0352562f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.68
cc_96 VPB N_VPWR_c_681_n 0.00895394f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.68
cc_97 VPB N_VPWR_c_682_n 0.00899828f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.68
cc_98 VPB N_VPWR_c_683_n 0.157251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_684_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.35
cc_100 VPB N_VPWR_c_685_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_101 VPB N_VPWR_c_686_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_102 VPB N_VPWR_c_680_n 0.0872008f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_103 VPB N_VPWR_c_688_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.515
cc_104 N_D_M1022_g N_C_M1014_g 0.0181303f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_105 N_D_M1006_g N_C_M1007_g 0.0148426f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_106 N_D_c_111_n N_C_M1007_g 2.7317e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_107 N_D_c_111_n N_C_c_168_n 0.0134722f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_D_c_106_n N_C_c_168_n 0.00153052f $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_109 N_D_c_111_n N_C_c_169_n 0.00133235f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_110 N_D_c_106_n N_C_c_169_n 0.0274741f $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_111 N_D_M1002_g N_A_27_368#_c_387_n 0.0150267f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_112 N_D_M1003_g N_A_27_368#_c_387_n 0.0140221f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_113 N_D_M1004_g N_A_27_368#_c_395_n 0.00867919f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_114 N_D_M1006_g N_A_27_368#_c_395_n 8.62308e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_115 N_D_M1004_g N_A_27_368#_c_389_n 0.0119307f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_116 N_D_M1006_g N_A_27_368#_c_389_n 0.0139978f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_117 N_D_M1006_g N_A_27_368#_c_390_n 4.63009e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_118 N_D_M1004_g N_A_27_368#_c_391_n 0.00194226f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_119 N_D_M1002_g N_Y_c_458_n 0.0162996f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_120 N_D_c_111_n N_Y_c_458_n 0.0065328f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_121 N_D_M1003_g N_Y_c_460_n 0.012931f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_122 N_D_M1004_g N_Y_c_460_n 0.0142562f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_123 N_D_c_111_n N_Y_c_460_n 0.0422425f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_124 N_D_c_106_n N_Y_c_460_n 4.90767e-19 $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_125 N_D_M1001_g N_Y_c_449_n 0.0162996f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_126 N_D_c_111_n N_Y_c_449_n 0.113145f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_127 N_D_M1001_g N_Y_c_450_n 0.00423262f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_128 N_D_M1022_g N_Y_c_450_n 0.00160267f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_129 N_D_c_106_n N_Y_c_450_n 0.0260064f $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_130 N_D_M1002_g N_Y_c_469_n 0.0147264f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_131 N_D_M1003_g N_Y_c_469_n 0.0106907f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_132 N_D_M1004_g N_Y_c_469_n 4.41999e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_133 N_D_c_111_n N_Y_c_469_n 0.0235495f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_134 N_D_c_106_n N_Y_c_469_n 5.54777e-19 $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_135 N_D_M1006_g N_Y_c_474_n 0.011604f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_136 N_D_c_111_n N_Y_c_474_n 0.023072f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_137 N_D_c_106_n N_Y_c_474_n 8.57329e-19 $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_138 N_D_M1022_g N_Y_c_451_n 0.0159102f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_139 N_D_c_106_n N_Y_c_451_n 0.00377017f $X=1.86 $Y=1.515 $X2=0 $Y2=0
cc_140 N_D_M1022_g N_Y_c_452_n 6.34175e-19 $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_141 N_D_M1001_g Y 0.024494f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_142 N_D_c_111_n Y 0.0349192f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_143 N_D_M1002_g N_VPWR_c_683_n 0.00333926f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_144 N_D_M1003_g N_VPWR_c_683_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_145 N_D_M1004_g N_VPWR_c_683_n 0.00333896f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_146 N_D_M1006_g N_VPWR_c_683_n 0.00333926f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_147 N_D_M1002_g N_VPWR_c_680_n 0.00426591f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_148 N_D_M1003_g N_VPWR_c_680_n 0.00422687f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_149 N_D_M1004_g N_VPWR_c_680_n 0.00423173f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_150 N_D_M1006_g N_VPWR_c_680_n 0.00423286f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_151 N_D_M1001_g N_VGND_c_761_n 0.00744799f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_152 N_D_M1022_g N_VGND_c_762_n 0.0136269f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_153 N_D_M1001_g N_VGND_c_772_n 0.00461464f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_154 N_D_M1022_g N_VGND_c_772_n 0.00383152f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_155 N_D_M1001_g N_VGND_c_773_n 0.00916349f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_156 N_D_M1022_g N_VGND_c_773_n 0.00762539f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_157 N_C_M1023_g N_B_M1009_g 0.0176979f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_158 N_C_c_168_n B 0.0364929f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_159 N_C_c_169_n B 0.00428128f $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_160 N_C_c_168_n N_B_c_238_n 3.01993e-19 $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_161 N_C_c_169_n N_B_c_238_n 0.0241886f $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_162 N_C_M1007_g N_A_27_368#_c_389_n 0.00100838f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_163 N_C_M1007_g N_A_27_368#_c_390_n 4.63009e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_164 N_C_M1007_g N_A_27_368#_c_403_n 0.0178906f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_165 N_C_M1012_g N_A_27_368#_c_403_n 0.0142175f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_166 N_C_c_168_n N_A_27_368#_c_403_n 0.0359263f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_167 N_C_c_169_n N_A_27_368#_c_403_n 4.90767e-19 $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_168 N_C_M1015_g N_A_27_368#_c_407_n 0.0142562f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_169 N_C_M1017_g N_A_27_368#_c_407_n 0.0158758f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_170 N_C_c_168_n N_A_27_368#_c_407_n 0.0403041f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_171 N_C_c_169_n N_A_27_368#_c_407_n 4.88651e-19 $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_172 N_C_c_168_n N_A_27_368#_c_411_n 0.016575f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_173 N_C_c_169_n N_A_27_368#_c_411_n 5.54777e-19 $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_174 N_C_M1023_g N_Y_c_446_n 0.0142504f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_175 N_C_c_169_n N_Y_c_446_n 0.00205646f $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_176 N_C_M1023_g N_Y_c_447_n 4.81487e-19 $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_177 N_C_M1014_g N_Y_c_451_n 0.0134054f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_178 N_C_M1014_g N_Y_c_452_n 0.0138796f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_179 N_C_M1023_g N_Y_c_452_n 0.00160267f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_180 N_C_c_168_n N_Y_c_452_n 0.113128f $X=3.62 $Y=1.515 $X2=0 $Y2=0
cc_181 N_C_c_169_n N_Y_c_452_n 0.0268231f $X=3.71 $Y=1.515 $X2=0 $Y2=0
cc_182 N_C_M1007_g N_A_499_368#_c_553_n 0.00828022f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_183 N_C_M1012_g N_A_499_368#_c_553_n 0.009254f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_184 N_C_M1015_g N_A_499_368#_c_553_n 5.56591e-19 $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_185 N_C_M1012_g N_A_499_368#_c_547_n 0.0116345f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_186 N_C_M1015_g N_A_499_368#_c_547_n 0.0116345f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_187 N_C_M1007_g N_A_499_368#_c_548_n 0.00348237f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_188 N_C_M1012_g N_A_499_368#_c_548_n 0.00194226f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_189 N_C_M1012_g N_A_499_368#_c_560_n 5.56591e-19 $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_190 N_C_M1015_g N_A_499_368#_c_560_n 0.009254f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_191 N_C_M1017_g N_A_499_368#_c_560_n 0.0140199f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_192 N_C_M1017_g N_A_499_368#_c_549_n 0.0137576f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_193 N_C_M1015_g N_A_499_368#_c_551_n 0.00194226f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_194 N_C_M1017_g N_A_499_368#_c_551_n 0.00194226f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_195 N_C_M1007_g N_VPWR_c_683_n 0.00517089f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_196 N_C_M1012_g N_VPWR_c_683_n 0.00333896f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_197 N_C_M1015_g N_VPWR_c_683_n 0.00333896f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_198 N_C_M1017_g N_VPWR_c_683_n 0.00333896f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_199 N_C_M1007_g N_VPWR_c_680_n 0.00978686f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_200 N_C_M1012_g N_VPWR_c_680_n 0.00422685f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_201 N_C_M1015_g N_VPWR_c_680_n 0.00422685f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_202 N_C_M1017_g N_VPWR_c_680_n 0.00427818f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_203 N_C_M1014_g N_VGND_c_762_n 0.00572988f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_204 N_C_M1023_g N_VGND_c_763_n 0.0136269f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_205 N_C_M1014_g N_VGND_c_767_n 0.00433162f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_206 N_C_M1023_g N_VGND_c_767_n 0.00383152f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_207 N_C_M1014_g N_VGND_c_773_n 0.00822119f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_208 N_C_M1023_g N_VGND_c_773_n 0.00762539f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B_M1013_g N_A_M1008_g 0.0120753f $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_210 B N_A_M1008_g 0.00715549f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_211 B N_A_c_312_n 0.00854105f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_212 N_B_c_238_n N_A_c_312_n 0.0120753f $X=6.135 $Y=1.515 $X2=0 $Y2=0
cc_213 B N_A_M1011_g 7.59625e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_214 B N_A_c_319_n 8.80022e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_215 B N_A_c_321_n 0.0112317f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_216 B N_A_27_368#_c_392_n 0.0159469f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_217 N_B_M1009_g N_Y_c_446_n 0.0114826f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_218 B N_Y_c_446_n 0.022854f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B_M1009_g N_Y_c_447_n 0.00856181f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B_M1020_g N_Y_c_447_n 0.0132207f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B_M1020_g N_Y_c_448_n 0.0134377f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_222 B N_Y_c_448_n 0.127864f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_223 N_B_c_238_n N_Y_c_448_n 0.0373023f $X=6.135 $Y=1.515 $X2=0 $Y2=0
cc_224 N_B_M1009_g N_Y_c_453_n 0.00257802f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B_M1020_g N_Y_c_453_n 0.00393109f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_226 B N_Y_c_453_n 0.0281223f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B_c_238_n N_Y_c_453_n 0.00232957f $X=6.135 $Y=1.515 $X2=0 $Y2=0
cc_228 N_B_M1000_g N_A_499_368#_c_549_n 0.0137576f $X=4.765 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B_M1000_g N_A_499_368#_c_567_n 0.0137902f $X=4.765 $Y=2.4 $X2=0 $Y2=0
cc_230 N_B_M1005_g N_A_499_368#_c_567_n 0.00922424f $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_231 N_B_M1010_g N_A_499_368#_c_567_n 5.5995e-19 $X=5.685 $Y=2.4 $X2=0 $Y2=0
cc_232 N_B_M1005_g N_A_499_368#_c_550_n 0.0117578f $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_233 N_B_M1010_g N_A_499_368#_c_550_n 0.0137f $X=5.685 $Y=2.4 $X2=0 $Y2=0
cc_234 N_B_M1013_g N_A_499_368#_c_550_n 0.00423362f $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_235 N_B_M1005_g N_A_499_368#_c_573_n 5.5995e-19 $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_236 N_B_M1010_g N_A_499_368#_c_573_n 0.00922424f $X=5.685 $Y=2.4 $X2=0 $Y2=0
cc_237 N_B_M1013_g N_A_499_368#_c_573_n 0.00777833f $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B_M1000_g N_A_499_368#_c_552_n 0.00194226f $X=4.765 $Y=2.4 $X2=0 $Y2=0
cc_239 N_B_M1005_g N_A_499_368#_c_552_n 0.00194226f $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_240 B N_A_879_368#_c_610_n 0.0218203f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B_c_238_n N_A_879_368#_c_610_n 0.00151288f $X=6.135 $Y=1.515 $X2=0
+ $Y2=0
cc_242 N_B_M1000_g N_A_879_368#_c_618_n 0.0142681f $X=4.765 $Y=2.4 $X2=0 $Y2=0
cc_243 N_B_M1005_g N_A_879_368#_c_618_n 0.0142681f $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_244 B N_A_879_368#_c_618_n 0.0472481f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_245 N_B_c_238_n N_A_879_368#_c_618_n 4.90767e-19 $X=6.135 $Y=1.515 $X2=0
+ $Y2=0
cc_246 N_B_M1010_g N_A_879_368#_c_622_n 0.0142681f $X=5.685 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B_M1013_g N_A_879_368#_c_622_n 0.0142681f $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_248 B N_A_879_368#_c_622_n 0.0463814f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_249 N_B_c_238_n N_A_879_368#_c_622_n 4.90767e-19 $X=6.135 $Y=1.515 $X2=0
+ $Y2=0
cc_250 N_B_M1013_g N_A_879_368#_c_612_n 2.4399e-19 $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_251 B N_A_879_368#_c_627_n 0.00507353f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_252 B N_A_879_368#_c_628_n 0.0174726f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_253 N_B_c_238_n N_A_879_368#_c_628_n 6.78061e-19 $X=6.135 $Y=1.515 $X2=0
+ $Y2=0
cc_254 B N_A_879_368#_c_630_n 0.0198447f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_255 N_B_M1000_g N_VPWR_c_683_n 0.00333896f $X=4.765 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B_M1005_g N_VPWR_c_683_n 0.00333896f $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B_M1010_g N_VPWR_c_683_n 0.00333896f $X=5.685 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B_M1013_g N_VPWR_c_683_n 0.00517089f $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_259 N_B_M1000_g N_VPWR_c_680_n 0.00427818f $X=4.765 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B_M1005_g N_VPWR_c_680_n 0.00422886f $X=5.215 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B_M1010_g N_VPWR_c_680_n 0.00422886f $X=5.685 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B_M1013_g N_VPWR_c_680_n 0.00978686f $X=6.135 $Y=2.4 $X2=0 $Y2=0
cc_263 N_B_M1009_g N_VGND_c_763_n 0.00432719f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_264 N_B_M1020_g N_VGND_c_765_n 0.00510848f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_265 N_B_M1009_g N_VGND_c_773_n 0.00820772f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B_M1020_g N_VGND_c_773_n 0.00825037f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B_M1009_g N_VGND_c_775_n 0.00434272f $X=4.21 $Y=0.74 $X2=0 $Y2=0
cc_268 N_B_M1020_g N_VGND_c_775_n 0.00434272f $X=4.64 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_c_312_n N_Y_c_448_n 0.0147383f $X=6.675 $Y=1.555 $X2=0 $Y2=0
cc_270 N_A_M1016_g N_Y_c_448_n 0.0146105f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_c_321_n N_Y_c_448_n 0.014057f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_272 N_A_M1016_g N_Y_c_454_n 9.31832e-19 $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_M1021_g N_Y_c_454_n 0.00330748f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_c_319_n N_Y_c_454_n 0.0132405f $X=7.98 $Y=1.465 $X2=0 $Y2=0
cc_275 N_A_c_320_n N_Y_c_454_n 0.00433553f $X=8.03 $Y=1.405 $X2=0 $Y2=0
cc_276 N_A_c_321_n N_Y_c_454_n 0.0406673f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_277 N_A_M1008_g N_A_499_368#_c_550_n 3.1137e-19 $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A_M1008_g N_A_879_368#_c_612_n 0.012057f $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A_M1011_g N_A_879_368#_c_612_n 4.10971e-19 $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_280 N_A_M1008_g N_A_879_368#_c_627_n 0.0157145f $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A_c_311_n N_A_879_368#_c_627_n 0.0055433f $X=7.045 $Y=1.555 $X2=0 $Y2=0
cc_282 N_A_M1011_g N_A_879_368#_c_627_n 0.014323f $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A_c_321_n N_A_879_368#_c_627_n 0.00643572f $X=7.805 $Y=1.405 $X2=0
+ $Y2=0
cc_284 N_A_M1008_g N_A_879_368#_c_613_n 4.09618e-19 $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_285 N_A_M1011_g N_A_879_368#_c_613_n 0.0121532f $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A_M1018_g N_A_879_368#_c_613_n 0.0121532f $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A_M1019_g N_A_879_368#_c_613_n 4.09618e-19 $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_288 N_A_M1018_g N_A_879_368#_c_641_n 0.014323f $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A_M1019_g N_A_879_368#_c_641_n 0.014323f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A_c_319_n N_A_879_368#_c_641_n 0.00430135f $X=7.98 $Y=1.465 $X2=0 $Y2=0
cc_291 N_A_c_321_n N_A_879_368#_c_641_n 0.027461f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_292 N_A_M1018_g N_A_879_368#_c_614_n 5.96661e-19 $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A_M1019_g N_A_879_368#_c_614_n 0.00399698f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_294 A N_A_879_368#_c_614_n 0.0264899f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_295 N_A_M1018_g N_A_879_368#_c_615_n 4.09618e-19 $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A_M1019_g N_A_879_368#_c_615_n 0.0130924f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A_M1008_g N_A_879_368#_c_630_n 8.84614e-19 $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A_M1011_g N_A_879_368#_c_651_n 0.00105868f $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A_M1018_g N_A_879_368#_c_651_n 0.00105868f $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A_c_319_n N_A_879_368#_c_651_n 0.00191987f $X=7.98 $Y=1.465 $X2=0 $Y2=0
cc_301 N_A_c_321_n N_A_879_368#_c_651_n 0.01334f $X=7.805 $Y=1.405 $X2=0 $Y2=0
cc_302 N_A_M1008_g N_VPWR_c_681_n 0.00246131f $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A_M1011_g N_VPWR_c_681_n 0.00233982f $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A_M1018_g N_VPWR_c_682_n 0.00233982f $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A_M1019_g N_VPWR_c_682_n 0.003737f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A_M1008_g N_VPWR_c_683_n 0.005209f $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_307 N_A_M1011_g N_VPWR_c_685_n 0.005209f $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_308 N_A_M1018_g N_VPWR_c_685_n 0.005209f $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_309 N_A_M1019_g N_VPWR_c_686_n 0.005209f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_310 N_A_M1008_g N_VPWR_c_680_n 0.00982636f $X=6.585 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A_M1011_g N_VPWR_c_680_n 0.00982526f $X=7.135 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A_M1018_g N_VPWR_c_680_n 0.00982526f $X=7.585 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A_M1019_g N_VPWR_c_680_n 0.00986267f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_314 N_A_M1021_g N_VGND_c_766_n 0.0151922f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_315 A N_VGND_c_766_n 0.026357f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_316 N_A_c_319_n N_VGND_c_766_n 5.98537e-19 $X=7.98 $Y=1.465 $X2=0 $Y2=0
cc_317 N_A_M1016_g N_VGND_c_770_n 0.00383152f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_M1021_g N_VGND_c_770_n 0.00383152f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_M1016_g N_VGND_c_773_n 0.00755866f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_M1021_g N_VGND_c_773_n 0.00760481f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_M1016_g N_VGND_c_776_n 0.0148268f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_27_368#_c_387_n N_Y_M1002_d 0.00165831f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_323 N_A_27_368#_c_389_n N_Y_M1004_d 0.00218982f $X=2.095 $Y=2.99 $X2=0 $Y2=0
cc_324 N_A_27_368#_M1002_s N_Y_c_458_n 0.00253686f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_325 N_A_27_368#_c_386_n N_Y_c_458_n 0.00427553f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_326 N_A_27_368#_M1002_s N_Y_c_456_n 0.00383494f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_327 N_A_27_368#_c_386_n N_Y_c_456_n 0.0206806f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_328 N_A_27_368#_M1003_s N_Y_c_460_n 0.00314376f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_329 N_A_27_368#_c_395_n N_Y_c_460_n 0.0148589f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_330 N_A_27_368#_c_387_n N_Y_c_469_n 0.0159318f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_331 N_A_27_368#_c_389_n N_Y_c_474_n 0.0177084f $X=2.095 $Y=2.99 $X2=0 $Y2=0
cc_332 N_A_27_368#_c_390_n N_Y_c_451_n 0.00568183f $X=2.18 $Y=2.12 $X2=0 $Y2=0
cc_333 N_A_27_368#_M1002_s Y 0.00217208f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_334 N_A_27_368#_c_403_n N_A_499_368#_M1007_d 0.00314376f $X=2.97 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_335 N_A_27_368#_c_407_n N_A_499_368#_M1015_d 0.00314376f $X=3.895 $Y=2.035
+ $X2=0 $Y2=0
cc_336 N_A_27_368#_c_403_n N_A_499_368#_c_553_n 0.0170259f $X=2.97 $Y=2.035
+ $X2=0 $Y2=0
cc_337 N_A_27_368#_M1012_s N_A_499_368#_c_547_n 0.00165831f $X=2.945 $Y=1.84
+ $X2=0 $Y2=0
cc_338 N_A_27_368#_c_430_p N_A_499_368#_c_547_n 0.0118736f $X=3.08 $Y=2.57 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_c_389_n N_A_499_368#_c_548_n 0.0110621f $X=2.095 $Y=2.99
+ $X2=0 $Y2=0
cc_340 N_A_27_368#_c_407_n N_A_499_368#_c_560_n 0.0170259f $X=3.895 $Y=2.035
+ $X2=0 $Y2=0
cc_341 N_A_27_368#_M1017_s N_A_499_368#_c_549_n 0.00266942f $X=3.845 $Y=1.84
+ $X2=0 $Y2=0
cc_342 N_A_27_368#_c_392_n N_A_499_368#_c_549_n 0.0184743f $X=3.98 $Y=2.115
+ $X2=0 $Y2=0
cc_343 N_A_27_368#_c_392_n N_A_879_368#_c_610_n 0.0128664f $X=3.98 $Y=2.115
+ $X2=0 $Y2=0
cc_344 N_A_27_368#_c_392_n N_A_879_368#_c_611_n 0.0396908f $X=3.98 $Y=2.115
+ $X2=0 $Y2=0
cc_345 N_A_27_368#_c_387_n N_VPWR_c_683_n 0.0439866f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_388_n N_VPWR_c_683_n 0.0236566f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_27_368#_c_389_n N_VPWR_c_683_n 0.0562636f $X=2.095 $Y=2.99 $X2=0
+ $Y2=0
cc_348 N_A_27_368#_c_391_n N_VPWR_c_683_n 0.0178163f $X=1.27 $Y=2.99 $X2=0 $Y2=0
cc_349 N_A_27_368#_c_387_n N_VPWR_c_680_n 0.0246722f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_350 N_A_27_368#_c_388_n N_VPWR_c_680_n 0.0128296f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_389_n N_VPWR_c_680_n 0.0314185f $X=2.095 $Y=2.99 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_391_n N_VPWR_c_680_n 0.00958215f $X=1.27 $Y=2.99 $X2=0
+ $Y2=0
cc_353 N_Y_c_445_n N_VGND_M1001_d 0.00326483f $X=0.355 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_354 N_Y_c_449_n N_VGND_M1001_d 5.5277e-19 $X=0.615 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_355 N_Y_c_451_n N_VGND_M1022_d 0.00250873f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_356 N_Y_c_446_n N_VGND_M1023_d 0.00250873f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_357 N_Y_c_448_n N_VGND_M1020_s 0.0398609f $X=7.24 $Y=1.045 $X2=0 $Y2=0
cc_358 N_Y_c_445_n N_VGND_c_761_n 0.0207726f $X=0.355 $Y=1.095 $X2=0 $Y2=0
cc_359 N_Y_c_449_n N_VGND_c_761_n 0.00427553f $X=0.615 $Y=0.765 $X2=0 $Y2=0
cc_360 N_Y_c_450_n N_VGND_c_761_n 0.0232074f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_361 N_Y_c_450_n N_VGND_c_762_n 0.0192747f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_362 N_Y_c_451_n N_VGND_c_762_n 0.0209867f $X=2.41 $Y=0.765 $X2=0 $Y2=0
cc_363 N_Y_c_452_n N_VGND_c_762_n 0.0213507f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_364 N_Y_c_446_n N_VGND_c_763_n 0.0209867f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_365 N_Y_c_447_n N_VGND_c_763_n 0.0191765f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_366 N_Y_c_452_n N_VGND_c_763_n 0.0192747f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_367 N_Y_c_447_n N_VGND_c_765_n 0.0174363f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_368 N_Y_c_448_n N_VGND_c_765_n 0.181264f $X=7.24 $Y=1.045 $X2=0 $Y2=0
cc_369 N_Y_c_454_n N_VGND_c_766_n 0.0265927f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_370 N_Y_c_452_n N_VGND_c_767_n 0.0523677f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_371 N_Y_c_454_n N_VGND_c_770_n 0.0288054f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_372 N_Y_c_450_n N_VGND_c_772_n 0.0499979f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_373 N_Y_c_447_n N_VGND_c_773_n 0.0118826f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_374 N_Y_c_450_n N_VGND_c_773_n 0.041525f $X=1.74 $Y=0.765 $X2=0 $Y2=0
cc_375 N_Y_c_452_n N_VGND_c_773_n 0.0434345f $X=3.59 $Y=0.765 $X2=0 $Y2=0
cc_376 N_Y_c_454_n N_VGND_c_773_n 0.02303f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_377 N_Y_c_447_n N_VGND_c_775_n 0.0144922f $X=4.425 $Y=0.515 $X2=0 $Y2=0
cc_378 N_Y_c_454_n N_VGND_c_776_n 0.0203431f $X=7.335 $Y=0.965 $X2=0 $Y2=0
cc_379 N_A_499_368#_c_549_n N_A_879_368#_M1000_s 0.00266942f $X=4.825 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_380 N_A_499_368#_c_550_n N_A_879_368#_M1005_s 0.00187091f $X=5.745 $Y=2.99
+ $X2=0 $Y2=0
cc_381 N_A_499_368#_c_549_n N_A_879_368#_c_611_n 0.0184743f $X=4.825 $Y=2.99
+ $X2=0 $Y2=0
cc_382 N_A_499_368#_M1000_d N_A_879_368#_c_618_n 0.00318402f $X=4.855 $Y=1.84
+ $X2=0 $Y2=0
cc_383 N_A_499_368#_c_567_n N_A_879_368#_c_618_n 0.0162994f $X=4.99 $Y=2.385
+ $X2=0 $Y2=0
cc_384 N_A_499_368#_c_550_n N_A_879_368#_c_662_n 0.0133959f $X=5.745 $Y=2.99
+ $X2=0 $Y2=0
cc_385 N_A_499_368#_M1010_d N_A_879_368#_c_622_n 0.00318402f $X=5.775 $Y=1.84
+ $X2=0 $Y2=0
cc_386 N_A_499_368#_c_573_n N_A_879_368#_c_622_n 0.0162994f $X=5.91 $Y=2.385
+ $X2=0 $Y2=0
cc_387 N_A_499_368#_c_550_n N_A_879_368#_c_612_n 0.00375633f $X=5.745 $Y=2.99
+ $X2=0 $Y2=0
cc_388 N_A_499_368#_c_550_n N_VPWR_c_681_n 0.00294199f $X=5.745 $Y=2.99 $X2=0
+ $Y2=0
cc_389 N_A_499_368#_c_547_n N_VPWR_c_683_n 0.0357927f $X=3.365 $Y=2.99 $X2=0
+ $Y2=0
cc_390 N_A_499_368#_c_548_n N_VPWR_c_683_n 0.0234458f $X=2.795 $Y=2.99 $X2=0
+ $Y2=0
cc_391 N_A_499_368#_c_549_n N_VPWR_c_683_n 0.0718669f $X=4.825 $Y=2.99 $X2=0
+ $Y2=0
cc_392 N_A_499_368#_c_550_n N_VPWR_c_683_n 0.0605268f $X=5.745 $Y=2.99 $X2=0
+ $Y2=0
cc_393 N_A_499_368#_c_551_n N_VPWR_c_683_n 0.0234458f $X=3.53 $Y=2.99 $X2=0
+ $Y2=0
cc_394 N_A_499_368#_c_552_n N_VPWR_c_683_n 0.0234458f $X=4.99 $Y=2.99 $X2=0
+ $Y2=0
cc_395 N_A_499_368#_c_547_n N_VPWR_c_680_n 0.0200586f $X=3.365 $Y=2.99 $X2=0
+ $Y2=0
cc_396 N_A_499_368#_c_548_n N_VPWR_c_680_n 0.0125551f $X=2.795 $Y=2.99 $X2=0
+ $Y2=0
cc_397 N_A_499_368#_c_549_n N_VPWR_c_680_n 0.0411134f $X=4.825 $Y=2.99 $X2=0
+ $Y2=0
cc_398 N_A_499_368#_c_550_n N_VPWR_c_680_n 0.0333657f $X=5.745 $Y=2.99 $X2=0
+ $Y2=0
cc_399 N_A_499_368#_c_551_n N_VPWR_c_680_n 0.0125551f $X=3.53 $Y=2.99 $X2=0
+ $Y2=0
cc_400 N_A_499_368#_c_552_n N_VPWR_c_680_n 0.0125551f $X=4.99 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_879_368#_c_627_n N_VPWR_M1008_s 0.00781989f $X=7.195 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_402 N_A_879_368#_c_641_n N_VPWR_M1018_s 0.00595031f $X=8.195 $Y=2.035 $X2=0
+ $Y2=0
cc_403 N_A_879_368#_c_612_n N_VPWR_c_681_n 0.0258971f $X=6.36 $Y=2.445 $X2=0
+ $Y2=0
cc_404 N_A_879_368#_c_627_n N_VPWR_c_681_n 0.0208278f $X=7.195 $Y=2.035 $X2=0
+ $Y2=0
cc_405 N_A_879_368#_c_613_n N_VPWR_c_681_n 0.0266809f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_406 N_A_879_368#_c_613_n N_VPWR_c_682_n 0.0266809f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_407 N_A_879_368#_c_641_n N_VPWR_c_682_n 0.0208278f $X=8.195 $Y=2.035 $X2=0
+ $Y2=0
cc_408 N_A_879_368#_c_615_n N_VPWR_c_682_n 0.0266809f $X=8.36 $Y=2.815 $X2=0
+ $Y2=0
cc_409 N_A_879_368#_c_612_n N_VPWR_c_683_n 0.0118717f $X=6.36 $Y=2.445 $X2=0
+ $Y2=0
cc_410 N_A_879_368#_c_613_n N_VPWR_c_685_n 0.0144623f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_411 N_A_879_368#_c_615_n N_VPWR_c_686_n 0.014549f $X=8.36 $Y=2.815 $X2=0
+ $Y2=0
cc_412 N_A_879_368#_c_612_n N_VPWR_c_680_n 0.00975826f $X=6.36 $Y=2.445 $X2=0
+ $Y2=0
cc_413 N_A_879_368#_c_613_n N_VPWR_c_680_n 0.0118344f $X=7.36 $Y=2.815 $X2=0
+ $Y2=0
cc_414 N_A_879_368#_c_615_n N_VPWR_c_680_n 0.0119743f $X=8.36 $Y=2.815 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o21a_2.pex.spice
* Created: Fri Aug 28 17:54:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21A_2%A1 1 3 6 8 9 10 11
c25 11 0 1.25174e-19 $X=0.72 $Y=1.295
c26 1 0 1.4014e-19 $X=0.7 $Y=1.22
r27 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r28 11 16 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r29 10 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r30 8 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.625 $Y=1.385
+ $X2=0.61 $Y2=1.385
r31 8 9 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.385
+ $X2=0.625 $Y2=1.22
r32 4 9 34.7346 $w=1.65e-07 $l=3.76696e-07 $layer=POLY_cond $X=0.725 $Y=1.55
+ $X2=0.625 $Y2=1.22
r33 4 6 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.725 $Y=1.55
+ $X2=0.725 $Y2=2.34
r34 1 9 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.625
+ $Y2=1.22
r35 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.7
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%A2 3 7 8 11 13
c31 13 0 1.25174e-19 $X=1.22 $Y=1.22
c32 8 0 1.79042e-19 $X=1.2 $Y=1.295
r33 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.385
+ $X2=1.22 $Y2=1.55
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.385
+ $X2=1.22 $Y2=1.22
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.385 $X2=1.22 $Y2=1.385
r36 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.22 $Y=1.295 $X2=1.22
+ $Y2=1.385
r37 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.31 $Y=0.74 $X2=1.31
+ $Y2=1.22
r38 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.145 $Y=2.34
+ $X2=1.145 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%B1 3 7 8 11 12 13
c39 13 0 3.89014e-20 $X=1.79 $Y=1.22
c40 3 0 9.62843e-20 $X=1.715 $Y=2.34
r41 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.385
+ $X2=1.79 $Y2=1.55
r42 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.385
+ $X2=1.79 $Y2=1.22
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.385 $X2=1.79 $Y2=1.385
r44 8 12 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.79 $Y2=1.365
r45 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.785 $Y=0.74
+ $X2=1.785 $Y2=1.22
r46 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.715 $Y=2.34
+ $X2=1.715 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%A_247_368# 1 2 9 13 15 17 18 19 20 22 25 29
+ 30 33 36 38 39 43
r78 48 49 8.48094 $w=3.41e-07 $l=6e-08 $layer=POLY_cond $X=2.855 $Y=1.415
+ $X2=2.915 $Y2=1.415
r79 44 48 53.0059 $w=3.41e-07 $l=3.75e-07 $layer=POLY_cond $X=2.48 $Y=1.415
+ $X2=2.855 $Y2=1.415
r80 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.385 $X2=2.48 $Y2=1.385
r81 40 43 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.21 $Y=1.385
+ $X2=2.48 $Y2=1.385
r82 37 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.55
+ $X2=2.21 $Y2=1.385
r83 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.21 $Y=1.55
+ $X2=2.21 $Y2=1.72
r84 36 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=1.22
+ $X2=2.21 $Y2=1.385
r85 36 39 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.21 $Y=1.22
+ $X2=2.21 $Y2=1.01
r86 31 39 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.1 $Y=0.815
+ $X2=2.1 $Y2=1.01
r87 31 33 9.16044 $w=3.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.1 $Y=0.815 $X2=2.1
+ $Y2=0.505
r88 29 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.125 $Y=1.805
+ $X2=2.21 $Y2=1.72
r89 29 30 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.125 $Y=1.805
+ $X2=1.655 $Y2=1.805
r90 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.49 $Y=1.985
+ $X2=1.49 $Y2=2.695
r91 23 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.49 $Y=1.89
+ $X2=1.655 $Y2=1.805
r92 23 25 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.49 $Y=1.89
+ $X2=1.49 $Y2=1.985
r93 20 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.345 $Y=1.22
+ $X2=3.345 $Y2=0.74
r94 19 49 25.9675 $w=3.41e-07 $l=1.52971e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.915 $Y2=1.415
r95 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.27 $Y=1.295
+ $X2=3.345 $Y2=1.22
r96 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.27 $Y=1.295
+ $X2=2.99 $Y2=1.295
r97 15 49 22.0049 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.915 $Y=1.22
+ $X2=2.915 $Y2=1.415
r98 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.915 $Y=1.22
+ $X2=2.915 $Y2=0.74
r99 11 48 17.6972 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=2.855 $Y=1.61
+ $X2=2.855 $Y2=1.415
r100 11 13 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.855 $Y=1.61
+ $X2=2.855 $Y2=2.4
r101 7 44 10.6012 $w=3.41e-07 $l=7.5e-08 $layer=POLY_cond $X=2.405 $Y=1.415
+ $X2=2.48 $Y2=1.415
r102 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.405 $Y=1.55
+ $X2=2.405 $Y2=2.4
r103 2 27 400 $w=1.7e-07 $l=9.74192e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.84 $X2=1.49 $Y2=2.695
r104 2 25 400 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.84 $X2=1.49 $Y2=1.985
r105 1 33 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.37 $X2=2 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%VPWR 1 2 3 12 18 24 27 28 29 35 42 49 50 53
+ 56
r42 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 50 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 47 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.13 $Y2=3.33
r47 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 46 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 43 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.13 $Y2=3.33
r52 43 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.13 $Y2=3.33
r54 42 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r58 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 35 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.13 $Y2=3.33
r60 35 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 33 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 29 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 29 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 27 32 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.335 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.335 $Y=3.33
+ $X2=0.5 $Y2=3.33
r67 26 37 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.665 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.665 $Y=3.33
+ $X2=0.5 $Y2=3.33
r69 22 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r70 22 24 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.225
r71 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.13 $Y=2.145
+ $X2=2.13 $Y2=2.825
r72 16 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=3.33
r73 16 21 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=2.825
r74 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.5 $Y=1.985 $X2=0.5
+ $Y2=2.695
r75 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.5 $Y=3.245 $X2=0.5
+ $Y2=3.33
r76 10 15 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.5 $Y=3.245 $X2=0.5
+ $Y2=2.695
r77 3 24 300 $w=1.7e-07 $l=4.68455e-07 $layer=licon1_PDIFF $count=2 $X=2.945
+ $Y=1.84 $X2=3.13 $Y2=2.225
r78 2 21 400 $w=1.7e-07 $l=1.13594e-06 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.84 $X2=2.13 $Y2=2.825
r79 2 18 400 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.84 $X2=2.13 $Y2=2.145
r80 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.5 $Y2=2.695
r81 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.84 $X2=0.5 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%X 1 2 9 13 14 15 16 22 33
c31 22 0 9.62843e-20 $X=3.13 $Y=1.72
r32 22 33 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=3.13 $Y=1.72
+ $X2=3.13 $Y2=1.665
r33 16 22 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.805
+ $X2=3.13 $Y2=1.805
r34 16 33 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.13 $Y=1.65
+ $X2=3.13 $Y2=1.665
r35 15 16 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.65
r36 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=0.925
+ $X2=3.13 $Y2=1.295
r37 13 14 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.13 $Y=0.515
+ $X2=3.13 $Y2=0.925
r38 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.63 $Y=1.985
+ $X2=2.63 $Y2=2.815
r39 7 16 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.63 $Y=1.805
+ $X2=3.12 $Y2=1.805
r40 7 9 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.63 $Y=1.89 $X2=2.63
+ $Y2=1.985
r41 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.815
r42 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=1.985
r43 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.99
+ $Y=0.37 $X2=3.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%A_54_74# 1 2 7 9 11 13 15
r26 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.84 $X2=1.57
+ $Y2=0.925
r27 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.57 $Y=0.84
+ $X2=1.57 $Y2=0.505
r28 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0.925
+ $X2=0.415 $Y2=0.925
r29 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.925
+ $X2=1.57 $Y2=0.925
r30 11 12 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.405 $Y=0.925
+ $X2=0.58 $Y2=0.925
r31 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=0.84 $X2=0.415
+ $Y2=0.925
r32 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.415 $Y=0.84
+ $X2=0.415 $Y2=0.505
r33 2 20 182 $w=1.7e-07 $l=6.40859e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.37 $X2=1.57 $Y2=0.925
r34 2 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.37 $X2=1.57 $Y2=0.505
r35 1 18 182 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.37 $X2=0.415 $Y2=0.925
r36 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.37 $X2=0.415 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__O21A_2%VGND 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r44 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r48 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r51 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.12
+ $Y2=0
r52 34 46 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.657
+ $Y2=0
r53 34 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.12
+ $Y2=0
r54 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r55 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 30 40 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=0.992
+ $Y2=0
r57 30 32 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=2.16
+ $Y2=0
r58 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r59 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.16
+ $Y2=0
r60 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r61 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r62 24 40 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.992
+ $Y2=0
r63 24 26 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.72
+ $Y2=0
r64 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r65 22 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r66 18 46 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.657 $Y2=0
r67 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=0.085 $X2=3.6
+ $Y2=0.515
r68 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r69 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.515
r70 10 40 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.992 $Y=0.085
+ $X2=0.992 $Y2=0
r71 10 12 10.6044 $w=4.83e-07 $l=4.3e-07 $layer=LI1_cond $X=0.992 $Y=0.085
+ $X2=0.992 $Y2=0.515
r72 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.515
r73 2 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.37 $X2=2.63 $Y2=0.515
r74 1 12 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.37 $X2=0.99 $Y2=0.515
.ends


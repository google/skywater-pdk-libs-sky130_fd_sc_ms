* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkinv_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X35 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X38 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

* File: sky130_fd_sc_ms__o21ai_2.pex.spice
* Created: Fri Aug 28 17:54:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21AI_2%A1 3 7 11 15 19 20 22 23 25 31 32
c79 32 0 1.62564e-19 $X=1.92 $Y=1.515
c80 31 0 1.76387e-19 $X=1.92 $Y=1.515
c81 20 0 1.66928e-19 $X=0.43 $Y=1.515
c82 15 0 1.83442e-19 $X=1.955 $Y=2.4
c83 11 0 1.73347e-19 $X=1.925 $Y=0.74
r84 31 34 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.515
+ $X2=1.92 $Y2=1.68
r85 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.515
+ $X2=1.92 $Y2=1.35
r86 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.515 $X2=1.92 $Y2=1.515
r87 25 32 3.45023 $w=5.18e-07 $l=1.5e-07 $layer=LI1_cond $X=2.015 $Y=1.665
+ $X2=2.015 $Y2=1.515
r88 24 25 6.55543 $w=5.18e-07 $l=2.85e-07 $layer=LI1_cond $X=2.015 $Y=1.95
+ $X2=2.015 $Y2=1.665
r89 22 24 9.39785 $w=1.7e-07 $l=2.995e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=2.015 $Y2=1.95
r90 22 23 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=0.595 $Y2=2.035
r91 20 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.515
+ $X2=0.43 $Y2=1.68
r92 20 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.515
+ $X2=0.43 $Y2=1.35
r93 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.515 $X2=0.43 $Y2=1.515
r94 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.43 $Y=1.95
+ $X2=0.595 $Y2=2.035
r95 17 19 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.43 $Y=1.95
+ $X2=0.43 $Y2=1.515
r96 15 34 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.955 $Y=2.4
+ $X2=1.955 $Y2=1.68
r97 11 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=0.74
+ $X2=1.925 $Y2=1.35
r98 7 28 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.35
r99 3 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%A2 3 7 11 15 17 23 24
c58 23 0 1.02944e-19 $X=1.35 $Y=1.515
r59 24 25 2.23839 $w=3.23e-07 $l=1.5e-08 $layer=POLY_cond $X=1.44 $Y=1.515
+ $X2=1.455 $Y2=1.515
r60 22 24 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=1.35 $Y=1.515
+ $X2=1.44 $Y2=1.515
r61 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.515 $X2=1.35 $Y2=1.515
r62 20 22 52.9752 $w=3.23e-07 $l=3.55e-07 $layer=POLY_cond $X=0.995 $Y=1.515
+ $X2=1.35 $Y2=1.515
r63 19 20 5.96904 $w=3.23e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.515
+ $X2=0.995 $Y2=1.515
r64 17 23 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.515
r65 13 25 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.515
r66 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r67 9 24 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.35
+ $X2=1.44 $Y2=1.515
r68 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.44 $Y=1.35 $X2=1.44
+ $Y2=0.74
r69 5 20 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r70 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r71 1 19 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.515
r72 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%B1 3 7 9 11 13 15 17 18 19
c50 19 0 1.98552e-19 $X=3.12 $Y=1.295
c51 3 0 1.89026e-19 $X=2.405 $Y=2.4
r52 22 24 12.518 $w=4.12e-07 $l=1.07e-07 $layer=POLY_cond $X=3 $Y=1.385 $X2=3
+ $Y2=1.492
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.385 $X2=3.07 $Y2=1.385
r54 19 23 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.07 $Y=1.295 $X2=3.07
+ $Y2=1.385
r55 15 22 39.8282 $w=4.12e-07 $l=2.22486e-07 $layer=POLY_cond $X=2.865 $Y=1.22
+ $X2=3 $Y2=1.385
r56 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.865 $Y=1.22
+ $X2=2.865 $Y2=0.74
r57 11 24 29.9374 $w=4.12e-07 $l=1.97129e-07 $layer=POLY_cond $X=2.855 $Y=1.615
+ $X2=3 $Y2=1.492
r58 11 13 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=2.855 $Y=1.615
+ $X2=2.855 $Y2=2.4
r59 10 18 0.134175 $w=2.45e-07 $l=1.93494e-07 $layer=POLY_cond $X=2.495 $Y=1.492
+ $X2=2.315 $Y2=1.52
r60 9 24 14.985 $w=2.45e-07 $l=2.35e-07 $layer=POLY_cond $X=2.765 $Y=1.492 $X2=3
+ $Y2=1.492
r61 9 10 68.4515 $w=2.45e-07 $l=2.7e-07 $layer=POLY_cond $X=2.765 $Y=1.492
+ $X2=2.495 $Y2=1.492
r62 5 18 27.9716 $w=1.65e-07 $l=1.8775e-07 $layer=POLY_cond $X=2.4 $Y=1.37
+ $X2=2.315 $Y2=1.52
r63 5 7 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.4 $Y=1.37 $X2=2.4
+ $Y2=0.74
r64 1 18 27.9716 $w=1.65e-07 $l=1.32571e-07 $layer=POLY_cond $X=2.405 $Y=1.615
+ $X2=2.315 $Y2=1.52
r65 1 3 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=2.405 $Y=1.615
+ $X2=2.405 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%VPWR 1 2 3 10 12 16 18 20 24 26 31 40 44
c49 2 0 1.62564e-19 $X=2.045 $Y=1.84
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 35 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 32 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.22 $Y2=3.33
r57 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 31 43 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r59 31 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 27 37 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r63 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 26 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.22 $Y2=3.33
r65 26 29 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r67 24 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 20 23 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=2.815
r69 18 43 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r70 18 23 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r71 14 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=3.245
+ $X2=2.22 $Y2=3.33
r72 14 16 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=2.22 $Y=3.245
+ $X2=2.22 $Y2=2.805
r73 10 37 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r74 10 12 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.455
r75 3 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.815
r76 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=1.985
r77 2 16 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.84 $X2=2.18 $Y2=2.805
r78 1 12 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%A_119_368# 1 2 9 11 12 14
c30 14 0 1.89026e-19 $X=1.73 $Y=2.805
c31 11 0 8.04979e-20 $X=1.565 $Y=2.99
r32 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.73 $Y=2.805
+ $X2=1.73 $Y2=2.99
r33 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=1.73 $Y2=2.99
r34 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=0.895 $Y2=2.99
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r36 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.73 $Y=2.905 $X2=0.73
+ $Y2=2.455
r37 2 14 600 $w=1.7e-07 $l=1.05345e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.73 $Y2=2.805
r38 1 9 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%Y 1 2 3 10 14 18 23 24 25 26 36 44
c43 44 0 1.76387e-19 $X=2.66 $Y=1.82
r44 32 36 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.66 $Y=1.955 $X2=2.66
+ $Y2=1.985
r45 25 33 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.375
+ $X2=2.66 $Y2=2.29
r46 25 38 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.375
+ $X2=2.66 $Y2=2.46
r47 25 26 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=2.66 $Y=2.475 $X2=2.66
+ $Y2=2.775
r48 25 38 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.66 $Y=2.475
+ $X2=2.66 $Y2=2.46
r49 24 32 0.128049 $w=2.68e-07 $l=3e-09 $layer=LI1_cond $X=2.66 $Y=1.952
+ $X2=2.66 $Y2=1.955
r50 24 44 6.23403 $w=2.68e-07 $l=1.32e-07 $layer=LI1_cond $X=2.66 $Y=1.952
+ $X2=2.66 $Y2=1.82
r51 24 33 10.7988 $w=2.68e-07 $l=2.53e-07 $layer=LI1_cond $X=2.66 $Y=2.037
+ $X2=2.66 $Y2=2.29
r52 24 36 2.21952 $w=2.68e-07 $l=5.2e-08 $layer=LI1_cond $X=2.66 $Y=2.037
+ $X2=2.66 $Y2=1.985
r53 23 44 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=2.63 $Y=1.13
+ $X2=2.63 $Y2=1.82
r54 18 21 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.23 $Y=2.375
+ $X2=1.23 $Y2=2.51
r55 12 23 6.22208 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.605 $Y=1 $X2=2.605
+ $Y2=1.13
r56 12 14 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=2.605 $Y=1 $X2=2.605
+ $Y2=0.88
r57 11 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.375
+ $X2=1.23 $Y2=2.375
r58 10 25 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=2.66 $Y2=2.375
r59 10 11 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=2.525 $Y=2.375
+ $X2=1.395 $Y2=2.375
r60 3 25 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.4
r61 3 36 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=1.985
r62 2 21 600 $w=1.7e-07 $l=7.56869e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.51
r63 1 14 182 $w=1.7e-07 $l=5.88897e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.37 $X2=2.645 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%A_27_74# 1 2 3 4 15 17 18 21 23 25 27 31 35
c60 27 0 1.98552e-19 $X=2.915 $Y=0.435
c61 25 0 1.73347e-19 $X=2.18 $Y=0.52
c62 17 0 1.66928e-19 $X=1.125 $Y=1.095
r63 28 33 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.305 $Y=0.435
+ $X2=2.18 $Y2=0.435
r64 27 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.435
+ $X2=3.08 $Y2=0.435
r65 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.435
+ $X2=2.305 $Y2=0.435
r66 25 33 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.52 $X2=2.18
+ $Y2=0.435
r67 25 26 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=2.18 $Y=0.52
+ $X2=2.18 $Y2=1.01
r68 24 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.095
+ $X2=1.25 $Y2=1.095
r69 23 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.18 $Y2=1.01
r70 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=1.375 $Y2=1.095
r71 19 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.01
+ $X2=1.25 $Y2=1.095
r72 19 21 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.25 $Y=1.01
+ $X2=1.25 $Y2=0.515
r73 17 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=1.25 $Y2=1.095
r74 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=0.445 $Y2=1.095
r75 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r76 13 15 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r77 4 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
r78 3 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r79 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r80 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r44 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r48 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r50 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.16
+ $Y2=0
r51 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r54 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r55 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r56 22 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r57 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r60 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r61 15 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r62 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 15 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r65 11 13 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.665
r66 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r67 7 9 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.665
r68 2 13 182 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.37 $X2=1.71 $Y2=0.665
r69 1 9 182 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.665
.ends


* File: sky130_fd_sc_ms__dlxtp_1.spice
* Created: Fri Aug 28 17:30:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlxtp_1.pex.spice"
.subckt sky130_fd_sc_ms__dlxtp_1  VNB VPB D GATE VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_A_119_88#_M1006_d N_D_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.1815 AS=0.1705 PD=1.76 PS=1.72 NRD=9.816 NRS=5.448 M=1 R=3.66667
+ SA=75000.2 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1001 N_VGND_M1001_d N_A_119_88#_M1001_g N_A_239_85#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.250643 AS=0.2238 PD=1.89466 PS=2.14 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1014 A_514_149# N_A_386_326#_M1014_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.142257 PD=0.66 PS=1.07534 NRD=18.564 NRS=125.712 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_592_149#_M1004_d N_A_562_123#_M1004_g A_514_149# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0996776 AS=0.0504 PD=0.872586 PS=0.66 NRD=24.276 NRS=18.564 M=1
+ R=2.8 SA=75001.5 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_239_85#_M1015_d N_A_685_59#_M1015_g N_A_592_149#_M1004_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.222 AS=0.175622 PD=2.08 PS=1.53741 NRD=0.804 NRS=16.212 M=1
+ R=4.93333 SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_592_149#_M1009_g N_A_386_326#_M1009_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.19615 AS=0.2109 PD=1.41 PS=2.05 NRD=34.056 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1003 N_A_685_59#_M1003_d N_A_562_123#_M1003_g N_VGND_M1009_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.19615 PD=2.05 PS=1.41 NRD=0 NRS=34.056 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_GATE_M1016_g N_A_562_123#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.261625 AS=0.222 PD=1.545 PS=2.08 NRD=48.408 NRS=1.62 M=1 R=4.93333
+ SA=75000.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1005 N_Q_M1005_d N_A_386_326#_M1005_g N_VGND_M1016_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.261625 PD=2.05 PS=1.545 NRD=0 NRS=48.408 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_119_88#_M1008_d N_D_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2352 AS=0.2352 PD=2.24 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1007 N_VPWR_M1007_d N_A_119_88#_M1007_g N_A_229_392#_M1007_s VPB PSHORT L=0.18
+ W=1 AD=0.257658 AS=0.28 PD=2.35211 PS=2.56 NRD=39.9122 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90000.4 A=0.18 P=2.36 MULT=1
MM1002 N_A_422_392#_M1002_d N_A_386_326#_M1002_g N_VPWR_M1007_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1176 AS=0.108217 PD=1.4 PS=0.987887 NRD=0 NRS=95.0525 M=1
+ R=2.33333 SA=90000.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1013 N_A_592_149#_M1013_d N_A_562_123#_M1013_g N_A_229_392#_M1013_s VPB PSHORT
+ L=0.18 W=1 AD=0.219366 AS=0.28 PD=1.90845 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90000.5 A=0.18 P=2.36 MULT=1
MM1017 N_A_422_392#_M1017_d N_A_685_59#_M1017_g N_A_592_149#_M1013_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.18665 AS=0.0921338 PD=1.8 PS=0.801549 NRD=39.8531
+ NRS=77.0861 M=1 R=2.33333 SA=90000.7 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_592_149#_M1010_g N_A_386_326#_M1010_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.3276 AS=0.3528 PD=2.18286 PS=2.87 NRD=41.764 NRS=2.6201 M=1
+ R=6.22222 SA=90000.2 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1011 N_A_685_59#_M1011_d N_A_562_123#_M1011_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2457 PD=2.24 PS=1.63714 NRD=0 NRS=55.6919 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1012 N_VPWR_M1012_d N_GATE_M1012_g N_A_562_123#_M1012_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1854 AS=0.2352 PD=1.30714 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1000 N_Q_M1000_d N_A_386_326#_M1000_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2472 PD=2.8 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=15.2636 P=20.15
c_81 VNB 0 7.64129e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dlxtp_1.pxi.spice"
*
.ends
*
*

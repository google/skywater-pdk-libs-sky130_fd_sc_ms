* File: sky130_fd_sc_ms__o31a_1.pxi.spice
* Created: Fri Aug 28 18:02:01 2020
* 
x_PM_SKY130_FD_SC_MS__O31A_1%A_84_48# N_A_84_48#_M1001_d N_A_84_48#_M1002_d
+ N_A_84_48#_M1008_g N_A_84_48#_M1006_g N_A_84_48#_c_67_n N_A_84_48#_c_83_p
+ N_A_84_48#_c_126_p N_A_84_48#_c_75_n N_A_84_48#_c_76_n N_A_84_48#_c_68_n
+ N_A_84_48#_c_69_n N_A_84_48#_c_70_n N_A_84_48#_c_71_n N_A_84_48#_c_99_p
+ N_A_84_48#_c_72_n PM_SKY130_FD_SC_MS__O31A_1%A_84_48#
x_PM_SKY130_FD_SC_MS__O31A_1%A1 N_A1_M1007_g N_A1_M1004_g A1 N_A1_c_151_n
+ N_A1_c_152_n PM_SKY130_FD_SC_MS__O31A_1%A1
x_PM_SKY130_FD_SC_MS__O31A_1%A2 N_A2_M1003_g N_A2_M1009_g A2 N_A2_c_192_n
+ N_A2_c_193_n PM_SKY130_FD_SC_MS__O31A_1%A2
x_PM_SKY130_FD_SC_MS__O31A_1%A3 N_A3_M1002_g N_A3_M1000_g A3 N_A3_c_226_n
+ N_A3_c_227_n PM_SKY130_FD_SC_MS__O31A_1%A3
x_PM_SKY130_FD_SC_MS__O31A_1%B1 N_B1_M1005_g N_B1_M1001_g B1 N_B1_c_264_n
+ N_B1_c_265_n PM_SKY130_FD_SC_MS__O31A_1%B1
x_PM_SKY130_FD_SC_MS__O31A_1%X N_X_M1008_s N_X_M1006_s N_X_c_295_n N_X_c_296_n X
+ X X X N_X_c_297_n PM_SKY130_FD_SC_MS__O31A_1%X
x_PM_SKY130_FD_SC_MS__O31A_1%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_321_n
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n VPWR N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_320_n N_VPWR_c_328_n PM_SKY130_FD_SC_MS__O31A_1%VPWR
x_PM_SKY130_FD_SC_MS__O31A_1%VGND N_VGND_M1008_d N_VGND_M1003_d N_VGND_c_360_n
+ N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n VGND N_VGND_c_364_n
+ N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n PM_SKY130_FD_SC_MS__O31A_1%VGND
x_PM_SKY130_FD_SC_MS__O31A_1%A_230_94# N_A_230_94#_M1007_d N_A_230_94#_M1000_d
+ N_A_230_94#_c_399_n N_A_230_94#_c_400_n N_A_230_94#_c_401_n
+ N_A_230_94#_c_402_n PM_SKY130_FD_SC_MS__O31A_1%A_230_94#
cc_1 VNB N_A_84_48#_M1008_g 0.030112f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_M1006_g 5.70835e-19 $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_3 VNB N_A_84_48#_c_67_n 2.46719e-19 $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.95
cc_4 VNB N_A_84_48#_c_68_n 0.0233423f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.615
cc_5 VNB N_A_84_48#_c_69_n 0.0253498f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=1.95
cc_6 VNB N_A_84_48#_c_70_n 0.0338659f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_7 VNB N_A_84_48#_c_71_n 0.0026276f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_8 VNB N_A_84_48#_c_72_n 0.0137511f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=1.13
cc_9 VNB N_A1_M1007_g 0.026484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_151_n 0.0243418f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_11 VNB N_A1_c_152_n 0.00495499f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_12 VNB N_A2_M1003_g 0.0247917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1009_g 0.00133404f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.32
cc_14 VNB N_A2_c_192_n 0.032497f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_15 VNB N_A2_c_193_n 0.00206174f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_16 VNB N_A3_M1000_g 0.0277067f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.32
cc_17 VNB N_A3_c_226_n 0.0263879f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_18 VNB N_A3_c_227_n 0.00182951f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_19 VNB N_B1_M1001_g 0.0287531f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.32
cc_20 VNB N_B1_c_264_n 0.0266136f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_21 VNB N_B1_c_265_n 0.00535768f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_22 VNB N_X_c_295_n 0.0265914f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_23 VNB N_X_c_296_n 0.0139041f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_24 VNB N_X_c_297_n 0.0249534f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=1.95
cc_25 VNB N_VPWR_c_320_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_26 VNB N_VGND_c_360_n 0.0212254f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_27 VNB N_VGND_c_361_n 0.0189386f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.65
cc_28 VNB N_VGND_c_362_n 0.023893f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.035
cc_29 VNB N_VGND_c_363_n 0.00702069f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.12
cc_30 VNB N_VGND_c_364_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.715
cc_31 VNB N_VGND_c_365_n 0.0370094f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_32 VNB N_VGND_c_366_n 0.227175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_367_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.035
cc_34 VNB N_A_230_94#_c_399_n 0.00335993f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_35 VNB N_A_230_94#_c_400_n 0.0191055f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.65
cc_36 VNB N_A_230_94#_c_401_n 0.0070898f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_37 VNB N_A_230_94#_c_402_n 0.00330195f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.65
cc_38 VPB N_A_84_48#_M1006_g 0.0306852f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_39 VPB N_A_84_48#_c_67_n 0.00287184f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.95
cc_40 VPB N_A_84_48#_c_75_n 0.00483137f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.375
cc_41 VPB N_A_84_48#_c_76_n 0.0082934f $X=-0.19 $Y=1.66 $X2=3.085 $Y2=2.035
cc_42 VPB N_A_84_48#_c_69_n 0.0125324f $X=-0.19 $Y=1.66 $X2=3.17 $Y2=1.95
cc_43 VPB N_A1_M1004_g 0.0220334f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.32
cc_44 VPB N_A1_c_151_n 0.00562917f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_45 VPB N_A1_c_152_n 0.00301265f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_46 VPB N_A2_M1009_g 0.021567f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.32
cc_47 VPB N_A2_c_193_n 0.00294484f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_48 VPB N_A3_M1002_g 0.0233132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A3_c_226_n 0.00570789f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_50 VPB N_A3_c_227_n 0.00200497f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_51 VPB N_B1_M1005_g 0.0248849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_B1_c_264_n 0.00564178f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_53 VPB N_B1_c_265_n 0.00346359f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_54 VPB X 0.0142465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB X 0.0419191f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.715
cc_56 VPB N_X_c_297_n 0.0075744f $X=-0.19 $Y=1.66 $X2=3.17 $Y2=1.95
cc_57 VPB N_VPWR_c_321_n 0.0165614f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_58 VPB N_VPWR_c_322_n 0.0292965f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_59 VPB N_VPWR_c_323_n 0.0501782f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.95
cc_60 VPB N_VPWR_c_324_n 0.00603306f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=2.035
cc_61 VPB N_VPWR_c_325_n 0.0191572f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.375
cc_62 VPB N_VPWR_c_326_n 0.0120081f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_63 VPB N_VPWR_c_320_n 0.0973629f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_64 VPB N_VPWR_c_328_n 0.00891827f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.485
cc_65 N_A_84_48#_M1008_g N_A1_M1007_g 0.0209698f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A_84_48#_c_70_n N_A1_M1007_g 0.00145529f $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_67 N_A_84_48#_c_71_n N_A1_M1007_g 6.58026e-19 $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_68 N_A_84_48#_M1006_g N_A1_M1004_g 0.0155963f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A_84_48#_c_67_n N_A1_M1004_g 0.00351106f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_70 N_A_84_48#_c_83_p N_A1_M1004_g 0.0178415f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_71 N_A_84_48#_M1006_g N_A1_c_151_n 7.81769e-19 $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A_84_48#_c_67_n N_A1_c_151_n 2.15441e-19 $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_73 N_A_84_48#_c_83_p N_A1_c_151_n 7.00522e-19 $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_74 N_A_84_48#_c_70_n N_A1_c_151_n 0.0187646f $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_75 N_A_84_48#_c_71_n N_A1_c_151_n 0.00170526f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_76 N_A_84_48#_c_67_n N_A1_c_152_n 0.0102298f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_77 N_A_84_48#_c_83_p N_A1_c_152_n 0.0238723f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A_84_48#_c_70_n N_A1_c_152_n 3.43766e-19 $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_79 N_A_84_48#_c_71_n N_A1_c_152_n 0.0240984f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_80 N_A_84_48#_c_83_p N_A2_M1009_g 0.0172246f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_84_48#_c_75_n N_A2_M1009_g 0.00353794f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_82 N_A_84_48#_c_83_p N_A2_c_192_n 4.87141e-19 $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_83 N_A_84_48#_c_83_p N_A2_c_193_n 0.022134f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_84 N_A_84_48#_c_83_p N_A3_M1002_g 0.0131671f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_84_48#_c_75_n N_A3_M1002_g 0.0162942f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_86 N_A_84_48#_c_99_p N_A3_M1002_g 8.8334e-19 $X=2.36 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_84_48#_c_99_p N_A3_c_226_n 7.63688e-19 $X=2.36 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_84_48#_c_83_p N_A3_c_227_n 0.0108932f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_89 N_A_84_48#_c_99_p N_A3_c_227_n 0.0130747f $X=2.36 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A_84_48#_c_75_n N_B1_M1005_g 0.00959126f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_91 N_A_84_48#_c_76_n N_B1_M1005_g 0.0185418f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_84_48#_c_69_n N_B1_M1005_g 0.00553924f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_93 N_A_84_48#_c_68_n N_B1_M1001_g 0.0132958f $X=3.08 $Y=0.615 $X2=0 $Y2=0
cc_94 N_A_84_48#_c_69_n N_B1_M1001_g 0.00714331f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_95 N_A_84_48#_c_76_n N_B1_c_264_n 7.01228e-19 $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_84_48#_c_69_n N_B1_c_264_n 0.00739878f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_97 N_A_84_48#_c_76_n N_B1_c_265_n 0.0247432f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_84_48#_c_69_n N_B1_c_265_n 0.0330212f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A_84_48#_M1008_g N_X_c_295_n 0.00805909f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_84_48#_M1008_g N_X_c_296_n 0.00278926f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_84_48#_c_71_n N_X_c_296_n 0.00138666f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_102 N_A_84_48#_M1006_g X 0.00293426f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_84_48#_c_67_n X 0.00567891f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_104 N_A_84_48#_c_70_n X 2.41927e-19 $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_105 N_A_84_48#_c_71_n X 0.00231492f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_106 N_A_84_48#_M1006_g X 0.0148712f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_84_48#_M1008_g N_X_c_297_n 0.0122939f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_84_48#_M1006_g N_X_c_297_n 0.00262394f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_84_48#_c_67_n N_X_c_297_n 0.00525749f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_110 N_A_84_48#_c_71_n N_X_c_297_n 0.0249901f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_111 N_A_84_48#_c_67_n N_VPWR_M1006_d 0.00221445f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_84_48#_c_83_p N_VPWR_M1006_d 0.0113618f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_84_48#_c_126_p N_VPWR_M1006_d 0.00269585f $X=0.795 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_84_48#_c_76_n N_VPWR_M1005_d 0.0199129f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_84_48#_c_69_n N_VPWR_M1005_d 0.00225668f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_116 N_A_84_48#_M1006_g N_VPWR_c_321_n 0.00799837f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_84_48#_c_83_p N_VPWR_c_321_n 0.0213608f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_118 N_A_84_48#_c_126_p N_VPWR_c_321_n 0.0116292f $X=0.795 $Y=2.035 $X2=0
+ $Y2=0
cc_119 N_A_84_48#_c_70_n N_VPWR_c_321_n 3.55059e-19 $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_120 N_A_84_48#_c_75_n N_VPWR_c_322_n 0.0394063f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_121 N_A_84_48#_c_76_n N_VPWR_c_322_n 0.0206354f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_122 N_A_84_48#_c_75_n N_VPWR_c_323_n 0.010336f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_123 N_A_84_48#_M1006_g N_VPWR_c_325_n 0.005209f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_84_48#_M1006_g N_VPWR_c_320_n 0.00990503f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_84_48#_c_75_n N_VPWR_c_320_n 0.0113305f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_126 N_A_84_48#_c_83_p A_259_368# 0.0096152f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_84_48#_c_83_p A_343_368# 0.0146661f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_84_48#_M1008_g N_VGND_c_360_n 0.00946427f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_84_48#_c_70_n N_VGND_c_360_n 0.00320573f $X=0.59 $Y=1.485 $X2=0 $Y2=0
cc_130 N_A_84_48#_c_71_n N_VGND_c_360_n 0.0140528f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_131 N_A_84_48#_M1008_g N_VGND_c_364_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_84_48#_c_68_n N_VGND_c_365_n 0.0107295f $X=3.08 $Y=0.615 $X2=0 $Y2=0
cc_133 N_A_84_48#_M1008_g N_VGND_c_366_n 0.00828717f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_134 N_A_84_48#_c_68_n N_VGND_c_366_n 0.0117056f $X=3.08 $Y=0.615 $X2=0 $Y2=0
cc_135 N_A_84_48#_c_72_n N_A_230_94#_c_400_n 0.00795851f $X=3.085 $Y=1.13 $X2=0
+ $Y2=0
cc_136 N_A_84_48#_c_68_n N_A_230_94#_c_402_n 0.019893f $X=3.08 $Y=0.615 $X2=0
+ $Y2=0
cc_137 N_A1_M1007_g N_A2_M1003_g 0.022073f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_138 N_A1_c_151_n N_A2_M1009_g 0.0757718f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_c_152_n N_A2_M1009_g 4.93984e-19 $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A1_c_151_n N_A2_c_192_n 0.0175581f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A1_c_152_n N_A2_c_192_n 0.00160123f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A1_M1007_g N_A2_c_193_n 2.93475e-19 $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_143 N_A1_c_151_n N_A2_c_193_n 8.38565e-19 $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A1_c_152_n N_A2_c_193_n 0.0320796f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_M1004_g X 6.43937e-19 $X=1.205 $Y=2.34 $X2=0 $Y2=0
cc_146 N_A1_M1004_g N_VPWR_c_321_n 0.00611549f $X=1.205 $Y=2.34 $X2=0 $Y2=0
cc_147 N_A1_M1004_g N_VPWR_c_323_n 0.0059286f $X=1.205 $Y=2.34 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_VPWR_c_320_n 0.00610055f $X=1.205 $Y=2.34 $X2=0 $Y2=0
cc_149 N_A1_M1007_g N_VGND_c_360_n 0.00744236f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_150 N_A1_M1007_g N_VGND_c_362_n 0.00485498f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_151 N_A1_M1007_g N_VGND_c_366_n 0.00514438f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_152 N_A1_M1007_g N_A_230_94#_c_399_n 0.00590569f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_153 N_A1_M1007_g N_A_230_94#_c_401_n 0.00247091f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_154 N_A1_c_151_n N_A_230_94#_c_401_n 0.00109337f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A1_c_152_n N_A_230_94#_c_401_n 0.0133988f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A2_M1003_g N_A3_M1000_g 0.0169838f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_157 N_A2_c_192_n N_A3_M1000_g 0.00168165f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_158 N_A2_c_193_n N_A3_M1000_g 2.86174e-19 $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_159 N_A2_M1009_g N_A3_c_226_n 0.0532073f $X=1.625 $Y=2.34 $X2=0 $Y2=0
cc_160 N_A2_c_192_n N_A3_c_226_n 0.0170634f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A2_c_193_n N_A3_c_226_n 0.00198873f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A2_c_192_n N_A3_c_227_n 9.75214e-19 $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_163 N_A2_c_193_n N_A3_c_227_n 0.0278487f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_164 N_A2_M1009_g N_VPWR_c_323_n 0.0059286f $X=1.625 $Y=2.34 $X2=0 $Y2=0
cc_165 N_A2_M1009_g N_VPWR_c_320_n 0.00610055f $X=1.625 $Y=2.34 $X2=0 $Y2=0
cc_166 N_A2_M1003_g N_VGND_c_361_n 0.0070805f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_167 N_A2_M1003_g N_VGND_c_362_n 0.00507111f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VGND_c_366_n 0.00514438f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_169 N_A2_M1003_g N_A_230_94#_c_399_n 0.00279704f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_170 N_A2_M1003_g N_A_230_94#_c_400_n 0.0163236f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_171 N_A2_c_192_n N_A_230_94#_c_400_n 0.00125621f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_172 N_A2_c_193_n N_A_230_94#_c_400_n 0.0249418f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_173 N_A3_M1002_g N_B1_M1005_g 0.019299f $X=2.135 $Y=2.34 $X2=0 $Y2=0
cc_174 N_A3_c_227_n N_B1_M1005_g 3.38956e-19 $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_175 N_A3_M1000_g N_B1_M1001_g 0.023509f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_176 N_A3_c_226_n N_B1_c_264_n 0.0206294f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A3_c_227_n N_B1_c_264_n 3.80681e-19 $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A3_M1002_g N_B1_c_265_n 2.6794e-19 $X=2.135 $Y=2.34 $X2=0 $Y2=0
cc_179 N_A3_c_226_n N_B1_c_265_n 0.00188197f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A3_c_227_n N_B1_c_265_n 0.0347534f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A3_M1002_g N_VPWR_c_322_n 0.00257616f $X=2.135 $Y=2.34 $X2=0 $Y2=0
cc_182 N_A3_M1002_g N_VPWR_c_323_n 0.0056753f $X=2.135 $Y=2.34 $X2=0 $Y2=0
cc_183 N_A3_M1002_g N_VPWR_c_320_n 0.00610055f $X=2.135 $Y=2.34 $X2=0 $Y2=0
cc_184 N_A3_M1000_g N_VGND_c_361_n 0.00716063f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_185 N_A3_M1000_g N_VGND_c_365_n 0.00507111f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_186 N_A3_M1000_g N_VGND_c_366_n 0.00514438f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_187 N_A3_M1000_g N_A_230_94#_c_400_n 0.0165716f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_188 N_A3_c_226_n N_A_230_94#_c_400_n 0.00118031f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A3_c_227_n N_A_230_94#_c_400_n 0.0202397f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A3_M1000_g N_A_230_94#_c_402_n 0.00275413f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_191 N_B1_M1005_g N_VPWR_c_322_n 0.0106618f $X=2.675 $Y=2.26 $X2=0 $Y2=0
cc_192 N_B1_M1005_g N_VPWR_c_323_n 0.00401533f $X=2.675 $Y=2.26 $X2=0 $Y2=0
cc_193 N_B1_M1005_g N_VPWR_c_320_n 0.00465661f $X=2.675 $Y=2.26 $X2=0 $Y2=0
cc_194 N_B1_M1001_g N_VGND_c_365_n 0.00485498f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_195 N_B1_M1001_g N_VGND_c_366_n 0.00514438f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_196 N_B1_M1001_g N_A_230_94#_c_400_n 0.00247983f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_197 N_B1_c_264_n N_A_230_94#_c_400_n 0.00101797f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_198 N_B1_c_265_n N_A_230_94#_c_400_n 0.0141977f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_199 N_B1_M1001_g N_A_230_94#_c_402_n 0.00594451f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_200 X N_VPWR_c_321_n 0.0271803f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_201 X N_VPWR_c_325_n 0.0163338f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_202 X N_VPWR_c_320_n 0.0134516f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_203 N_X_c_295_n N_VGND_c_360_n 0.0312028f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_204 N_X_c_295_n N_VGND_c_364_n 0.0159025f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_205 N_X_c_295_n N_VGND_c_366_n 0.0131064f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_206 N_VGND_c_360_n N_A_230_94#_c_399_n 0.0190445f $X=0.78 $Y=0.515 $X2=0
+ $Y2=0
cc_207 N_VGND_c_361_n N_A_230_94#_c_399_n 0.00929705f $X=1.945 $Y=0.615 $X2=0
+ $Y2=0
cc_208 N_VGND_c_362_n N_A_230_94#_c_399_n 0.0105078f $X=1.765 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_366_n N_A_230_94#_c_399_n 0.0115086f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_M1003_d N_A_230_94#_c_400_n 0.00923283f $X=1.655 $Y=0.47 $X2=0
+ $Y2=0
cc_211 N_VGND_c_361_n N_A_230_94#_c_400_n 0.0282971f $X=1.945 $Y=0.615 $X2=0
+ $Y2=0
cc_212 N_VGND_c_360_n N_A_230_94#_c_401_n 0.00760062f $X=0.78 $Y=0.515 $X2=0
+ $Y2=0
cc_213 N_VGND_c_361_n N_A_230_94#_c_402_n 0.00976671f $X=1.945 $Y=0.615 $X2=0
+ $Y2=0
cc_214 N_VGND_c_365_n N_A_230_94#_c_402_n 0.0103491f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_366_n N_A_230_94#_c_402_n 0.0113354f $X=3.12 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__xnor3_1.spice
* Created: Fri Aug 28 18:18:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xnor3_1.pex.spice"
.subckt sky130_fd_sc_ms__xnor3_1  VNB VPB C B A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_81_268#_M1003_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.24975 AS=0.2109 PD=1.90103 PS=2.05 NRD=45.804 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_232_162#_M1013_d N_C_M1013_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.1575 AS=0.14175 PD=1.59 PS=1.07897 NRD=0 NRS=80.712 M=1 R=2.8 SA=75000.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 N_A_81_268#_M1008_d N_C_M1008_g N_A_371_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1006 N_A_363_394#_M1006_d N_A_232_162#_M1006_g N_A_81_268#_M1008_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=6.552 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1001 N_A_786_100#_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.36 PD=2.05 PS=2.83 NRD=0 NRS=69.96 M=1 R=4.93333 SA=75000.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_371_74#_M1007_d N_A_786_100#_M1007_g N_A_897_54#_M1007_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1328 AS=0.374625 PD=1.055 PS=2.77 NRD=12.18 NRS=99.432 M=1
+ R=4.26667 SA=75000.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_1116_383#_M1004_d N_B_M1004_g N_A_371_74#_M1007_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.137177 AS=0.1328 PD=1.26792 PS=1.055 NRD=20.616 NRS=13.116 M=1
+ R=4.26667 SA=75000.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_363_394#_M1021_d N_A_786_100#_M1021_g N_A_1116_383#_M1004_d VNB
+ NLOWVT L=0.15 W=0.42 AD=0.0792057 AS=0.0900226 PD=0.780566 PS=0.832075
+ NRD=18.564 NRS=5.712 M=1 R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1014 N_A_897_54#_M1014_d N_B_M1014_g N_A_363_394#_M1021_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1104 AS=0.120694 PD=0.985 PS=1.18943 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A_M1017_g N_A_897_54#_M1014_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1376 AS=0.1104 PD=1.07 PS=0.985 NRD=20.616 NRS=0 M=1 R=4.26667 SA=75001.8
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_1116_383#_M1005_d N_A_897_54#_M1005_g N_VGND_M1017_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1376 PD=1.85 PS=1.07 NRD=0 NRS=7.488 M=1
+ R=4.26667 SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_A_81_268#_M1016_g N_X_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.289164 AS=0.3024 PD=2.06182 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1018 N_A_232_162#_M1018_d N_C_M1018_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.165236 PD=1.84 PS=1.17818 NRD=0 NRS=70.7821 M=1 R=3.55556
+ SA=90000.9 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1000 N_A_81_268#_M1000_d N_C_M1000_g N_A_363_394#_M1000_s VPB PSHORT L=0.18
+ W=0.84 AD=0.196375 AS=0.2352 PD=1.395 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1019 N_A_371_74#_M1019_d N_A_232_162#_M1019_g N_A_81_268#_M1000_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.231 AS=0.196375 PD=2.23 PS=1.395 NRD=0 NRS=17.5724 M=1
+ R=4.66667 SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1002 N_A_786_100#_M1002_d N_B_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.4026 PD=2.78 PS=3.05 NRD=0 NRS=13.1793 M=1 R=6.22222 SA=90000.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1009 N_A_363_394#_M1009_d N_A_786_100#_M1009_g N_A_897_54#_M1009_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.160735 AS=0.35325 PD=1.35649 PS=2.84 NRD=0 NRS=85.7147 M=1
+ R=4.66667 SA=90000.3 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1010 N_A_1116_383#_M1010_d N_B_M1010_g N_A_363_394#_M1009_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.122465 PD=0.91 PS=1.03351 NRD=0 NRS=24.6053 M=1
+ R=3.55556 SA=90000.8 SB=90002.4 A=0.1152 P=1.64 MULT=1
MM1012 N_A_371_74#_M1012_d N_A_786_100#_M1012_g N_A_1116_383#_M1010_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.150573 AS=0.0864 PD=1.12 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90001.2 SB=90001.9 A=0.1152 P=1.64 MULT=1
MM1015 N_A_897_54#_M1015_d N_B_M1015_g N_A_371_74#_M1012_d VPB PSHORT L=0.18
+ W=0.84 AD=0.157043 AS=0.197627 PD=1.24174 PS=1.47 NRD=18.7544 NRS=42.1974 M=1
+ R=4.66667 SA=90001.5 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_A_897_54#_M1015_d VPB PSHORT L=0.18 W=1
+ AD=0.1775 AS=0.186957 PD=1.355 PS=1.47826 NRD=15.7403 NRS=0 M=1 R=5.55556
+ SA=90001.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_A_1116_383#_M1011_d N_A_897_54#_M1011_g N_VPWR_M1020_d VPB PSHORT
+ L=0.18 W=1 AD=0.285 AS=0.1775 PD=2.57 PS=1.355 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90002.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__xnor3_1.pxi.spice"
*
.ends
*
*

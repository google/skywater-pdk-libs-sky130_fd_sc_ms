* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_136_392# C a_220_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VGND a_44_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND B a_44_392# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X3 a_220_392# B a_334_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 VPWR a_44_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_334_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 a_44_392# D a_136_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 a_44_392# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X8 VGND D a_44_392# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X9 a_44_392# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends

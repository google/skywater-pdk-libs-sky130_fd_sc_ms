* File: sky130_fd_sc_ms__a211o_1.pex.spice
* Created: Wed Sep  2 11:49:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A211O_1%A_81_264# 1 2 3 12 16 18 19 20 25 27 29 31
+ 35 40
c77 27 0 3.92783e-20 $X=3.125 $Y=1.18
c78 25 0 1.62677e-19 $X=2.28 $Y=1.195
c79 19 0 1.71301e-19 $X=1.13 $Y=1.485
r80 42 43 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.445 $Y=1.18
+ $X2=2.445 $Y2=1.195
r81 40 42 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.445 $Y=1.02
+ $X2=2.445 $Y2=1.18
r82 31 33 19.7165 $w=4.13e-07 $l=7.1e-07 $layer=LI1_cond $X=3.332 $Y=2.105
+ $X2=3.332 $Y2=2.815
r83 29 46 2.59301 $w=4.15e-07 $l=1e-07 $layer=LI1_cond $X=3.332 $Y=1.28
+ $X2=3.332 $Y2=1.18
r84 29 31 22.91 $w=4.13e-07 $l=8.25e-07 $layer=LI1_cond $X=3.332 $Y=1.28
+ $X2=3.332 $Y2=2.105
r85 28 42 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.18 $X2=2.445
+ $Y2=1.18
r86 27 46 5.36752 $w=2e-07 $l=2.07e-07 $layer=LI1_cond $X=3.125 $Y=1.18
+ $X2=3.332 $Y2=1.18
r87 27 28 28.5591 $w=1.98e-07 $l=5.15e-07 $layer=LI1_cond $X=3.125 $Y=1.18
+ $X2=2.61 $Y2=1.18
r88 26 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=1.195
+ $X2=1.33 $Y2=1.195
r89 25 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=1.195
+ $X2=2.445 $Y2=1.195
r90 25 26 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.28 $Y=1.195
+ $X2=1.415 $Y2=1.195
r91 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.115
+ $Y=1.485 $X2=1.115 $Y2=1.485
r92 20 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.33 $Y=1.525
+ $X2=1.33 $Y2=1.195
r93 20 22 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.245 $Y=1.525
+ $X2=1.115 $Y2=1.525
r94 19 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.13 $Y=1.485
+ $X2=1.115 $Y2=1.485
r95 18 23 92.6765 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=0.585 $Y=1.485
+ $X2=1.115 $Y2=1.485
r96 14 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.205 $Y=1.32
+ $X2=1.13 $Y2=1.485
r97 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.205 $Y=1.32
+ $X2=1.205 $Y2=0.74
r98 10 18 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.495 $Y=1.65
+ $X2=0.585 $Y2=1.485
r99 10 12 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.495 $Y=1.65
+ $X2=0.495 $Y2=2.4
r100 3 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.96 $X2=3.29 $Y2=2.815
r101 3 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=1.96 $X2=3.29 $Y2=2.105
r102 2 46 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.68 $X2=3.375 $Y2=1.17
r103 1 40 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.68 $X2=2.445 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%A2 3 7 9 12
c35 9 0 1.71301e-19 $X=1.68 $Y=1.665
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.615
+ $X2=1.67 $Y2=1.78
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.615
+ $X2=1.67 $Y2=1.45
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.615 $X2=1.67 $Y2=1.615
r39 7 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.755 $Y=1 $X2=1.755
+ $Y2=1.45
r40 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.745 $Y=2.46
+ $X2=1.745 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%A1 3 7 9 10 14
c42 7 0 3.92783e-20 $X=2.23 $Y=1
r43 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.615
+ $X2=2.21 $Y2=1.78
r44 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.615
+ $X2=2.21 $Y2=1.45
r45 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=2.64 $Y2=1.615
r46 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.615 $X2=2.21 $Y2=1.615
r47 7 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.23 $Y=1 $X2=2.23
+ $Y2=1.45
r48 3 17 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.225 $Y=2.46
+ $X2=2.225 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%B1 4 5 7 12 13 15 23
c43 12 0 1.23467e-19 $X=2.71 $Y=0.405
c44 4 0 3.92096e-20 $X=2.66 $Y=1
r45 15 23 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=2.275 $Y2=0.462
r46 13 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.405
+ $X2=2.71 $Y2=0.57
r47 12 23 15.9147 $w=3.13e-07 $l=4.35e-07 $layer=LI1_cond $X=2.71 $Y=0.412
+ $X2=2.275 $Y2=0.412
r48 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=0.405 $X2=2.71 $Y2=0.405
r49 5 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.675 $Y=1.485 $X2=2.675
+ $Y2=1.395
r50 5 7 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=2.675 $Y=1.485
+ $X2=2.675 $Y2=2.46
r51 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.66 $Y=1 $X2=2.66
+ $Y2=1.395
r52 4 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.66 $Y=1 $X2=2.66
+ $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%C1 3 8 10 11 12 15 16
r35 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=0.405 $X2=3.55 $Y2=0.405
r36 12 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.55 $Y=0.555
+ $X2=3.55 $Y2=0.405
r37 11 15 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=3.235 $Y=0.405
+ $X2=3.55 $Y2=0.405
r38 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.105 $Y=1.395
+ $X2=3.105 $Y2=1.545
r39 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.16 $Y=1 $X2=3.16
+ $Y2=1.395
r40 5 11 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.16 $Y=0.57
+ $X2=3.235 $Y2=0.405
r41 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.16 $Y=0.57 $X2=3.16
+ $Y2=1
r42 3 10 355.669 $w=1.8e-07 $l=9.15e-07 $layer=POLY_cond $X=3.065 $Y=2.46
+ $X2=3.065 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%X 1 2 9 12 13 14 21 30
r20 19 21 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.26 $Y=1.995 $X2=0.26
+ $Y2=2.035
r21 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r22 12 19 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.995
r23 12 30 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=0.26 $Y=1.972
+ $X2=0.26 $Y2=1.82
r24 12 13 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.405
r25 12 21 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.26 $Y=2.057
+ $X2=0.26 $Y2=2.035
r26 9 11 13.9526 $w=7.17e-07 $l=8.2e-07 $layer=LI1_cond $X=0.17 $Y=0.737
+ $X2=0.99 $Y2=0.737
r27 7 9 9.47984 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=0.737
r28 7 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r29 2 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r30 2 14 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r31 1 11 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.865
+ $Y=0.37 $X2=0.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r41 33 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 30 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 27 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.76 $Y2=3.33
r47 27 29 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 22 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.76 $Y2=3.33
r51 22 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 20 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 18 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 18 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.885 $Y=3.33 $X2=1.985
+ $Y2=3.33
r56 17 32 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 17 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.085 $Y=3.33 $X2=1.985
+ $Y2=3.33
r58 13 19 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=3.33
r59 13 15 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=2.455
r60 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.76 $Y=1.985
+ $X2=0.76 $Y2=2.815
r61 7 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r62 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=2.815
r63 2 15 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=1.835
+ $Y=1.96 $X2=1.985 $Y2=2.455
r64 1 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.815
r65 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%A_279_392# 1 2 7 9 11 13 15
r39 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=2.12 $X2=2.45
+ $Y2=2.035
r40 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.45 $Y=2.12
+ $X2=2.45 $Y2=2.815
r41 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.035
+ $X2=1.52 $Y2=2.035
r42 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=2.035
+ $X2=2.45 $Y2=2.035
r43 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.285 $Y=2.035
+ $X2=1.685 $Y2=2.035
r44 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.12 $X2=1.52
+ $Y2=2.035
r45 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.52 $Y=2.12 $X2=1.52
+ $Y2=2.815
r46 2 20 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.96 $X2=2.45 $Y2=2.115
r47 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.96 $X2=2.45 $Y2=2.815
r48 1 18 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.115
r49 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.96 $X2=1.52 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_1%VGND 1 2 9 13 16 20 22 24 34 35 38 41
r46 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r49 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 32 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.13
+ $Y2=0
r51 32 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r52 31 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r53 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 27 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r55 26 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r56 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 24 38 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.48
+ $Y2=0
r58 24 30 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r59 22 42 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r60 22 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r61 18 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.945 $Y=0.825
+ $X2=3.13 $Y2=0.825
r62 16 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.74
+ $X2=3.13 $Y2=0.825
r63 15 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r64 15 16 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.74
r65 14 38 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.48
+ $Y2=0
r66 13 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.13
+ $Y2=0
r67 13 14 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=1.705 $Y2=0
r68 9 11 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.48 $Y=0.495
+ $X2=1.48 $Y2=0.835
r69 7 38 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=0.085 $X2=1.48
+ $Y2=0
r70 7 9 10.8976 $w=4.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.48 $Y=0.085 $X2=1.48
+ $Y2=0.495
r71 2 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.68 $X2=2.945 $Y2=0.825
r72 1 11 182 $w=1.7e-07 $l=5.80625e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.37 $X2=1.54 $Y2=0.835
r73 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.28
+ $Y=0.37 $X2=1.42 $Y2=0.495
.ends


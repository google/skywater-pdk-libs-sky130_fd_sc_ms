* NGSPICE file created from sky130_fd_sc_ms__o311a_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_219_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.958e+11p pd=4.3e+06u as=1.1042e+12p ps=7.58e+06u
M1001 a_135_74# C1 a_32_74# VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=2.701e+11p ps=2.21e+06u
M1002 VGND A3 a_219_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_447_368# A2 a_363_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=2.688e+11p ps=2.72e+06u
M1004 VPWR A1 a_447_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.2132e+12p pd=8.73e+06u as=0p ps=0u
M1005 X a_32_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1006 a_32_74# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=6.736e+11p pd=5.52e+06u as=0p ps=0u
M1007 VPWR C1 a_32_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A1 a_219_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_32_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_363_368# A3 a_32_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_32_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1012 VPWR a_32_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_219_74# B1 a_135_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


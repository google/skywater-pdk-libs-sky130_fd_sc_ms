* File: sky130_fd_sc_ms__a21bo_1.pex.spice
* Created: Wed Sep  2 11:50:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21BO_1%A2 1 3 8 10 11 15
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.405 $X2=0.27 $Y2=0.405
r31 11 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.405
r32 10 14 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.46 $Y=0.405
+ $X2=0.27 $Y2=0.405
r33 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.535 $Y=1 $X2=0.535
+ $Y2=1.395
r34 5 10 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.535 $Y=0.57
+ $X2=0.46 $Y2=0.405
r35 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.535 $Y=0.57
+ $X2=0.535 $Y2=1
r36 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.485 $X2=0.52
+ $Y2=1.395
r37 1 3 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=0.52 $Y=1.485
+ $X2=0.52 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%A1 3 7 9 12
c37 12 0 6.82625e-20 $X=0.985 $Y=1.615
c38 7 0 4.71918e-20 $X=1 $Y=2.46
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.615
+ $X2=0.985 $Y2=1.78
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.615
+ $X2=0.985 $Y2=1.45
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.615 $X2=0.985 $Y2=1.615
r42 9 13 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=0.985 $Y2=1.615
r43 7 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1 $Y=2.46 $X2=1
+ $Y2=1.78
r44 3 14 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.895 $Y=1 $X2=0.895
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%A_272_110# 1 2 7 9 12 14 16 18 20 21 26 28
+ 33
r65 30 33 8.00764 $w=5.88e-07 $l=3.95e-07 $layer=LI1_cond $X=2.16 $Y=0.645
+ $X2=2.555 $Y2=0.645
r66 24 29 0.0912679 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=1.945
+ $X2=2.08 $Y2=1.945
r67 24 26 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=1.945
+ $X2=2.53 $Y2=1.945
r68 22 30 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.16 $Y=0.94
+ $X2=2.16 $Y2=0.645
r69 22 28 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=0.94
+ $X2=2.16 $Y2=1.1
r70 21 37 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.08 $Y=1.265
+ $X2=2.08 $Y2=1.47
r71 20 28 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=1.265
+ $X2=2.08 $Y2=1.1
r72 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.08
+ $Y=1.265 $X2=2.08 $Y2=1.265
r73 18 29 13.7904 $w=3.3e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=1.605
+ $X2=2.08 $Y2=1.945
r74 18 20 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=1.605
+ $X2=2.08 $Y2=1.265
r75 15 16 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.54 $Y=1.47 $X2=1.45
+ $Y2=1.47
r76 14 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.47
+ $X2=2.08 $Y2=1.47
r77 14 15 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.915 $Y=1.47
+ $X2=1.54 $Y2=1.47
r78 10 16 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.545
+ $X2=1.45 $Y2=1.47
r79 10 12 355.669 $w=1.8e-07 $l=9.15e-07 $layer=POLY_cond $X=1.45 $Y=1.545
+ $X2=1.45 $Y2=2.46
r80 7 16 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.435 $Y=1.395
+ $X2=1.45 $Y2=1.47
r81 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.435 $Y=1.395
+ $X2=1.435 $Y2=1
r82 2 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.84 $X2=2.53 $Y2=1.985
r83 1 33 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.37 $X2=2.555 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%B1_N 3 7 9 12
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.55
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.22
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.385 $X2=2.68 $Y2=1.385
r39 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.68 $Y=1.295 $X2=2.68
+ $Y2=1.385
r40 7 14 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.77 $Y=0.645
+ $X2=2.77 $Y2=1.22
r41 3 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=2.755 $Y=2.26
+ $X2=2.755 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%A_194_136# 1 2 9 13 17 19 20 23 29 31 34 35
+ 38 39
c84 39 0 1.9051e-19 $X=3.25 $Y=1.485
c85 35 0 6.82625e-20 $X=1.667 $Y=1.94
c86 34 0 9.10919e-20 $X=3.17 $Y=2.24
r87 39 44 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.485
+ $X2=3.25 $Y2=1.65
r88 39 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.485
+ $X2=3.25 $Y2=1.32
r89 38 41 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=1.485
+ $X2=3.25 $Y2=1.65
r90 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.485 $X2=3.25 $Y2=1.485
r91 34 41 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.17 $Y=2.24 $X2=3.17
+ $Y2=1.65
r92 32 36 1.64875 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=1.76 $Y=2.325
+ $X2=1.667 $Y2=2.325
r93 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=2.325
+ $X2=3.17 $Y2=2.24
r94 31 32 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.085 $Y=2.325
+ $X2=1.76 $Y2=2.325
r95 27 36 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.667 $Y=2.41
+ $X2=1.667 $Y2=2.325
r96 27 29 2.99754 $w=1.83e-07 $l=5e-08 $layer=LI1_cond $X=1.667 $Y=2.41
+ $X2=1.667 $Y2=2.46
r97 24 36 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.667 $Y=2.24
+ $X2=1.667 $Y2=2.325
r98 24 26 8.09337 $w=1.83e-07 $l=1.35e-07 $layer=LI1_cond $X=1.667 $Y=2.24
+ $X2=1.667 $Y2=2.105
r99 23 35 5.60801 $w=1.83e-07 $l=9.2e-08 $layer=LI1_cond $X=1.667 $Y=2.032
+ $X2=1.667 $Y2=1.94
r100 23 26 4.37641 $w=1.83e-07 $l=7.3e-08 $layer=LI1_cond $X=1.667 $Y=2.032
+ $X2=1.667 $Y2=2.105
r101 21 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.66 $Y=1.28
+ $X2=1.66 $Y2=1.94
r102 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.575 $Y=1.195
+ $X2=1.66 $Y2=1.28
r103 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.575 $Y=1.195
+ $X2=1.315 $Y2=1.195
r104 15 20 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.13 $Y=1.11
+ $X2=1.315 $Y2=1.195
r105 15 17 9.49987 $w=3.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.13 $Y=1.11
+ $X2=1.13 $Y2=0.805
r106 13 44 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.29 $Y=2.4
+ $X2=3.29 $Y2=1.65
r107 9 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.245 $Y=0.74
+ $X2=3.245 $Y2=1.32
r108 2 29 300 $w=1.7e-07 $l=5.63471e-07 $layer=licon1_PDIFF $count=2 $X=1.54
+ $Y=1.96 $X2=1.675 $Y2=2.46
r109 2 26 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.96 $X2=1.675 $Y2=2.105
r110 1 17 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.97
+ $Y=0.68 $X2=1.13 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%A_34_392# 1 2 7 9 11 13 15
c32 7 0 4.71918e-20 $X=0.295 $Y=2.12
r33 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.12
+ $X2=1.225 $Y2=2.035
r34 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.225 $Y=2.12
+ $X2=1.225 $Y2=2.815
r35 12 18 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.46 $Y=2.035
+ $X2=0.295 $Y2=2.03
r36 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=2.035
+ $X2=1.225 $Y2=2.035
r37 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.06 $Y=2.035 $X2=0.46
+ $Y2=2.035
r38 7 18 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.295 $Y=2.12 $X2=0.295
+ $Y2=2.03
r39 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.295 $Y=2.12
+ $X2=0.295 $Y2=2.815
r40 2 20 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.96 $X2=1.225 $Y2=2.115
r41 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.96 $X2=1.225 $Y2=2.815
r42 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.96 $X2=0.295 $Y2=2.105
r43 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.96 $X2=0.295 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%VPWR 1 2 11 15 17 19 29 30 33 36
r38 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=3.33
+ $X2=3.065 $Y2=3.33
r43 27 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.23 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 20 33 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.86 $Y=3.33 $X2=0.76
+ $Y2=3.33
r50 20 22 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=3.065 $Y2=3.33
r52 19 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=2.64
+ $Y2=3.33
r53 17 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=3.33
r56 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=2.745
r57 9 33 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=3.33
r58 9 11 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.455
r59 2 15 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=3.065 $Y2=2.745
r60 1 11 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.96 $X2=0.76 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%X 1 2 9 13 14 15 16 24 33
r25 21 24 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=3.592 $Y=1.982
+ $X2=3.592 $Y2=1.985
r26 15 16 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=3.592 $Y=2.405
+ $X2=3.592 $Y2=2.775
r27 14 21 0.567357 $w=3.23e-07 $l=1.6e-08 $layer=LI1_cond $X=3.592 $Y=1.966
+ $X2=3.592 $Y2=1.982
r28 14 33 7.78643 $w=3.23e-07 $l=1.46e-07 $layer=LI1_cond $X=3.592 $Y=1.966
+ $X2=3.592 $Y2=1.82
r29 14 15 12.5528 $w=3.23e-07 $l=3.54e-07 $layer=LI1_cond $X=3.592 $Y=2.051
+ $X2=3.592 $Y2=2.405
r30 14 24 2.34035 $w=3.23e-07 $l=6.6e-08 $layer=LI1_cond $X=3.592 $Y=2.051
+ $X2=3.592 $Y2=1.985
r31 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.13 $X2=3.67
+ $Y2=1.82
r32 7 13 10.9702 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=3.525 $Y=0.9
+ $X2=3.525 $Y2=1.13
r33 7 9 10.0107 $w=4.58e-07 $l=3.85e-07 $layer=LI1_cond $X=3.525 $Y=0.9
+ $X2=3.525 $Y2=0.515
r34 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.515 $Y2=2.815
r35 2 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.515 $Y2=1.985
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.32
+ $Y=0.37 $X2=3.46 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_1%VGND 1 2 3 11 14 18 21 24 25 27 28 29 35 44
+ 45 48
c59 18 0 1.9051e-19 $X=3.005 $Y=0.665
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r63 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.65
+ $Y2=0
r65 39 41 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.64
+ $Y2=0
r66 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r67 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.65
+ $Y2=0
r69 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.2
+ $Y2=0
r70 33 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r71 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 29 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r73 29 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r74 27 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.64
+ $Y2=0
r75 27 28 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.007
+ $Y2=0
r76 26 44 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.6
+ $Y2=0
r77 26 28 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.007
+ $Y2=0
r78 24 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r79 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.69
+ $Y2=0
r80 23 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=1.2
+ $Y2=0
r81 23 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.69
+ $Y2=0
r82 21 22 11.7247 $w=3.85e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.09
+ $X2=0.69 $Y2=1.09
r83 16 28 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.007 $Y=0.085
+ $X2=3.007 $Y2=0
r84 16 18 31.0892 $w=2.13e-07 $l=5.8e-07 $layer=LI1_cond $X=3.007 $Y=0.085
+ $X2=3.007 $Y2=0.665
r85 12 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0
r86 12 14 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0.835
r87 11 22 5.54671 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=0.84 $X2=0.69
+ $Y2=1.09
r88 10 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r89 10 11 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.84
r90 3 18 182 $w=1.7e-07 $l=3.66367e-07 $layer=licon1_NDIFF $count=1 $X=2.845
+ $Y=0.37 $X2=3.005 $Y2=0.665
r91 2 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.68 $X2=1.65 $Y2=0.835
r92 1 21 182 $w=1.7e-07 $l=4.68348e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.68 $X2=0.32 $Y2=1.09
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__nor4b_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__nor4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.350000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.350000 1.855000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.395000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.110000 0.815000 1.440000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.862400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.290000 0.350000 1.620000 1.010000 ;
        RECT 1.290000 1.010000 3.275000 1.180000 ;
        RECT 2.300000 0.350000 2.630000 1.010000 ;
        RECT 2.905000 1.850000 3.275000 2.980000 ;
        RECT 3.105000 1.180000 3.275000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
        RECT 0.790000  0.085000 1.120000 0.940000 ;
        RECT 1.790000  0.085000 2.120000 0.840000 ;
        RECT 2.800000  0.085000 3.130000 0.840000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.360000 3.415000 ;
        RECT 0.835000 2.290000 1.165000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105000 0.350000 0.620000 0.940000 ;
      RECT 0.105000 0.940000 0.275000 1.820000 ;
      RECT 0.105000 1.820000 0.595000 1.950000 ;
      RECT 0.105000 1.950000 2.735000 2.120000 ;
      RECT 0.105000 2.120000 0.595000 2.700000 ;
      RECT 2.565000 1.350000 2.935000 1.680000 ;
      RECT 2.565000 1.680000 2.735000 1.950000 ;
  END
END sky130_fd_sc_ms__nor4b_1

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a221o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__a221o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.255000 1.765000 0.565000 ;
        RECT 1.595000 0.565000 1.765000 1.040000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 0.255000 2.755000 0.505000 ;
        RECT 2.525000 0.505000 2.755000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.615000 1.300000 9.495000 1.750000 ;
        RECT 9.095000 1.210000 9.495000 1.300000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.470000 0.255000 7.045000 0.505000 ;
        RECT 6.845000 0.505000 7.045000 0.670000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.470000 5.735000 2.150000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.355000 1.920000 ;
        RECT 0.125000 1.920000 4.525000 2.090000 ;
        RECT 2.850000 2.090000 4.525000 2.190000 ;
        RECT 3.005000 1.010000 4.540000 1.180000 ;
        RECT 3.005000 1.180000 3.235000 1.410000 ;
        RECT 3.430000 0.440000 3.760000 1.010000 ;
        RECT 4.290000 0.480000 4.540000 1.010000 ;
      LAYER mcon ;
        RECT 0.155000 1.210000 0.325000 1.380000 ;
        RECT 3.035000 1.210000 3.205000 1.380000 ;
      LAYER met1 ;
        RECT 0.095000 1.180000 0.385000 1.225000 ;
        RECT 0.095000 1.225000 3.265000 1.365000 ;
        RECT 0.095000 1.365000 0.385000 1.410000 ;
        RECT 2.975000 1.180000 3.265000 1.225000 ;
        RECT 2.975000 1.365000 3.265000 1.410000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
        RECT 1.935000  0.085000 2.105000 0.675000 ;
        RECT 1.935000  0.675000 2.330000 1.070000 ;
        RECT 3.000000  0.085000 3.250000 0.840000 ;
        RECT 3.940000  0.085000 4.110000 0.840000 ;
        RECT 4.720000  0.085000 5.440000 0.960000 ;
        RECT 6.130000  0.085000 6.300000 0.675000 ;
        RECT 6.130000  0.675000 6.525000 0.960000 ;
        RECT 6.275000  0.960000 6.525000 1.280000 ;
        RECT 7.215000  0.085000 7.465000 1.090000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.600000 3.415000 ;
        RECT 0.320000 2.260000 0.650000 3.245000 ;
        RECT 1.395000 2.600000 2.065000 3.245000 ;
        RECT 2.845000 2.700000 3.175000 3.245000 ;
        RECT 3.745000 2.700000 4.075000 3.245000 ;
        RECT 4.645000 2.700000 4.975000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.315000 0.655000 0.565000 0.735000 ;
      RECT 0.315000 0.735000 1.425000 0.905000 ;
      RECT 0.315000 0.905000 0.565000 1.010000 ;
      RECT 0.745000 1.075000 1.075000 1.580000 ;
      RECT 0.745000 1.580000 4.880000 1.750000 ;
      RECT 0.890000 2.260000 2.565000 2.360000 ;
      RECT 0.890000 2.360000 7.150000 2.430000 ;
      RECT 0.890000 2.430000 1.220000 2.900000 ;
      RECT 1.255000 0.905000 1.425000 1.240000 ;
      RECT 1.255000 1.240000 2.760000 1.410000 ;
      RECT 2.235000 2.430000 7.150000 2.530000 ;
      RECT 2.235000 2.530000 2.565000 2.900000 ;
      RECT 2.510000 0.840000 2.760000 1.240000 ;
      RECT 3.595000 1.350000 4.880000 1.580000 ;
      RECT 4.710000 1.130000 6.090000 1.300000 ;
      RECT 4.710000 1.300000 4.880000 1.350000 ;
      RECT 5.470000 2.700000 6.700000 2.905000 ;
      RECT 5.470000 2.905000 8.830000 3.075000 ;
      RECT 5.610000 0.580000 5.940000 1.130000 ;
      RECT 5.920000 1.300000 6.090000 1.600000 ;
      RECT 5.920000 1.600000 8.445000 1.770000 ;
      RECT 5.920000 1.770000 6.250000 2.190000 ;
      RECT 6.705000 0.840000 7.035000 1.260000 ;
      RECT 6.705000 1.260000 7.935000 1.430000 ;
      RECT 6.820000 1.940000 8.380000 2.110000 ;
      RECT 6.820000 2.110000 7.150000 2.360000 ;
      RECT 6.870000 2.530000 7.150000 2.735000 ;
      RECT 7.425000 2.280000 7.755000 2.905000 ;
      RECT 7.685000 0.255000 8.925000 0.425000 ;
      RECT 7.685000 0.425000 7.935000 1.260000 ;
      RECT 8.010000 2.110000 8.380000 2.735000 ;
      RECT 8.115000 0.595000 8.445000 1.600000 ;
      RECT 8.580000 1.940000 8.830000 2.905000 ;
      RECT 8.625000 0.425000 8.925000 1.040000 ;
  END
END sky130_fd_sc_ms__a221o_4

* File: sky130_fd_sc_ms__o2111ai_2.pxi.spice
* Created: Fri Aug 28 17:52:06 2020
* 
x_PM_SKY130_FD_SC_MS__O2111AI_2%D1 N_D1_M1011_g N_D1_c_103_n N_D1_M1014_g
+ N_D1_M1012_g N_D1_c_105_n N_D1_M1016_g N_D1_c_106_n N_D1_c_107_n D1
+ PM_SKY130_FD_SC_MS__O2111AI_2%D1
x_PM_SKY130_FD_SC_MS__O2111AI_2%C1 N_C1_M1001_g N_C1_M1013_g N_C1_M1002_g
+ N_C1_M1015_g C1 N_C1_c_155_n PM_SKY130_FD_SC_MS__O2111AI_2%C1
x_PM_SKY130_FD_SC_MS__O2111AI_2%B1 N_B1_M1017_g N_B1_c_211_n N_B1_c_212_n
+ N_B1_M1018_g N_B1_M1007_g N_B1_M1009_g N_B1_c_215_n N_B1_c_216_n B1 B1 B1
+ PM_SKY130_FD_SC_MS__O2111AI_2%B1
x_PM_SKY130_FD_SC_MS__O2111AI_2%A2 N_A2_M1000_g N_A2_M1003_g N_A2_M1019_g
+ N_A2_M1005_g A2 A2 N_A2_c_277_n PM_SKY130_FD_SC_MS__O2111AI_2%A2
x_PM_SKY130_FD_SC_MS__O2111AI_2%A1 N_A1_M1004_g N_A1_M1006_g N_A1_M1010_g
+ N_A1_M1008_g A1 A1 N_A1_c_325_n PM_SKY130_FD_SC_MS__O2111AI_2%A1
x_PM_SKY130_FD_SC_MS__O2111AI_2%VPWR N_VPWR_M1011_s N_VPWR_M1012_s
+ N_VPWR_M1015_s N_VPWR_M1018_s N_VPWR_M1006_d N_VPWR_c_368_n N_VPWR_c_369_n
+ N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n
+ VPWR N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n
+ N_VPWR_c_367_n N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n
+ PM_SKY130_FD_SC_MS__O2111AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O2111AI_2%Y N_Y_M1014_s N_Y_M1011_d N_Y_M1013_d
+ N_Y_M1017_d N_Y_M1003_d N_Y_c_453_n N_Y_c_447_n N_Y_c_448_n N_Y_c_473_n
+ N_Y_c_449_n N_Y_c_450_n N_Y_c_451_n N_Y_c_493_n N_Y_c_498_n Y Y Y Y Y
+ N_Y_c_446_n Y Y PM_SKY130_FD_SC_MS__O2111AI_2%Y
x_PM_SKY130_FD_SC_MS__O2111AI_2%A_697_368# N_A_697_368#_M1003_s
+ N_A_697_368#_M1005_s N_A_697_368#_M1008_s N_A_697_368#_c_529_n
+ N_A_697_368#_c_530_n N_A_697_368#_c_531_n N_A_697_368#_c_536_n
+ N_A_697_368#_c_537_n N_A_697_368#_c_532_n N_A_697_368#_c_533_n
+ PM_SKY130_FD_SC_MS__O2111AI_2%A_697_368#
x_PM_SKY130_FD_SC_MS__O2111AI_2%A_40_74# N_A_40_74#_M1014_d N_A_40_74#_M1016_d
+ N_A_40_74#_M1002_d N_A_40_74#_c_564_n N_A_40_74#_c_565_n N_A_40_74#_c_566_n
+ N_A_40_74#_c_567_n N_A_40_74#_c_568_n N_A_40_74#_c_582_n
+ PM_SKY130_FD_SC_MS__O2111AI_2%A_40_74#
x_PM_SKY130_FD_SC_MS__O2111AI_2%A_299_74# N_A_299_74#_M1001_s
+ N_A_299_74#_M1007_s N_A_299_74#_c_604_n N_A_299_74#_c_611_n
+ N_A_299_74#_c_605_n PM_SKY130_FD_SC_MS__O2111AI_2%A_299_74#
x_PM_SKY130_FD_SC_MS__O2111AI_2%A_510_74# N_A_510_74#_M1007_d
+ N_A_510_74#_M1009_d N_A_510_74#_M1019_d N_A_510_74#_M1010_d
+ N_A_510_74#_c_630_n N_A_510_74#_c_631_n N_A_510_74#_c_632_n
+ N_A_510_74#_c_633_n N_A_510_74#_c_634_n N_A_510_74#_c_635_n
+ N_A_510_74#_c_636_n N_A_510_74#_c_637_n N_A_510_74#_c_638_n
+ N_A_510_74#_c_639_n PM_SKY130_FD_SC_MS__O2111AI_2%A_510_74#
x_PM_SKY130_FD_SC_MS__O2111AI_2%VGND N_VGND_M1000_s N_VGND_M1004_s
+ N_VGND_c_693_n N_VGND_c_694_n VGND N_VGND_c_695_n N_VGND_c_696_n
+ N_VGND_c_697_n N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n
+ PM_SKY130_FD_SC_MS__O2111AI_2%VGND
cc_1 VNB N_D1_M1011_g 0.00871317f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_2 VNB N_D1_c_103_n 0.0204008f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.22
cc_3 VNB N_D1_M1012_g 0.00555556f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_4 VNB N_D1_c_105_n 0.0159551f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_5 VNB N_D1_c_106_n 0.0507325f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_6 VNB N_D1_c_107_n 0.0357086f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.385
cc_7 VNB D1 0.0126727f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_C1_M1001_g 0.0219968f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_9 VNB N_C1_M1013_g 0.00164866f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_10 VNB N_C1_M1002_g 0.0275487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C1_M1015_g 0.00159486f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_12 VNB C1 0.00888795f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.385
cc_13 VNB N_C1_c_155_n 0.0491382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_211_n 0.0123976f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.22
cc_15 VNB N_B1_c_212_n 0.0149711f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_16 VNB N_B1_M1007_g 0.0314339f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.74
cc_17 VNB N_B1_M1009_g 0.024203f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.385
cc_18 VNB N_B1_c_215_n 0.0142667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_216_n 0.024603f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB B1 0.00931452f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_21 VNB N_A2_M1000_g 0.0232975f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_22 VNB N_A2_M1019_g 0.0232975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB A2 0.00232957f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.385
cc_24 VNB N_A2_c_277_n 0.0343868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_M1004_g 0.0245199f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_26 VNB N_A1_M1010_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A1 0.0161791f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.385
cc_28 VNB N_A1_c_325_n 0.045324f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_29 VNB N_VPWR_c_367_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_446_n 0.00289639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_40_74#_c_564_n 0.0222939f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_32 VNB N_A_40_74#_c_565_n 0.00448726f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.74
cc_33 VNB N_A_40_74#_c_566_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_34 VNB N_A_40_74#_c_567_n 0.00325f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.385
cc_35 VNB N_A_40_74#_c_568_n 0.0157968f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_36 VNB N_A_299_74#_c_604_n 0.0199129f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_37 VNB N_A_299_74#_c_605_n 0.00240543f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.74
cc_38 VNB N_A_510_74#_c_630_n 0.00380647f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_39 VNB N_A_510_74#_c_631_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.385
cc_40 VNB N_A_510_74#_c_632_n 0.00417749f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.385
cc_41 VNB N_A_510_74#_c_633_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_42 VNB N_A_510_74#_c_634_n 0.00575126f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_43 VNB N_A_510_74#_c_635_n 0.00207041f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_44 VNB N_A_510_74#_c_636_n 0.0148256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_510_74#_c_637_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_510_74#_c_638_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_510_74#_c_639_n 0.00211286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_693_n 0.00335558f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_49 VNB N_VGND_c_694_n 0.00562151f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.74
cc_50 VNB N_VGND_c_695_n 0.095433f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.385
cc_51 VNB N_VGND_c_696_n 0.0175706f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_52 VNB N_VGND_c_697_n 0.0188229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_698_n 0.32741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_699_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_700_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_D1_M1011_g 0.0274077f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_57 VPB N_D1_M1012_g 0.0225188f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_58 VPB N_C1_M1013_g 0.0230883f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_59 VPB N_C1_M1015_g 0.0227912f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.385
cc_60 VPB N_B1_M1017_g 0.0218051f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_61 VPB N_B1_c_211_n 0.00314639f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.22
cc_62 VPB N_B1_c_212_n 7.74996e-19 $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_63 VPB N_B1_M1018_g 0.0246451f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_64 VPB N_B1_c_215_n 0.00191514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B1_c_216_n 0.0155439f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_66 VPB B1 0.0114786f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_67 VPB N_A2_M1003_g 0.0247875f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_68 VPB N_A2_M1005_g 0.0197873f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.385
cc_69 VPB A2 0.00696541f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.385
cc_70 VPB N_A2_c_277_n 0.00456027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A1_M1006_g 0.0218877f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_72 VPB N_A1_M1008_g 0.0281514f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.385
cc_73 VPB A1 0.0107587f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.385
cc_74 VPB N_A1_c_325_n 0.0127586f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_75 VPB N_VPWR_c_368_n 0.011928f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.385
cc_76 VPB N_VPWR_c_369_n 0.0563264f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.385
cc_77 VPB N_VPWR_c_370_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_78 VPB N_VPWR_c_371_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_372_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_80 VPB N_VPWR_c_373_n 0.0148873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_374_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_375_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_376_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_377_n 0.0389588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_378_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_367_n 0.0846271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_380_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_381_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_382_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_383_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_Y_c_447_n 0.00630481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_Y_c_448_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_93 VPB N_Y_c_449_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_94 VPB N_Y_c_450_n 0.0117034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_Y_c_451_n 0.00223855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB Y 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_697_368#_c_529_n 0.00554152f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.22
cc_98 VPB N_A_697_368#_c_530_n 0.00473643f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=0.74
cc_99 VPB N_A_697_368#_c_531_n 0.00376758f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.385
cc_100 VPB N_A_697_368#_c_532_n 0.0075506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_697_368#_c_533_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_102 N_D1_c_105_n N_C1_M1001_g 0.0120716f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_103 N_D1_c_107_n N_C1_M1001_g 0.0103282f $X=0.995 $Y=1.385 $X2=0 $Y2=0
cc_104 N_D1_M1012_g N_C1_M1013_g 0.0259151f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_105 N_D1_c_107_n C1 0.00147127f $X=0.995 $Y=1.385 $X2=0 $Y2=0
cc_106 N_D1_M1012_g N_C1_c_155_n 0.0103282f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_107 N_D1_M1011_g N_VPWR_c_369_n 0.00649184f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_108 N_D1_c_106_n N_VPWR_c_369_n 0.00185549f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_109 D1 N_VPWR_c_369_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_110 N_D1_M1012_g N_VPWR_c_370_n 0.0038215f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_111 N_D1_M1011_g N_VPWR_c_375_n 0.005209f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_112 N_D1_M1012_g N_VPWR_c_375_n 0.005209f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_113 N_D1_M1011_g N_VPWR_c_367_n 0.00986139f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_114 N_D1_M1012_g N_VPWR_c_367_n 0.0098216f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_115 N_D1_c_105_n N_Y_c_453_n 0.00519789f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_116 N_D1_M1012_g N_Y_c_447_n 0.0175141f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_117 N_D1_M1012_g N_Y_c_451_n 7.56966e-19 $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_118 N_D1_M1011_g Y 0.0138377f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_119 N_D1_M1012_g Y 0.00753353f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_120 N_D1_c_107_n Y 0.0141808f $X=0.995 $Y=1.385 $X2=0 $Y2=0
cc_121 D1 Y 0.0153466f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_122 N_D1_M1011_g Y 0.00329777f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_123 N_D1_M1012_g Y 9.19315e-19 $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_124 N_D1_c_103_n N_Y_c_446_n 0.00446631f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_125 N_D1_c_105_n N_Y_c_446_n 0.0046202f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_126 N_D1_c_107_n N_Y_c_446_n 0.00997992f $X=0.995 $Y=1.385 $X2=0 $Y2=0
cc_127 D1 N_Y_c_446_n 0.0125724f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_128 N_D1_M1011_g Y 0.0137261f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_129 N_D1_M1012_g Y 0.0139698f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_130 N_D1_c_103_n N_A_40_74#_c_564_n 0.00904821f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_131 N_D1_c_105_n N_A_40_74#_c_564_n 6.7158e-19 $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_132 N_D1_c_106_n N_A_40_74#_c_564_n 0.00177966f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_133 D1 N_A_40_74#_c_564_n 0.0219843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_134 N_D1_c_103_n N_A_40_74#_c_565_n 0.0100245f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_135 N_D1_c_105_n N_A_40_74#_c_565_n 0.0120041f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_136 N_D1_c_103_n N_A_40_74#_c_566_n 0.00282152f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_137 N_D1_c_103_n N_VGND_c_695_n 0.00278247f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_138 N_D1_c_105_n N_VGND_c_695_n 0.00278271f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_139 N_D1_c_103_n N_VGND_c_698_n 0.00357287f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_140 N_D1_c_105_n N_VGND_c_698_n 0.00353526f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_141 N_C1_M1015_g N_B1_M1017_g 0.0202992f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_142 C1 N_B1_c_212_n 4.71864e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_143 N_C1_c_155_n N_B1_c_212_n 0.0202992f $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_144 C1 B1 0.0103841f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_145 N_C1_c_155_n B1 0.00440251f $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_146 N_C1_M1013_g N_VPWR_c_370_n 0.00366558f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_147 N_C1_M1013_g N_VPWR_c_371_n 0.005209f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_148 N_C1_M1015_g N_VPWR_c_371_n 0.005209f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_149 N_C1_M1015_g N_VPWR_c_372_n 0.0027763f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_150 N_C1_M1013_g N_VPWR_c_367_n 0.00982832f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_151 N_C1_M1015_g N_VPWR_c_367_n 0.00982376f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_152 N_C1_M1013_g N_Y_c_447_n 0.0141693f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_153 C1 N_Y_c_447_n 0.0152996f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_C1_c_155_n N_Y_c_447_n 4.1732e-19 $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_155 N_C1_M1013_g N_Y_c_448_n 0.0115311f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_156 N_C1_M1015_g N_Y_c_448_n 0.0125215f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_157 N_C1_M1015_g N_Y_c_473_n 0.0151969f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_158 C1 N_Y_c_473_n 0.00561225f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_C1_M1015_g N_Y_c_449_n 6.50516e-19 $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_160 N_C1_M1013_g N_Y_c_451_n 0.00486388f $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_161 N_C1_M1015_g N_Y_c_451_n 0.00469835f $X=1.945 $Y=2.4 $X2=0 $Y2=0
cc_162 C1 N_Y_c_451_n 0.0279601f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_C1_c_155_n N_Y_c_451_n 7.11382e-19 $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_164 N_C1_M1013_g Y 7.90299e-19 $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_165 C1 Y 0.0111018f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_166 N_C1_c_155_n Y 2.90167e-19 $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_167 N_C1_M1001_g N_Y_c_446_n 5.93224e-19 $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_168 C1 N_Y_c_446_n 0.00514333f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_169 N_C1_M1013_g Y 6.46654e-19 $X=1.495 $Y=2.4 $X2=0 $Y2=0
cc_170 N_C1_M1001_g N_A_40_74#_c_565_n 9.48753e-19 $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_171 N_C1_M1001_g N_A_40_74#_c_567_n 2.64945e-19 $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_172 N_C1_M1001_g N_A_40_74#_c_568_n 0.00100394f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_173 N_C1_M1002_g N_A_40_74#_c_568_n 0.0104532f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_174 C1 N_A_40_74#_c_568_n 0.003612f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_175 N_C1_c_155_n N_A_40_74#_c_568_n 0.00108687f $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_176 N_C1_M1001_g N_A_40_74#_c_582_n 0.0106874f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_177 N_C1_M1002_g N_A_40_74#_c_582_n 0.00854195f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_178 C1 N_A_40_74#_c_582_n 0.0319834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_179 N_C1_c_155_n N_A_40_74#_c_582_n 8.78523e-19 $X=1.945 $Y=1.465 $X2=0 $Y2=0
cc_180 N_C1_M1002_g N_A_299_74#_c_604_n 0.0112994f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_181 N_C1_M1001_g N_A_299_74#_c_605_n 0.00608065f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_182 N_C1_M1002_g N_A_299_74#_c_605_n 4.46617e-19 $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_183 N_C1_M1002_g N_A_510_74#_c_630_n 8.65009e-19 $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_184 N_C1_M1002_g N_A_510_74#_c_632_n 0.00183941f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_185 N_C1_M1001_g N_VGND_c_695_n 0.0043213f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_186 N_C1_M1002_g N_VGND_c_695_n 0.00278271f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_187 N_C1_M1001_g N_VGND_c_698_n 0.00447557f $X=1.42 $Y=0.74 $X2=0 $Y2=0
cc_188 N_C1_M1002_g N_VGND_c_698_n 0.00359085f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B1_M1009_g N_A2_M1000_g 0.0169057f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B1_c_216_n A2 2.25782e-19 $X=3.335 $Y=1.515 $X2=0 $Y2=0
cc_191 B1 A2 0.0290777f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_192 N_B1_c_216_n N_A2_c_277_n 0.0169057f $X=3.335 $Y=1.515 $X2=0 $Y2=0
cc_193 B1 N_A2_c_277_n 0.00627403f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_194 N_B1_M1017_g N_VPWR_c_372_n 0.0027763f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_195 N_B1_M1018_g N_VPWR_c_373_n 0.00501904f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_196 N_B1_M1017_g N_VPWR_c_376_n 0.005209f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_197 N_B1_M1018_g N_VPWR_c_376_n 0.005209f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_198 N_B1_M1017_g N_VPWR_c_367_n 0.00982376f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_199 N_B1_M1018_g N_VPWR_c_367_n 0.00987399f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_200 N_B1_M1017_g N_Y_c_473_n 0.0169825f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_201 N_B1_M1017_g N_Y_c_449_n 0.0119382f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_202 N_B1_M1018_g N_Y_c_449_n 0.0166062f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_203 N_B1_M1018_g N_Y_c_450_n 0.0150541f $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_204 N_B1_c_215_n N_Y_c_450_n 0.00286223f $X=2.755 $Y=1.53 $X2=0 $Y2=0
cc_205 B1 N_Y_c_450_n 0.0710723f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B1_M1017_g N_Y_c_451_n 0.0014449f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_207 N_B1_M1017_g N_Y_c_493_n 0.00186015f $X=2.395 $Y=2.4 $X2=0 $Y2=0
cc_208 N_B1_c_211_n N_Y_c_493_n 5.61336e-19 $X=2.755 $Y=1.605 $X2=0 $Y2=0
cc_209 N_B1_M1018_g N_Y_c_493_n 8.84614e-19 $X=2.845 $Y=2.4 $X2=0 $Y2=0
cc_210 B1 N_Y_c_493_n 0.0194095f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_211 N_B1_M1007_g N_A_40_74#_c_568_n 0.00129437f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B1_M1007_g N_A_299_74#_c_604_n 0.0132622f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B1_M1009_g N_A_299_74#_c_604_n 0.00500371f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B1_M1009_g N_A_299_74#_c_611_n 0.00491451f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B1_M1007_g N_A_510_74#_c_630_n 0.00750528f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B1_M1009_g N_A_510_74#_c_630_n 8.63392e-19 $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B1_M1007_g N_A_510_74#_c_631_n 0.0093986f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_218 N_B1_M1009_g N_A_510_74#_c_631_n 0.0134662f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B1_c_216_n N_A_510_74#_c_631_n 0.00381149f $X=3.335 $Y=1.515 $X2=0
+ $Y2=0
cc_220 B1 N_A_510_74#_c_631_n 0.0512198f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_221 N_B1_c_211_n N_A_510_74#_c_632_n 0.0012943f $X=2.755 $Y=1.605 $X2=0 $Y2=0
cc_222 N_B1_M1007_g N_A_510_74#_c_632_n 0.00326704f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B1_c_215_n N_A_510_74#_c_632_n 0.00135494f $X=2.755 $Y=1.53 $X2=0 $Y2=0
cc_224 B1 N_A_510_74#_c_632_n 0.0289808f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B1_M1009_g N_A_510_74#_c_633_n 3.92031e-19 $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_226 B1 N_A_510_74#_c_634_n 3.67275e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_227 B1 N_A_510_74#_c_638_n 0.0153286f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_M1009_g N_VGND_c_693_n 5.13093e-19 $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_M1007_g N_VGND_c_695_n 0.00278271f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B1_M1009_g N_VGND_c_695_n 0.00430908f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B1_M1007_g N_VGND_c_698_n 0.00359085f $X=2.91 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B1_M1009_g N_VGND_c_698_n 0.00817424f $X=3.41 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A2_M1019_g N_A1_M1004_g 0.0195237f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A2_M1005_g N_A1_M1006_g 0.0132434f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_235 A2 N_A1_M1006_g 0.00276109f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_236 A2 A1 0.0272178f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_237 A2 N_A1_c_325_n 0.0105349f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_238 N_A2_c_277_n N_A1_c_325_n 0.0211634f $X=4.305 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A2_M1003_g N_VPWR_c_373_n 8.64401e-19 $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A2_M1003_g N_VPWR_c_377_n 0.00333926f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A2_M1005_g N_VPWR_c_377_n 0.00333926f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A2_M1003_g N_VPWR_c_367_n 0.0042782f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A2_M1005_g N_VPWR_c_367_n 0.00422798f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A2_M1003_g N_Y_c_450_n 0.0196047f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A2_M1003_g N_Y_c_498_n 0.0161585f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A2_M1005_g N_Y_c_498_n 0.0108737f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_247 A2 N_Y_c_498_n 0.0202798f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_248 N_A2_c_277_n N_Y_c_498_n 5.54777e-19 $X=4.305 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A2_M1003_g N_A_697_368#_c_530_n 0.0149058f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A2_M1005_g N_A_697_368#_c_530_n 0.0137017f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_251 A2 N_A_697_368#_c_536_n 0.0143992f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_252 A2 N_A_697_368#_c_537_n 0.00286247f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_253 N_A2_M1000_g N_A_299_74#_c_604_n 3.00542e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1000_g N_A_510_74#_c_633_n 3.92313e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A2_M1000_g N_A_510_74#_c_634_n 0.0177742f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_M1019_g N_A_510_74#_c_634_n 0.0136953f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_257 A2 N_A_510_74#_c_634_n 0.0344116f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_258 N_A2_c_277_n N_A_510_74#_c_634_n 0.00359948f $X=4.305 $Y=1.515 $X2=0
+ $Y2=0
cc_259 N_A2_M1019_g N_A_510_74#_c_635_n 4.03583e-19 $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_260 A2 N_A_510_74#_c_636_n 3.30926e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_261 A2 N_A_510_74#_c_639_n 0.0223224f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_262 N_A2_M1000_g N_VGND_c_693_n 0.0105278f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_M1019_g N_VGND_c_693_n 0.0091926f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A2_M1000_g N_VGND_c_695_n 0.00383152f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_M1019_g N_VGND_c_696_n 0.00444681f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A2_M1000_g N_VGND_c_698_n 0.00757637f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A2_M1019_g N_VGND_c_698_n 0.00877616f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A1_M1006_g N_VPWR_c_374_n 0.0120713f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A1_M1008_g N_VPWR_c_374_n 0.00334717f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A1_M1006_g N_VPWR_c_377_n 0.00460063f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A1_M1008_g N_VPWR_c_378_n 0.005209f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A1_M1006_g N_VPWR_c_367_n 0.00908665f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A1_M1008_g N_VPWR_c_367_n 0.00985824f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_274 N_A1_M1006_g N_A_697_368#_c_530_n 0.00101073f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A1_M1006_g N_A_697_368#_c_537_n 0.0197444f $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A1_M1008_g N_A_697_368#_c_537_n 0.0132272f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_277 A1 N_A_697_368#_c_537_n 0.0279568f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_278 N_A1_c_325_n N_A_697_368#_c_537_n 0.00308477f $X=5.25 $Y=1.515 $X2=0
+ $Y2=0
cc_279 N_A1_M1008_g N_A_697_368#_c_532_n 8.84614e-19 $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_280 A1 N_A_697_368#_c_532_n 0.0254941f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_281 N_A1_c_325_n N_A_697_368#_c_532_n 2.88522e-19 $X=5.25 $Y=1.515 $X2=0
+ $Y2=0
cc_282 N_A1_M1006_g N_A_697_368#_c_533_n 8.97786e-19 $X=4.755 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A1_M1008_g N_A_697_368#_c_533_n 0.0117965f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A1_M1004_g N_A_510_74#_c_635_n 0.00913563f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A1_M1010_g N_A_510_74#_c_635_n 9.66583e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A1_M1004_g N_A_510_74#_c_636_n 0.0151535f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A1_M1010_g N_A_510_74#_c_636_n 0.0140467f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_288 A1 N_A_510_74#_c_636_n 0.0542669f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_289 N_A1_c_325_n N_A_510_74#_c_636_n 0.00732318f $X=5.25 $Y=1.515 $X2=0 $Y2=0
cc_290 N_A1_M1010_g N_A_510_74#_c_637_n 0.00159319f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A1_M1004_g N_A_510_74#_c_639_n 0.00155819f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A1_M1004_g N_VGND_c_693_n 5.12014e-19 $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A1_M1004_g N_VGND_c_694_n 0.00426511f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A1_M1010_g N_VGND_c_694_n 0.013385f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A1_M1004_g N_VGND_c_696_n 0.00434272f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A1_M1010_g N_VGND_c_697_n 0.00383152f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A1_M1004_g N_VGND_c_698_n 0.00820816f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A1_M1010_g N_VGND_c_698_n 0.00761342f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_299 N_VPWR_M1012_s N_Y_c_447_n 0.00218982f $X=1.085 $Y=1.84 $X2=0 $Y2=0
cc_300 N_VPWR_c_370_n N_Y_c_447_n 0.0167599f $X=1.27 $Y=2.305 $X2=0 $Y2=0
cc_301 N_VPWR_c_370_n N_Y_c_448_n 0.0283501f $X=1.27 $Y=2.305 $X2=0 $Y2=0
cc_302 N_VPWR_c_371_n N_Y_c_448_n 0.0144623f $X=2.085 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_c_372_n N_Y_c_448_n 0.0233699f $X=2.17 $Y=2.455 $X2=0 $Y2=0
cc_304 N_VPWR_c_367_n N_Y_c_448_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_305 N_VPWR_M1015_s N_Y_c_473_n 0.00761058f $X=2.035 $Y=1.84 $X2=0 $Y2=0
cc_306 N_VPWR_c_372_n N_Y_c_473_n 0.0126919f $X=2.17 $Y=2.455 $X2=0 $Y2=0
cc_307 N_VPWR_c_372_n N_Y_c_449_n 0.0233699f $X=2.17 $Y=2.455 $X2=0 $Y2=0
cc_308 N_VPWR_c_373_n N_Y_c_449_n 0.0234083f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_309 N_VPWR_c_376_n N_Y_c_449_n 0.0144623f $X=2.985 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_c_367_n N_Y_c_449_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_M1018_s N_Y_c_450_n 0.0052384f $X=2.935 $Y=1.84 $X2=0 $Y2=0
cc_312 N_VPWR_c_373_n N_Y_c_450_n 0.0197477f $X=3.07 $Y=2.455 $X2=0 $Y2=0
cc_313 N_VPWR_c_369_n Y 0.0062222f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_314 N_VPWR_c_369_n Y 0.0339179f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_315 N_VPWR_c_370_n Y 0.0322767f $X=1.27 $Y=2.305 $X2=0 $Y2=0
cc_316 N_VPWR_c_375_n Y 0.0144623f $X=1.105 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_367_n Y 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_c_373_n N_A_697_368#_c_529_n 0.0397231f $X=3.07 $Y=2.455 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_374_n N_A_697_368#_c_530_n 0.0103602f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_377_n N_A_697_368#_c_530_n 0.0581059f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_367_n N_A_697_368#_c_530_n 0.0324093f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_373_n N_A_697_368#_c_531_n 0.011925f $X=3.07 $Y=2.455 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_377_n N_A_697_368#_c_531_n 0.0179217f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_367_n N_A_697_368#_c_531_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_325 N_VPWR_M1006_d N_A_697_368#_c_537_n 0.00408051f $X=4.845 $Y=1.84 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_374_n N_A_697_368#_c_537_n 0.0189268f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_374_n N_A_697_368#_c_533_n 0.0266809f $X=4.98 $Y=2.455 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_378_n N_A_697_368#_c_533_n 0.014549f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_329 N_VPWR_c_367_n N_A_697_368#_c_533_n 0.0119743f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_Y_c_450_n N_A_697_368#_M1003_s 0.00567673f $X=3.915 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_331 N_Y_c_450_n N_A_697_368#_c_529_n 0.0197477f $X=3.915 $Y=2.035 $X2=0 $Y2=0
cc_332 N_Y_M1003_d N_A_697_368#_c_530_n 0.00165831f $X=3.945 $Y=1.84 $X2=0 $Y2=0
cc_333 N_Y_c_498_n N_A_697_368#_c_530_n 0.0159318f $X=4.08 $Y=2.115 $X2=0 $Y2=0
cc_334 N_Y_M1014_s N_A_40_74#_c_565_n 0.00176461f $X=0.635 $Y=0.37 $X2=0 $Y2=0
cc_335 N_Y_c_453_n N_A_40_74#_c_565_n 0.0143448f $X=0.775 $Y=0.86 $X2=0 $Y2=0
cc_336 N_Y_c_447_n N_A_40_74#_c_567_n 0.00549175f $X=1.555 $Y=1.885 $X2=0 $Y2=0
cc_337 N_Y_c_446_n N_A_40_74#_c_567_n 0.00503069f $X=0.77 $Y=1.345 $X2=0 $Y2=0
cc_338 N_A_40_74#_c_582_n N_A_299_74#_M1001_s 0.00470069f $X=1.97 $Y=0.862
+ $X2=-0.19 $Y2=-0.245
cc_339 N_A_40_74#_M1002_d N_A_299_74#_c_604_n 0.00274343f $X=1.995 $Y=0.37 $X2=0
+ $Y2=0
cc_340 N_A_40_74#_c_568_n N_A_299_74#_c_604_n 0.0202288f $X=2.135 $Y=0.86 $X2=0
+ $Y2=0
cc_341 N_A_40_74#_c_582_n N_A_299_74#_c_604_n 0.00364964f $X=1.97 $Y=0.862 $X2=0
+ $Y2=0
cc_342 N_A_40_74#_c_565_n N_A_299_74#_c_605_n 0.0112234f $X=1.12 $Y=0.34 $X2=0
+ $Y2=0
cc_343 N_A_40_74#_c_582_n N_A_299_74#_c_605_n 0.0197079f $X=1.97 $Y=0.862 $X2=0
+ $Y2=0
cc_344 N_A_40_74#_c_568_n N_A_510_74#_c_630_n 0.0286351f $X=2.135 $Y=0.86 $X2=0
+ $Y2=0
cc_345 N_A_40_74#_c_568_n N_A_510_74#_c_632_n 0.00854265f $X=2.135 $Y=0.86 $X2=0
+ $Y2=0
cc_346 N_A_40_74#_c_565_n N_VGND_c_695_n 0.050626f $X=1.12 $Y=0.34 $X2=0 $Y2=0
cc_347 N_A_40_74#_c_566_n N_VGND_c_695_n 0.0235688f $X=0.51 $Y=0.34 $X2=0 $Y2=0
cc_348 N_A_40_74#_c_565_n N_VGND_c_698_n 0.028285f $X=1.12 $Y=0.34 $X2=0 $Y2=0
cc_349 N_A_40_74#_c_566_n N_VGND_c_698_n 0.0127152f $X=0.51 $Y=0.34 $X2=0 $Y2=0
cc_350 N_A_40_74#_c_582_n N_VGND_c_698_n 0.00653179f $X=1.97 $Y=0.862 $X2=0
+ $Y2=0
cc_351 N_A_299_74#_c_604_n N_A_510_74#_M1007_d 0.00273752f $X=3.03 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_352 N_A_299_74#_c_604_n N_A_510_74#_c_630_n 0.0203278f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_353 N_A_299_74#_M1007_s N_A_510_74#_c_631_n 0.00250873f $X=2.985 $Y=0.37
+ $X2=0 $Y2=0
cc_354 N_A_299_74#_c_604_n N_A_510_74#_c_631_n 0.00304353f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_355 N_A_299_74#_c_611_n N_A_510_74#_c_631_n 0.0207721f $X=3.195 $Y=0.635
+ $X2=0 $Y2=0
cc_356 N_A_299_74#_c_604_n N_A_510_74#_c_633_n 0.00370621f $X=3.03 $Y=0.34 $X2=0
+ $Y2=0
cc_357 N_A_299_74#_c_604_n N_VGND_c_693_n 0.0029789f $X=3.03 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_299_74#_c_604_n N_VGND_c_695_n 0.101637f $X=3.03 $Y=0.34 $X2=0 $Y2=0
cc_359 N_A_299_74#_c_605_n N_VGND_c_695_n 0.0225845f $X=1.635 $Y=0.34 $X2=0
+ $Y2=0
cc_360 N_A_299_74#_c_604_n N_VGND_c_698_n 0.0575414f $X=3.03 $Y=0.34 $X2=0 $Y2=0
cc_361 N_A_299_74#_c_605_n N_VGND_c_698_n 0.0124836f $X=1.635 $Y=0.34 $X2=0
+ $Y2=0
cc_362 N_A_510_74#_c_634_n N_VGND_M1000_s 0.00197722f $X=4.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_363 N_A_510_74#_c_636_n N_VGND_M1004_s 0.00250873f $X=5.35 $Y=1.095 $X2=0
+ $Y2=0
cc_364 N_A_510_74#_c_633_n N_VGND_c_693_n 0.0182488f $X=3.625 $Y=0.515 $X2=0
+ $Y2=0
cc_365 N_A_510_74#_c_634_n N_VGND_c_693_n 0.0172656f $X=4.42 $Y=1.095 $X2=0
+ $Y2=0
cc_366 N_A_510_74#_c_635_n N_VGND_c_693_n 0.0168193f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_510_74#_c_635_n N_VGND_c_694_n 0.0184106f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_368 N_A_510_74#_c_636_n N_VGND_c_694_n 0.0210288f $X=5.35 $Y=1.095 $X2=0
+ $Y2=0
cc_369 N_A_510_74#_c_637_n N_VGND_c_694_n 0.0182902f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_370 N_A_510_74#_c_633_n N_VGND_c_695_n 0.00749631f $X=3.625 $Y=0.515 $X2=0
+ $Y2=0
cc_371 N_A_510_74#_c_635_n N_VGND_c_696_n 0.0109942f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_372 N_A_510_74#_c_637_n N_VGND_c_697_n 0.011066f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_373 N_A_510_74#_c_633_n N_VGND_c_698_n 0.0062048f $X=3.625 $Y=0.515 $X2=0
+ $Y2=0
cc_374 N_A_510_74#_c_635_n N_VGND_c_698_n 0.00904371f $X=4.505 $Y=0.515 $X2=0
+ $Y2=0
cc_375 N_A_510_74#_c_637_n N_VGND_c_698_n 0.00915947f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__dlrtp_2.pex.spice
* Created: Wed Sep  2 12:05:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRTP_2%D 3 7 9 12 13
c28 7 0 1.60049e-19 $X=0.52 $Y=0.835
r29 12 15 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.78
r30 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.45
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r32 9 13 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r33 7 14 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.52 $Y=0.835
+ $X2=0.52 $Y2=1.45
r34 3 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=0.505 $Y=2.38 $X2=0.505
+ $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%GATE 3 6 8 11 13
c39 8 0 2.85504e-19 $X=1.2 $Y=1.295
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.385
+ $X2=1.155 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.385
+ $X2=1.155 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.385 $X2=1.155 $Y2=1.385
r43 8 12 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.385
r44 6 14 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=1.125 $Y=2.38
+ $X2=1.125 $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.1 $Y=0.74 $X2=1.1
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%A_235_74# 1 2 9 13 17 19 20 23 25 26 28 30
+ 31 34 35 36 40 47 52 56 57 58
c151 35 0 1.78997e-19 $X=3.92 $Y=0.34
c152 26 0 1.86781e-19 $X=2.045 $Y=1.42
c153 25 0 1.25456e-19 $X=2.045 $Y=1.585
c154 23 0 1.18818e-19 $X=3.845 $Y=0.615
c155 20 0 2.9829e-19 $X=3.26 $Y=1.735
c156 19 0 1.64562e-19 $X=3.76 $Y=1.735
r157 56 58 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.957 $Y=1.425
+ $X2=3.957 $Y2=1.26
r158 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.425 $X2=3.925 $Y2=1.425
r159 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.585 $X2=1.725 $Y2=1.585
r160 49 52 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.54 $Y=1.585
+ $X2=1.725 $Y2=1.585
r161 45 47 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.35 $Y=2.105
+ $X2=1.54 $Y2=2.105
r162 42 43 13.8993 $w=4.73e-07 $l=3.45e-07 $layer=LI1_cond $X=1.387 $Y=0.665
+ $X2=1.387 $Y2=1.01
r163 40 42 3.77709 $w=4.73e-07 $l=1.5e-07 $layer=LI1_cond $X=1.387 $Y=0.515
+ $X2=1.387 $Y2=0.665
r164 37 58 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.005 $Y=0.425
+ $X2=4.005 $Y2=1.26
r165 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=0.34
+ $X2=4.005 $Y2=0.425
r166 35 36 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.92 $Y=0.34
+ $X2=2.975 $Y2=0.34
r167 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.89 $Y=0.425
+ $X2=2.975 $Y2=0.34
r168 33 34 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.89 $Y=0.425
+ $X2=2.89 $Y2=0.58
r169 32 42 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=1.625 $Y=0.665
+ $X2=1.387 $Y2=0.665
r170 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.805 $Y=0.665
+ $X2=2.89 $Y2=0.58
r171 31 32 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.805 $Y=0.665
+ $X2=1.625 $Y2=0.665
r172 30 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.94
+ $X2=1.54 $Y2=2.105
r173 29 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.75
+ $X2=1.54 $Y2=1.585
r174 29 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=1.75
+ $X2=1.54 $Y2=1.94
r175 28 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.42
+ $X2=1.54 $Y2=1.585
r176 28 43 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.54 $Y=1.42
+ $X2=1.54 $Y2=1.01
r177 25 53 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=2.045 $Y=1.585
+ $X2=1.725 $Y2=1.585
r178 25 26 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.045 $Y=1.585
+ $X2=2.045 $Y2=1.42
r179 21 57 39.2009 $w=2.58e-07 $l=2.0106e-07 $layer=POLY_cond $X=3.845 $Y=1.26
+ $X2=3.925 $Y2=1.425
r180 21 23 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.845 $Y=1.26
+ $X2=3.845 $Y2=0.615
r181 19 57 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=3.76 $Y=1.735
+ $X2=3.925 $Y2=1.425
r182 19 20 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.76 $Y=1.735
+ $X2=3.26 $Y2=1.735
r183 15 20 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.17 $Y=1.81
+ $X2=3.26 $Y2=1.735
r184 15 17 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=3.17 $Y=1.81
+ $X2=3.17 $Y2=2.46
r185 11 26 34.7346 $w=1.65e-07 $l=1.3e-07 $layer=POLY_cond $X=2.175 $Y=1.42
+ $X2=2.045 $Y2=1.42
r186 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.175 $Y=1.42
+ $X2=2.175 $Y2=0.86
r187 7 26 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=2.135 $Y=1.75
+ $X2=2.045 $Y2=1.42
r188 7 9 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.135 $Y=1.75
+ $X2=2.135 $Y2=2.38
r189 2 45 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.96 $X2=1.35 $Y2=2.105
r190 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.175
+ $Y=0.37 $X2=1.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%A_27_392# 1 2 9 13 17 19 20 22 23 26 28 31
+ 32
c96 31 0 1.66318e-19 $X=2.675 $Y=1.605
c97 26 0 1.66802e-19 $X=2.595 $Y=2.44
r98 32 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.605
+ $X2=2.675 $Y2=1.77
r99 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.605
+ $X2=2.675 $Y2=1.44
r100 31 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=1.605
+ $X2=2.675 $Y2=1.77
r101 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.605 $X2=2.675 $Y2=1.605
r102 28 29 7.80343 $w=6.41e-07 $l=4.1e-07 $layer=LI1_cond $X=0.485 $Y=2.115
+ $X2=0.485 $Y2=2.525
r103 26 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.595 $Y=2.44
+ $X2=2.595 $Y2=1.77
r104 24 29 8.74498 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.855 $Y=2.525
+ $X2=0.485 $Y2=2.525
r105 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.51 $Y=2.525
+ $X2=2.595 $Y2=2.44
r106 23 24 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=2.51 $Y=2.525
+ $X2=0.855 $Y2=2.525
r107 22 28 10.6318 $w=6.41e-07 $l=3.5812e-07 $layer=LI1_cond $X=0.77 $Y=1.95
+ $X2=0.485 $Y2=2.115
r108 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.77 $Y=1.28
+ $X2=0.77 $Y2=1.95
r109 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.77 $Y2=1.28
r110 19 20 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.685 $Y=1.195
+ $X2=0.47 $Y2=1.195
r111 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.305 $Y=1.11
+ $X2=0.47 $Y2=1.195
r112 15 17 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.305 $Y=1.11
+ $X2=0.305 $Y2=0.835
r113 13 36 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.765 $Y=0.69
+ $X2=2.765 $Y2=1.44
r114 9 37 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=2.75 $Y=2.46 $X2=2.75
+ $Y2=1.77
r115 2 28 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r116 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.56 $X2=0.305 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%A_347_98# 1 2 9 12 15 16 19 21 22 23 26 27
+ 33 37 41 47 50
c112 47 0 3.48291e-20 $X=3.215 $Y=1.285
c113 33 0 1.86781e-19 $X=2.23 $Y=1.085
c114 26 0 1.64562e-19 $X=3.895 $Y=2.215
r115 47 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.285
+ $X2=3.215 $Y2=1.12
r116 46 48 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.182 $Y=1.285
+ $X2=3.182 $Y2=1.45
r117 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.285 $X2=3.215 $Y2=1.285
r118 39 41 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.975 $Y=2.025
+ $X2=3.135 $Y2=2.025
r119 35 37 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.91 $Y=2.105
+ $X2=2.145 $Y2=2.105
r120 32 33 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.085
+ $X2=2.23 $Y2=1.085
r121 30 32 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.88 $Y=1.085
+ $X2=2.145 $Y2=1.085
r122 27 52 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.895 $Y=2.215
+ $X2=3.705 $Y2=2.215
r123 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=2.215 $X2=3.895 $Y2=2.215
r124 24 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.895 $Y=2.905
+ $X2=3.895 $Y2=2.215
r125 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.73 $Y=2.99
+ $X2=3.895 $Y2=2.905
r126 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.73 $Y=2.99
+ $X2=3.06 $Y2=2.99
r127 21 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=1.94
+ $X2=3.135 $Y2=2.025
r128 21 48 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.135 $Y=1.94
+ $X2=3.135 $Y2=1.45
r129 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.975 $Y=2.905
+ $X2=3.06 $Y2=2.99
r130 18 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.11
+ $X2=2.975 $Y2=2.025
r131 18 19 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.975 $Y=2.11
+ $X2=2.975 $Y2=2.905
r132 16 46 5.21861 $w=2.63e-07 $l=1.2e-07 $layer=LI1_cond $X=3.182 $Y=1.165
+ $X2=3.182 $Y2=1.285
r133 16 33 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.05 $Y=1.165
+ $X2=2.23 $Y2=1.165
r134 15 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.94
+ $X2=2.145 $Y2=2.105
r135 14 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.25
+ $X2=2.145 $Y2=1.085
r136 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.145 $Y=1.25
+ $X2=2.145 $Y2=1.94
r137 10 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=2.38
+ $X2=3.705 $Y2=2.215
r138 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.705 $Y=2.38
+ $X2=3.705 $Y2=2.75
r139 9 50 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.155 $Y=0.69
+ $X2=3.155 $Y2=1.12
r140 2 35 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.96 $X2=1.91 $Y2=2.105
r141 1 30 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.49 $X2=1.88 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%A_832_55# 1 2 7 9 14 18 22 26 30 34 36 39 43
+ 49 51 53 55 58 59 60 70 75
c138 60 0 3.83707e-20 $X=5.34 $Y=1.72
c139 51 0 7.10122e-20 $X=6.05 $Y=1.805
r140 75 76 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=6.645 $Y=1.465
+ $X2=6.66 $Y2=1.465
r141 72 73 1.49689 $w=3.22e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.465
+ $X2=6.205 $Y2=1.465
r142 63 64 4.69791 $w=4.88e-07 $l=1.4e-07 $layer=LI1_cond $X=5.34 $Y=2.24
+ $X2=5.34 $Y2=2.38
r143 62 63 6.22449 $w=4.88e-07 $l=2.55e-07 $layer=LI1_cond $X=5.34 $Y=1.985
+ $X2=5.34 $Y2=2.24
r144 59 62 4.39376 $w=4.88e-07 $l=1.8e-07 $layer=LI1_cond $X=5.34 $Y=1.805
+ $X2=5.34 $Y2=1.985
r145 59 60 7.50345 $w=4.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=1.805
+ $X2=5.34 $Y2=1.72
r146 58 60 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.18 $Y=1.13
+ $X2=5.18 $Y2=1.72
r147 56 75 13.472 $w=3.22e-07 $l=9e-08 $layer=POLY_cond $X=6.555 $Y=1.465
+ $X2=6.645 $Y2=1.465
r148 56 73 52.3913 $w=3.22e-07 $l=3.5e-07 $layer=POLY_cond $X=6.555 $Y=1.465
+ $X2=6.205 $Y2=1.465
r149 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.555
+ $Y=1.465 $X2=6.555 $Y2=1.465
r150 53 67 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.135 $Y=1.465
+ $X2=6.135 $Y2=1.805
r151 53 55 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.22 $Y=1.465
+ $X2=6.555 $Y2=1.465
r152 52 59 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=5.585 $Y=1.805
+ $X2=5.34 $Y2=1.805
r153 51 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.05 $Y=1.805
+ $X2=6.135 $Y2=1.805
r154 51 52 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.05 $Y=1.805
+ $X2=5.585 $Y2=1.805
r155 49 64 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.42 $Y=2.815
+ $X2=5.42 $Y2=2.38
r156 41 58 9.97136 $w=4.18e-07 $l=2.1e-07 $layer=LI1_cond $X=5.055 $Y=0.92
+ $X2=5.055 $Y2=1.13
r157 41 43 11.1128 $w=4.18e-07 $l=4.05e-07 $layer=LI1_cond $X=5.055 $Y=0.92
+ $X2=5.055 $Y2=0.515
r158 39 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=2.215
+ $X2=4.465 $Y2=2.38
r159 39 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=2.215
+ $X2=4.465 $Y2=2.05
r160 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.465
+ $Y=2.215 $X2=4.465 $Y2=2.215
r161 36 63 4.01183 $w=2.8e-07 $l=2.45e-07 $layer=LI1_cond $X=5.095 $Y=2.24
+ $X2=5.34 $Y2=2.24
r162 36 38 25.93 $w=2.78e-07 $l=6.3e-07 $layer=LI1_cond $X=5.095 $Y=2.24
+ $X2=4.465 $Y2=2.24
r163 32 34 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.235 $Y=0.975
+ $X2=4.375 $Y2=0.975
r164 28 76 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.63
+ $X2=6.66 $Y2=1.465
r165 28 30 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.66 $Y=1.63
+ $X2=6.66 $Y2=2.4
r166 24 75 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.3
+ $X2=6.645 $Y2=1.465
r167 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.645 $Y=1.3
+ $X2=6.645 $Y2=0.74
r168 20 73 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=1.465
r169 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.205 $Y=1.3
+ $X2=6.205 $Y2=0.74
r170 16 72 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=1.465
r171 16 18 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=2.4
r172 14 71 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.39 $Y=2.75
+ $X2=4.39 $Y2=2.38
r173 10 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.375 $Y=1.05
+ $X2=4.375 $Y2=0.975
r174 10 70 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.375 $Y=1.05
+ $X2=4.375 $Y2=2.05
r175 7 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.235 $Y=0.9
+ $X2=4.235 $Y2=0.975
r176 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.235 $Y=0.9 $X2=4.235
+ $Y2=0.615
r177 2 62 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.84 $X2=5.42 $Y2=1.985
r178 2 49 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.84 $X2=5.42 $Y2=2.815
r179 1 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.37 $X2=5.01 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%A_646_74# 1 2 9 13 15 16 17 23 24 28 32 33
+ 35
c89 9 0 7.10122e-20 $X=5.195 $Y=2.4
r90 32 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=2.57
+ $X2=3.395 $Y2=2.405
r91 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.515 $X2=4.825 $Y2=1.515
r92 26 28 10.6547 $w=2.63e-07 $l=2.45e-07 $layer=LI1_cond $X=4.792 $Y=1.76
+ $X2=4.792 $Y2=1.515
r93 25 35 1.34256 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.655 $Y=1.845
+ $X2=3.522 $Y2=1.845
r94 24 26 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=4.66 $Y=1.845
+ $X2=4.792 $Y2=1.76
r95 24 25 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.66 $Y=1.845
+ $X2=3.655 $Y2=1.845
r96 23 35 5.16603 $w=1.7e-07 $l=1.06325e-07 $layer=LI1_cond $X=3.57 $Y=1.76
+ $X2=3.522 $Y2=1.845
r97 22 23 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.57 $Y=0.845
+ $X2=3.57 $Y2=1.76
r98 20 35 5.16603 $w=1.7e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.475 $Y=1.93
+ $X2=3.522 $Y2=1.845
r99 20 33 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.475 $Y=1.93
+ $X2=3.475 $Y2=2.405
r100 17 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.485 $Y=0.72
+ $X2=3.57 $Y2=0.845
r101 17 19 1.22 $w=2.5e-07 $l=2.5e-08 $layer=LI1_cond $X=3.485 $Y=0.72 $X2=3.46
+ $Y2=0.72
r102 15 29 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.105 $Y=1.515
+ $X2=4.825 $Y2=1.515
r103 15 16 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=1.515
+ $X2=5.105 $Y2=1.35
r104 11 16 34.7346 $w=1.65e-07 $l=1.2e-07 $layer=POLY_cond $X=5.225 $Y=1.35
+ $X2=5.105 $Y2=1.35
r105 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.225 $Y=1.35
+ $X2=5.225 $Y2=0.74
r106 7 16 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=5.195 $Y=1.68
+ $X2=5.105 $Y2=1.35
r107 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.195 $Y=1.68
+ $X2=5.195 $Y2=2.4
r108 2 32 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.96 $X2=3.395 $Y2=2.57
r109 1 19 182 $w=1.7e-07 $l=4.09145e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.37 $X2=3.46 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%RESET_B 3 6 8 11 12 13
c41 13 0 3.83707e-20 $X=5.675 $Y=1.22
r42 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.385
+ $X2=5.675 $Y2=1.55
r43 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.385
+ $X2=5.675 $Y2=1.22
r44 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.675
+ $Y=1.385 $X2=5.675 $Y2=1.385
r45 8 12 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.52 $Y=1.365
+ $X2=5.675 $Y2=1.365
r46 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.645 $Y=2.4
+ $X2=5.645 $Y2=1.55
r47 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.615 $Y=0.74
+ $X2=5.615 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%VPWR 1 2 3 4 5 20 24 28 32 34 37 38 39 48 55
+ 60 66 69 76 80
r82 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r83 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r84 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 64 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r87 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r88 61 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=5.92 $Y2=3.33
r89 61 63 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=6.48 $Y2=3.33
r90 60 79 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.977 $Y2=3.33
r91 60 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 59 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r93 59 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r95 56 58 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.085 $Y=3.33
+ $X2=5.52 $Y2=3.33
r96 55 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.92 $Y2=3.33
r97 55 58 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r100 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r101 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 48 56 8.68381 $w=1.7e-07 $l=3.18e-07 $layer=LI1_cond $X=4.767 $Y=3.33
+ $X2=5.085 $Y2=3.33
r103 48 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 48 69 9.70048 $w=6.33e-07 $l=5.15e-07 $layer=LI1_cond $X=4.767 $Y=3.33
+ $X2=4.767 $Y2=2.815
r105 48 53 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.45 $Y=3.33
+ $X2=4.08 $Y2=3.33
r106 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 44 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r111 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r113 41 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 39 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r115 39 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 37 46 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.445 $Y2=3.33
r118 36 50 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.61 $Y=3.33 $X2=2.64
+ $Y2=3.33
r119 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.445 $Y2=3.33
r120 32 79 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.977 $Y2=3.33
r121 32 34 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.305
r122 28 31 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.92 $Y=2.145
+ $X2=5.92 $Y2=2.825
r123 26 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=3.33
r124 26 31 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=2.825
r125 22 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=3.33
r126 22 24 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=2.945
r127 18 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r128 18 20 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.945
r129 5 34 300 $w=1.7e-07 $l=5.43392e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=1.84 $X2=6.92 $Y2=2.305
r130 4 31 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.84 $X2=5.92 $Y2=2.825
r131 4 28 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.84 $X2=5.92 $Y2=2.145
r132 3 69 600 $w=1.7e-07 $l=3.995e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=2.54 $X2=4.765 $Y2=2.815
r133 2 24 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.96 $X2=2.445 $Y2=2.945
r134 1 20 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.815 $Y2=2.945
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%Q 1 2 9 11 13 15 16 17 24
r43 23 24 25.3036 $w=2.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.96 $Y=1.8
+ $X2=6.96 $Y2=1.295
r44 22 24 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.96 $Y=1.13
+ $X2=6.96 $Y2=1.295
r45 19 21 13.6724 $w=2.32e-07 $l=2.6e-07 $layer=LI1_cond $X=6.42 $Y=1.885
+ $X2=6.42 $Y2=2.145
r46 18 19 2.55969 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=1.885
+ $X2=6.42 $Y2=1.885
r47 17 23 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.96 $Y2=1.8
r48 17 18 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.585 $Y2=1.885
r49 15 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.96 $Y2=1.13
r50 15 16 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.585 $Y2=1.045
r51 11 21 4.04823 $w=3.3e-07 $l=8e-08 $layer=LI1_cond $X=6.42 $Y=2.225 $X2=6.42
+ $Y2=2.145
r52 11 13 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=6.42 $Y=2.225 $X2=6.42
+ $Y2=2.825
r53 7 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.42 $Y=0.96
+ $X2=6.585 $Y2=1.045
r54 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.42 $Y=0.96 $X2=6.42
+ $Y2=0.515
r55 2 21 400 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=2.145
r56 2 13 400 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=2.825
r57 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.37 $X2=6.42 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_2%VGND 1 2 3 4 5 20 24 28 30 32 34 35 41 50 57
+ 62 68 71 74 78
c80 24 0 1.18818e-19 $X=4.45 $Y=0.615
r81 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r82 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r83 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r85 66 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r86 66 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r87 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r88 63 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=5.92
+ $Y2=0
r89 63 65 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=6.48
+ $Y2=0
r90 62 77 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r91 62 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r92 61 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r93 61 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r94 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 58 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=4.45
+ $Y2=0
r96 58 60 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=5.52
+ $Y2=0
r97 57 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.92
+ $Y2=0
r98 57 60 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.52
+ $Y2=0
r99 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r101 52 55 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r102 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r103 50 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.45
+ $Y2=0
r104 50 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=0
+ $X2=4.08 $Y2=0
r105 49 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r106 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r107 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r108 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r110 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r111 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r112 43 45 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r113 41 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r114 41 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r115 37 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.64
+ $Y2=0
r116 35 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.16 $Y2=0
r117 34 39 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.47
+ $Y2=0.325
r118 34 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.635
+ $Y2=0
r119 34 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.305
+ $Y2=0
r120 30 77 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r121 30 32 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.625
r122 26 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r123 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.515
r124 22 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r125 22 24 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.615
r126 18 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r127 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.515
r128 5 32 182 $w=1.7e-07 $l=3.40624e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.37 $X2=6.92 $Y2=0.625
r129 4 28 91 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=2 $X=5.69
+ $Y=0.37 $X2=5.92 $Y2=0.515
r130 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.31
+ $Y=0.405 $X2=4.45 $Y2=0.615
r131 2 39 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.49 $X2=2.47 $Y2=0.325
r132 1 20 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.56 $X2=0.815 $Y2=0.515
.ends


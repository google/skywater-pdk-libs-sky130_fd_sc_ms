* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor2_4 A B VGND VNB VPB VPWR Y
X0 a_27_74# B a_119_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_511_74# a_119_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 Y B a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 Y a_119_368# a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_511_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_950_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_119_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X7 Y a_119_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_511_74# a_119_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 Y a_119_368# a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_119_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X11 a_511_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND B a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_950_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_950_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_511_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_950_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VPWR A a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 VGND A a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR A a_119_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X20 VGND A a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR a_119_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 VGND B a_511_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR B a_119_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X24 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X25 a_119_368# B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 a_511_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VPWR A a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 Y B a_950_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__a222oi_1.pxi.spice
* Created: Fri Aug 28 17:02:12 2020
* 
x_PM_SKY130_FD_SC_MS__A222OI_1%C1 N_C1_M1001_g N_C1_M1003_g C1 N_C1_c_73_n
+ N_C1_c_74_n N_C1_c_75_n PM_SKY130_FD_SC_MS__A222OI_1%C1
x_PM_SKY130_FD_SC_MS__A222OI_1%C2 N_C2_M1000_g N_C2_M1011_g C2 C2 N_C2_c_103_n
+ N_C2_c_104_n PM_SKY130_FD_SC_MS__A222OI_1%C2
x_PM_SKY130_FD_SC_MS__A222OI_1%B2 N_B2_M1009_g N_B2_M1002_g N_B2_c_137_n
+ N_B2_c_138_n N_B2_c_139_n B2 B2 N_B2_c_141_n PM_SKY130_FD_SC_MS__A222OI_1%B2
x_PM_SKY130_FD_SC_MS__A222OI_1%B1 N_B1_M1004_g N_B1_M1010_g N_B1_c_176_n
+ N_B1_c_177_n N_B1_c_178_n B1 B1 N_B1_c_180_n PM_SKY130_FD_SC_MS__A222OI_1%B1
x_PM_SKY130_FD_SC_MS__A222OI_1%A1 N_A1_c_216_n N_A1_M1008_g N_A1_M1006_g
+ N_A1_c_217_n A1 A1 N_A1_c_218_n N_A1_c_219_n N_A1_c_220_n
+ PM_SKY130_FD_SC_MS__A222OI_1%A1
x_PM_SKY130_FD_SC_MS__A222OI_1%A2 N_A2_M1005_g N_A2_M1007_g A2 A2 N_A2_c_258_n
+ PM_SKY130_FD_SC_MS__A222OI_1%A2
x_PM_SKY130_FD_SC_MS__A222OI_1%Y N_Y_M1003_s N_Y_M1004_d N_Y_M1001_s N_Y_M1011_d
+ N_Y_c_288_n N_Y_c_289_n N_Y_c_283_n N_Y_c_298_n N_Y_c_300_n N_Y_c_284_n
+ N_Y_c_290_n N_Y_c_291_n N_Y_c_285_n N_Y_c_323_n Y Y Y Y
+ PM_SKY130_FD_SC_MS__A222OI_1%Y
x_PM_SKY130_FD_SC_MS__A222OI_1%A_119_392# N_A_119_392#_M1001_d
+ N_A_119_392#_M1009_d N_A_119_392#_c_366_n N_A_119_392#_c_363_n
+ N_A_119_392#_c_364_n N_A_119_392#_c_371_n
+ PM_SKY130_FD_SC_MS__A222OI_1%A_119_392#
x_PM_SKY130_FD_SC_MS__A222OI_1%A_369_392# N_A_369_392#_M1009_s
+ N_A_369_392#_M1010_d N_A_369_392#_M1007_d N_A_369_392#_c_393_n
+ N_A_369_392#_c_388_n N_A_369_392#_c_405_n N_A_369_392#_c_389_n
+ N_A_369_392#_c_390_n N_A_369_392#_c_391_n N_A_369_392#_c_392_n
+ PM_SKY130_FD_SC_MS__A222OI_1%A_369_392#
x_PM_SKY130_FD_SC_MS__A222OI_1%VPWR N_VPWR_M1008_d N_VPWR_c_431_n N_VPWR_c_432_n
+ N_VPWR_c_433_n VPWR N_VPWR_c_434_n N_VPWR_c_430_n
+ PM_SKY130_FD_SC_MS__A222OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A222OI_1%VGND N_VGND_M1000_d N_VGND_M1005_d N_VGND_c_466_n
+ N_VGND_c_467_n VGND N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n
+ N_VGND_c_471_n PM_SKY130_FD_SC_MS__A222OI_1%VGND
cc_1 VNB N_C1_M1001_g 0.0124041f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_2 VNB N_C1_c_73_n 0.0334751f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_3 VNB N_C1_c_74_n 0.0274553f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_4 VNB N_C1_c_75_n 0.023864f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.12
cc_5 VNB C2 0.0030793f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C2_c_103_n 0.0628469f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.12
cc_7 VNB N_C2_c_104_n 0.0197172f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.455
cc_8 VNB N_B2_c_137_n 0.0194107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B2_c_138_n 0.0279322f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_10 VNB N_B2_c_139_n 0.00289239f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_11 VNB B2 0.00168047f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_12 VNB N_B2_c_141_n 0.0187447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_176_n 0.0196919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_177_n 0.0219347f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_15 VNB N_B1_c_178_n 0.00227135f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_16 VNB B1 0.00551108f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_17 VNB N_B1_c_180_n 0.0158166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_216_n 0.0209748f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_19 VNB N_A1_c_217_n 0.00340501f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.285
cc_20 VNB N_A1_c_218_n 0.018178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_219_n 0.0152451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_220_n 0.0199469f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.455
cc_23 VNB N_A2_M1005_g 0.0265625f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_24 VNB N_A2_M1007_g 0.00970738f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_25 VNB A2 0.0100538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_258_n 0.0591204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_283_n 0.0189692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_284_n 0.0072208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_285_n 0.00618121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.0158532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB Y 8.17974e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_430_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_466_n 0.0128247f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.69
cc_34 VNB N_VGND_c_467_n 0.0321458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_468_n 0.0459918f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.455
cc_36 VNB N_VGND_c_469_n 0.0299712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_470_n 0.0355947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_471_n 0.253868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_C1_M1001_g 0.039542f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_40 VPB N_C1_c_74_n 0.00936426f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_41 VPB N_C2_M1011_g 0.0256615f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_42 VPB C2 0.0020523f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB N_C2_c_103_n 0.0212071f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.12
cc_44 VPB N_B2_M1009_g 0.0259391f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_45 VPB N_B2_c_139_n 0.015002f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_46 VPB B2 0.00139606f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_47 VPB N_B1_M1010_g 0.0234341f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_48 VPB N_B1_c_178_n 0.0126891f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_49 VPB B1 0.00245553f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_50 VPB N_A1_M1008_g 0.0249188f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.12
cc_51 VPB N_A1_c_217_n 0.0139902f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_52 VPB N_A1_c_219_n 0.00483286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A2_M1007_g 0.0414634f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_54 VPB A2 0.00812361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_Y_c_288_n 0.0094557f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.12
cc_56 VPB N_Y_c_289_n 0.0348765f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.455
cc_57 VPB N_Y_c_290_n 0.00524858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_Y_c_291_n 0.021965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB Y 0.0084656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_119_392#_c_363_n 0.0214994f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_61 VPB N_A_119_392#_c_364_n 0.00378342f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_62 VPB N_A_369_392#_c_388_n 0.00275585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_369_392#_c_389_n 0.00881223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_369_392#_c_390_n 0.0348765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_369_392#_c_391_n 0.0146198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_369_392#_c_392_n 0.00797468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_431_n 0.00976602f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.69
cc_68 VPB N_VPWR_c_432_n 0.0832085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_433_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.285
cc_70 VPB N_VPWR_c_434_n 0.0207426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_430_n 0.0704432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_C1_M1001_g N_C2_M1011_g 0.023964f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_73 N_C1_c_73_n C2 6.88337e-19 $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_74 N_C1_c_74_n C2 0.0264482f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_75 N_C1_c_73_n N_C2_c_103_n 0.041753f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_76 N_C1_c_74_n N_C2_c_103_n 0.00286882f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_77 N_C1_c_75_n N_C2_c_104_n 0.041753f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_78 N_C1_M1001_g N_Y_c_288_n 8.84614e-19 $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_79 N_C1_c_73_n N_Y_c_288_n 4.87918e-19 $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_80 N_C1_c_74_n N_Y_c_288_n 0.0264502f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_81 N_C1_M1001_g N_Y_c_289_n 0.0118657f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_82 N_C1_c_75_n N_Y_c_283_n 0.00793201f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_83 N_C1_M1001_g N_Y_c_298_n 0.0131783f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_84 N_C1_c_74_n N_Y_c_298_n 0.0113214f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_85 N_C1_c_74_n N_Y_c_300_n 0.00942884f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_86 N_C1_c_75_n N_Y_c_300_n 0.00806212f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_87 N_C1_c_73_n N_Y_c_284_n 0.00412259f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_88 N_C1_c_74_n N_Y_c_284_n 0.026382f $X=0.43 $Y=1.285 $X2=0 $Y2=0
cc_89 N_C1_c_75_n N_Y_c_284_n 7.15802e-19 $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_90 N_C1_M1001_g N_A_119_392#_c_364_n 0.003398f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_91 N_C1_M1001_g N_VPWR_c_432_n 0.005209f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_92 N_C1_M1001_g N_VPWR_c_430_n 0.00987672f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_93 N_C1_c_75_n N_VGND_c_469_n 0.00434272f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_94 N_C1_c_75_n N_VGND_c_470_n 0.00126064f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_95 N_C1_c_75_n N_VGND_c_471_n 0.00437003f $X=0.43 $Y=1.12 $X2=0 $Y2=0
cc_96 N_C2_c_103_n N_B2_c_141_n 0.00733596f $X=1.15 $Y=1.285 $X2=0 $Y2=0
cc_97 N_C2_M1011_g N_Y_c_289_n 6.25319e-19 $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_98 N_C2_c_104_n N_Y_c_283_n 0.00159871f $X=1.075 $Y=1.12 $X2=0 $Y2=0
cc_99 N_C2_M1011_g N_Y_c_298_n 0.0166675f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_100 C2 N_Y_c_298_n 0.0090993f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_C2_c_103_n N_Y_c_298_n 0.00233214f $X=1.15 $Y=1.285 $X2=0 $Y2=0
cc_102 C2 N_Y_c_300_n 0.0237068f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_C2_c_103_n N_Y_c_300_n 0.00216104f $X=1.15 $Y=1.285 $X2=0 $Y2=0
cc_104 N_C2_c_104_n N_Y_c_300_n 0.0178302f $X=1.075 $Y=1.12 $X2=0 $Y2=0
cc_105 N_C2_M1011_g N_Y_c_290_n 0.00466492f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_106 C2 N_Y_c_291_n 0.0157066f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_C2_c_103_n N_Y_c_291_n 0.00144582f $X=1.15 $Y=1.285 $X2=0 $Y2=0
cc_108 C2 Y 0.0526461f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_C2_c_103_n Y 0.00765712f $X=1.15 $Y=1.285 $X2=0 $Y2=0
cc_110 N_C2_c_104_n Y 0.00440102f $X=1.075 $Y=1.12 $X2=0 $Y2=0
cc_111 N_C2_M1011_g N_A_119_392#_c_366_n 0.0129722f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_112 N_C2_M1011_g N_A_119_392#_c_363_n 0.0137576f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_113 N_C2_M1011_g N_A_119_392#_c_364_n 0.0019123f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_114 N_C2_M1011_g N_VPWR_c_432_n 0.00333896f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_115 N_C2_M1011_g N_VPWR_c_430_n 0.00428385f $X=1.005 $Y=2.46 $X2=0 $Y2=0
cc_116 N_C2_c_104_n N_VGND_c_469_n 0.00383152f $X=1.075 $Y=1.12 $X2=0 $Y2=0
cc_117 N_C2_c_104_n N_VGND_c_470_n 0.0102512f $X=1.075 $Y=1.12 $X2=0 $Y2=0
cc_118 N_C2_c_104_n N_VGND_c_471_n 0.00369533f $X=1.075 $Y=1.12 $X2=0 $Y2=0
cc_119 N_B2_M1009_g N_B1_M1010_g 0.0244331f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_120 N_B2_c_137_n N_B1_c_176_n 0.0205102f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_121 N_B2_c_138_n N_B1_c_177_n 0.0205102f $X=2.14 $Y=1.625 $X2=0 $Y2=0
cc_122 N_B2_c_139_n N_B1_c_178_n 0.0205102f $X=2.14 $Y=1.79 $X2=0 $Y2=0
cc_123 B2 B1 0.0438819f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B2_c_141_n B1 0.00410205f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_125 B2 N_B1_c_180_n 8.23261e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B2_c_141_n N_B1_c_180_n 0.0205102f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_127 N_B2_M1009_g N_Y_c_290_n 0.00429611f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_128 B2 N_Y_c_290_n 4.44645e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B2_M1009_g N_Y_c_291_n 0.00112371f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_130 N_B2_c_137_n N_Y_c_285_n 0.0013851f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_131 N_B2_c_137_n N_Y_c_323_n 0.0132291f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_132 B2 N_Y_c_323_n 0.0233092f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_133 N_B2_c_141_n N_Y_c_323_n 0.00112191f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_134 N_B2_c_137_n Y 0.00508329f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_135 B2 Y 0.0496775f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B2_c_141_n Y 0.00350374f $X=2.14 $Y=1.285 $X2=0 $Y2=0
cc_137 N_B2_c_138_n Y 0.00350374f $X=2.14 $Y=1.625 $X2=0 $Y2=0
cc_138 N_B2_M1009_g N_A_119_392#_c_363_n 0.0163065f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_139 N_B2_M1009_g N_A_369_392#_c_393_n 0.0131585f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_140 B2 N_A_369_392#_c_393_n 0.0113019f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B2_M1009_g N_A_369_392#_c_391_n 0.0108312f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_142 N_B2_c_139_n N_A_369_392#_c_391_n 9.9377e-19 $X=2.14 $Y=1.79 $X2=0 $Y2=0
cc_143 B2 N_A_369_392#_c_391_n 0.0129339f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_144 N_B2_M1009_g N_VPWR_c_432_n 0.00333926f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_145 N_B2_M1009_g N_VPWR_c_430_n 0.00428387f $X=2.215 $Y=2.46 $X2=0 $Y2=0
cc_146 N_B2_c_137_n N_VGND_c_468_n 0.00383152f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_147 N_B2_c_137_n N_VGND_c_470_n 0.00946983f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_148 N_B2_c_137_n N_VGND_c_471_n 0.00369533f $X=2.14 $Y=1.12 $X2=0 $Y2=0
cc_149 N_B1_c_177_n N_A1_c_216_n 0.0111092f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_150 N_B1_M1010_g N_A1_M1008_g 0.0125401f $X=2.715 $Y=2.46 $X2=0 $Y2=0
cc_151 N_B1_c_178_n N_A1_c_217_n 0.0111092f $X=2.71 $Y=1.79 $X2=0 $Y2=0
cc_152 B1 N_A1_c_218_n 0.00258451f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B1_c_180_n N_A1_c_218_n 0.0111092f $X=2.71 $Y=1.285 $X2=0 $Y2=0
cc_154 B1 N_A1_c_219_n 0.0352122f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_c_180_n N_A1_c_219_n 0.00237949f $X=2.71 $Y=1.285 $X2=0 $Y2=0
cc_156 N_B1_c_176_n N_A1_c_220_n 0.00516683f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_157 N_B1_c_176_n N_Y_c_285_n 0.0157946f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_158 B1 N_Y_c_285_n 0.0262962f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_159 N_B1_c_180_n N_Y_c_285_n 0.00121333f $X=2.71 $Y=1.285 $X2=0 $Y2=0
cc_160 N_B1_M1010_g N_A_119_392#_c_363_n 0.00448675f $X=2.715 $Y=2.46 $X2=0
+ $Y2=0
cc_161 N_B1_M1010_g N_A_119_392#_c_371_n 0.00721229f $X=2.715 $Y=2.46 $X2=0
+ $Y2=0
cc_162 N_B1_M1010_g N_A_369_392#_c_393_n 0.0144961f $X=2.715 $Y=2.46 $X2=0 $Y2=0
cc_163 N_B1_c_178_n N_A_369_392#_c_393_n 4.32055e-19 $X=2.71 $Y=1.79 $X2=0 $Y2=0
cc_164 B1 N_A_369_392#_c_393_n 0.0202798f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B1_M1010_g N_A_369_392#_c_391_n 4.54422e-19 $X=2.715 $Y=2.46 $X2=0
+ $Y2=0
cc_166 N_B1_c_178_n N_A_369_392#_c_392_n 2.71489e-19 $X=2.71 $Y=1.79 $X2=0 $Y2=0
cc_167 B1 N_A_369_392#_c_392_n 0.00261022f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_168 N_B1_M1010_g N_VPWR_c_432_n 0.00517089f $X=2.715 $Y=2.46 $X2=0 $Y2=0
cc_169 N_B1_M1010_g N_VPWR_c_430_n 0.00979708f $X=2.715 $Y=2.46 $X2=0 $Y2=0
cc_170 N_B1_c_176_n N_VGND_c_468_n 0.00288916f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_171 N_B1_c_176_n N_VGND_c_470_n 7.41728e-19 $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_172 N_B1_c_176_n N_VGND_c_471_n 0.00359465f $X=2.71 $Y=1.12 $X2=0 $Y2=0
cc_173 N_A1_c_219_n N_A2_M1005_g 0.0074729f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_174 N_A1_c_220_n N_A2_M1005_g 0.0263949f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_175 N_A1_c_216_n N_A2_M1007_g 0.0263949f $X=3.305 $Y=1.61 $X2=0 $Y2=0
cc_176 N_A1_M1008_g N_A2_M1007_g 0.023632f $X=3.215 $Y=2.46 $X2=0 $Y2=0
cc_177 N_A1_c_218_n A2 4.05463e-19 $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_178 N_A1_c_219_n A2 0.0495144f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_179 N_A1_c_218_n N_A2_c_258_n 0.0263949f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_180 N_A1_c_218_n N_Y_c_285_n 0.00268566f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_181 N_A1_c_219_n N_Y_c_285_n 0.0149686f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_182 N_A1_c_220_n N_Y_c_285_n 0.0116062f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_183 N_A1_M1008_g N_A_119_392#_c_363_n 3.17612e-19 $X=3.215 $Y=2.46 $X2=0
+ $Y2=0
cc_184 N_A1_M1008_g N_A_369_392#_c_388_n 0.0118701f $X=3.215 $Y=2.46 $X2=0 $Y2=0
cc_185 N_A1_M1008_g N_A_369_392#_c_405_n 0.0136434f $X=3.215 $Y=2.46 $X2=0 $Y2=0
cc_186 N_A1_c_217_n N_A_369_392#_c_405_n 0.00112785f $X=3.305 $Y=1.79 $X2=0
+ $Y2=0
cc_187 N_A1_c_219_n N_A_369_392#_c_405_n 0.0407226f $X=3.32 $Y=1.285 $X2=0 $Y2=0
cc_188 N_A1_M1008_g N_A_369_392#_c_390_n 8.48253e-19 $X=3.215 $Y=2.46 $X2=0
+ $Y2=0
cc_189 N_A1_M1008_g N_A_369_392#_c_392_n 0.00196977f $X=3.215 $Y=2.46 $X2=0
+ $Y2=0
cc_190 N_A1_M1008_g N_VPWR_c_431_n 0.00230487f $X=3.215 $Y=2.46 $X2=0 $Y2=0
cc_191 N_A1_M1008_g N_VPWR_c_432_n 0.005209f $X=3.215 $Y=2.46 $X2=0 $Y2=0
cc_192 N_A1_M1008_g N_VPWR_c_430_n 0.00983523f $X=3.215 $Y=2.46 $X2=0 $Y2=0
cc_193 N_A1_c_220_n N_VGND_c_467_n 0.00222027f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_194 N_A1_c_220_n N_VGND_c_468_n 0.00432706f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_195 N_A1_c_220_n N_VGND_c_471_n 0.00819572f $X=3.305 $Y=1.12 $X2=0 $Y2=0
cc_196 N_A2_M1005_g N_Y_c_285_n 0.00174219f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_197 N_A2_M1007_g N_A_369_392#_c_388_n 8.8709e-19 $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_198 N_A2_M1007_g N_A_369_392#_c_405_n 0.0182002f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_199 N_A2_M1007_g N_A_369_392#_c_389_n 0.0013033f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_200 A2 N_A_369_392#_c_389_n 0.0252512f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_201 N_A2_c_258_n N_A_369_392#_c_389_n 0.00121003f $X=4.05 $Y=1.345 $X2=0
+ $Y2=0
cc_202 N_A2_M1007_g N_A_369_392#_c_390_n 0.0128569f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_203 N_A2_M1007_g N_VPWR_c_431_n 0.00989997f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_204 N_A2_M1007_g N_VPWR_c_434_n 0.005209f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_205 N_A2_M1007_g N_VPWR_c_430_n 0.00987818f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_206 N_A2_M1005_g N_VGND_c_467_n 0.0161695f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_207 A2 N_VGND_c_467_n 0.0184523f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A2_c_258_n N_VGND_c_467_n 0.00206909f $X=4.05 $Y=1.345 $X2=0 $Y2=0
cc_209 N_A2_M1005_g N_VGND_c_468_n 0.00383152f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_210 N_A2_M1005_g N_VGND_c_471_n 0.0075725f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_211 N_Y_c_298_n N_A_119_392#_M1001_d 0.00943905f $X=1.115 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_212 N_Y_c_298_n N_A_119_392#_c_366_n 0.0189268f $X=1.115 $Y=2.045 $X2=0 $Y2=0
cc_213 N_Y_M1011_d N_A_119_392#_c_363_n 0.00335038f $X=1.095 $Y=1.96 $X2=0 $Y2=0
cc_214 N_Y_c_291_n N_A_119_392#_c_363_n 0.0388717f $X=1.28 $Y=2.125 $X2=0 $Y2=0
cc_215 N_Y_c_289_n N_A_119_392#_c_364_n 0.0037133f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_216 N_Y_c_291_n N_A_369_392#_c_391_n 0.0681652f $X=1.28 $Y=2.125 $X2=0 $Y2=0
cc_217 N_Y_c_289_n N_VPWR_c_432_n 0.014549f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_218 N_Y_c_289_n N_VPWR_c_430_n 0.0119743f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_219 N_Y_c_300_n A_119_74# 0.0072096f $X=1.485 $Y=0.865 $X2=-0.19 $Y2=-0.245
cc_220 N_Y_c_300_n N_VGND_M1000_d 0.0162958f $X=1.485 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_221 N_Y_c_323_n N_VGND_M1000_d 0.0126943f $X=2.525 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_222 Y N_VGND_M1000_d 0.00918472f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_223 N_Y_c_285_n N_VGND_c_467_n 0.0207642f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_224 N_Y_c_285_n N_VGND_c_468_n 0.0395123f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_225 N_Y_c_283_n N_VGND_c_469_n 0.0144324f $X=0.305 $Y=0.515 $X2=0 $Y2=0
cc_226 N_Y_c_283_n N_VGND_c_470_n 0.00836615f $X=0.305 $Y=0.515 $X2=0 $Y2=0
cc_227 N_Y_c_300_n N_VGND_c_470_n 0.0349649f $X=1.485 $Y=0.865 $X2=0 $Y2=0
cc_228 N_Y_c_285_n N_VGND_c_470_n 0.00748454f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_229 N_Y_c_323_n N_VGND_c_470_n 0.024446f $X=2.525 $Y=0.64 $X2=0 $Y2=0
cc_230 Y N_VGND_c_470_n 0.0257144f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_231 N_Y_c_283_n N_VGND_c_471_n 0.0119472f $X=0.305 $Y=0.515 $X2=0 $Y2=0
cc_232 N_Y_c_300_n N_VGND_c_471_n 0.0179064f $X=1.485 $Y=0.865 $X2=0 $Y2=0
cc_233 N_Y_c_285_n N_VGND_c_471_n 0.0302537f $X=3.195 $Y=0.495 $X2=0 $Y2=0
cc_234 N_Y_c_323_n N_VGND_c_471_n 0.0130236f $X=2.525 $Y=0.64 $X2=0 $Y2=0
cc_235 Y N_VGND_c_471_n 0.00127411f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_236 N_Y_c_323_n A_461_74# 0.0072096f $X=2.525 $Y=0.64 $X2=-0.19 $Y2=-0.245
cc_237 N_A_119_392#_c_363_n N_A_369_392#_M1009_s 0.00266942f $X=2.325 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_238 N_A_119_392#_M1009_d N_A_369_392#_c_393_n 0.00884137f $X=2.305 $Y=1.96
+ $X2=0 $Y2=0
cc_239 N_A_119_392#_c_371_n N_A_369_392#_c_393_n 0.0189268f $X=2.49 $Y=2.465
+ $X2=0 $Y2=0
cc_240 N_A_119_392#_c_363_n N_A_369_392#_c_388_n 0.0039531f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_241 N_A_119_392#_c_363_n N_A_369_392#_c_391_n 0.0205035f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_242 N_A_119_392#_c_363_n N_VPWR_c_431_n 0.00275197f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_243 N_A_119_392#_c_363_n N_VPWR_c_432_n 0.111406f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_244 N_A_119_392#_c_364_n N_VPWR_c_432_n 0.0235512f $X=0.945 $Y=2.99 $X2=0
+ $Y2=0
cc_245 N_A_119_392#_c_363_n N_VPWR_c_430_n 0.0630647f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_246 N_A_119_392#_c_364_n N_VPWR_c_430_n 0.0126924f $X=0.945 $Y=2.99 $X2=0
+ $Y2=0
cc_247 N_A_369_392#_c_405_n N_VPWR_M1008_d 0.0071387f $X=3.875 $Y=2.045
+ $X2=-0.19 $Y2=1.66
cc_248 N_A_369_392#_c_388_n N_VPWR_c_431_n 0.0263057f $X=2.99 $Y=2.815 $X2=0
+ $Y2=0
cc_249 N_A_369_392#_c_405_n N_VPWR_c_431_n 0.0237567f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_250 N_A_369_392#_c_390_n N_VPWR_c_431_n 0.0433291f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_369_392#_c_388_n N_VPWR_c_432_n 0.014549f $X=2.99 $Y=2.815 $X2=0
+ $Y2=0
cc_252 N_A_369_392#_c_390_n N_VPWR_c_434_n 0.014549f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_253 N_A_369_392#_c_388_n N_VPWR_c_430_n 0.0119743f $X=2.99 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_A_369_392#_c_390_n N_VPWR_c_430_n 0.0119743f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0

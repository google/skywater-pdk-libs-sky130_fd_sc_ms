* File: sky130_fd_sc_ms__o41a_2.spice
* Created: Wed Sep  2 12:26:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o41a_2.pex.spice"
.subckt sky130_fd_sc_ms__o41a_2  VNB VPB A1 A2 A3 A4 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A1_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_27_74#_M1013_d N_A2_M1013_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A3_M1003_g N_A_27_74#_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.21645 AS=0.1036 PD=1.325 PS=1.02 NRD=25.944 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1000 N_A_27_74#_M1000_d N_A4_M1000_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.21645 PD=1.035 PS=1.325 NRD=2.424 NRS=23.508 M=1 R=4.93333
+ SA=75001.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_A_431_368#_M1009_d N_B1_M1009_g N_A_27_74#_M1000_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.10915 PD=2.19 PS=1.035 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_431_368#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1001_d N_A_431_368#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1002 A_119_368# N_A1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90003.7
+ A=0.2016 P=2.6 MULT=1
MM1005 A_203_368# N_A2_M1005_g A_119_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1008 A_317_368# N_A3_M1008_g A_203_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=24.6053 M=1 R=6.22222 SA=90001.2
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1006 N_A_431_368#_M1006_d N_A4_M1006_g A_317_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.223789 AS=0.2184 PD=1.59547 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222
+ SA=90001.8 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_A_431_368#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.5 AS=0.199811 PD=2.0283 PS=1.42453 NRD=0 NRS=22.9702 M=1 R=5.55556
+ SA=90002.3 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1010_d N_A_431_368#_M1010_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.56 PD=1.39 PS=2.2717 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1010_d N_A_431_368#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__o41a_2.pxi.spice"
*
.ends
*
*

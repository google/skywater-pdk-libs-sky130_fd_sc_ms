* NGSPICE file created from sky130_fd_sc_ms__nor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nor3_2 A B C VGND VNB VPB VPWR Y
M1000 a_27_368# C Y VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=8.38e+06u as=3.584e+11p ps=2.88e+06u
M1001 a_309_368# B a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.384e+11p pd=5.62e+06u as=0p ps=0u
M1002 Y C a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_309_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.248e+11p ps=2.82e+06u
M1004 a_27_368# B a_309_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_309_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C Y VNB nlowvt w=740000u l=150000u
+  ad=9.176e+11p pd=5.44e+06u as=4.699e+11p ps=4.23e+06u
M1007 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* NGSPICE file created from sky130_fd_sc_ms__dlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_84_48# a_334_338# a_286_392# VPB pshort w=1e+06u l=180000u
+  ad=3.991e+11p pd=3.21e+06u as=2.4e+11p ps=2.48e+06u
M1001 VGND a_27_74# a_491_124# VNB nlowvt w=420000u l=150000u
+  ad=1.78525e+12p pd=1.468e+07u as=2.3775e+11p ps=2.39e+06u
M1002 VPWR a_27_74# a_527_508# VPB pshort w=420000u l=180000u
+  ad=3.0253e+12p pd=1.906e+07u as=1.008e+11p ps=1.32e+06u
M1003 VPWR a_84_48# a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 GCLK a_1047_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.216e+11p pd=5.59e+06u as=0p ps=0u
M1005 a_1047_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1006 GCLK a_1047_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 GCLK a_1047_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1047_368# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.416e+11p pd=2.85e+06u as=0p ps=0u
M1009 VGND a_1047_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_1047_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_491_124# a_334_338# a_84_48# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.587e+11p ps=2.25e+06u
M1012 VPWR CLK a_334_54# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 VGND a_1047_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_27_74# a_1047_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_334_338# a_334_54# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 GCLK a_1047_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_286_80# GATE VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 a_84_48# a_334_54# a_286_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND CLK a_334_54# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.333e+11p ps=2.19e+06u
M1020 VGND a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1021 a_1047_368# a_27_74# a_1047_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 VPWR a_1047_368# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_286_392# GATE VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_527_508# a_334_54# a_84_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_334_338# a_334_54# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.675e+11p pd=2.66e+06u as=0p ps=0u
.ends


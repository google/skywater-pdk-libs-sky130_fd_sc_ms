* File: sky130_fd_sc_ms__a2111oi_1.spice
* Created: Wed Sep  2 11:49:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2111oi_1.pex.spice"
.subckt sky130_fd_sc_ms__a2111oi_1  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_D1_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_C1_M1006_g N_Y_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.185
+ AS=0.1036 PD=1.24 PS=1.02 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.185 PD=1.02 PS=1.24 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 A_461_74# N_A1_M1002_g N_Y_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.7 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_461_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75002.2 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1007 A_159_368# N_D1_M1007_g N_Y_M1007_s VPB PSHORT L=0.18 W=1.12 AD=0.1176
+ AS=0.2912 PD=1.33 PS=2.76 NRD=8.7862 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90002.2
+ A=0.2016 P=2.6 MULT=1
MM1004 A_237_368# N_C1_M1004_g A_159_368# VPB PSHORT L=0.18 W=1.12 AD=0.2016
+ AS=0.1176 PD=1.48 PS=1.33 NRD=21.9852 NRS=8.7862 M=1 R=6.22222 SA=90000.6
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1005 N_A_345_368#_M1005_d N_B1_M1005_g A_237_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.2016 PD=1.48 PS=1.48 NRD=2.6201 NRS=21.9852 M=1 R=6.22222
+ SA=90001.1 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_345_368#_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.2016 PD=1.48 PS=1.48 NRD=2.6201 NRS=11.426 M=1 R=6.22222
+ SA=90001.6 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1000 N_A_345_368#_M1000_d N_A2_M1000_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2016 PD=2.76 PS=1.48 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90002.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__a2111oi_1.pxi.spice"
*
.ends
*
*

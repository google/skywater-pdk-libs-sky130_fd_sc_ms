* File: sky130_fd_sc_ms__o221ai_1.spice
* Created: Wed Sep  2 12:23:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o221ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o221ai_1  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1009 N_A_114_74#_M1009_d N_C1_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 N_A_114_74#_M1003_d N_B1_M1003_g N_A_239_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1001 N_A_239_74#_M1001_d N_B2_M1001_g N_A_114_74#_M1003_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_239_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2368 AS=0.1295 PD=1.38 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1006 N_A_239_74#_M1006_d N_A1_M1006_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2368 PD=2.05 PS=1.38 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_C1_M1002_g N_Y_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.4088 AS=0.3136 PD=1.85 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1004 A_327_368# N_B1_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.4088 PD=1.36 PS=1.85 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90001.8
+ A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1007_d N_B2_M1007_g A_327_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90001.5 SB=90001.3
+ A=0.2016 P=2.6 MULT=1
MM1005 A_525_368# N_A2_M1005_g N_Y_M1007_d VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=20.2122 M=1 R=6.22222 SA=90002.1
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_525_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90002.7 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o221ai_1.pxi.spice"
*
.ends
*
*

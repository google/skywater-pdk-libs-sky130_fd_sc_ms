* File: sky130_fd_sc_ms__nor3_4.pxi.spice
* Created: Wed Sep  2 12:16:11 2020
* 
x_PM_SKY130_FD_SC_MS__NOR3_4%A N_A_M1008_g N_A_M1004_g N_A_M1016_g N_A_M1009_g
+ N_A_c_115_n N_A_M1012_g N_A_c_116_n N_A_M1014_g N_A_c_163_p N_A_c_108_n
+ N_A_c_140_p N_A_c_124_p N_A_c_109_n N_A_c_110_n N_A_c_111_n N_A_c_125_p A A A
+ N_A_c_112_n N_A_c_122_p PM_SKY130_FD_SC_MS__NOR3_4%A
x_PM_SKY130_FD_SC_MS__NOR3_4%B N_B_M1003_g N_B_c_238_n N_B_M1006_g N_B_c_239_n
+ N_B_c_240_n N_B_M1013_g N_B_M1005_g N_B_M1010_g N_B_M1011_g N_B_c_244_n
+ N_B_c_245_n N_B_c_257_n N_B_c_246_n B B N_B_c_247_n N_B_c_248_n N_B_c_249_n
+ N_B_c_250_n N_B_c_251_n B B N_B_c_252_n PM_SKY130_FD_SC_MS__NOR3_4%B
x_PM_SKY130_FD_SC_MS__NOR3_4%C N_C_M1000_g N_C_c_356_n N_C_c_357_n N_C_M1002_g
+ N_C_M1001_g N_C_c_359_n N_C_M1007_g N_C_M1015_g N_C_c_361_n N_C_c_362_n
+ N_C_M1017_g N_C_c_363_n N_C_c_364_n N_C_c_365_n N_C_c_366_n C C C C
+ N_C_c_368_n PM_SKY130_FD_SC_MS__NOR3_4%C
x_PM_SKY130_FD_SC_MS__NOR3_4%A_27_368# N_A_27_368#_M1008_d N_A_27_368#_M1009_d
+ N_A_27_368#_M1005_d N_A_27_368#_M1011_d N_A_27_368#_M1014_d
+ N_A_27_368#_c_461_n N_A_27_368#_c_462_n N_A_27_368#_c_475_n
+ N_A_27_368#_c_463_n N_A_27_368#_c_480_n N_A_27_368#_c_485_n
+ N_A_27_368#_c_464_n N_A_27_368#_c_487_n N_A_27_368#_c_465_n
+ N_A_27_368#_c_466_n N_A_27_368#_c_467_n N_A_27_368#_c_494_n
+ N_A_27_368#_c_495_n N_A_27_368#_c_496_n N_A_27_368#_c_468_n
+ PM_SKY130_FD_SC_MS__NOR3_4%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR3_4%VPWR N_VPWR_M1008_s N_VPWR_M1012_s N_VPWR_c_548_n
+ N_VPWR_c_549_n VPWR N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_547_n N_VPWR_c_554_n N_VPWR_c_555_n PM_SKY130_FD_SC_MS__NOR3_4%VPWR
x_PM_SKY130_FD_SC_MS__NOR3_4%A_298_368# N_A_298_368#_M1003_s
+ N_A_298_368#_M1001_s N_A_298_368#_M1017_s N_A_298_368#_M1010_s
+ N_A_298_368#_c_616_n N_A_298_368#_c_617_n N_A_298_368#_c_618_n
+ PM_SKY130_FD_SC_MS__NOR3_4%A_298_368#
x_PM_SKY130_FD_SC_MS__NOR3_4%Y N_Y_M1004_s N_Y_M1006_d N_Y_M1002_d N_Y_M1000_d
+ N_Y_M1015_d N_Y_c_660_n N_Y_c_661_n N_Y_c_662_n N_Y_c_698_n N_Y_c_663_n
+ N_Y_c_664_n N_Y_c_668_n N_Y_c_665_n N_Y_c_666_n N_Y_c_717_n N_Y_c_669_n
+ N_Y_c_670_n Y PM_SKY130_FD_SC_MS__NOR3_4%Y
x_PM_SKY130_FD_SC_MS__NOR3_4%VGND N_VGND_M1004_d N_VGND_M1016_d N_VGND_M1013_s
+ N_VGND_M1007_s N_VGND_c_772_n N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n
+ N_VGND_c_776_n N_VGND_c_777_n VGND N_VGND_c_778_n N_VGND_c_779_n
+ N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n N_VGND_c_784_n
+ PM_SKY130_FD_SC_MS__NOR3_4%VGND
cc_1 VNB N_A_M1004_g 0.0307057f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1016_g 0.024721f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.74
cc_3 VNB N_A_c_108_n 0.00103091f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_4 VNB N_A_c_109_n 0.0027193f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_5 VNB N_A_c_110_n 0.16813f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_6 VNB N_A_c_111_n 0.0357942f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_7 VNB N_A_c_112_n 0.0479327f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.515
cc_8 VNB N_B_c_238_n 0.0156992f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_9 VNB N_B_c_239_n 0.0193149f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.74
cc_10 VNB N_B_c_240_n 0.0161096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_M1005_g 0.00903762f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=1.77
cc_12 VNB N_B_M1010_g 0.00789458f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.4
cc_13 VNB N_B_M1011_g 0.00773158f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_14 VNB N_B_c_244_n 0.0111069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_245_n 0.0256494f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=2.02
cc_16 VNB N_B_c_246_n 0.0147148f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_17 VNB N_B_c_247_n 0.0114101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_248_n 0.0861994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_249_n 0.0037819f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.515
cc_20 VNB N_B_c_250_n 0.00684755f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_21 VNB N_B_c_251_n 0.00930406f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=2.045
cc_22 VNB N_B_c_252_n 0.00306353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_356_n 0.00870882f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_24 VNB N_C_c_357_n 0.0055414f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_C_M1002_g 0.0363229f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.35
cc_26 VNB N_C_c_359_n 0.00232143f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_27 VNB N_C_M1007_g 0.0396304f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=2.4
cc_28 VNB N_C_c_361_n 0.0100449f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_29 VNB N_C_c_362_n 0.00752287f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_30 VNB N_C_c_363_n 0.0732211f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=2.02
cc_31 VNB N_C_c_364_n 0.0021832f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_32 VNB N_C_c_365_n 0.00435531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_C_c_366_n 0.0194928f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_34 VNB C 0.00924763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C_c_368_n 0.14102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_547_n 0.283096f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_37 VNB N_Y_c_660_n 0.0103011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_661_n 0.00348993f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=1.77
cc_39 VNB N_Y_c_662_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=1.77
cc_40 VNB N_Y_c_663_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=5.805 $Y2=2.105
cc_41 VNB N_Y_c_664_n 0.0314239f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=2.02
cc_42 VNB N_Y_c_665_n 0.00896499f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_43 VNB N_Y_c_666_n 0.00226854f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_44 VNB Y 0.00248769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_772_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.68
cc_46 VNB N_VGND_c_773_n 0.0505972f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_47 VNB N_VGND_c_774_n 0.00900483f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=2.4
cc_48 VNB N_VGND_c_775_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.92
cc_49 VNB N_VGND_c_776_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_50 VNB N_VGND_c_777_n 0.0120529f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.255
cc_51 VNB N_VGND_c_778_n 0.019013f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_52 VNB N_VGND_c_779_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_53 VNB N_VGND_c_780_n 0.0915322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_781_n 0.388363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_782_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.515
cc_56 VNB N_VGND_c_783_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_57 VNB N_VGND_c_784_n 0.00596278f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.045
cc_58 VPB N_A_M1008_g 0.0285106f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.4
cc_59 VPB N_A_M1009_g 0.0205508f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_60 VPB N_A_c_115_n 0.0159622f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=1.77
cc_61 VPB N_A_c_116_n 0.0209495f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=1.77
cc_62 VPB N_A_c_108_n 0.0014948f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_63 VPB N_A_c_109_n 0.00149128f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_64 VPB N_A_c_111_n 0.0206988f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=1.515
cc_65 VPB N_A_c_112_n 0.00538875f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=1.515
cc_66 VPB N_B_M1003_g 0.0238324f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_67 VPB N_B_M1005_g 0.0219647f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=1.77
cc_68 VPB N_B_M1010_g 0.0201742f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=2.4
cc_69 VPB N_B_M1011_g 0.0218281f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_70 VPB N_B_c_257_n 0.00155728f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_71 VPB N_B_c_247_n 0.00569486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_C_M1000_g 0.0228832f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.4
cc_73 VPB N_C_c_356_n 0.00857758f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_74 VPB N_C_c_357_n 0.00415775f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_75 VPB N_C_M1001_g 0.0218674f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.68
cc_76 VPB N_C_c_359_n 0.00330321f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_77 VPB N_C_M1015_g 0.0218304f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.92
cc_78 VPB N_C_c_361_n 0.0115314f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_79 VPB N_C_c_362_n 0.00969026f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_80 VPB N_C_M1017_g 0.0214009f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=2.255
cc_81 VPB N_C_c_364_n 0.00318934f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_82 VPB N_C_c_365_n 0.00224265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_27_368#_c_461_n 0.0295461f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=2.4
cc_84 VPB N_A_27_368#_c_462_n 0.0197196f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=2.4
cc_85 VPB N_A_27_368#_c_463_n 0.00202145f $X=-0.19 $Y=1.66 $X2=3.85 $Y2=2.255
cc_86 VPB N_A_27_368#_c_464_n 0.00211347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_27_368#_c_465_n 0.0303776f $X=-0.19 $Y=1.66 $X2=3.935 $Y2=2.255
cc_88 VPB N_A_27_368#_c_466_n 0.0190607f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.95
cc_89 VPB N_A_27_368#_c_467_n 0.00708086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_368#_c_468_n 0.0071123f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=2.045
cc_91 VPB N_VPWR_c_548_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=1.35
cc_92 VPB N_VPWR_c_549_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.68
cc_93 VPB N_VPWR_c_550_n 0.0178682f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=1.77
cc_94 VPB N_VPWR_c_551_n 0.116778f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=2.4
cc_95 VPB N_VPWR_c_552_n 0.0177091f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=2.02
cc_96 VPB N_VPWR_c_547_n 0.0745626f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_97 VPB N_VPWR_c_554_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_555_n 0.00601813f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=1.515
cc_99 VPB N_A_298_368#_c_616_n 0.00997561f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.68
cc_100 VPB N_A_298_368#_c_617_n 0.00227131f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=2.4
cc_101 VPB N_A_298_368#_c_618_n 0.00194561f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_102 VPB N_Y_c_668_n 0.00849352f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_103 VPB N_Y_c_669_n 0.00828589f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.95
cc_104 VPB N_Y_c_670_n 5.90677e-19 $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.95
cc_105 A N_B_M1003_g 0.00440718f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_106 N_A_c_122_p N_B_M1003_g 0.0159278f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_107 N_A_M1016_g N_B_c_238_n 0.0209692f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_c_124_p N_B_M1005_g 0.0128424f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_109 N_A_c_125_p N_B_M1005_g 0.0029722f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_110 N_A_c_124_p N_B_M1010_g 0.0116635f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_111 N_A_c_124_p N_B_M1011_g 0.0149678f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_112 N_A_c_111_n N_B_M1011_g 0.0434836f $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_113 N_A_M1016_g N_B_c_244_n 0.00879955f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_c_108_n N_B_c_257_n 0.0130906f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_115 A N_B_c_257_n 7.95053e-19 $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_116 N_A_c_112_n N_B_c_257_n 0.00150439f $X=0.935 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A_c_122_p N_B_c_257_n 0.0162196f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_118 N_A_c_108_n N_B_c_246_n 0.00231165f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A_c_112_n N_B_c_246_n 0.0240797f $X=0.935 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A_M1009_g N_B_c_247_n 0.0240797f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_c_122_p N_B_c_247_n 7.44609e-19 $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_122 N_A_c_109_n N_B_c_248_n 0.00328264f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_123 N_A_c_110_n N_B_c_248_n 0.0110664f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_124 N_A_c_140_p N_B_c_251_n 0.00799671f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_125 A N_B_c_251_n 0.00663543f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_126 N_A_c_140_p N_C_M1000_g 0.0144158f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_127 A N_C_M1000_g 0.0051931f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_128 N_A_c_140_p N_C_M1001_g 0.0132684f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_129 N_A_c_140_p N_C_M1015_g 0.0132684f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_130 N_A_c_125_p N_C_M1015_g 7.87653e-19 $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_131 N_A_c_140_p N_C_c_361_n 8.81995e-19 $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_132 N_A_c_140_p N_C_M1017_g 0.00934032f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_133 N_A_c_124_p N_C_M1017_g 3.15447e-19 $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_134 N_A_c_125_p N_C_M1017_g 0.00923418f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_135 N_A_c_109_n C 0.0276579f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_136 N_A_c_110_n C 0.00275385f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_137 N_A_c_109_n N_C_c_368_n 2.67785e-19 $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_138 N_A_c_110_n N_C_c_368_n 0.0179842f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_139 N_A_c_122_p N_A_27_368#_M1009_d 0.00791461f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_140 N_A_c_124_p N_A_27_368#_M1005_d 0.00321662f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_141 N_A_c_124_p N_A_27_368#_M1011_d 0.00761058f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_142 N_A_M1008_g N_A_27_368#_c_461_n 9.84618e-19 $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_c_108_n N_A_27_368#_c_461_n 0.00119904f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A_M1008_g N_A_27_368#_c_462_n 9.71144e-19 $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_M1008_g N_A_27_368#_c_475_n 0.0164451f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_M1009_g N_A_27_368#_c_475_n 0.0110002f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_c_163_p N_A_27_368#_c_475_n 0.018363f $X=0.77 $Y=1.92 $X2=0 $Y2=0
cc_148 N_A_c_112_n N_A_27_368#_c_475_n 2.39739e-19 $X=0.935 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A_c_122_p N_A_27_368#_c_475_n 0.00726436f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_150 N_A_c_140_p N_A_27_368#_c_480_n 0.117054f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_151 N_A_c_124_p N_A_27_368#_c_480_n 0.0179f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_152 N_A_c_125_p N_A_27_368#_c_480_n 0.0082338f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_153 A N_A_27_368#_c_480_n 0.0131482f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_154 N_A_c_122_p N_A_27_368#_c_480_n 0.00951666f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_155 N_A_c_124_p N_A_27_368#_c_485_n 0.0356639f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_156 N_A_c_115_n N_A_27_368#_c_464_n 2.98687e-19 $X=5.775 $Y=1.77 $X2=0 $Y2=0
cc_157 N_A_c_115_n N_A_27_368#_c_487_n 0.0109315f $X=5.775 $Y=1.77 $X2=0 $Y2=0
cc_158 N_A_c_116_n N_A_27_368#_c_487_n 0.0164145f $X=6.225 $Y=1.77 $X2=0 $Y2=0
cc_159 N_A_c_124_p N_A_27_368#_c_487_n 0.0252862f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_160 N_A_c_111_n N_A_27_368#_c_487_n 2.29439e-19 $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A_c_116_n N_A_27_368#_c_465_n 9.80186e-19 $X=6.225 $Y=1.77 $X2=0 $Y2=0
cc_162 N_A_c_109_n N_A_27_368#_c_465_n 0.00125279f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_163 N_A_c_116_n N_A_27_368#_c_466_n 9.71144e-19 $X=6.225 $Y=1.77 $X2=0 $Y2=0
cc_164 N_A_c_122_p N_A_27_368#_c_494_n 0.0151841f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_165 N_A_c_124_p N_A_27_368#_c_495_n 0.0141652f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_166 N_A_c_124_p N_A_27_368#_c_496_n 0.0126293f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_167 N_A_c_163_p N_VPWR_M1008_s 0.00217078f $X=0.77 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A_c_124_p N_VPWR_M1012_s 0.00202466f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_169 N_A_c_109_n N_VPWR_M1012_s 2.90423e-19 $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_170 N_A_M1008_g N_VPWR_c_548_n 0.0110077f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_M1009_g N_VPWR_c_548_n 0.00829914f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_c_115_n N_VPWR_c_549_n 0.00780794f $X=5.775 $Y=1.77 $X2=0 $Y2=0
cc_173 N_A_c_116_n N_VPWR_c_549_n 0.0107582f $X=6.225 $Y=1.77 $X2=0 $Y2=0
cc_174 N_A_M1008_g N_VPWR_c_550_n 0.00460063f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_M1009_g N_VPWR_c_551_n 0.00460063f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A_c_115_n N_VPWR_c_551_n 0.00460063f $X=5.775 $Y=1.77 $X2=0 $Y2=0
cc_177 N_A_c_116_n N_VPWR_c_552_n 0.00460063f $X=6.225 $Y=1.77 $X2=0 $Y2=0
cc_178 N_A_M1008_g N_VPWR_c_547_n 0.00459562f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_M1009_g N_VPWR_c_547_n 0.00455949f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_c_115_n N_VPWR_c_547_n 0.00450916f $X=5.775 $Y=1.77 $X2=0 $Y2=0
cc_181 N_A_c_116_n N_VPWR_c_547_n 0.00454512f $X=6.225 $Y=1.77 $X2=0 $Y2=0
cc_182 N_A_c_140_p N_A_298_368#_M1003_s 0.00240508f $X=3.85 $Y=2.255 $X2=-0.19
+ $Y2=-0.245
cc_183 A N_A_298_368#_M1003_s 0.0116967f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_184 N_A_c_122_p N_A_298_368#_M1003_s 0.0025653f $X=1.625 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_c_140_p N_A_298_368#_M1001_s 0.0070381f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_186 N_A_c_124_p N_A_298_368#_M1017_s 0.00748795f $X=5.805 $Y=2.105 $X2=0
+ $Y2=0
cc_187 N_A_c_125_p N_A_298_368#_M1017_s 0.00363072f $X=3.935 $Y=2.105 $X2=0
+ $Y2=0
cc_188 N_A_c_124_p N_A_298_368#_M1010_s 0.00321012f $X=5.805 $Y=2.105 $X2=0
+ $Y2=0
cc_189 N_A_c_115_n N_A_298_368#_c_618_n 3.14035e-19 $X=5.775 $Y=1.77 $X2=0 $Y2=0
cc_190 N_A_c_140_p N_Y_M1000_d 0.00677658f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_191 N_A_c_140_p N_Y_M1015_d 0.00677658f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_192 N_A_M1016_g N_Y_c_660_n 0.0148128f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_c_108_n N_Y_c_660_n 0.00446029f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A_c_112_n N_Y_c_660_n 0.00124519f $X=0.935 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A_M1004_g N_Y_c_661_n 0.00582181f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_M1016_g N_Y_c_661_n 0.00129659f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_c_108_n N_Y_c_661_n 0.0239178f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A_c_112_n N_Y_c_661_n 8.68732e-19 $X=0.935 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A_M1016_g N_Y_c_662_n 6.36864e-19 $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_c_109_n N_Y_c_664_n 0.00639395f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_201 N_A_c_110_n N_Y_c_664_n 0.00389741f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_202 N_A_c_140_p N_Y_c_668_n 0.00510648f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_203 N_A_c_124_p N_Y_c_668_n 0.0714309f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_204 N_A_c_109_n N_Y_c_668_n 0.00559649f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_205 N_A_c_111_n N_Y_c_668_n 5.18582e-19 $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A_c_125_p N_Y_c_668_n 0.0082338f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_207 N_A_c_109_n N_Y_c_665_n 0.0204255f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_208 N_A_c_110_n N_Y_c_665_n 0.00556001f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_209 N_A_c_140_p N_Y_c_669_n 0.0949959f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_210 N_A_M1004_g Y 0.00840664f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_M1016_g Y 0.00914611f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_M1004_g N_VGND_c_773_n 0.00647381f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_M1016_g N_VGND_c_774_n 0.00625757f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_M1004_g N_VGND_c_778_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_M1016_g N_VGND_c_778_n 0.00445602f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_c_109_n N_VGND_c_780_n 0.0148959f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_217 N_A_c_110_n N_VGND_c_780_n 0.0101867f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_218 N_A_M1004_g N_VGND_c_781_n 0.00824041f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_M1016_g N_VGND_c_781_n 0.00857802f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_c_109_n N_VGND_c_781_n 0.0120047f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_221 N_A_c_110_n N_VGND_c_781_n 0.00834893f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_222 N_B_c_250_n N_C_c_356_n 0.00686768f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_223 N_B_M1003_g N_C_c_357_n 0.0375592f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_224 N_B_c_239_n N_C_c_357_n 0.00558626f $X=1.85 $Y=1.26 $X2=0 $Y2=0
cc_225 N_B_c_257_n N_C_c_357_n 0.00100564f $X=1.475 $Y=1.435 $X2=0 $Y2=0
cc_226 N_B_c_247_n N_C_c_357_n 0.007253f $X=1.475 $Y=1.68 $X2=0 $Y2=0
cc_227 N_B_c_251_n N_C_c_357_n 0.00686768f $X=2.045 $Y=1.35 $X2=0 $Y2=0
cc_228 N_B_c_240_n N_C_M1002_g 0.0257968f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_229 N_B_c_249_n N_C_M1002_g 0.019948f $X=2.585 $Y=1.35 $X2=0 $Y2=0
cc_230 N_B_c_245_n N_C_M1007_g 0.0203249f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_231 N_B_c_252_n N_C_M1007_g 2.71203e-19 $X=2.755 $Y=1.35 $X2=0 $Y2=0
cc_232 N_B_c_245_n N_C_c_362_n 0.0163161f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_233 N_B_M1005_g N_C_c_363_n 0.0449663f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_234 N_B_c_245_n N_C_c_363_n 0.0216801f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_235 N_B_c_248_n N_C_c_363_n 0.00958311f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_236 N_B_c_252_n N_C_c_364_n 0.00309543f $X=2.755 $Y=1.35 $X2=0 $Y2=0
cc_237 N_B_c_248_n C 0.00105275f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_238 N_B_c_248_n N_C_c_368_n 0.0205126f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_239 N_B_M1003_g N_A_27_368#_c_463_n 0.00554736f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_240 N_B_M1003_g N_A_27_368#_c_480_n 0.011853f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B_M1005_g N_A_27_368#_c_480_n 0.0112434f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_242 N_B_M1010_g N_A_27_368#_c_485_n 0.010732f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_243 N_B_M1011_g N_A_27_368#_c_485_n 0.0108952f $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_244 N_B_M1011_g N_A_27_368#_c_464_n 2.98687e-19 $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B_M1003_g N_A_27_368#_c_494_n 0.00493036f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B_M1005_g N_A_27_368#_c_495_n 0.0060734f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B_M1003_g N_VPWR_c_548_n 4.76121e-19 $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_248 N_B_M1011_g N_VPWR_c_549_n 3.9902e-19 $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_249 N_B_M1003_g N_VPWR_c_551_n 0.00387245f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_250 N_B_M1005_g N_VPWR_c_551_n 0.00333926f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_251 N_B_M1010_g N_VPWR_c_551_n 0.00335119f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_252 N_B_M1011_g N_VPWR_c_551_n 0.00518311f $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_253 N_B_M1003_g N_VPWR_c_547_n 0.00488273f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_254 N_B_M1005_g N_VPWR_c_547_n 0.00423213f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_255 N_B_M1010_g N_VPWR_c_547_n 0.00421776f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B_M1011_g N_VPWR_c_547_n 0.00524643f $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B_M1003_g N_A_298_368#_c_616_n 0.00264208f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B_M1005_g N_A_298_368#_c_617_n 0.0111696f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_259 N_B_M1010_g N_A_298_368#_c_617_n 0.00920596f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B_M1005_g N_A_298_368#_c_618_n 7.79815e-19 $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B_M1010_g N_A_298_368#_c_618_n 0.00655172f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B_M1011_g N_A_298_368#_c_618_n 0.00685613f $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_263 N_B_c_238_n N_Y_c_660_n 0.0128008f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_264 N_B_c_244_n N_Y_c_660_n 0.00354091f $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_265 N_B_c_257_n N_Y_c_660_n 0.0172045f $X=1.475 $Y=1.435 $X2=0 $Y2=0
cc_266 N_B_c_238_n N_Y_c_662_n 0.00622488f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_267 N_B_c_240_n N_Y_c_662_n 0.0079293f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_268 N_B_c_240_n N_Y_c_698_n 0.0105176f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_269 N_B_c_250_n N_Y_c_698_n 0.035669f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_270 N_B_c_251_n N_Y_c_698_n 0.00635832f $X=2.045 $Y=1.35 $X2=0 $Y2=0
cc_271 N_B_c_240_n N_Y_c_663_n 5.95058e-19 $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_272 N_B_c_245_n N_Y_c_664_n 0.157951f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_273 N_B_c_248_n N_Y_c_664_n 0.00910698f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_274 N_B_M1005_g N_Y_c_668_n 0.0124091f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_275 N_B_M1010_g N_Y_c_668_n 0.0116635f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_276 N_B_M1011_g N_Y_c_668_n 0.00651638f $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_277 N_B_c_248_n N_Y_c_668_n 0.00509515f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_278 N_B_M1010_g N_Y_c_665_n 0.00349992f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_279 N_B_M1011_g N_Y_c_665_n 0.00450306f $X=5.325 $Y=2.4 $X2=0 $Y2=0
cc_280 N_B_c_245_n N_Y_c_665_n 0.0249855f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_281 N_B_c_248_n N_Y_c_665_n 0.0172245f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_282 N_B_c_238_n N_Y_c_666_n 0.00551466f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_283 N_B_c_239_n N_Y_c_666_n 0.00245638f $X=1.85 $Y=1.26 $X2=0 $Y2=0
cc_284 N_B_c_240_n N_Y_c_666_n 0.00540275f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_285 N_B_c_257_n N_Y_c_666_n 0.00777454f $X=1.475 $Y=1.435 $X2=0 $Y2=0
cc_286 N_B_c_251_n N_Y_c_666_n 0.0196452f $X=2.045 $Y=1.35 $X2=0 $Y2=0
cc_287 N_B_c_249_n N_Y_c_717_n 0.0229777f $X=2.585 $Y=1.35 $X2=0 $Y2=0
cc_288 N_B_c_245_n N_Y_c_669_n 0.0366882f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_289 N_B_c_250_n N_Y_c_669_n 0.0392333f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_290 N_B_c_245_n N_Y_c_670_n 0.122294f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_291 N_B_c_238_n Y 6.20067e-19 $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_292 N_B_c_238_n N_VGND_c_774_n 0.00477239f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_293 N_B_c_240_n N_VGND_c_775_n 0.00381161f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_294 N_B_c_238_n N_VGND_c_779_n 0.00434272f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_295 N_B_c_240_n N_VGND_c_779_n 0.00434272f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_296 N_B_c_238_n N_VGND_c_781_n 0.00821239f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_297 N_B_c_240_n N_VGND_c_781_n 0.0044609f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_298 N_C_M1000_g N_A_27_368#_c_480_n 0.0131577f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_299 N_C_M1001_g N_A_27_368#_c_480_n 0.0132419f $X=2.605 $Y=2.4 $X2=0 $Y2=0
cc_300 N_C_M1015_g N_A_27_368#_c_480_n 0.0132419f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_301 N_C_M1017_g N_A_27_368#_c_480_n 0.013162f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_302 N_C_M1000_g N_A_27_368#_c_494_n 0.00160878f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_303 N_C_M1017_g N_A_27_368#_c_495_n 9.98792e-19 $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_304 N_C_M1000_g N_VPWR_c_551_n 0.00333926f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_305 N_C_M1001_g N_VPWR_c_551_n 0.00333926f $X=2.605 $Y=2.4 $X2=0 $Y2=0
cc_306 N_C_M1015_g N_VPWR_c_551_n 0.00333926f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_307 N_C_M1017_g N_VPWR_c_551_n 0.00333926f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_308 N_C_M1000_g N_VPWR_c_547_n 0.00425421f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_309 N_C_M1001_g N_VPWR_c_547_n 0.00425433f $X=2.605 $Y=2.4 $X2=0 $Y2=0
cc_310 N_C_M1015_g N_VPWR_c_547_n 0.00425433f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_311 N_C_M1017_g N_VPWR_c_547_n 0.00425457f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_312 N_C_M1000_g N_A_298_368#_c_616_n 0.0140067f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_313 N_C_M1001_g N_A_298_368#_c_616_n 0.0144631f $X=2.605 $Y=2.4 $X2=0 $Y2=0
cc_314 N_C_M1015_g N_A_298_368#_c_616_n 0.0144631f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_315 N_C_M1017_g N_A_298_368#_c_616_n 0.0142824f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_316 N_C_M1002_g N_Y_c_662_n 5.99621e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_317 N_C_M1002_g N_Y_c_698_n 0.00917824f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_318 N_C_M1002_g N_Y_c_663_n 0.00744777f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_319 N_C_M1007_g N_Y_c_663_n 0.0115222f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_320 N_C_M1007_g N_Y_c_664_n 0.0105704f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_321 N_C_c_363_n N_Y_c_664_n 0.0148401f $X=3.83 $Y=1.545 $X2=0 $Y2=0
cc_322 C N_Y_c_664_n 0.112382f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_323 N_C_c_368_n N_Y_c_664_n 0.0178347f $X=5.31 $Y=0.505 $X2=0 $Y2=0
cc_324 N_C_c_361_n N_Y_c_668_n 6.45276e-19 $X=3.725 $Y=1.62 $X2=0 $Y2=0
cc_325 N_C_M1017_g N_Y_c_668_n 0.010586f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_326 N_C_c_365_n N_Y_c_668_n 0.00293152f $X=3.815 $Y=1.62 $X2=0 $Y2=0
cc_327 N_C_M1002_g N_Y_c_666_n 8.58155e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_328 N_C_M1002_g N_Y_c_717_n 7.17169e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_329 N_C_M1007_g N_Y_c_717_n 7.17169e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_330 N_C_M1000_g N_Y_c_669_n 0.00401358f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_331 N_C_c_356_n N_Y_c_669_n 0.00557729f $X=2.42 $Y=1.62 $X2=0 $Y2=0
cc_332 N_C_M1001_g N_Y_c_669_n 0.0171368f $X=2.605 $Y=2.4 $X2=0 $Y2=0
cc_333 N_C_c_359_n N_Y_c_669_n 0.00785813f $X=2.85 $Y=1.62 $X2=0 $Y2=0
cc_334 N_C_M1015_g N_Y_c_669_n 0.0167274f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_335 N_C_M1015_g N_Y_c_670_n 0.00186773f $X=3.215 $Y=2.4 $X2=0 $Y2=0
cc_336 N_C_c_361_n N_Y_c_670_n 0.00897092f $X=3.725 $Y=1.62 $X2=0 $Y2=0
cc_337 N_C_M1002_g N_VGND_c_775_n 0.00519354f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_338 N_C_M1002_g N_VGND_c_776_n 0.00434272f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_339 N_C_M1007_g N_VGND_c_776_n 0.00434272f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_340 N_C_M1007_g N_VGND_c_777_n 0.00500066f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_341 N_C_c_366_n N_VGND_c_777_n 0.00758204f $X=3.905 $Y=0.505 $X2=0 $Y2=0
cc_342 C N_VGND_c_777_n 0.0133731f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_343 N_C_c_366_n N_VGND_c_780_n 0.0360112f $X=3.905 $Y=0.505 $X2=0 $Y2=0
cc_344 C N_VGND_c_780_n 0.0766498f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_345 N_C_M1002_g N_VGND_c_781_n 0.0044609f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_346 N_C_M1007_g N_VGND_c_781_n 0.0045006f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_347 N_C_c_366_n N_VGND_c_781_n 0.0528683f $X=3.905 $Y=0.505 $X2=0 $Y2=0
cc_348 C N_VGND_c_781_n 0.0658172f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_349 N_A_27_368#_c_475_n N_VPWR_M1008_s 0.00322221f $X=1.09 $Y=2.425 $X2=-0.19
+ $Y2=1.66
cc_350 N_A_27_368#_c_487_n N_VPWR_M1012_s 0.00322315f $X=6.365 $Y=2.445 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_462_n N_VPWR_c_548_n 0.0105596f $X=0.275 $Y=2.815 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_475_n N_VPWR_c_548_n 0.0166216f $X=1.09 $Y=2.425 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_463_n N_VPWR_c_548_n 0.0105596f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_464_n N_VPWR_c_549_n 0.0111923f $X=5.55 $Y=2.835 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_487_n N_VPWR_c_549_n 0.0166604f $X=6.365 $Y=2.445 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_466_n N_VPWR_c_549_n 0.00990073f $X=6.45 $Y=2.815 $X2=0
+ $Y2=0
cc_357 N_A_27_368#_c_462_n N_VPWR_c_550_n 0.011066f $X=0.275 $Y=2.815 $X2=0
+ $Y2=0
cc_358 N_A_27_368#_c_463_n N_VPWR_c_551_n 0.0109126f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_359 N_A_27_368#_c_480_n N_VPWR_c_551_n 0.00283666f $X=4.485 $Y=2.595 $X2=0
+ $Y2=0
cc_360 N_A_27_368#_c_464_n N_VPWR_c_551_n 0.00811275f $X=5.55 $Y=2.835 $X2=0
+ $Y2=0
cc_361 N_A_27_368#_c_466_n N_VPWR_c_552_n 0.011066f $X=6.45 $Y=2.815 $X2=0 $Y2=0
cc_362 N_A_27_368#_c_462_n N_VPWR_c_547_n 0.00915947f $X=0.275 $Y=2.815 $X2=0
+ $Y2=0
cc_363 N_A_27_368#_c_475_n N_VPWR_c_547_n 0.0129559f $X=1.09 $Y=2.425 $X2=0
+ $Y2=0
cc_364 N_A_27_368#_c_463_n N_VPWR_c_547_n 0.00899513f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_365 N_A_27_368#_c_480_n N_VPWR_c_547_n 0.0103153f $X=4.485 $Y=2.595 $X2=0
+ $Y2=0
cc_366 N_A_27_368#_c_485_n N_VPWR_c_547_n 0.00707445f $X=5.465 $Y=2.445 $X2=0
+ $Y2=0
cc_367 N_A_27_368#_c_464_n N_VPWR_c_547_n 0.006266f $X=5.55 $Y=2.835 $X2=0 $Y2=0
cc_368 N_A_27_368#_c_487_n N_VPWR_c_547_n 0.013213f $X=6.365 $Y=2.445 $X2=0
+ $Y2=0
cc_369 N_A_27_368#_c_466_n N_VPWR_c_547_n 0.00915947f $X=6.45 $Y=2.815 $X2=0
+ $Y2=0
cc_370 N_A_27_368#_c_480_n N_A_298_368#_M1003_s 0.00740542f $X=4.485 $Y=2.595
+ $X2=-0.19 $Y2=1.66
cc_371 N_A_27_368#_c_480_n N_A_298_368#_M1001_s 0.00726344f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_372 N_A_27_368#_c_480_n N_A_298_368#_M1017_s 0.00818977f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_373 N_A_27_368#_c_485_n N_A_298_368#_M1010_s 0.00329277f $X=5.465 $Y=2.445
+ $X2=0 $Y2=0
cc_374 N_A_27_368#_c_463_n N_A_298_368#_c_616_n 0.00487876f $X=1.175 $Y=2.815
+ $X2=0 $Y2=0
cc_375 N_A_27_368#_c_480_n N_A_298_368#_c_616_n 0.157228f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_376 N_A_27_368#_M1005_d N_A_298_368#_c_617_n 0.00165831f $X=4.515 $Y=1.84
+ $X2=0 $Y2=0
cc_377 N_A_27_368#_c_480_n N_A_298_368#_c_617_n 0.00742366f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_378 N_A_27_368#_c_485_n N_A_298_368#_c_617_n 0.00463687f $X=5.465 $Y=2.445
+ $X2=0 $Y2=0
cc_379 N_A_27_368#_c_495_n N_A_298_368#_c_617_n 0.0132901f $X=4.61 $Y=2.445
+ $X2=0 $Y2=0
cc_380 N_A_27_368#_c_485_n N_A_298_368#_c_618_n 0.0157942f $X=5.465 $Y=2.445
+ $X2=0 $Y2=0
cc_381 N_A_27_368#_c_464_n N_A_298_368#_c_618_n 0.0111923f $X=5.55 $Y=2.835
+ $X2=0 $Y2=0
cc_382 N_A_27_368#_c_480_n N_Y_M1000_d 0.0069612f $X=4.485 $Y=2.595 $X2=0 $Y2=0
cc_383 N_A_27_368#_c_480_n N_Y_M1015_d 0.0069612f $X=4.485 $Y=2.595 $X2=0 $Y2=0
cc_384 N_A_27_368#_M1005_d N_Y_c_668_n 0.00166235f $X=4.515 $Y=1.84 $X2=0 $Y2=0
cc_385 N_VPWR_c_548_n N_A_298_368#_c_616_n 0.0028351f $X=0.725 $Y=2.79 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_551_n N_A_298_368#_c_616_n 0.218071f $X=5.835 $Y=3.33 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_547_n N_A_298_368#_c_616_n 0.12348f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_c_549_n N_A_298_368#_c_618_n 0.00207737f $X=6 $Y=2.8 $X2=0 $Y2=0
cc_389 N_VPWR_c_551_n N_A_298_368#_c_618_n 0.0223085f $X=5.835 $Y=3.33 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_547_n N_A_298_368#_c_618_n 0.0122976f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_A_298_368#_c_616_n N_Y_M1000_d 0.00365107f $X=4.173 $Y=2.962 $X2=0
+ $Y2=0
cc_392 N_A_298_368#_c_616_n N_Y_M1015_d 0.00365107f $X=4.173 $Y=2.962 $X2=0
+ $Y2=0
cc_393 N_A_298_368#_M1017_s N_Y_c_668_n 0.00339007f $X=3.905 $Y=1.84 $X2=0 $Y2=0
cc_394 N_A_298_368#_M1010_s N_Y_c_668_n 0.0016705f $X=4.965 $Y=1.84 $X2=0 $Y2=0
cc_395 N_A_298_368#_M1001_s N_Y_c_669_n 0.00402365f $X=2.695 $Y=1.84 $X2=0 $Y2=0
cc_396 N_Y_c_660_n N_VGND_M1016_d 0.00342052f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_397 N_Y_c_698_n N_VGND_M1013_s 0.00669573f $X=2.545 $Y=0.925 $X2=0 $Y2=0
cc_398 N_Y_c_664_n N_VGND_M1007_s 0.0147644f $X=5.135 $Y=0.925 $X2=0 $Y2=0
cc_399 N_Y_c_661_n N_VGND_c_773_n 0.00555794f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_400 Y N_VGND_c_773_n 0.0243474f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_401 N_Y_c_660_n N_VGND_c_774_n 0.0240821f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_402 N_Y_c_662_n N_VGND_c_774_n 0.0191389f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_403 Y N_VGND_c_774_n 0.0191765f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_404 N_Y_c_662_n N_VGND_c_775_n 0.0127977f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_405 N_Y_c_698_n N_VGND_c_775_n 0.0243503f $X=2.545 $Y=0.925 $X2=0 $Y2=0
cc_406 N_Y_c_663_n N_VGND_c_775_n 0.0127977f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_407 N_Y_c_663_n N_VGND_c_776_n 0.0144609f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_408 N_Y_c_663_n N_VGND_c_777_n 0.0122213f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_409 N_Y_c_664_n N_VGND_c_777_n 0.0244298f $X=5.135 $Y=0.925 $X2=0 $Y2=0
cc_410 Y N_VGND_c_778_n 0.0145221f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_411 N_Y_c_662_n N_VGND_c_779_n 0.0144922f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_412 N_Y_c_662_n N_VGND_c_781_n 0.0118826f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_413 N_Y_c_698_n N_VGND_c_781_n 0.0110662f $X=2.545 $Y=0.925 $X2=0 $Y2=0
cc_414 N_Y_c_663_n N_VGND_c_781_n 0.0118703f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_415 N_Y_c_664_n N_VGND_c_781_n 0.0226485f $X=5.135 $Y=0.925 $X2=0 $Y2=0
cc_416 Y N_VGND_c_781_n 0.0119308f $X=0.635 $Y=0.47 $X2=0 $Y2=0

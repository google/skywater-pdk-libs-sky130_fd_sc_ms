* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_29_368# B2 a_297_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_293_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_29_368# B1 a_297_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_675_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR A1 a_297_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 VPWR A2 a_297_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_297_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 Y A1 a_675_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_297_368# B2 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 Y C1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Y B1 a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_297_368# B1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_297_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_293_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND B2 a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_675_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND A2 a_675_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_29_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_139_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=6.14e+06u as=6.608e+11p ps=5.66e+06u
M1001 a_139_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y B1 a_139_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1003 Y A1 a_223_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=3.108e+11p ps=2.32e+06u
M1004 a_223_74# A2 a_145_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1005 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.291e+11p pd=4.39e+06u as=0p ps=0u
M1006 a_145_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_139_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__a2bb2oi_2.pxi.spice
* Created: Fri Aug 28 17:04:42 2020
* 
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%A1_N N_A1_N_c_94_n N_A1_N_c_95_n N_A1_N_M1001_g
+ N_A1_N_M1011_g A1_N N_A1_N_c_98_n N_A1_N_c_99_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_2%A1_N
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%A2_N N_A2_N_M1015_g N_A2_N_M1007_g A2_N
+ N_A2_N_c_122_n N_A2_N_c_123_n PM_SKY130_FD_SC_MS__A2BB2OI_2%A2_N
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%A_212_102# N_A_212_102#_M1011_d
+ N_A_212_102#_M1015_d N_A_212_102#_M1002_g N_A_212_102#_M1012_g
+ N_A_212_102#_M1003_g N_A_212_102#_c_159_n N_A_212_102#_c_160_n
+ N_A_212_102#_M1004_g N_A_212_102#_c_162_n N_A_212_102#_c_163_n
+ N_A_212_102#_c_164_n N_A_212_102#_c_168_n N_A_212_102#_c_165_n
+ N_A_212_102#_c_169_n N_A_212_102#_c_170_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_2%A_212_102#
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%B2 N_B2_M1008_g N_B2_M1000_g N_B2_M1009_g
+ N_B2_M1006_g B2 N_B2_c_251_n N_B2_c_252_n PM_SKY130_FD_SC_MS__A2BB2OI_2%B2
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%B1 N_B1_M1010_g N_B1_M1005_g N_B1_M1014_g
+ N_B1_M1013_g B1 B1 N_B1_c_302_n PM_SKY130_FD_SC_MS__A2BB2OI_2%B1
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%VPWR N_VPWR_M1001_s N_VPWR_M1008_d
+ N_VPWR_M1010_d N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n VPWR
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_340_n
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%A_424_368# N_A_424_368#_M1003_s
+ N_A_424_368#_M1004_s N_A_424_368#_M1009_s N_A_424_368#_M1013_s
+ N_A_424_368#_c_396_n N_A_424_368#_c_397_n N_A_424_368#_c_398_n
+ N_A_424_368#_c_399_n N_A_424_368#_c_413_n N_A_424_368#_c_417_n
+ N_A_424_368#_c_400_n N_A_424_368#_c_421_n N_A_424_368#_c_401_n
+ N_A_424_368#_c_402_n N_A_424_368#_c_427_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_2%A_424_368#
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%Y N_Y_M1002_d N_Y_M1000_d N_Y_M1003_d
+ N_Y_c_452_n N_Y_c_463_n N_Y_c_453_n N_Y_c_454_n N_Y_c_455_n N_Y_c_456_n
+ N_Y_c_457_n Y Y N_Y_c_459_n PM_SKY130_FD_SC_MS__A2BB2OI_2%Y
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%VGND N_VGND_M1011_s N_VGND_M1007_d
+ N_VGND_M1012_s N_VGND_M1005_s N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n VGND N_VGND_c_515_n
+ N_VGND_c_516_n N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n
+ N_VGND_c_521_n N_VGND_c_522_n PM_SKY130_FD_SC_MS__A2BB2OI_2%VGND
x_PM_SKY130_FD_SC_MS__A2BB2OI_2%A_615_74# N_A_615_74#_M1000_s
+ N_A_615_74#_M1006_s N_A_615_74#_M1014_d N_A_615_74#_c_586_n
+ N_A_615_74#_c_587_n N_A_615_74#_c_588_n N_A_615_74#_c_589_n
+ N_A_615_74#_c_590_n PM_SKY130_FD_SC_MS__A2BB2OI_2%A_615_74#
cc_1 VNB N_A1_N_c_94_n 0.0481442f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.36
cc_2 VNB N_A1_N_c_95_n 0.00925795f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.315
cc_3 VNB N_A1_N_M1001_g 0.0292726f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.46
cc_4 VNB N_A1_N_M1011_g 0.00957864f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.83
cc_5 VNB N_A1_N_c_98_n 0.0520748f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.36
cc_6 VNB N_A1_N_c_99_n 0.0173999f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_7 VNB N_A2_N_M1007_g 0.0275221f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.435
cc_8 VNB N_A2_N_c_122_n 0.0181234f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_9 VNB N_A2_N_c_123_n 0.00389989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_212_102#_M1002_g 0.0199064f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.83
cc_11 VNB N_A_212_102#_M1012_g 0.0212056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_212_102#_M1003_g 5.41114e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_13 VNB N_A_212_102#_c_159_n 0.0246498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_212_102#_c_160_n 0.052356f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_15 VNB N_A_212_102#_M1004_g 4.91966e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_212_102#_c_162_n 0.00309191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_212_102#_c_163_n 0.00291468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_212_102#_c_164_n 0.00312382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_212_102#_c_165_n 0.0113965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_M1008_g 4.57279e-19 $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.315
cc_21 VNB N_B2_M1000_g 0.0246759f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.435
cc_22 VNB N_B2_M1009_g 4.54698e-19 $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.225
cc_23 VNB N_B2_M1006_g 0.0224057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B2_c_251_n 9.30952e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B2_c_252_n 0.0439207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_M1005_g 0.023004f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.435
cc_27 VNB N_B1_M1014_g 0.0326336f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.225
cc_28 VNB B1 0.00470982f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_29 VNB N_B1_c_302_n 0.0453065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_340_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_452_n 0.00188975f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_32 VNB N_Y_c_453_n 0.0015351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_454_n 0.00179199f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_34 VNB N_Y_c_455_n 0.0147551f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_35 VNB N_Y_c_456_n 0.00208742f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.555
cc_36 VNB N_Y_c_457_n 0.00330895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB Y 0.00478477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_459_n 0.00839017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_509_n 0.0384995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_510_n 0.00956096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_511_n 0.0132072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_512_n 0.00559476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_513_n 0.0409229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_514_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_515_n 0.0184856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_516_n 0.0209509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_517_n 0.0155887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_518_n 0.0220155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_519_n 0.324227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_520_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_521_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_522_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_615_74#_c_586_n 0.0085563f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.83
cc_54 VNB N_A_615_74#_c_587_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.36
cc_55 VNB N_A_615_74#_c_588_n 0.0162677f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.45
cc_56 VNB N_A_615_74#_c_589_n 0.00225785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_615_74#_c_590_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.555
cc_58 VPB N_A1_N_M1001_g 0.0388248f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.46
cc_59 VPB N_A2_N_M1015_g 0.0256517f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.315
cc_60 VPB N_A2_N_c_122_n 0.0120608f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_61 VPB N_A2_N_c_123_n 0.00813645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_212_102#_M1003_g 0.0249008f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.45
cc_63 VPB N_A_212_102#_M1004_g 0.0217327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_212_102#_c_168_n 0.0153951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_212_102#_c_169_n 0.00668605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_212_102#_c_170_n 0.00593631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_B2_M1008_g 0.0218378f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.315
cc_68 VPB N_B2_M1009_g 0.0218481f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.225
cc_69 VPB N_B2_c_251_n 0.00251854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_B1_M1010_g 0.0202406f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.315
cc_71 VPB N_B1_M1013_g 0.0281481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB B1 0.00544426f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.45
cc_73 VPB N_B1_c_302_n 0.00525849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_341_n 0.0616596f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_75 VPB N_VPWR_c_342_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.45
cc_76 VPB N_VPWR_c_343_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.555
cc_77 VPB N_VPWR_c_344_n 0.0206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_345_n 0.0648853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_346_n 0.0164265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_347_n 0.0197776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_340_n 0.103585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_349_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_350_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_351_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_424_368#_c_396_n 0.0120542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_424_368#_c_397_n 0.00475153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_424_368#_c_398_n 0.00460831f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.45
cc_88 VPB N_A_424_368#_c_399_n 0.00315626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_424_368#_c_400_n 0.00176163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_424_368#_c_401_n 0.0171219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_424_368#_c_402_n 0.0345796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_Y_c_454_n 0.00163227f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.45
cc_93 N_A1_N_c_94_n N_A2_N_M1007_g 0.0165728f $X=0.91 $Y=0.36 $X2=0 $Y2=0
cc_94 N_A1_N_M1001_g N_A2_N_c_122_n 0.098121f $X=0.97 $Y=2.46 $X2=0 $Y2=0
cc_95 N_A1_N_M1001_g N_A2_N_c_123_n 0.00968467f $X=0.97 $Y=2.46 $X2=0 $Y2=0
cc_96 N_A1_N_M1011_g N_A_212_102#_c_162_n 0.00729347f $X=0.985 $Y=0.83 $X2=0
+ $Y2=0
cc_97 N_A1_N_c_95_n N_A_212_102#_c_164_n 0.00464063f $X=0.97 $Y=1.315 $X2=0
+ $Y2=0
cc_98 N_A1_N_M1011_g N_A_212_102#_c_164_n 0.00416728f $X=0.985 $Y=0.83 $X2=0
+ $Y2=0
cc_99 N_A1_N_M1001_g N_A_212_102#_c_169_n 0.00280028f $X=0.97 $Y=2.46 $X2=0
+ $Y2=0
cc_100 N_A1_N_M1001_g N_VPWR_c_341_n 0.0257097f $X=0.97 $Y=2.46 $X2=0 $Y2=0
cc_101 N_A1_N_M1001_g N_VPWR_c_345_n 0.00460063f $X=0.97 $Y=2.46 $X2=0 $Y2=0
cc_102 N_A1_N_M1001_g N_VPWR_c_340_n 0.00908061f $X=0.97 $Y=2.46 $X2=0 $Y2=0
cc_103 N_A1_N_c_94_n N_VGND_c_509_n 0.0216612f $X=0.91 $Y=0.36 $X2=0 $Y2=0
cc_104 N_A1_N_M1011_g N_VGND_c_509_n 0.00217288f $X=0.985 $Y=0.83 $X2=0 $Y2=0
cc_105 N_A1_N_c_98_n N_VGND_c_509_n 0.00156654f $X=0.27 $Y=0.36 $X2=0 $Y2=0
cc_106 N_A1_N_c_99_n N_VGND_c_509_n 0.0294445f $X=0.27 $Y=0.45 $X2=0 $Y2=0
cc_107 N_A1_N_c_94_n N_VGND_c_510_n 0.0032259f $X=0.91 $Y=0.36 $X2=0 $Y2=0
cc_108 N_A1_N_c_98_n N_VGND_c_515_n 0.00703799f $X=0.27 $Y=0.36 $X2=0 $Y2=0
cc_109 N_A1_N_c_99_n N_VGND_c_515_n 0.0179317f $X=0.27 $Y=0.45 $X2=0 $Y2=0
cc_110 N_A1_N_c_94_n N_VGND_c_516_n 0.00680549f $X=0.91 $Y=0.36 $X2=0 $Y2=0
cc_111 N_A1_N_c_98_n N_VGND_c_519_n 0.0117623f $X=0.27 $Y=0.36 $X2=0 $Y2=0
cc_112 N_A1_N_c_99_n N_VGND_c_519_n 0.0121515f $X=0.27 $Y=0.45 $X2=0 $Y2=0
cc_113 N_A2_N_M1007_g N_A_212_102#_M1002_g 0.0272428f $X=1.46 $Y=0.83 $X2=0
+ $Y2=0
cc_114 N_A2_N_c_122_n N_A_212_102#_c_160_n 0.00880632f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_115 N_A2_N_M1007_g N_A_212_102#_c_163_n 0.0149733f $X=1.46 $Y=0.83 $X2=0
+ $Y2=0
cc_116 N_A2_N_c_122_n N_A_212_102#_c_163_n 0.00305246f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_117 N_A2_N_c_123_n N_A_212_102#_c_163_n 0.0174383f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_118 N_A2_N_c_122_n N_A_212_102#_c_164_n 0.00163439f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_119 N_A2_N_c_123_n N_A_212_102#_c_164_n 0.0214254f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_120 N_A2_N_M1015_g N_A_212_102#_c_168_n 0.0147227f $X=1.36 $Y=2.46 $X2=0
+ $Y2=0
cc_121 N_A2_N_M1007_g N_A_212_102#_c_165_n 0.00403933f $X=1.46 $Y=0.83 $X2=0
+ $Y2=0
cc_122 N_A2_N_c_122_n N_A_212_102#_c_165_n 0.00143871f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_123 N_A2_N_c_123_n N_A_212_102#_c_165_n 0.0168013f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_124 N_A2_N_M1015_g N_A_212_102#_c_169_n 0.00500006f $X=1.36 $Y=2.46 $X2=0
+ $Y2=0
cc_125 N_A2_N_c_122_n N_A_212_102#_c_169_n 0.00403602f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_126 N_A2_N_c_123_n N_A_212_102#_c_169_n 0.0124349f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_127 N_A2_N_M1015_g N_A_212_102#_c_170_n 0.00519584f $X=1.36 $Y=2.46 $X2=0
+ $Y2=0
cc_128 N_A2_N_c_122_n N_A_212_102#_c_170_n 0.00303087f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_129 N_A2_N_c_123_n N_A_212_102#_c_170_n 0.00999859f $X=1.435 $Y=1.615 $X2=0
+ $Y2=0
cc_130 N_A2_N_M1015_g N_VPWR_c_341_n 0.00340742f $X=1.36 $Y=2.46 $X2=0 $Y2=0
cc_131 N_A2_N_M1015_g N_VPWR_c_345_n 0.005209f $X=1.36 $Y=2.46 $X2=0 $Y2=0
cc_132 N_A2_N_M1015_g N_VPWR_c_340_n 0.00988003f $X=1.36 $Y=2.46 $X2=0 $Y2=0
cc_133 N_A2_N_M1015_g N_A_424_368#_c_396_n 0.00101941f $X=1.36 $Y=2.46 $X2=0
+ $Y2=0
cc_134 N_A2_N_M1015_g N_A_424_368#_c_398_n 0.00260566f $X=1.36 $Y=2.46 $X2=0
+ $Y2=0
cc_135 N_A2_N_M1007_g N_VGND_c_509_n 2.29767e-19 $X=1.46 $Y=0.83 $X2=0 $Y2=0
cc_136 N_A2_N_M1007_g N_VGND_c_510_n 0.00556969f $X=1.46 $Y=0.83 $X2=0 $Y2=0
cc_137 N_A2_N_M1007_g N_VGND_c_516_n 0.00481372f $X=1.46 $Y=0.83 $X2=0 $Y2=0
cc_138 N_A2_N_M1007_g N_VGND_c_519_n 0.00502397f $X=1.46 $Y=0.83 $X2=0 $Y2=0
cc_139 N_A_212_102#_M1004_g N_B2_M1008_g 0.0122285f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_212_102#_c_159_n N_B2_c_251_n 9.99339e-19 $X=2.83 $Y=1.575 $X2=0
+ $Y2=0
cc_141 N_A_212_102#_c_159_n N_B2_c_252_n 0.0122285f $X=2.83 $Y=1.575 $X2=0 $Y2=0
cc_142 N_A_212_102#_c_169_n N_VPWR_c_341_n 0.0324718f $X=1.585 $Y=2.115 $X2=0
+ $Y2=0
cc_143 N_A_212_102#_M1004_g N_VPWR_c_342_n 3.91772e-19 $X=2.92 $Y=2.4 $X2=0
+ $Y2=0
cc_144 N_A_212_102#_M1003_g N_VPWR_c_345_n 0.00333926f $X=2.47 $Y=2.4 $X2=0
+ $Y2=0
cc_145 N_A_212_102#_M1004_g N_VPWR_c_345_n 0.00333896f $X=2.92 $Y=2.4 $X2=0
+ $Y2=0
cc_146 N_A_212_102#_c_168_n N_VPWR_c_345_n 0.0216883f $X=1.585 $Y=2.815 $X2=0
+ $Y2=0
cc_147 N_A_212_102#_M1003_g N_VPWR_c_340_n 0.0042782f $X=2.47 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_212_102#_M1004_g N_VPWR_c_340_n 0.00422796f $X=2.92 $Y=2.4 $X2=0
+ $Y2=0
cc_149 N_A_212_102#_c_168_n N_VPWR_c_340_n 0.0178836f $X=1.585 $Y=2.815 $X2=0
+ $Y2=0
cc_150 N_A_212_102#_M1003_g N_A_424_368#_c_396_n 0.00147158f $X=2.47 $Y=2.4
+ $X2=0 $Y2=0
cc_151 N_A_212_102#_c_160_n N_A_424_368#_c_396_n 0.0051692f $X=2.56 $Y=1.575
+ $X2=0 $Y2=0
cc_152 N_A_212_102#_c_165_n N_A_424_368#_c_396_n 0.0105084f $X=1.825 $Y=1.65
+ $X2=0 $Y2=0
cc_153 N_A_212_102#_c_170_n N_A_424_368#_c_396_n 0.0902949f $X=1.665 $Y=1.95
+ $X2=0 $Y2=0
cc_154 N_A_212_102#_M1003_g N_A_424_368#_c_397_n 0.0147971f $X=2.47 $Y=2.4 $X2=0
+ $Y2=0
cc_155 N_A_212_102#_M1004_g N_A_424_368#_c_397_n 0.0132535f $X=2.92 $Y=2.4 $X2=0
+ $Y2=0
cc_156 N_A_212_102#_c_168_n N_A_424_368#_c_398_n 0.00682755f $X=1.585 $Y=2.815
+ $X2=0 $Y2=0
cc_157 N_A_212_102#_M1004_g N_A_424_368#_c_399_n 0.00429672f $X=2.92 $Y=2.4
+ $X2=0 $Y2=0
cc_158 N_A_212_102#_M1003_g N_A_424_368#_c_413_n 7.26148e-19 $X=2.47 $Y=2.4
+ $X2=0 $Y2=0
cc_159 N_A_212_102#_M1004_g N_A_424_368#_c_413_n 0.0111671f $X=2.92 $Y=2.4 $X2=0
+ $Y2=0
cc_160 N_A_212_102#_M1002_g N_Y_c_452_n 3.0814e-19 $X=1.95 $Y=0.78 $X2=0 $Y2=0
cc_161 N_A_212_102#_M1012_g N_Y_c_452_n 3.0814e-19 $X=2.38 $Y=0.78 $X2=0 $Y2=0
cc_162 N_A_212_102#_M1012_g N_Y_c_463_n 0.0183036f $X=2.38 $Y=0.78 $X2=0 $Y2=0
cc_163 N_A_212_102#_c_160_n N_Y_c_463_n 0.00156873f $X=2.56 $Y=1.575 $X2=0 $Y2=0
cc_164 N_A_212_102#_c_160_n N_Y_c_453_n 0.00101398f $X=2.56 $Y=1.575 $X2=0 $Y2=0
cc_165 N_A_212_102#_c_165_n N_Y_c_453_n 0.0102843f $X=1.825 $Y=1.65 $X2=0 $Y2=0
cc_166 N_A_212_102#_M1003_g N_Y_c_454_n 0.0193352f $X=2.47 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A_212_102#_c_159_n N_Y_c_454_n 0.013082f $X=2.83 $Y=1.575 $X2=0 $Y2=0
cc_168 N_A_212_102#_c_160_n N_Y_c_454_n 0.00696484f $X=2.56 $Y=1.575 $X2=0 $Y2=0
cc_169 N_A_212_102#_M1004_g N_Y_c_454_n 0.00379157f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A_212_102#_c_165_n N_Y_c_454_n 0.0113048f $X=1.825 $Y=1.65 $X2=0 $Y2=0
cc_171 N_A_212_102#_c_170_n N_Y_c_454_n 0.00469336f $X=1.665 $Y=1.95 $X2=0 $Y2=0
cc_172 N_A_212_102#_c_159_n N_Y_c_455_n 0.0109044f $X=2.83 $Y=1.575 $X2=0 $Y2=0
cc_173 N_A_212_102#_M1012_g Y 0.00798713f $X=2.38 $Y=0.78 $X2=0 $Y2=0
cc_174 N_A_212_102#_c_165_n Y 0.0104157f $X=1.825 $Y=1.65 $X2=0 $Y2=0
cc_175 N_A_212_102#_c_163_n N_VGND_M1007_d 0.00156264f $X=1.74 $Y=1.195 $X2=0
+ $Y2=0
cc_176 N_A_212_102#_c_165_n N_VGND_M1007_d 8.63167e-19 $X=1.825 $Y=1.65 $X2=0
+ $Y2=0
cc_177 N_A_212_102#_c_162_n N_VGND_c_509_n 0.022536f $X=1.22 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_A_212_102#_c_164_n N_VGND_c_509_n 0.00314439f $X=1.33 $Y=1.195 $X2=0
+ $Y2=0
cc_179 N_A_212_102#_M1002_g N_VGND_c_510_n 0.0124909f $X=1.95 $Y=0.78 $X2=0
+ $Y2=0
cc_180 N_A_212_102#_M1012_g N_VGND_c_510_n 4.87951e-19 $X=2.38 $Y=0.78 $X2=0
+ $Y2=0
cc_181 N_A_212_102#_c_162_n N_VGND_c_510_n 0.00123145f $X=1.22 $Y=0.655 $X2=0
+ $Y2=0
cc_182 N_A_212_102#_c_163_n N_VGND_c_510_n 0.0120046f $X=1.74 $Y=1.195 $X2=0
+ $Y2=0
cc_183 N_A_212_102#_c_165_n N_VGND_c_510_n 0.00902191f $X=1.825 $Y=1.65 $X2=0
+ $Y2=0
cc_184 N_A_212_102#_M1002_g N_VGND_c_511_n 4.49156e-19 $X=1.95 $Y=0.78 $X2=0
+ $Y2=0
cc_185 N_A_212_102#_M1012_g N_VGND_c_511_n 0.0105465f $X=2.38 $Y=0.78 $X2=0
+ $Y2=0
cc_186 N_A_212_102#_c_160_n N_VGND_c_511_n 6.99248e-19 $X=2.56 $Y=1.575 $X2=0
+ $Y2=0
cc_187 N_A_212_102#_c_162_n N_VGND_c_516_n 0.00825865f $X=1.22 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_212_102#_M1002_g N_VGND_c_517_n 0.00455951f $X=1.95 $Y=0.78 $X2=0
+ $Y2=0
cc_189 N_A_212_102#_M1012_g N_VGND_c_517_n 0.00455951f $X=2.38 $Y=0.78 $X2=0
+ $Y2=0
cc_190 N_A_212_102#_M1002_g N_VGND_c_519_n 0.00447788f $X=1.95 $Y=0.78 $X2=0
+ $Y2=0
cc_191 N_A_212_102#_M1012_g N_VGND_c_519_n 0.00447788f $X=2.38 $Y=0.78 $X2=0
+ $Y2=0
cc_192 N_A_212_102#_c_162_n N_VGND_c_519_n 0.0098462f $X=1.22 $Y=0.655 $X2=0
+ $Y2=0
cc_193 N_A_212_102#_M1012_g N_A_615_74#_c_586_n 7.64007e-19 $X=2.38 $Y=0.78
+ $X2=0 $Y2=0
cc_194 N_B2_M1009_g N_B1_M1010_g 0.0135543f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_195 N_B2_M1006_g N_B1_M1005_g 0.0193758f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_196 N_B2_c_251_n B1 0.0288576f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_197 N_B2_c_252_n B1 0.0044137f $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_198 N_B2_c_251_n N_B1_c_302_n 3.05931e-19 $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_199 N_B2_c_252_n N_B1_c_302_n 0.0194779f $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_200 N_B2_M1008_g N_VPWR_c_342_n 0.0121257f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_201 N_B2_M1009_g N_VPWR_c_342_n 0.01274f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_202 N_B2_M1009_g N_VPWR_c_343_n 5.41206e-19 $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_203 N_B2_M1008_g N_VPWR_c_345_n 0.00460063f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_204 N_B2_M1009_g N_VPWR_c_346_n 0.00460063f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_205 N_B2_M1008_g N_VPWR_c_340_n 0.00908665f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_206 N_B2_M1009_g N_VPWR_c_340_n 0.00908665f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_207 N_B2_M1008_g N_A_424_368#_c_397_n 0.00101073f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_208 N_B2_M1008_g N_A_424_368#_c_399_n 4.97677e-19 $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_209 N_B2_M1008_g N_A_424_368#_c_417_n 0.0179786f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_210 N_B2_M1009_g N_A_424_368#_c_417_n 0.0194916f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B2_c_251_n N_A_424_368#_c_417_n 0.0218447f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_212 N_B2_c_252_n N_A_424_368#_c_417_n 4.5617e-19 $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_213 N_B2_c_251_n N_Y_c_454_n 0.0100292f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_214 N_B2_c_252_n N_Y_c_454_n 0.00234545f $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_215 N_B2_M1000_g N_Y_c_456_n 0.0133827f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B2_c_251_n N_Y_c_456_n 0.00435083f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_217 N_B2_c_252_n N_Y_c_456_n 0.00249037f $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_218 N_B2_M1000_g N_Y_c_457_n 0.0111719f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B2_M1006_g N_Y_c_457_n 0.0058626f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B2_c_251_n N_Y_c_457_n 0.0220896f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_221 N_B2_c_252_n N_Y_c_457_n 7.46584e-19 $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_222 N_B2_M1000_g N_Y_c_459_n 0.00746753f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B2_c_251_n N_Y_c_459_n 0.00753152f $X=3.57 $Y=1.485 $X2=0 $Y2=0
cc_224 N_B2_c_252_n N_Y_c_459_n 0.00275234f $X=3.82 $Y=1.485 $X2=0 $Y2=0
cc_225 N_B2_M1000_g N_VGND_c_511_n 0.00702892f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B2_M1006_g N_VGND_c_512_n 6.37019e-19 $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B2_M1000_g N_VGND_c_513_n 0.00291649f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B2_M1006_g N_VGND_c_513_n 0.00291649f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B2_M1000_g N_VGND_c_519_n 0.0036412f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B2_M1006_g N_VGND_c_519_n 0.00359219f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B2_M1000_g N_A_615_74#_c_586_n 0.01124f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B2_M1006_g N_A_615_74#_c_586_n 0.0142063f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B2_M1006_g N_A_615_74#_c_589_n 0.00127665f $X=3.845 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B1_M1010_g N_VPWR_c_342_n 5.41206e-19 $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_235 N_B1_M1010_g N_VPWR_c_343_n 0.0127835f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_236 N_B1_M1013_g N_VPWR_c_343_n 0.0158915f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_237 N_B1_M1010_g N_VPWR_c_346_n 0.00460063f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B1_M1013_g N_VPWR_c_347_n 0.00460063f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_239 N_B1_M1010_g N_VPWR_c_340_n 0.00908665f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_240 N_B1_M1013_g N_VPWR_c_340_n 0.00912473f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B1_M1010_g N_A_424_368#_c_421_n 0.0142562f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_242 N_B1_M1013_g N_A_424_368#_c_421_n 0.0182976f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_243 B1 N_A_424_368#_c_421_n 0.0359152f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_244 N_B1_c_302_n N_A_424_368#_c_421_n 4.90767e-19 $X=4.72 $Y=1.515 $X2=0
+ $Y2=0
cc_245 N_B1_M1013_g N_A_424_368#_c_401_n 8.13654e-19 $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B1_M1013_g N_A_424_368#_c_402_n 0.00147311f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_247 B1 N_A_424_368#_c_427_n 0.0141817f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_248 N_B1_M1005_g N_VGND_c_512_n 0.00977449f $X=4.275 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B1_M1014_g N_VGND_c_512_n 0.00328502f $X=4.705 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B1_M1005_g N_VGND_c_513_n 0.00383152f $X=4.275 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B1_M1014_g N_VGND_c_518_n 0.00434272f $X=4.705 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B1_M1005_g N_VGND_c_519_n 0.00757637f $X=4.275 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B1_M1014_g N_VGND_c_519_n 0.00824186f $X=4.705 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B1_M1005_g N_A_615_74#_c_588_n 0.0128967f $X=4.275 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B1_M1014_g N_A_615_74#_c_588_n 0.0165989f $X=4.705 $Y=0.74 $X2=0 $Y2=0
cc_256 B1 N_A_615_74#_c_588_n 0.0400398f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_257 N_B1_c_302_n N_A_615_74#_c_588_n 0.00426023f $X=4.72 $Y=1.515 $X2=0 $Y2=0
cc_258 B1 N_A_615_74#_c_589_n 0.0153286f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_259 N_B1_M1005_g N_A_615_74#_c_590_n 7.07591e-19 $X=4.275 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B1_M1014_g N_A_615_74#_c_590_n 0.0100626f $X=4.705 $Y=0.74 $X2=0 $Y2=0
cc_261 N_VPWR_c_342_n N_A_424_368#_c_397_n 0.0103602f $X=3.595 $Y=2.455 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_345_n N_A_424_368#_c_397_n 0.0586721f $X=3.43 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_340_n N_A_424_368#_c_397_n 0.0325115f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_345_n N_A_424_368#_c_398_n 0.0179217f $X=3.43 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_340_n N_A_424_368#_c_398_n 0.00971942f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_266 N_VPWR_M1008_d N_A_424_368#_c_417_n 0.0031498f $X=3.46 $Y=1.84 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_342_n N_A_424_368#_c_417_n 0.0170259f $X=3.595 $Y=2.455 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_342_n N_A_424_368#_c_400_n 0.0233699f $X=3.595 $Y=2.455 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_343_n N_A_424_368#_c_400_n 0.0233699f $X=4.495 $Y=2.455 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_346_n N_A_424_368#_c_400_n 0.00749631f $X=4.33 $Y=3.33 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_340_n N_A_424_368#_c_400_n 0.0062048f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_272 N_VPWR_M1010_d N_A_424_368#_c_421_n 0.00314376f $X=4.36 $Y=1.84 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_343_n N_A_424_368#_c_421_n 0.0170259f $X=4.495 $Y=2.455 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_343_n N_A_424_368#_c_402_n 0.0234083f $X=4.495 $Y=2.455 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_347_n N_A_424_368#_c_402_n 0.011066f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_276 N_VPWR_c_340_n N_A_424_368#_c_402_n 0.00915947f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_277 N_A_424_368#_c_397_n N_Y_M1003_d 0.00165831f $X=2.98 $Y=2.99 $X2=0 $Y2=0
cc_278 N_A_424_368#_c_396_n N_Y_c_463_n 0.00163427f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_279 N_A_424_368#_c_396_n N_Y_c_453_n 0.00147466f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A_424_368#_c_396_n N_Y_c_454_n 0.0302573f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_424_368#_c_397_n N_Y_c_454_n 0.014259f $X=2.98 $Y=2.99 $X2=0 $Y2=0
cc_282 N_A_424_368#_c_399_n N_Y_c_454_n 0.0110894f $X=3.105 $Y=2.12 $X2=0 $Y2=0
cc_283 N_A_424_368#_c_399_n N_Y_c_455_n 0.0120729f $X=3.105 $Y=2.12 $X2=0 $Y2=0
cc_284 N_A_424_368#_c_401_n N_A_615_74#_c_588_n 0.00831718f $X=4.985 $Y=2.12
+ $X2=0 $Y2=0
cc_285 N_Y_c_463_n N_VGND_M1012_s 2.88975e-19 $X=2.525 $Y=1.065 $X2=0 $Y2=0
cc_286 Y N_VGND_M1012_s 0.00295773f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_287 N_Y_c_452_n N_VGND_c_510_n 0.0203993f $X=2.165 $Y=0.555 $X2=0 $Y2=0
cc_288 N_Y_c_452_n N_VGND_c_511_n 0.0157399f $X=2.165 $Y=0.555 $X2=0 $Y2=0
cc_289 N_Y_c_463_n N_VGND_c_511_n 0.00280727f $X=2.525 $Y=1.065 $X2=0 $Y2=0
cc_290 Y N_VGND_c_511_n 0.0212357f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_291 N_Y_c_452_n N_VGND_c_517_n 0.00645633f $X=2.165 $Y=0.555 $X2=0 $Y2=0
cc_292 N_Y_c_452_n N_VGND_c_519_n 0.00605288f $X=2.165 $Y=0.555 $X2=0 $Y2=0
cc_293 N_Y_c_456_n N_A_615_74#_M1000_s 7.34034e-19 $X=3.465 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_294 N_Y_c_459_n N_A_615_74#_M1000_s 0.00318338f $X=3.235 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_295 N_Y_M1000_d N_A_615_74#_c_586_n 0.00178571f $X=3.49 $Y=0.37 $X2=0 $Y2=0
cc_296 N_Y_c_457_n N_A_615_74#_c_586_n 0.0162079f $X=3.63 $Y=0.95 $X2=0 $Y2=0
cc_297 N_Y_c_459_n N_A_615_74#_c_586_n 0.0155322f $X=3.235 $Y=1.195 $X2=0 $Y2=0
cc_298 N_Y_c_457_n N_A_615_74#_c_589_n 0.00678603f $X=3.63 $Y=0.95 $X2=0 $Y2=0
cc_299 N_VGND_c_511_n N_A_615_74#_c_586_n 0.0156798f $X=2.595 $Y=0.645 $X2=0
+ $Y2=0
cc_300 N_VGND_c_513_n N_A_615_74#_c_586_n 0.038121f $X=4.325 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_c_519_n N_A_615_74#_c_586_n 0.0321651f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_512_n N_A_615_74#_c_587_n 0.00947603f $X=4.49 $Y=0.595 $X2=0
+ $Y2=0
cc_303 N_VGND_c_513_n N_A_615_74#_c_587_n 0.00758556f $X=4.325 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_519_n N_A_615_74#_c_587_n 0.00627867f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_M1005_s N_A_615_74#_c_588_n 0.00176461f $X=4.35 $Y=0.37 $X2=0
+ $Y2=0
cc_306 N_VGND_c_512_n N_A_615_74#_c_588_n 0.0153337f $X=4.49 $Y=0.595 $X2=0
+ $Y2=0
cc_307 N_VGND_c_512_n N_A_615_74#_c_590_n 0.0182902f $X=4.49 $Y=0.595 $X2=0
+ $Y2=0
cc_308 N_VGND_c_518_n N_A_615_74#_c_590_n 0.0145639f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_519_n N_A_615_74#_c_590_n 0.0119984f $X=5.04 $Y=0 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__ebufn_8.ext - technology: sky130A

.subckt sky130_fd_sc_ms__ebufn_8 A TE_B VGND VNB VPB VPWR Z
M1000 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.0054e+12p pd=1.874e+07u as=1.2506e+12p ps=1.226e+07u
M1001 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.3048e+12p pd=1.129e+07u as=2.8168e+12p ps=2.519e+07u
M1002 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.213e+11p ps=8.41e+06u
M1008 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.4573e+12p ps=1.808e+07u
M1010 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_84_48# A VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 Z a_84_48# a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_28_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR TE_B a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A a_84_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_833_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_84_48# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR TE_B a_833_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.544e+11p ps=3.23e+06u
M1029 VGND TE_B a_833_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1030 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR A a_84_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_28_368# a_84_48# Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_27_74# a_833_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


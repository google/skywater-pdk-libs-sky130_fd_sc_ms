* File: sky130_fd_sc_ms__a2bb2o_1.pxi.spice
* Created: Fri Aug 28 17:04:06 2020
* 
x_PM_SKY130_FD_SC_MS__A2BB2O_1%A_93_264# N_A_93_264#_M1002_d N_A_93_264#_M1009_s
+ N_A_93_264#_M1000_g N_A_93_264#_M1006_g N_A_93_264#_c_85_n N_A_93_264#_c_92_n
+ N_A_93_264#_c_153_p N_A_93_264#_c_174_p N_A_93_264#_c_93_n N_A_93_264#_c_94_n
+ N_A_93_264#_c_95_n N_A_93_264#_c_86_n N_A_93_264#_c_97_n N_A_93_264#_c_87_n
+ N_A_93_264#_c_126_p N_A_93_264#_c_88_n N_A_93_264#_c_89_n N_A_93_264#_c_98_n
+ PM_SKY130_FD_SC_MS__A2BB2O_1%A_93_264#
x_PM_SKY130_FD_SC_MS__A2BB2O_1%A1_N N_A1_N_M1001_g N_A1_N_M1004_g A1_N
+ N_A1_N_c_189_n N_A1_N_c_190_n PM_SKY130_FD_SC_MS__A2BB2O_1%A1_N
x_PM_SKY130_FD_SC_MS__A2BB2O_1%A2_N N_A2_N_c_226_n N_A2_N_M1007_g N_A2_N_c_227_n
+ N_A2_N_M1005_g A2_N PM_SKY130_FD_SC_MS__A2BB2O_1%A2_N
x_PM_SKY130_FD_SC_MS__A2BB2O_1%A_257_126# N_A_257_126#_M1004_d
+ N_A_257_126#_M1007_d N_A_257_126#_M1002_g N_A_257_126#_M1009_g
+ N_A_257_126#_c_268_n N_A_257_126#_c_269_n N_A_257_126#_c_270_n
+ N_A_257_126#_c_271_n N_A_257_126#_c_275_n N_A_257_126#_c_276_n
+ N_A_257_126#_c_277_n N_A_257_126#_c_272_n N_A_257_126#_c_273_n
+ PM_SKY130_FD_SC_MS__A2BB2O_1%A_257_126#
x_PM_SKY130_FD_SC_MS__A2BB2O_1%B2 N_B2_M1003_g N_B2_M1011_g B2 N_B2_c_340_n
+ PM_SKY130_FD_SC_MS__A2BB2O_1%B2
x_PM_SKY130_FD_SC_MS__A2BB2O_1%B1 N_B1_M1008_g N_B1_c_377_n N_B1_M1010_g B1 B1
+ N_B1_c_380_n PM_SKY130_FD_SC_MS__A2BB2O_1%B1
x_PM_SKY130_FD_SC_MS__A2BB2O_1%X N_X_M1006_s N_X_M1000_s N_X_c_406_n N_X_c_407_n
+ X X X N_X_c_410_n N_X_c_408_n X PM_SKY130_FD_SC_MS__A2BB2O_1%X
x_PM_SKY130_FD_SC_MS__A2BB2O_1%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_c_431_n
+ N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n VPWR N_VPWR_c_435_n
+ N_VPWR_c_436_n N_VPWR_c_430_n N_VPWR_c_438_n PM_SKY130_FD_SC_MS__A2BB2O_1%VPWR
x_PM_SKY130_FD_SC_MS__A2BB2O_1%A_533_392# N_A_533_392#_M1009_d
+ N_A_533_392#_M1010_d N_A_533_392#_c_478_n N_A_533_392#_c_479_n
+ N_A_533_392#_c_480_n N_A_533_392#_c_481_n N_A_533_392#_c_482_n
+ PM_SKY130_FD_SC_MS__A2BB2O_1%A_533_392#
x_PM_SKY130_FD_SC_MS__A2BB2O_1%VGND N_VGND_M1006_d N_VGND_M1005_d N_VGND_M1008_d
+ N_VGND_c_503_n N_VGND_c_519_n N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_562_n
+ N_VGND_c_553_n N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n VGND N_VGND_c_513_n
+ N_VGND_c_514_n PM_SKY130_FD_SC_MS__A2BB2O_1%VGND
cc_1 VNB N_A_93_264#_M1000_g 5.3677e-19 $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_2 VNB N_A_93_264#_M1006_g 0.024394f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_3 VNB N_A_93_264#_c_85_n 3.96917e-19 $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.79
cc_4 VNB N_A_93_264#_c_86_n 0.00914112f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.79
cc_5 VNB N_A_93_264#_c_87_n 3.76316e-19 $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.12
cc_6 VNB N_A_93_264#_c_88_n 0.0354364f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.485
cc_7 VNB N_A_93_264#_c_89_n 0.00668603f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.485
cc_8 VNB N_A1_N_M1001_g 0.00222805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A1_N 0.00271775f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_10 VNB N_A1_N_c_189_n 0.0313834f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.32
cc_11 VNB N_A1_N_c_190_n 0.0166691f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_12 VNB N_A2_N_c_226_n 0.0384047f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=0.63
cc_13 VNB N_A2_N_c_227_n 0.0199265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2_N 0.00300577f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_15 VNB N_A_257_126#_M1002_g 0.020051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_257_126#_c_268_n 0.00104163f $X=-0.19 $Y=-0.245 $X2=1.325
+ $Y2=1.875
cc_17 VNB N_A_257_126#_c_269_n 0.00564675f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.96
cc_18 VNB N_A_257_126#_c_270_n 0.0152508f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.875
cc_19 VNB N_A_257_126#_c_271_n 0.0462783f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.875
cc_20 VNB N_A_257_126#_c_272_n 0.00162172f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_21 VNB N_A_257_126#_c_273_n 0.021289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B2_M1003_g 0.0216081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B2 0.00401095f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_24 VNB N_B2_c_340_n 0.0198707f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_25 VNB N_B1_M1008_g 0.013239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_377_n 0.00887504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_M1010_g 0.0187569f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_28 VNB B1 0.0355701f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.32
cc_29 VNB N_B1_c_380_n 0.0531247f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.875
cc_30 VNB N_X_c_406_n 0.02872f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.4
cc_31 VNB N_X_c_407_n 0.0124546f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_32 VNB N_X_c_408_n 0.0241894f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_33 VNB N_VPWR_c_430_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.12
cc_34 VNB N_VGND_c_503_n 0.0122286f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.81
cc_35 VNB N_VGND_c_504_n 0.00822066f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.96
cc_36 VNB N_VGND_c_505_n 0.0102407f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.875
cc_37 VNB N_VGND_c_506_n 0.0234937f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.21
cc_38 VNB N_VGND_c_507_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.79
cc_39 VNB N_VGND_c_508_n 0.0397362f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=2.635
cc_40 VNB N_VGND_c_509_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=2.635
cc_41 VNB N_VGND_c_510_n 0.00661898f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.12
cc_42 VNB N_VGND_c_511_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_43 VNB N_VGND_c_512_n 0.022756f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.12
cc_44 VNB N_VGND_c_513_n 0.0272571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_514_n 0.263154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A_93_264#_M1000_g 0.0278178f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_47 VPB N_A_93_264#_c_85_n 0.00128976f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.79
cc_48 VPB N_A_93_264#_c_92_n 0.00689106f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.875
cc_49 VPB N_A_93_264#_c_93_n 0.0149438f $X=-0.19 $Y=1.66 $X2=2.02 $Y2=1.875
cc_50 VPB N_A_93_264#_c_94_n 0.0114911f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.99
cc_51 VPB N_A_93_264#_c_95_n 0.00202512f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=2.99
cc_52 VPB N_A_93_264#_c_86_n 0.0028976f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.79
cc_53 VPB N_A_93_264#_c_97_n 0.00527363f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=2.635
cc_54 VPB N_A_93_264#_c_98_n 0.00661228f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.875
cc_55 VPB N_A1_N_M1001_g 0.0283851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A2_N_c_226_n 0.0116045f $X=-0.19 $Y=1.66 $X2=2.595 $Y2=0.63
cc_57 VPB N_A2_N_M1007_g 0.0219185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_257_126#_M1009_g 0.0268165f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.81
cc_59 VPB N_A_257_126#_c_275_n 0.00773021f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=1.79
cc_60 VPB N_A_257_126#_c_276_n 0.00135977f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=2.635
cc_61 VPB N_A_257_126#_c_277_n 0.0058758f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.12
cc_62 VPB N_A_257_126#_c_273_n 0.0139187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B2_M1011_g 0.0228498f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.65
cc_64 VPB B2 0.00232698f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_65 VPB N_B2_c_340_n 0.0103695f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.81
cc_66 VPB N_B1_M1010_g 0.0409432f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.65
cc_67 VPB X 0.0481048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_410_n 0.0134913f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.12
cc_69 VPB N_X_c_408_n 0.00770854f $X=-0.19 $Y=1.66 $X2=2.735 $Y2=1.12
cc_70 VPB N_VPWR_c_431_n 0.00610667f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_71 VPB N_VPWR_c_432_n 0.00396743f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.81
cc_72 VPB N_VPWR_c_433_n 0.0227874f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.79
cc_73 VPB N_VPWR_c_434_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.875
cc_74 VPB N_VPWR_c_435_n 0.0504652f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=2.99
cc_75 VPB N_VPWR_c_436_n 0.0278922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_430_n 0.0837069f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.12
cc_77 VPB N_VPWR_c_438_n 0.00656574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_533_392#_c_478_n 0.00663239f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.65
cc_79 VPB N_A_533_392#_c_479_n 0.00179576f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.4
cc_80 VPB N_A_533_392#_c_480_n 0.00811042f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.32
cc_81 VPB N_A_533_392#_c_481_n 0.0125858f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.81
cc_82 VPB N_A_533_392#_c_482_n 0.0345796f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=1.65
cc_83 N_A_93_264#_M1000_g N_A1_N_M1001_g 0.033983f $X=0.7 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_93_264#_c_85_n N_A1_N_M1001_g 0.00278599f $X=0.815 $Y=1.79 $X2=0 $Y2=0
cc_85 N_A_93_264#_c_92_n N_A1_N_M1001_g 0.0170446f $X=1.325 $Y=1.875 $X2=0 $Y2=0
cc_86 N_A_93_264#_c_95_n N_A1_N_M1001_g 0.00125801f $X=1.495 $Y=2.99 $X2=0 $Y2=0
cc_87 N_A_93_264#_c_88_n N_A1_N_M1001_g 0.00100023f $X=0.63 $Y=1.485 $X2=0 $Y2=0
cc_88 N_A_93_264#_c_89_n N_A1_N_M1001_g 6.91159e-19 $X=0.815 $Y=1.485 $X2=0
+ $Y2=0
cc_89 N_A_93_264#_M1006_g A1_N 0.00242144f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_90 N_A_93_264#_c_92_n A1_N 0.0189017f $X=1.325 $Y=1.875 $X2=0 $Y2=0
cc_91 N_A_93_264#_c_88_n A1_N 2.74196e-19 $X=0.63 $Y=1.485 $X2=0 $Y2=0
cc_92 N_A_93_264#_c_89_n A1_N 0.0239351f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_93 N_A_93_264#_c_98_n A1_N 7.77974e-19 $X=1.41 $Y=1.875 $X2=0 $Y2=0
cc_94 N_A_93_264#_M1006_g N_A1_N_c_189_n 0.0205191f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_95 N_A_93_264#_c_92_n N_A1_N_c_189_n 0.00299885f $X=1.325 $Y=1.875 $X2=0
+ $Y2=0
cc_96 N_A_93_264#_c_89_n N_A1_N_c_189_n 0.00197815f $X=0.815 $Y=1.485 $X2=0
+ $Y2=0
cc_97 N_A_93_264#_M1006_g N_A1_N_c_190_n 0.0144354f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_98 N_A_93_264#_c_93_n N_A2_N_c_226_n 0.00661567f $X=2.02 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_93_264#_c_86_n N_A2_N_c_226_n 0.00653657f $X=2.105 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_93_264#_c_93_n N_A2_N_M1007_g 0.0137243f $X=2.02 $Y=1.875 $X2=0 $Y2=0
cc_101 N_A_93_264#_c_94_n N_A2_N_M1007_g 0.0159911f $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_102 N_A_93_264#_c_97_n N_A2_N_M1007_g 0.00319512f $X=2.35 $Y=2.635 $X2=0
+ $Y2=0
cc_103 N_A_93_264#_c_86_n N_A2_N_c_227_n 4.03823e-19 $X=2.105 $Y=1.79 $X2=0
+ $Y2=0
cc_104 N_A_93_264#_c_87_n N_A2_N_c_227_n 0.00551149f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_105 N_A_93_264#_c_93_n A2_N 0.022839f $X=2.02 $Y=1.875 $X2=0 $Y2=0
cc_106 N_A_93_264#_c_86_n A2_N 0.0309176f $X=2.105 $Y=1.79 $X2=0 $Y2=0
cc_107 N_A_93_264#_c_87_n A2_N 0.00263878f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_108 N_A_93_264#_c_94_n N_A_257_126#_M1007_d 0.00239704f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_109 N_A_93_264#_c_86_n N_A_257_126#_M1002_g 0.00584824f $X=2.105 $Y=1.79
+ $X2=0 $Y2=0
cc_110 N_A_93_264#_c_126_p N_A_257_126#_M1002_g 0.0108693f $X=2.735 $Y=1.12
+ $X2=0 $Y2=0
cc_111 N_A_93_264#_c_93_n N_A_257_126#_M1009_g 0.00100065f $X=2.02 $Y=1.875
+ $X2=0 $Y2=0
cc_112 N_A_93_264#_c_94_n N_A_257_126#_M1009_g 0.00699354f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_113 N_A_93_264#_c_97_n N_A_257_126#_M1009_g 0.00705138f $X=2.35 $Y=2.635
+ $X2=0 $Y2=0
cc_114 N_A_93_264#_M1006_g N_A_257_126#_c_269_n 6.54731e-19 $X=0.72 $Y=0.81
+ $X2=0 $Y2=0
cc_115 N_A_93_264#_M1009_s N_A_257_126#_c_275_n 0.00742973f $X=2.225 $Y=1.96
+ $X2=0 $Y2=0
cc_116 N_A_93_264#_c_93_n N_A_257_126#_c_275_n 0.0160722f $X=2.02 $Y=1.875 $X2=0
+ $Y2=0
cc_117 N_A_93_264#_c_94_n N_A_257_126#_c_275_n 0.00588659f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_118 N_A_93_264#_c_97_n N_A_257_126#_c_275_n 0.02253f $X=2.35 $Y=2.635 $X2=0
+ $Y2=0
cc_119 N_A_93_264#_M1009_s N_A_257_126#_c_276_n 0.00298247f $X=2.225 $Y=1.96
+ $X2=0 $Y2=0
cc_120 N_A_93_264#_c_93_n N_A_257_126#_c_276_n 0.014357f $X=2.02 $Y=1.875 $X2=0
+ $Y2=0
cc_121 N_A_93_264#_c_93_n N_A_257_126#_c_277_n 0.0243536f $X=2.02 $Y=1.875 $X2=0
+ $Y2=0
cc_122 N_A_93_264#_c_94_n N_A_257_126#_c_277_n 0.0203767f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_123 N_A_93_264#_c_97_n N_A_257_126#_c_277_n 0.0204056f $X=2.35 $Y=2.635 $X2=0
+ $Y2=0
cc_124 N_A_93_264#_c_86_n N_A_257_126#_c_272_n 0.02533f $X=2.105 $Y=1.79 $X2=0
+ $Y2=0
cc_125 N_A_93_264#_c_126_p N_A_257_126#_c_272_n 0.0142216f $X=2.735 $Y=1.12
+ $X2=0 $Y2=0
cc_126 N_A_93_264#_c_86_n N_A_257_126#_c_273_n 0.00319608f $X=2.105 $Y=1.79
+ $X2=0 $Y2=0
cc_127 N_A_93_264#_c_97_n N_A_257_126#_c_273_n 3.26401e-19 $X=2.35 $Y=2.635
+ $X2=0 $Y2=0
cc_128 N_A_93_264#_c_126_p N_A_257_126#_c_273_n 0.00161255f $X=2.735 $Y=1.12
+ $X2=0 $Y2=0
cc_129 N_A_93_264#_c_126_p N_B2_M1003_g 0.00425018f $X=2.735 $Y=1.12 $X2=0 $Y2=0
cc_130 N_A_93_264#_c_94_n N_B2_M1011_g 2.99783e-19 $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_131 N_A_93_264#_c_126_p B2 0.00133508f $X=2.735 $Y=1.12 $X2=0 $Y2=0
cc_132 N_A_93_264#_c_126_p N_B1_M1008_g 5.52341e-19 $X=2.735 $Y=1.12 $X2=0 $Y2=0
cc_133 N_A_93_264#_M1006_g N_X_c_406_n 6.44746e-19 $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_134 N_A_93_264#_c_88_n N_X_c_407_n 0.00288561f $X=0.63 $Y=1.485 $X2=0 $Y2=0
cc_135 N_A_93_264#_c_89_n N_X_c_407_n 0.0101951f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_136 N_A_93_264#_M1000_g N_X_c_410_n 0.00194972f $X=0.7 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_93_264#_c_153_p N_X_c_410_n 0.00672505f $X=0.9 $Y=1.875 $X2=0 $Y2=0
cc_138 N_A_93_264#_c_88_n N_X_c_410_n 0.00218979f $X=0.63 $Y=1.485 $X2=0 $Y2=0
cc_139 N_A_93_264#_c_89_n N_X_c_410_n 0.00792733f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_140 N_A_93_264#_M1000_g N_X_c_408_n 0.00225904f $X=0.7 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_93_264#_M1006_g N_X_c_408_n 0.00337861f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_142 N_A_93_264#_c_85_n N_X_c_408_n 0.00424168f $X=0.815 $Y=1.79 $X2=0 $Y2=0
cc_143 N_A_93_264#_c_88_n N_X_c_408_n 0.00231223f $X=0.63 $Y=1.485 $X2=0 $Y2=0
cc_144 N_A_93_264#_c_89_n N_X_c_408_n 0.0253043f $X=0.815 $Y=1.485 $X2=0 $Y2=0
cc_145 N_A_93_264#_c_92_n N_VPWR_M1000_d 0.0015839f $X=1.325 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_93_264#_c_153_p N_VPWR_M1000_d 5.61821e-19 $X=0.9 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_93_264#_M1000_g N_VPWR_c_431_n 0.0197727f $X=0.7 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_93_264#_c_92_n N_VPWR_c_431_n 0.0144497f $X=1.325 $Y=1.875 $X2=0
+ $Y2=0
cc_149 N_A_93_264#_c_153_p N_VPWR_c_431_n 0.00679503f $X=0.9 $Y=1.875 $X2=0
+ $Y2=0
cc_150 N_A_93_264#_c_95_n N_VPWR_c_431_n 0.00802251f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_151 N_A_93_264#_c_94_n N_VPWR_c_432_n 0.00280782f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_152 N_A_93_264#_M1000_g N_VPWR_c_433_n 0.00460063f $X=0.7 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_93_264#_c_94_n N_VPWR_c_435_n 0.0672123f $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_154 N_A_93_264#_c_95_n N_VPWR_c_435_n 0.0121867f $X=1.495 $Y=2.99 $X2=0 $Y2=0
cc_155 N_A_93_264#_M1000_g N_VPWR_c_430_n 0.00912809f $X=0.7 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_93_264#_c_94_n N_VPWR_c_430_n 0.0377688f $X=2.185 $Y=2.99 $X2=0 $Y2=0
cc_157 N_A_93_264#_c_95_n N_VPWR_c_430_n 0.00660921f $X=1.495 $Y=2.99 $X2=0
+ $Y2=0
cc_158 N_A_93_264#_c_174_p A_261_392# 0.0031191f $X=1.41 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_93_264#_c_94_n N_A_533_392#_c_479_n 0.00341172f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_160 N_A_93_264#_c_87_n N_VGND_M1005_d 0.00555114f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_161 N_A_93_264#_c_126_p N_VGND_M1005_d 0.00864797f $X=2.735 $Y=1.12 $X2=0
+ $Y2=0
cc_162 N_A_93_264#_M1006_g N_VGND_c_503_n 0.0147184f $X=0.72 $Y=0.81 $X2=0 $Y2=0
cc_163 N_A_93_264#_c_89_n N_VGND_c_503_n 0.00542821f $X=0.815 $Y=1.485 $X2=0
+ $Y2=0
cc_164 N_A_93_264#_M1002_d N_VGND_c_519_n 0.00370806f $X=2.595 $Y=0.63 $X2=0
+ $Y2=0
cc_165 N_A_93_264#_c_87_n N_VGND_c_519_n 0.013831f $X=2.19 $Y=1.12 $X2=0 $Y2=0
cc_166 N_A_93_264#_c_126_p N_VGND_c_519_n 0.0389185f $X=2.735 $Y=1.12 $X2=0
+ $Y2=0
cc_167 N_A_93_264#_M1002_d N_VGND_c_504_n 6.84302e-19 $X=2.595 $Y=0.63 $X2=0
+ $Y2=0
cc_168 N_A_93_264#_M1006_g N_VGND_c_506_n 0.00438299f $X=0.72 $Y=0.81 $X2=0
+ $Y2=0
cc_169 N_A_93_264#_c_126_p N_VGND_c_512_n 0.00469776f $X=2.735 $Y=1.12 $X2=0
+ $Y2=0
cc_170 N_A_93_264#_M1006_g N_VGND_c_514_n 0.00439883f $X=0.72 $Y=0.81 $X2=0
+ $Y2=0
cc_171 N_A1_N_M1001_g N_A2_N_c_226_n 0.0824247f $X=1.215 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_172 A1_N N_A2_N_c_226_n 0.00115052f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_173 N_A1_N_c_189_n N_A2_N_c_226_n 0.0201104f $X=1.17 $Y=1.455 $X2=-0.19
+ $Y2=-0.245
cc_174 A1_N N_A2_N_c_227_n 3.7319e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A1_N_c_190_n N_A2_N_c_227_n 0.0181059f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_176 A1_N A2_N 0.0281622f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_N_c_189_n A2_N 0.00114978f $X=1.17 $Y=1.455 $X2=0 $Y2=0
cc_178 N_A1_N_c_190_n A2_N 3.57707e-19 $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_179 A1_N N_A_257_126#_M1004_d 5.24173e-19 $X=1.115 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A1_N_c_190_n N_A_257_126#_c_268_n 0.00103147f $X=1.17 $Y=1.29 $X2=0
+ $Y2=0
cc_181 N_A1_N_M1001_g N_VPWR_c_431_n 0.00596796f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_182 N_A1_N_M1001_g N_VPWR_c_435_n 0.00553757f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_183 N_A1_N_M1001_g N_VPWR_c_430_n 0.0108852f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_184 A1_N N_VGND_M1006_d 0.00184725f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_185 A1_N N_VGND_c_503_n 0.0014989f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A1_N_c_189_n N_VGND_c_503_n 0.0027243f $X=1.17 $Y=1.455 $X2=0 $Y2=0
cc_187 N_A1_N_c_190_n N_VGND_c_503_n 0.0031179f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_188 N_A1_N_c_190_n N_VGND_c_508_n 0.00412698f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_189 N_A1_N_c_190_n N_VGND_c_514_n 0.00468052f $X=1.17 $Y=1.29 $X2=0 $Y2=0
cc_190 A2_N N_A_257_126#_M1004_d 2.07485e-19 $X=1.595 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_191 N_A2_N_c_226_n N_A_257_126#_M1002_g 0.00209308f $X=1.605 $Y=1.82 $X2=0
+ $Y2=0
cc_192 N_A2_N_c_227_n N_A_257_126#_c_268_n 0.0172182f $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_193 A2_N N_A_257_126#_c_268_n 0.00272717f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A2_N_c_227_n N_A_257_126#_c_269_n 7.6083e-19 $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_195 N_A2_N_c_227_n N_A_257_126#_c_270_n 0.00657983f $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_196 A2_N N_A_257_126#_c_270_n 0.0044198f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A2_N_c_227_n N_A_257_126#_c_271_n 3.36612e-19 $X=1.64 $Y=1.29 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_226_n N_A_257_126#_c_276_n 4.66378e-19 $X=1.605 $Y=1.82 $X2=0
+ $Y2=0
cc_199 N_A2_N_M1007_g N_A_257_126#_c_276_n 0.00240499f $X=1.605 $Y=2.46 $X2=0
+ $Y2=0
cc_200 N_A2_N_M1007_g N_A_257_126#_c_277_n 0.00840368f $X=1.605 $Y=2.46 $X2=0
+ $Y2=0
cc_201 N_A2_N_c_226_n N_A_257_126#_c_273_n 0.00502857f $X=1.605 $Y=1.82 $X2=0
+ $Y2=0
cc_202 N_A2_N_M1007_g N_VPWR_c_435_n 0.00333926f $X=1.605 $Y=2.46 $X2=0 $Y2=0
cc_203 N_A2_N_M1007_g N_VPWR_c_430_n 0.00427327f $X=1.605 $Y=2.46 $X2=0 $Y2=0
cc_204 A2_N N_VGND_M1005_d 0.00228426f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_205 N_A2_N_c_226_n N_VGND_c_519_n 0.00115762f $X=1.605 $Y=1.82 $X2=0 $Y2=0
cc_206 A2_N N_VGND_c_519_n 0.0041082f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_207 N_A2_N_c_227_n N_VGND_c_508_n 5.45085e-19 $X=1.64 $Y=1.29 $X2=0 $Y2=0
cc_208 N_A_257_126#_c_271_n N_B2_M1003_g 0.0270626f $X=2.43 $Y=0.355 $X2=0 $Y2=0
cc_209 N_A_257_126#_M1009_g N_B2_M1011_g 0.0143419f $X=2.575 $Y=2.46 $X2=0 $Y2=0
cc_210 N_A_257_126#_c_276_n N_B2_M1011_g 8.93354e-19 $X=2.445 $Y=2.13 $X2=0
+ $Y2=0
cc_211 N_A_257_126#_c_272_n B2 0.0208896f $X=2.5 $Y=1.615 $X2=0 $Y2=0
cc_212 N_A_257_126#_c_273_n B2 0.00114361f $X=2.5 $Y=1.615 $X2=0 $Y2=0
cc_213 N_A_257_126#_c_272_n N_B2_c_340_n 4.14706e-19 $X=2.5 $Y=1.615 $X2=0 $Y2=0
cc_214 N_A_257_126#_c_273_n N_B2_c_340_n 0.0207787f $X=2.5 $Y=1.615 $X2=0 $Y2=0
cc_215 N_A_257_126#_M1009_g N_VPWR_c_432_n 5.80216e-19 $X=2.575 $Y=2.46 $X2=0
+ $Y2=0
cc_216 N_A_257_126#_M1009_g N_VPWR_c_435_n 0.00517089f $X=2.575 $Y=2.46 $X2=0
+ $Y2=0
cc_217 N_A_257_126#_M1009_g N_VPWR_c_430_n 0.00983819f $X=2.575 $Y=2.46 $X2=0
+ $Y2=0
cc_218 N_A_257_126#_c_276_n N_A_533_392#_c_478_n 0.00580234f $X=2.445 $Y=2.13
+ $X2=0 $Y2=0
cc_219 N_A_257_126#_c_268_n N_VGND_c_503_n 0.0223974f $X=1.425 $Y=0.845 $X2=0
+ $Y2=0
cc_220 N_A_257_126#_c_269_n N_VGND_c_503_n 0.0219867f $X=1.59 $Y=0.387 $X2=0
+ $Y2=0
cc_221 N_A_257_126#_M1002_g N_VGND_c_519_n 0.00837945f $X=2.52 $Y=0.95 $X2=0
+ $Y2=0
cc_222 N_A_257_126#_c_270_n N_VGND_c_519_n 0.0573731f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_223 N_A_257_126#_c_271_n N_VGND_c_519_n 0.00391065f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_224 N_A_257_126#_c_270_n N_VGND_c_504_n 0.0210179f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_225 N_A_257_126#_c_271_n N_VGND_c_504_n 0.00727503f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_226 N_A_257_126#_c_269_n N_VGND_c_508_n 0.0218645f $X=1.59 $Y=0.387 $X2=0
+ $Y2=0
cc_227 N_A_257_126#_c_270_n N_VGND_c_508_n 0.0657312f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_228 N_A_257_126#_c_271_n N_VGND_c_508_n 0.00641604f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_229 N_A_257_126#_c_269_n N_VGND_c_514_n 0.0118577f $X=1.59 $Y=0.387 $X2=0
+ $Y2=0
cc_230 N_A_257_126#_c_270_n N_VGND_c_514_n 0.0366452f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_231 N_A_257_126#_c_271_n N_VGND_c_514_n 0.00987452f $X=2.43 $Y=0.355 $X2=0
+ $Y2=0
cc_232 N_B2_M1011_g N_B1_M1010_g 0.0263066f $X=3.025 $Y=2.46 $X2=0 $Y2=0
cc_233 B2 N_B1_M1010_g 0.00756601f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B2_c_340_n N_B1_M1010_g 0.0198084f $X=3.04 $Y=1.615 $X2=0 $Y2=0
cc_235 N_B2_M1003_g N_B1_c_380_n 0.0258771f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_236 N_B2_M1011_g N_VPWR_c_432_n 0.0129269f $X=3.025 $Y=2.46 $X2=0 $Y2=0
cc_237 N_B2_M1011_g N_VPWR_c_435_n 0.00460063f $X=3.025 $Y=2.46 $X2=0 $Y2=0
cc_238 N_B2_M1011_g N_VPWR_c_430_n 0.00908665f $X=3.025 $Y=2.46 $X2=0 $Y2=0
cc_239 B2 N_A_533_392#_c_478_n 8.43333e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B2_c_340_n N_A_533_392#_c_478_n 2.72398e-19 $X=3.04 $Y=1.615 $X2=0
+ $Y2=0
cc_241 N_B2_M1011_g N_A_533_392#_c_480_n 0.014478f $X=3.025 $Y=2.46 $X2=0 $Y2=0
cc_242 B2 N_A_533_392#_c_480_n 0.0257171f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B2_c_340_n N_A_533_392#_c_480_n 0.00333368f $X=3.04 $Y=1.615 $X2=0
+ $Y2=0
cc_244 N_B2_M1003_g N_VGND_c_519_n 0.00564957f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_245 B2 N_VGND_c_519_n 9.81631e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_246 N_B2_M1003_g N_VGND_c_504_n 0.00515291f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_247 N_B2_M1003_g N_VGND_c_505_n 0.00266787f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_248 N_B2_M1003_g N_VGND_c_553_n 0.00425334f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_249 B2 N_VGND_c_553_n 0.00366871f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_250 N_B2_c_340_n N_VGND_c_553_n 0.00117163f $X=3.04 $Y=1.615 $X2=0 $Y2=0
cc_251 N_B2_M1003_g N_VGND_c_510_n 0.00246733f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_252 N_B2_M1003_g N_VGND_c_512_n 0.00102955f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_253 N_B2_M1003_g N_VGND_c_514_n 0.00283952f $X=2.95 $Y=0.95 $X2=0 $Y2=0
cc_254 N_B1_M1010_g N_VPWR_c_432_n 0.0160415f $X=3.505 $Y=2.46 $X2=0 $Y2=0
cc_255 N_B1_M1010_g N_VPWR_c_436_n 0.00460063f $X=3.505 $Y=2.46 $X2=0 $Y2=0
cc_256 N_B1_M1010_g N_VPWR_c_430_n 0.00913687f $X=3.505 $Y=2.46 $X2=0 $Y2=0
cc_257 N_B1_M1010_g N_A_533_392#_c_480_n 0.0191613f $X=3.505 $Y=2.46 $X2=0 $Y2=0
cc_258 N_B1_M1010_g N_A_533_392#_c_481_n 4.17659e-19 $X=3.505 $Y=2.46 $X2=0
+ $Y2=0
cc_259 N_B1_M1010_g N_A_533_392#_c_482_n 4.69176e-19 $X=3.505 $Y=2.46 $X2=0
+ $Y2=0
cc_260 B1 N_VGND_M1008_d 0.0022726f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_261 B1 N_VGND_c_505_n 0.0330236f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_262 N_B1_c_380_n N_VGND_c_505_n 0.0137935f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_263 N_B1_M1008_g N_VGND_c_562_n 0.0124674f $X=3.49 $Y=0.95 $X2=0 $Y2=0
cc_264 B1 N_VGND_c_562_n 0.00390864f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_265 N_B1_M1008_g N_VGND_c_512_n 0.00872234f $X=3.49 $Y=0.95 $X2=0 $Y2=0
cc_266 N_B1_c_377_n N_VGND_c_512_n 0.00115069f $X=3.505 $Y=1.435 $X2=0 $Y2=0
cc_267 B1 N_VGND_c_512_n 0.0221741f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_268 N_B1_c_380_n N_VGND_c_512_n 0.00120812f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_269 B1 N_VGND_c_513_n 0.0476503f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_270 N_B1_c_380_n N_VGND_c_513_n 0.00865075f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_271 B1 N_VGND_c_514_n 0.0257336f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_272 N_B1_c_380_n N_VGND_c_514_n 0.0119279f $X=3.65 $Y=0.355 $X2=0 $Y2=0
cc_273 X N_VPWR_c_431_n 0.0287387f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_274 X N_VPWR_c_433_n 0.0193209f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_275 X N_VPWR_c_430_n 0.0159921f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_276 N_X_c_406_n N_VGND_c_503_n 0.021946f $X=0.505 $Y=0.585 $X2=0 $Y2=0
cc_277 N_X_c_406_n N_VGND_c_506_n 0.0161045f $X=0.505 $Y=0.585 $X2=0 $Y2=0
cc_278 N_X_c_406_n N_VGND_c_514_n 0.0163598f $X=0.505 $Y=0.585 $X2=0 $Y2=0
cc_279 N_VPWR_c_432_n N_A_533_392#_c_479_n 0.0236746f $X=3.265 $Y=2.455 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_435_n N_A_533_392#_c_479_n 0.00749631f $X=3.085 $Y=3.33 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_430_n N_A_533_392#_c_479_n 0.0062048f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_282 N_VPWR_M1011_d N_A_533_392#_c_480_n 0.00197722f $X=3.115 $Y=1.96 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_432_n N_A_533_392#_c_480_n 0.0194666f $X=3.265 $Y=2.455 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_432_n N_A_533_392#_c_482_n 0.0237131f $X=3.265 $Y=2.455 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_436_n N_A_533_392#_c_482_n 0.011066f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VPWR_c_430_n N_A_533_392#_c_482_n 0.00915947f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_287 N_A_533_392#_c_480_n N_VGND_c_512_n 0.00295854f $X=3.645 $Y=2.035 $X2=0
+ $Y2=0
cc_288 N_A_533_392#_c_481_n N_VGND_c_512_n 0.00793931f $X=3.77 $Y=2.12 $X2=0
+ $Y2=0
cc_289 N_VGND_c_505_n A_605_126# 0.00487694f $X=3.23 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_290 N_VGND_c_562_n A_605_126# 0.00244694f $X=3.54 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_291 N_VGND_c_553_n A_605_126# 0.00779459f $X=3.315 $Y=0.925 $X2=-0.19
+ $Y2=-0.245

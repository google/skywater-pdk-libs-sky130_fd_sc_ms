* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_685_140# a_27_74# a_412_140# VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=5.888e+11p ps=5.68e+06u
M1001 a_685_140# C a_882_137# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.888e+11p ps=5.68e+06u
M1002 a_412_140# a_27_74# a_685_140# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=3.5296e+12p pd=2.358e+07u as=2.8e+11p ps=2.56e+06u
M1004 a_475_388# D VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.3525e+12p pd=1.087e+07u as=0p ps=0u
M1005 X a_475_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1006 VPWR a_475_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_475_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_475_388# X VNB nlowvt w=740000u l=150000u
+  ad=1.1064e+12p pd=1.017e+07u as=4.44e+11p ps=4.16e+06u
M1009 a_475_388# a_200_74# a_412_140# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1010 VGND D a_882_137# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_475_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_475_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_475_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR D a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_475_388# a_200_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_475_388# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_200_74# a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR C a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_27_74# a_475_388# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_475_388# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_475_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_200_74# A_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1023 VGND B_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1024 a_200_74# A_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.915e+11p pd=1.99e+06u as=0p ps=0u
M1025 a_882_137# C a_685_140# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_882_137# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_412_140# a_200_74# a_475_388# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__nand4_1.pex.spice
* Created: Fri Aug 28 17:44:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4_1%D 3 7 8 11 13
r30 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=1.385
+ $X2=0.74 $Y2=1.55
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=1.385
+ $X2=0.74 $Y2=1.22
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.385 $X2=0.74 $Y2=1.385
r33 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.74 $Y=1.295 $X2=0.74
+ $Y2=1.385
r34 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.83 $Y=0.74 $X2=0.83
+ $Y2=1.22
r35 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.815 $Y=2.4
+ $X2=0.815 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_1%C 3 6 8 11 12 13
c34 13 0 3.78555e-20 $X=1.31 $Y=1.22
c35 12 0 1.64093e-19 $X=1.31 $Y=1.385
r36 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.385
+ $X2=1.31 $Y2=1.55
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.385
+ $X2=1.31 $Y2=1.22
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.385 $X2=1.31 $Y2=1.385
r39 8 12 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=1.365 $X2=1.31
+ $Y2=1.365
r40 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.265 $Y=2.4
+ $X2=1.265 $Y2=1.55
r41 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.22 $Y=0.74 $X2=1.22
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_1%B 3 6 8 11 13
c36 13 0 1.64093e-19 $X=1.88 $Y=1.22
c37 8 0 3.78555e-20 $X=2.16 $Y=1.295
r38 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.385
+ $X2=1.88 $Y2=1.55
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.385
+ $X2=1.88 $Y2=1.22
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.385 $X2=1.88 $Y2=1.385
r41 8 12 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=1.88 $Y2=1.365
r42 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.875 $Y=2.4
+ $X2=1.875 $Y2=1.55
r43 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.79 $Y=0.74 $X2=1.79
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_1%A 1 3 6 8 14
c23 6 0 1.85286e-19 $X=2.375 $Y=2.4
r24 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r25 12 14 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.375 $Y=1.385
+ $X2=2.61 $Y2=1.385
r26 10 12 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.36 $Y=1.385
+ $X2=2.375 $Y2=1.385
r27 8 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.385
r28 4 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.55
+ $X2=2.375 $Y2=1.385
r29 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.375 $Y=1.55
+ $X2=2.375 $Y2=2.4
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.22
+ $X2=2.36 $Y2=1.385
r31 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.36 $Y=1.22 $X2=2.36
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_1%VPWR 1 2 3 12 18 20 22 27 28 30 31 32 41 47
c40 1 0 1.38338e-19 $X=0.395 $Y=1.84
r41 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 41 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.657 $Y2=3.33
r45 41 43 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 36 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 32 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 32 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 30 39 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.565 $Y2=3.33
r53 29 43 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=1.565 $Y2=3.33
r55 27 35 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.54 $Y2=3.33
r57 26 39 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.705 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=3.33
+ $X2=0.54 $Y2=3.33
r59 22 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.6 $Y=1.985 $X2=2.6
+ $Y2=2.815
r60 20 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.6 $Y=3.245
+ $X2=2.657 $Y2=3.33
r61 20 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.6 $Y=3.245 $X2=2.6
+ $Y2=2.815
r62 16 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=3.245
+ $X2=1.565 $Y2=3.33
r63 16 18 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.565 $Y=3.245
+ $X2=1.565 $Y2=2.405
r64 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.54 $Y=2.145
+ $X2=0.54 $Y2=2.825
r65 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.54 $Y=3.245
+ $X2=0.54 $Y2=3.33
r66 10 15 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.54 $Y=3.245
+ $X2=0.54 $Y2=2.825
r67 3 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=2.815
r68 3 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=1.985
r69 2 18 300 $w=1.7e-07 $l=6.61721e-07 $layer=licon1_PDIFF $count=2 $X=1.355
+ $Y=1.84 $X2=1.565 $Y2=2.405
r70 1 15 400 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.84 $X2=0.54 $Y2=2.825
r71 1 12 400 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.84 $X2=0.54 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_1%Y 1 2 3 11 12 13 14 15 18 20 22 26 30 31 34
c78 20 0 1.85286e-19 $X=2.1 $Y=2.15
c79 15 0 1.38338e-19 $X=0.405 $Y=1.805
r80 31 34 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=1.985
+ $X2=1.68 $Y2=1.985
r81 31 33 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=1.985
+ $X2=2.1 $Y2=1.985
r82 28 34 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.205 $Y=1.985
+ $X2=1.68 $Y2=1.985
r83 28 30 6.46576 $w=2.5e-07 $l=1.88348e-07 $layer=LI1_cond $X=1.205 $Y=1.985
+ $X2=1.04 $Y2=1.935
r84 24 26 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.575 $Y=0.84
+ $X2=2.575 $Y2=0.515
r85 20 33 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=2.15 $X2=2.1
+ $Y2=1.985
r86 20 22 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.1 $Y=2.15 $X2=2.1
+ $Y2=2.815
r87 16 30 0.364692 $w=3.3e-07 $l=2.15e-07 $layer=LI1_cond $X=1.04 $Y=2.15
+ $X2=1.04 $Y2=1.935
r88 16 18 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.04 $Y=2.15
+ $X2=1.04 $Y2=2.815
r89 14 30 6.46576 $w=2.5e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.875 $Y=1.805
+ $X2=1.04 $Y2=1.935
r90 14 15 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=0.875 $Y=1.805
+ $X2=0.405 $Y2=1.805
r91 12 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.41 $Y=0.925
+ $X2=2.575 $Y2=0.84
r92 12 13 130.807 $w=1.68e-07 $l=2.005e-06 $layer=LI1_cond $X=2.41 $Y=0.925
+ $X2=0.405 $Y2=0.925
r93 11 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.72
+ $X2=0.405 $Y2=1.805
r94 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.32 $Y=1.01
+ $X2=0.405 $Y2=0.925
r95 10 11 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.32 $Y=1.01
+ $X2=0.32 $Y2=1.72
r96 3 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.84 $X2=2.1 $Y2=1.985
r97 3 22 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.84 $X2=2.1 $Y2=2.815
r98 2 30 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.84 $X2=1.04 $Y2=1.985
r99 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.84 $X2=1.04 $Y2=2.815
r100 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.435
+ $Y=0.37 $X2=2.575 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_1%VGND 1 4 8 9 12
r20 13 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r21 12 17 8.95014 $w=7.02e-07 $l=5.15e-07 $layer=LI1_cond $X=0.392 $Y=0
+ $X2=0.392 $Y2=0.515
r22 12 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r23 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 8 9 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r25 6 12 9.34032 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.392
+ $Y2=0
r26 6 8 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=0.785 $Y=0 $X2=2.64
+ $Y2=0
r27 4 9 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r28 4 15 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r29 1 17 91 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.615 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__clkinv_1.spice
* Created: Fri Aug 28 17:19:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkinv_1.pex.spice"
.subckt sky130_fd_sc_ms__clkinv_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.22535 AS=0.1491 PD=2.17 PS=1.55 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.3
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=0.84 AD=0.1134
+ AS=0.2268 PD=1.11 PS=2.22 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2 SB=90000.6
+ A=0.1512 P=2.04 MULT=1
MM1002 N_Y_M1001_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=0.84 AD=0.1134
+ AS=0.2268 PD=1.11 PS=2.22 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.6 SB=90000.2
+ A=0.1512 P=2.04 MULT=1
DX3_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_ms__clkinv_1.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__fah_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_416_392# A VGND VNB nlowvt w=640000u l=150000u
+  ad=4.247e+11p pd=4.22e+06u as=1.82425e+12p ps=1.593e+07u
M1001 COUT a_1454_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=2.404e+12p ps=1.999e+07u
M1002 a_852_424# a_481_379# a_117_368# VPB pshort w=840000u l=180000u
+  ad=1.1046e+12p pd=4.31e+06u as=6.58e+11p ps=5.31e+06u
M1003 a_517_424# B a_416_392# VNB nlowvt w=640000u l=150000u
+  ad=3.904e+11p pd=2.5e+06u as=0p ps=0u
M1004 a_852_424# B a_117_368# VNB nlowvt w=640000u l=150000u
+  ad=4.448e+11p pd=2.67e+06u as=7.401e+11p ps=4.99e+06u
M1005 a_117_368# a_481_379# a_517_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_1454_424# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_1898_424# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 a_1898_424# a_852_424# a_1692_424# VNB nlowvt w=640000u l=150000u
+  ad=4.729e+11p pd=2.9e+06u as=6.112e+11p ps=4.47e+06u
M1009 SUM a_1898_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_1692_424# a_2055_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1011 COUT a_1454_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 VGND A a_81_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.272e+11p ps=1.99e+06u
M1013 a_1454_424# a_852_424# a_481_379# VNB nlowvt w=640000u l=150000u
+  ad=5.6e+11p pd=3.03e+06u as=2.33e+11p ps=2.13e+06u
M1014 a_416_392# B a_852_424# VPB pshort w=840000u l=180000u
+  ad=5.398e+11p pd=4.87e+06u as=0p ps=0u
M1015 a_1692_424# a_517_424# a_1454_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1898_424# a_517_424# a_1692_424# VPB pshort w=840000u l=180000u
+  ad=5.082e+11p pd=2.89e+06u as=9.84e+11p ps=5.92e+06u
M1017 a_1692_424# CI VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1898_424# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.146e+11p ps=2.06e+06u
M1019 a_416_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1692_424# a_2055_424# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.642e+11p ps=3.01e+06u
M1021 a_1454_424# a_517_424# a_481_379# VPB pshort w=840000u l=180000u
+  ad=8.484e+11p pd=3.7e+06u as=3.654e+11p ps=2.93e+06u
M1022 a_2055_424# a_852_424# a_1898_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1692_424# CI VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_117_368# a_81_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_481_379# B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1692_424# a_852_424# a_1454_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_416_392# a_481_379# a_852_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_2055_424# a_517_424# a_1898_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A a_81_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1030 a_517_424# a_481_379# a_416_392# VPB pshort w=840000u l=180000u
+  ad=7.434e+11p pd=3.45e+06u as=0p ps=0u
M1031 SUM a_1898_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_117_368# B a_517_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_481_379# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_117_368# a_81_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_1454_424# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__a222o_1.pex.spice
* Created: Wed Sep  2 11:52:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A222O_1%C1 3 7 8 9 13 14 15
c29 14 0 1.41241e-19 $X=0.385 $Y=1.285
r30 13 16 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.285
+ $X2=0.407 $Y2=1.45
r31 13 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.285
+ $X2=0.407 $Y2=1.12
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.285 $X2=0.385 $Y2=1.285
r33 8 9 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r34 8 14 0.271163 $w=4.23e-07 $l=1e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.285
r35 7 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.52 $Y=0.69 $X2=0.52
+ $Y2=1.12
r36 3 16 388.71 $w=1.8e-07 $l=1e-06 $layer=POLY_cond $X=0.505 $Y=2.45 $X2=0.505
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%C2 1 3 6 8 11
c38 11 0 1.41241e-19 $X=1.11 $Y=1.285
c39 6 0 1.72297e-19 $X=1.11 $Y=2.45
r40 11 13 20.5296 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=1.11 $Y=1.285
+ $X2=1.225 $Y2=1.285
r41 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.285 $X2=1.225 $Y2=1.285
r42 4 11 12.2893 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.45
+ $X2=1.11 $Y2=1.285
r43 4 6 388.71 $w=1.8e-07 $l=1e-06 $layer=POLY_cond $X=1.11 $Y=1.45 $X2=1.11
+ $Y2=2.45
r44 1 11 35.7037 $w=2.7e-07 $l=2.70185e-07 $layer=POLY_cond $X=0.91 $Y=1.12
+ $X2=1.11 $Y2=1.285
r45 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.91 $Y=1.12 $X2=0.91
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%B2 3 8 10 11 12 15
c45 11 0 3.57238e-19 $X=1.635 $Y=1.84
r46 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r47 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.18
r48 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.345 $X2=1.765 $Y2=1.345
r49 10 11 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.635 $Y=1.69
+ $X2=1.635 $Y2=1.84
r50 10 18 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.675 $Y=1.69
+ $X2=1.675 $Y2=1.51
r51 8 17 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.855 $Y=0.69
+ $X2=1.855 $Y2=1.18
r52 3 11 163.344 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.61 $Y=2.45 $X2=1.61
+ $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%B1 1 3 8 9 10 11 15 16 17
c41 16 0 1.60193e-19 $X=2.385 $Y=1.285
r42 15 18 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=1.285
+ $X2=2.345 $Y2=1.45
r43 15 17 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=2.345 $Y=1.285
+ $X2=2.345 $Y2=1.12
r44 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.285 $X2=2.385 $Y2=1.285
r45 10 11 8.27194 $w=5.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.487 $Y=1.295
+ $X2=2.487 $Y2=1.665
r46 10 16 0.223566 $w=5.33e-07 $l=1e-08 $layer=LI1_cond $X=2.487 $Y=1.295
+ $X2=2.487 $Y2=1.285
r47 9 18 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.215 $Y=1.79
+ $X2=2.215 $Y2=1.45
r48 8 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.245 $Y=0.69
+ $X2=2.245 $Y2=1.12
r49 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.2 $Y=1.88 $X2=2.2
+ $Y2=1.79
r50 1 3 152.633 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=2.2 $Y=1.88 $X2=2.2
+ $Y2=2.45
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%A1 3 8 9 10 11 14 16
c34 11 0 7.1933e-20 $X=3.12 $Y=1.295
r35 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.285
+ $X2=3.09 $Y2=1.45
r36 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.285
+ $X2=3.09 $Y2=1.12
r37 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.285 $X2=3.09 $Y2=1.285
r38 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.227 $Y=1.69
+ $X2=3.227 $Y2=1.84
r39 9 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.18 $Y=1.69 $X2=3.18
+ $Y2=1.45
r40 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.26 $Y=2.415
+ $X2=3.26 $Y2=1.84
r41 3 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.18 $Y=0.69 $X2=3.18
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%A2 3 6 8 11 13
c39 6 0 7.1933e-20 $X=3.71 $Y=2.415
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.285
+ $X2=3.66 $Y2=1.45
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.285
+ $X2=3.66 $Y2=1.12
r42 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.285 $X2=3.66 $Y2=1.285
r43 6 14 375.105 $w=1.8e-07 $l=9.65e-07 $layer=POLY_cond $X=3.71 $Y=2.415
+ $X2=3.71 $Y2=1.45
r44 3 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.57 $Y=0.69 $X2=3.57
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%A_32_74# 1 2 3 12 16 20 22 23 28 32 35 36 37
+ 40 41 45 46
r106 46 50 40.7387 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.212 $Y=1.465
+ $X2=4.212 $Y2=1.63
r107 46 49 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.212 $Y=1.465
+ $X2=4.212 $Y2=1.3
r108 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.465 $X2=4.205 $Y2=1.465
r109 42 45 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.1 $Y=1.465
+ $X2=4.205 $Y2=1.465
r110 39 41 10.2865 $w=6.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.64
+ $X2=3.13 $Y2=0.64
r111 39 40 20.0288 $w=6.18e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=0.64
+ $X2=2.295 $Y2=0.64
r112 35 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=1.3 $X2=4.1
+ $Y2=1.465
r113 34 35 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.1 $Y=0.95 $X2=4.1
+ $Y2=1.3
r114 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=0.865
+ $X2=4.1 $Y2=0.95
r115 32 41 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.015 $Y=0.865
+ $X2=3.13 $Y2=0.865
r116 31 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=0.865
+ $X2=0.805 $Y2=0.865
r117 31 40 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=0.89 $Y=0.865
+ $X2=2.295 $Y2=0.865
r118 28 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=2.095
+ $X2=0.885 $Y2=1.93
r119 24 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.95
+ $X2=0.805 $Y2=0.865
r120 24 37 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.805 $Y=0.95
+ $X2=0.805 $Y2=1.93
r121 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.865
+ $X2=0.805 $Y2=0.865
r122 22 23 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.72 $Y=0.865
+ $X2=0.47 $Y2=0.865
r123 18 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.47 $Y2=0.865
r124 18 20 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.305 $Y2=0.515
r125 16 49 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.305 $Y=0.74
+ $X2=4.305 $Y2=1.3
r126 12 50 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.295 $Y=2.4
+ $X2=4.295 $Y2=1.63
r127 3 28 300 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.95 $X2=0.885 $Y2=2.095
r128 2 39 45.5 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_NDIFF $count=4 $X=2.32
+ $Y=0.37 $X2=2.965 $Y2=0.495
r129 1 20 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.37 $X2=0.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%A_27_390# 1 2 3 12 16 17 20 24 28 30
c43 20 0 1.72297e-19 $X=1.385 $Y=2.095
r44 26 28 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.425 $Y=2.905
+ $X2=2.425 $Y2=2.465
r45 25 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=2.99
+ $X2=1.385 $Y2=2.99
r46 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.26 $Y=2.99
+ $X2=2.425 $Y2=2.905
r47 24 25 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.26 $Y=2.99
+ $X2=1.55 $Y2=2.99
r48 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.385 $Y=2.095
+ $X2=1.385 $Y2=2.805
r49 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=2.905
+ $X2=1.385 $Y2=2.99
r50 18 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.385 $Y=2.905
+ $X2=1.385 $Y2=2.805
r51 16 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=2.99
+ $X2=1.385 $Y2=2.99
r52 16 17 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.22 $Y=2.99
+ $X2=0.445 $Y2=2.99
r53 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.125
+ $X2=0.28 $Y2=2.805
r54 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r55 10 15 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.805
r56 3 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.95 $X2=2.425 $Y2=2.465
r57 2 23 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.95 $X2=1.385 $Y2=2.805
r58 2 20 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.95 $X2=1.385 $Y2=2.095
r59 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.95 $X2=0.28 $Y2=2.805
r60 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.95 $X2=0.28 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%A_340_390# 1 2 9 11 13 16
c33 16 0 1.97045e-19 $X=1.885 $Y=2.095
r34 11 18 2.90003 $w=3.3e-07 $l=1.18e-07 $layer=LI1_cond $X=3.485 $Y=2.13
+ $X2=3.485 $Y2=2.012
r35 11 13 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=3.485 $Y=2.13
+ $X2=3.485 $Y2=2.77
r36 10 16 4.99254 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.05 $Y=2.045
+ $X2=1.885 $Y2=2.03
r37 9 18 4.86615 $w=1.7e-07 $l=1.80748e-07 $layer=LI1_cond $X=3.32 $Y=2.045
+ $X2=3.485 $Y2=2.012
r38 9 10 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=3.32 $Y=2.045
+ $X2=2.05 $Y2=2.045
r39 2 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=1.915 $X2=3.485 $Y2=2.06
r40 2 13 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=1.915 $X2=3.485 $Y2=2.77
r41 1 16 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=1.7
+ $Y=1.95 $X2=1.885 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%VPWR 1 2 9 13 18 19 20 29 35 36 39
r49 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 36 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r52 33 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.02 $Y2=3.33
r53 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r54 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 29 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.02 $Y2=3.33
r57 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 28 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 23 27 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 20 24 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 18 27 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.985 $Y2=3.33
r66 17 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.15 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=2.985 $Y2=3.33
r68 13 16 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=4.02 $Y=2.06
+ $X2=4.02 $Y2=2.815
r69 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.33
r70 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=2.815
r71 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=3.245
+ $X2=2.985 $Y2=3.33
r72 7 9 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.985 $Y=3.245
+ $X2=2.985 $Y2=2.385
r73 2 16 400 $w=1.7e-07 $l=1.00399e-06 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=1.915 $X2=4.02 $Y2=2.815
r74 2 13 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=1.915 $X2=4.02 $Y2=2.06
r75 1 9 300 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_PDIFF $count=2 $X=2.84
+ $Y=1.915 $X2=2.985 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%X 1 2 9 13 14 15 16 23 32
r25 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=4.532 $Y=1.997
+ $X2=4.532 $Y2=2.035
r26 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=4.532 $Y=2.405
+ $X2=4.532 $Y2=2.775
r27 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=4.532 $Y=1.973
+ $X2=4.532 $Y2=1.997
r28 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=4.532 $Y=1.973
+ $X2=4.532 $Y2=1.82
r29 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=4.532 $Y=2.058
+ $X2=4.532 $Y2=2.405
r30 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=4.532 $Y=2.058
+ $X2=4.532 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.625 $Y=1.13
+ $X2=4.625 $Y2=1.82
r32 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=4.532 $Y=0.953
+ $X2=4.532 $Y2=1.13
r33 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=4.532 $Y=0.953
+ $X2=4.532 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.38
+ $Y=0.37 $X2=4.52 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_1%VGND 1 2 7 14 24 25 30 36
r43 34 36 10.0102 $w=6.83e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=1.805 $Y2=0.257
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 32 34 0.69844 $w=6.83e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=0.257 $X2=1.68
+ $Y2=0.257
r46 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r47 28 32 7.68284 $w=6.83e-07 $l=4.4e-07 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=1.64 $Y2=0.257
r48 28 30 12.0182 $w=6.83e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=0.96 $Y2=0.257
r49 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r51 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r52 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.56
+ $Y2=0
r53 21 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r54 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r56 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r57 17 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.805
+ $Y2=0
r58 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 14 42 10.9023 $w=5.63e-07 $l=5.15e-07 $layer=LI1_cond $X=3.902 $Y=0
+ $X2=3.902 $Y2=0.515
r60 14 22 7.93092 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=3.902 $Y=0 $X2=4.185
+ $Y2=0
r61 14 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 14 20 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.6
+ $Y2=0
r63 12 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 11 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.96
+ $Y2=0
r65 11 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 7 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.6
+ $Y2=0
r67 7 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r68 2 42 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=3.645
+ $Y=0.37 $X2=3.9 $Y2=0.515
r69 1 32 91 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.37 $X2=1.64 $Y2=0.515
.ends


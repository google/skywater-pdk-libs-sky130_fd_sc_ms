* File: sky130_fd_sc_ms__dfxbp_1.pxi.spice
* Created: Fri Aug 28 17:24:30 2020
* 
x_PM_SKY130_FD_SC_MS__DFXBP_1%CLK N_CLK_M1015_g N_CLK_c_208_n N_CLK_M1025_g CLK
+ N_CLK_c_209_n N_CLK_c_210_n PM_SKY130_FD_SC_MS__DFXBP_1%CLK
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_27_74# N_A_27_74#_M1025_s N_A_27_74#_M1015_s
+ N_A_27_74#_M1014_g N_A_27_74#_c_241_n N_A_27_74#_M1017_g N_A_27_74#_M1002_g
+ N_A_27_74#_M1003_g N_A_27_74#_c_264_n N_A_27_74#_M1023_g N_A_27_74#_c_243_n
+ N_A_27_74#_M1020_g N_A_27_74#_c_266_n N_A_27_74#_c_245_n N_A_27_74#_c_267_n
+ N_A_27_74#_c_246_n N_A_27_74#_c_268_n N_A_27_74#_c_269_n N_A_27_74#_c_283_n
+ N_A_27_74#_c_247_n N_A_27_74#_c_248_n N_A_27_74#_c_249_n N_A_27_74#_c_250_n
+ N_A_27_74#_c_251_n N_A_27_74#_c_252_n N_A_27_74#_c_253_n N_A_27_74#_c_271_n
+ N_A_27_74#_c_272_n N_A_27_74#_c_254_n N_A_27_74#_c_255_n N_A_27_74#_c_256_n
+ N_A_27_74#_c_257_n N_A_27_74#_c_438_p N_A_27_74#_c_258_n N_A_27_74#_c_318_p
+ N_A_27_74#_c_366_p N_A_27_74#_c_259_n N_A_27_74#_c_260_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_27_74#
x_PM_SKY130_FD_SC_MS__DFXBP_1%D N_D_M1021_g N_D_c_481_n N_D_c_482_n N_D_M1009_g
+ N_D_c_487_n N_D_c_488_n D D N_D_c_489_n N_D_c_484_n D
+ PM_SKY130_FD_SC_MS__DFXBP_1%D
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_208_368# N_A_208_368#_M1017_d
+ N_A_208_368#_M1014_d N_A_208_368#_c_543_n N_A_208_368#_c_544_n
+ N_A_208_368#_c_555_n N_A_208_368#_M1026_g N_A_208_368#_M1012_g
+ N_A_208_368#_M1010_g N_A_208_368#_M1016_g N_A_208_368#_c_558_n
+ N_A_208_368#_c_547_n N_A_208_368#_c_559_n N_A_208_368#_c_560_n
+ N_A_208_368#_c_660_p N_A_208_368#_c_561_n N_A_208_368#_c_562_n
+ N_A_208_368#_c_563_n N_A_208_368#_c_564_n N_A_208_368#_c_548_n
+ N_A_208_368#_c_549_n N_A_208_368#_c_567_n N_A_208_368#_c_653_n
+ N_A_208_368#_c_618_n N_A_208_368#_c_568_n N_A_208_368#_c_550_n
+ N_A_208_368#_c_551_n N_A_208_368#_c_571_n N_A_208_368#_c_552_n
+ N_A_208_368#_c_553_n N_A_208_368#_c_554_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_208_368#
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_701_463# N_A_701_463#_M1008_d
+ N_A_701_463#_M1011_d N_A_701_463#_c_778_n N_A_701_463#_M1019_g
+ N_A_701_463#_c_771_n N_A_701_463#_c_772_n N_A_701_463#_M1005_g
+ N_A_701_463#_c_780_n N_A_701_463#_c_773_n N_A_701_463#_c_774_n
+ N_A_701_463#_c_775_n N_A_701_463#_c_782_n N_A_701_463#_c_776_n
+ N_A_701_463#_c_783_n N_A_701_463#_c_777_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_701_463#
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_546_447# N_A_546_447#_M1002_d
+ N_A_546_447#_M1026_d N_A_546_447#_M1011_g N_A_546_447#_M1008_g
+ N_A_546_447#_c_861_n N_A_546_447#_c_868_n N_A_546_447#_c_862_n
+ N_A_546_447#_c_863_n N_A_546_447#_c_864_n N_A_546_447#_c_865_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_546_447#
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_1191_120# N_A_1191_120#_M1018_s
+ N_A_1191_120#_M1001_s N_A_1191_120#_c_948_n N_A_1191_120#_M1013_g
+ N_A_1191_120#_c_963_n N_A_1191_120#_M1004_g N_A_1191_120#_M1006_g
+ N_A_1191_120#_M1024_g N_A_1191_120#_c_950_n N_A_1191_120#_M1022_g
+ N_A_1191_120#_M1007_g N_A_1191_120#_c_952_n N_A_1191_120#_c_967_n
+ N_A_1191_120#_c_953_n N_A_1191_120#_c_954_n N_A_1191_120#_c_955_n
+ N_A_1191_120#_c_969_n N_A_1191_120#_c_956_n N_A_1191_120#_c_957_n
+ N_A_1191_120#_c_970_n N_A_1191_120#_c_958_n N_A_1191_120#_c_959_n
+ N_A_1191_120#_c_960_n N_A_1191_120#_c_961_n N_A_1191_120#_c_962_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_1191_120#
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_1005_120# N_A_1005_120#_M1010_d
+ N_A_1005_120#_M1023_d N_A_1005_120#_M1018_g N_A_1005_120#_c_1091_n
+ N_A_1005_120#_M1001_g N_A_1005_120#_c_1093_n N_A_1005_120#_c_1098_n
+ N_A_1005_120#_c_1099_n N_A_1005_120#_c_1094_n N_A_1005_120#_c_1095_n
+ N_A_1005_120#_c_1096_n PM_SKY130_FD_SC_MS__DFXBP_1%A_1005_120#
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_1644_112# N_A_1644_112#_M1022_s
+ N_A_1644_112#_M1007_s N_A_1644_112#_M1000_g N_A_1644_112#_M1027_g
+ N_A_1644_112#_c_1175_n N_A_1644_112#_c_1180_n N_A_1644_112#_c_1176_n
+ N_A_1644_112#_c_1177_n N_A_1644_112#_c_1178_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_1644_112#
x_PM_SKY130_FD_SC_MS__DFXBP_1%VPWR N_VPWR_M1015_d N_VPWR_M1021_s N_VPWR_M1019_d
+ N_VPWR_M1004_d N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_c_1227_n N_VPWR_c_1228_n
+ N_VPWR_c_1229_n N_VPWR_c_1230_n N_VPWR_c_1231_n N_VPWR_c_1232_n
+ N_VPWR_c_1233_n VPWR N_VPWR_c_1234_n N_VPWR_c_1235_n N_VPWR_c_1236_n
+ N_VPWR_c_1237_n N_VPWR_c_1238_n N_VPWR_c_1239_n N_VPWR_c_1226_n
+ N_VPWR_c_1241_n N_VPWR_c_1242_n N_VPWR_c_1243_n N_VPWR_c_1244_n
+ N_VPWR_c_1245_n PM_SKY130_FD_SC_MS__DFXBP_1%VPWR
x_PM_SKY130_FD_SC_MS__DFXBP_1%A_423_503# N_A_423_503#_M1009_d
+ N_A_423_503#_M1021_d N_A_423_503#_c_1346_n N_A_423_503#_c_1347_n
+ N_A_423_503#_c_1350_n N_A_423_503#_c_1348_n
+ PM_SKY130_FD_SC_MS__DFXBP_1%A_423_503#
x_PM_SKY130_FD_SC_MS__DFXBP_1%Q N_Q_M1006_d N_Q_M1024_d N_Q_c_1387_n
+ N_Q_c_1388_n N_Q_c_1390_n N_Q_c_1389_n Q Q PM_SKY130_FD_SC_MS__DFXBP_1%Q
x_PM_SKY130_FD_SC_MS__DFXBP_1%Q_N N_Q_N_M1027_d N_Q_N_M1000_d N_Q_N_c_1422_n
+ N_Q_N_c_1423_n Q_N Q_N Q_N Q_N N_Q_N_c_1424_n PM_SKY130_FD_SC_MS__DFXBP_1%Q_N
x_PM_SKY130_FD_SC_MS__DFXBP_1%VGND N_VGND_M1025_d N_VGND_M1009_s N_VGND_M1005_d
+ N_VGND_M1013_d N_VGND_M1018_d N_VGND_M1022_d N_VGND_c_1447_n N_VGND_c_1448_n
+ N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n N_VGND_c_1452_n
+ N_VGND_c_1453_n N_VGND_c_1454_n N_VGND_c_1455_n VGND N_VGND_c_1456_n
+ N_VGND_c_1457_n N_VGND_c_1458_n N_VGND_c_1459_n N_VGND_c_1460_n
+ N_VGND_c_1461_n N_VGND_c_1462_n N_VGND_c_1463_n N_VGND_c_1464_n
+ N_VGND_c_1465_n PM_SKY130_FD_SC_MS__DFXBP_1%VGND
cc_1 VNB N_CLK_M1015_g 0.00933516f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.4
cc_2 VNB N_CLK_c_208_n 0.0249846f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_3 VNB N_CLK_c_209_n 0.0170997f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.385
cc_4 VNB N_CLK_c_210_n 0.043127f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.385
cc_5 VNB N_A_27_74#_M1014_g 0.00671647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_74#_c_241_n 0.0200827f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.385
cc_7 VNB N_A_27_74#_M1002_g 0.0501254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_243_n 0.0162777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_M1020_g 0.0105944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_245_n 0.025869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_246_n 0.0170752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_247_n 0.0116924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_248_n 0.00166535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_249_n 0.00186241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_250_n 0.00540141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_251_n 0.00281369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_252_n 0.0221511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_253_n 0.00163039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_254_n 7.82432e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_255_n 0.0118083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_256_n 0.0105648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_257_n 0.0414841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_258_n 0.00259079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_259_n 0.00103934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_260_n 0.0392937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_D_c_481_n 0.017978f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_27 VNB N_D_c_482_n 0.016457f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_28 VNB D 0.00823049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_D_c_484_n 0.0330064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB D 0.0010259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_208_368#_c_543_n 0.124043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_208_368#_c_544_n 0.0124378f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.385
cc_33 VNB N_A_208_368#_M1012_g 0.0273053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_208_368#_M1010_g 0.0222798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_208_368#_c_547_n 0.00597788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_208_368#_c_548_n 0.00235398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_208_368#_c_549_n 0.0161929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_208_368#_c_550_n 0.0239766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_208_368#_c_551_n 0.0046762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_208_368#_c_552_n 0.00313964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_208_368#_c_553_n 0.0118286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_208_368#_c_554_n 0.0763825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_701_463#_c_771_n 0.0165524f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.385
cc_44 VNB N_A_701_463#_c_772_n 0.0176421f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.385
cc_45 VNB N_A_701_463#_c_773_n 0.00671037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_701_463#_c_774_n 0.00169046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_701_463#_c_775_n 0.00267832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_701_463#_c_776_n 0.00358633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_701_463#_c_777_n 0.0561054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_546_447#_M1008_g 0.0470947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_546_447#_c_861_n 0.00118604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_546_447#_c_862_n 0.00823929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_546_447#_c_863_n 0.00382818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_546_447#_c_864_n 0.00233106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_546_447#_c_865_n 0.00956301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1191_120#_c_948_n 0.0180835f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_57 VNB N_A_1191_120#_M1006_g 0.0308613f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_58 VNB N_A_1191_120#_c_950_n 0.0496885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1191_120#_M1022_g 0.028129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1191_120#_c_952_n 0.0263396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1191_120#_c_953_n 0.0109904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1191_120#_c_954_n 0.00994684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1191_120#_c_955_n 0.0041626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1191_120#_c_956_n 0.00194748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1191_120#_c_957_n 0.00430774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1191_120#_c_958_n 0.00589238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1191_120#_c_959_n 0.0134552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1191_120#_c_960_n 0.00424067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1191_120#_c_961_n 0.0163416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1191_120#_c_962_n 0.0039729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1005_120#_M1018_g 0.0344116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1005_120#_c_1091_n 0.0422748f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.385
cc_73 VNB N_A_1005_120#_M1001_g 0.00295455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1005_120#_c_1093_n 0.00478673f $X=-0.19 $Y=-0.245 $X2=0.5
+ $Y2=1.385
cc_75 VNB N_A_1005_120#_c_1094_n 0.00830518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1005_120#_c_1095_n 0.00210839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1005_120#_c_1096_n 0.0367433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1644_112#_M1000_g 0.00181363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1644_112#_M1027_g 0.0283734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1644_112#_c_1175_n 0.00163563f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.365
cc_81 VNB N_A_1644_112#_c_1176_n 0.00581718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1644_112#_c_1177_n 0.033278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1644_112#_c_1178_n 4.13327e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VPWR_c_1226_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_423_503#_c_1346_n 0.00580587f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_86 VNB N_A_423_503#_c_1347_n 0.00234657f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.385
cc_87 VNB N_A_423_503#_c_1348_n 0.00770442f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.365
cc_88 VNB N_Q_c_1387_n 0.0118205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_Q_c_1388_n 0.00607215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_Q_c_1389_n 0.00334031f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_91 VNB N_Q_N_c_1422_n 0.0268838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_Q_N_c_1423_n 0.0131134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_Q_N_c_1424_n 0.0249582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1447_n 0.00896842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1448_n 0.00500733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1449_n 0.0221779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1450_n 0.00980886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1451_n 0.0167052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1452_n 0.0446216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1453_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1454_n 0.0349259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1455_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1456_n 0.0187989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1457_n 0.0228203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1458_n 0.0409948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1459_n 0.0210192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1460_n 0.0195955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1461_n 0.523824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1462_n 0.00728126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1463_n 0.00463313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1464_n 0.0144866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1465_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VPB N_CLK_M1015_g 0.028083f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.4
cc_114 VPB N_A_27_74#_M1014_g 0.0259311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_74#_M1002_g 0.00462901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_74#_M1003_g 0.0435067f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.365
cc_117 VPB N_A_27_74#_c_264_n 0.0199887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_74#_c_243_n 0.0110118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_74#_c_266_n 0.0235385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_74#_c_267_n 0.0426033f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_74#_c_268_n 0.00416746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_27_74#_c_269_n 0.00966261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_27_74#_c_249_n 0.00100809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_27_74#_c_271_n 0.00475834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_27_74#_c_272_n 0.044779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_27_74#_c_255_n 0.00162615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_D_M1021_g 0.0277866f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.4
cc_128 VPB N_D_c_487_n 0.00490033f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.385
cc_129 VPB N_D_c_488_n 0.00296382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_D_c_489_n 0.0417709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_208_368#_c_555_n 0.0557223f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.385
cc_132 VPB N_A_208_368#_M1026_g 0.038237f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.385
cc_133 VPB N_A_208_368#_M1016_g 0.0393201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_208_368#_c_558_n 0.00749605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_208_368#_c_559_n 0.00752859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_208_368#_c_560_n 0.00907849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_208_368#_c_561_n 0.00423784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_208_368#_c_562_n 0.00491526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_208_368#_c_563_n 0.0094181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_208_368#_c_564_n 0.0097708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_208_368#_c_548_n 0.0194931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_208_368#_c_549_n 0.0162754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_208_368#_c_567_n 0.00829109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_208_368#_c_568_n 0.00110644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_208_368#_c_550_n 0.0148529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_208_368#_c_551_n 3.5904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_208_368#_c_571_n 8.00764e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_208_368#_c_552_n 5.59442e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_208_368#_c_553_n 0.0261169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_701_463#_c_778_n 0.0195677f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_151 VPB N_A_701_463#_c_771_n 0.0369573f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.385
cc_152 VPB N_A_701_463#_c_780_n 0.0179854f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_153 VPB N_A_701_463#_c_774_n 0.00214217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_701_463#_c_782_n 0.00214694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_701_463#_c_783_n 0.00918998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_546_447#_M1011_g 0.025681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_546_447#_c_861_n 0.00483153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_546_447#_c_868_n 0.0171655f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_159 VPB N_A_546_447#_c_864_n 0.0040038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_546_447#_c_865_n 0.0376501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_1191_120#_c_963_n 0.0180762f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.385
cc_162 VPB N_A_1191_120#_M1024_g 0.0271348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_1191_120#_c_950_n 0.0243168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_1191_120#_M1007_g 0.0231255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_1191_120#_c_967_n 0.0679897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_1191_120#_c_954_n 8.17895e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_1191_120#_c_969_n 0.00925603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1191_120#_c_970_n 0.00196713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_1191_120#_c_958_n 0.0141289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_1191_120#_c_959_n 0.00360691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_1191_120#_c_960_n 0.00208859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_1191_120#_c_961_n 0.0041169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_1005_120#_M1001_g 0.0237159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_1005_120#_c_1098_n 0.00401672f $X=-0.19 $Y=1.66 $X2=0.24
+ $Y2=1.365
cc_175 VPB N_A_1005_120#_c_1099_n 0.0012271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_1005_120#_c_1094_n 0.00333943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1644_112#_M1000_g 0.0298295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_1644_112#_c_1180_n 0.00534596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1227_n 0.0055443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1228_n 0.00962306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1229_n 0.0201407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1230_n 0.0131829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1231_n 0.01786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1232_n 0.0476377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1233_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1234_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1235_n 0.0200756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1236_n 0.047945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1237_n 0.0216197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1238_n 0.0330829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1239_n 0.0189562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1226_n 0.125205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1241_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1242_n 0.00631318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1243_n 0.0152284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1244_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1245_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_423_503#_c_1346_n 0.00315188f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_199 VPB N_A_423_503#_c_1350_n 0.00241878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_Q_c_1390_n 0.00229785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_Q_c_1389_n 0.00422386f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_202 VPB Q 0.0136179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB Q_N 0.0123377f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_204 VPB Q_N 0.0415558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_Q_N_c_1424_n 0.00766684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 N_CLK_M1015_g N_A_27_74#_M1014_g 0.0339293f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_207 N_CLK_c_208_n N_A_27_74#_c_241_n 0.0181404f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_208 N_CLK_M1015_g N_A_27_74#_c_267_n 0.00147311f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_209 N_CLK_c_208_n N_A_27_74#_c_246_n 0.00882722f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_210 N_CLK_M1015_g N_A_27_74#_c_268_n 0.0189754f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_211 N_CLK_c_209_n N_A_27_74#_c_268_n 0.0102401f $X=0.335 $Y=1.385 $X2=0 $Y2=0
cc_212 N_CLK_c_210_n N_A_27_74#_c_268_n 0.00111883f $X=0.5 $Y=1.385 $X2=0 $Y2=0
cc_213 N_CLK_c_209_n N_A_27_74#_c_269_n 0.0201635f $X=0.335 $Y=1.385 $X2=0 $Y2=0
cc_214 N_CLK_c_210_n N_A_27_74#_c_269_n 0.00442617f $X=0.5 $Y=1.385 $X2=0 $Y2=0
cc_215 N_CLK_c_208_n N_A_27_74#_c_283_n 0.0119752f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_216 N_CLK_c_209_n N_A_27_74#_c_283_n 0.00263778f $X=0.335 $Y=1.385 $X2=0
+ $Y2=0
cc_217 N_CLK_c_208_n N_A_27_74#_c_247_n 0.00476731f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_218 N_CLK_c_209_n N_A_27_74#_c_247_n 0.0252086f $X=0.335 $Y=1.385 $X2=0 $Y2=0
cc_219 N_CLK_c_210_n N_A_27_74#_c_247_n 0.00160701f $X=0.5 $Y=1.385 $X2=0 $Y2=0
cc_220 N_CLK_c_208_n N_A_27_74#_c_248_n 0.00646623f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_221 N_CLK_c_209_n N_A_27_74#_c_248_n 0.0300243f $X=0.335 $Y=1.385 $X2=0 $Y2=0
cc_222 N_CLK_c_210_n N_A_27_74#_c_248_n 0.00313275f $X=0.5 $Y=1.385 $X2=0 $Y2=0
cc_223 N_CLK_M1015_g N_A_27_74#_c_258_n 0.00313275f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_224 N_CLK_c_209_n N_A_27_74#_c_260_n 2.79433e-19 $X=0.335 $Y=1.385 $X2=0
+ $Y2=0
cc_225 N_CLK_c_210_n N_A_27_74#_c_260_n 0.0207929f $X=0.5 $Y=1.385 $X2=0 $Y2=0
cc_226 N_CLK_M1015_g N_A_208_368#_c_558_n 2.39284e-19 $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_227 N_CLK_M1015_g N_A_208_368#_c_548_n 4.66032e-19 $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_228 N_CLK_M1015_g N_VPWR_c_1227_n 0.0200267f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_229 N_CLK_M1015_g N_VPWR_c_1234_n 0.00460063f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_230 N_CLK_M1015_g N_VPWR_c_1226_n 0.00912278f $X=0.5 $Y=2.4 $X2=0 $Y2=0
cc_231 N_CLK_c_208_n N_VGND_c_1447_n 0.0047967f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_232 N_CLK_c_208_n N_VGND_c_1456_n 0.00329783f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_233 N_CLK_c_208_n N_VGND_c_1461_n 0.00427533f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_234 N_A_27_74#_c_250_n N_D_c_481_n 0.00278405f $X=2.375 $Y=0.815 $X2=0 $Y2=0
cc_235 N_A_27_74#_M1002_g N_D_c_482_n 0.0172805f $X=3.015 $Y=0.805 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_250_n N_D_c_482_n 0.00588103f $X=2.375 $Y=0.815 $X2=0 $Y2=0
cc_237 N_A_27_74#_c_251_n N_D_c_482_n 0.00772943f $X=2.46 $Y=0.73 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_252_n N_D_c_482_n 0.00155847f $X=3.485 $Y=0.34 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_250_n D 0.0230701f $X=2.375 $Y=0.815 $X2=0 $Y2=0
cc_240 N_A_27_74#_M1014_g N_D_c_489_n 0.00199396f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_27_74#_M1002_g N_D_c_484_n 0.00223115f $X=3.015 $Y=0.805 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_250_n N_D_c_484_n 0.00533187f $X=2.375 $Y=0.815 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_250_n N_A_208_368#_M1017_d 0.00985275f $X=2.375 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_244 N_A_27_74#_M1002_g N_A_208_368#_c_543_n 0.00882199f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_245 N_A_27_74#_c_250_n N_A_208_368#_c_543_n 0.00395094f $X=2.375 $Y=0.815
+ $X2=0 $Y2=0
cc_246 N_A_27_74#_c_252_n N_A_208_368#_c_543_n 0.0145743f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_247 N_A_27_74#_c_253_n N_A_208_368#_c_543_n 0.0035998f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_248 N_A_27_74#_c_241_n N_A_208_368#_c_544_n 0.0153188f $X=1.135 $Y=1.22 $X2=0
+ $Y2=0
cc_249 N_A_27_74#_M1002_g N_A_208_368#_c_555_n 0.0125777f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_250 N_A_27_74#_M1003_g N_A_208_368#_M1026_g 0.0167452f $X=3.175 $Y=2.75 $X2=0
+ $Y2=0
cc_251 N_A_27_74#_c_272_n N_A_208_368#_M1026_g 0.0125777f $X=3.285 $Y=1.91 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_M1002_g N_A_208_368#_M1012_g 0.00817548f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_253 N_A_27_74#_c_252_n N_A_208_368#_M1012_g 0.0121187f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_254 N_A_27_74#_c_271_n N_A_208_368#_M1012_g 0.001104f $X=3.485 $Y=1.912 $X2=0
+ $Y2=0
cc_255 N_A_27_74#_c_272_n N_A_208_368#_M1012_g 7.27492e-19 $X=3.285 $Y=1.91
+ $X2=0 $Y2=0
cc_256 N_A_27_74#_c_254_n N_A_208_368#_M1012_g 0.00486574f $X=3.57 $Y=0.58 $X2=0
+ $Y2=0
cc_257 N_A_27_74#_c_255_n N_A_208_368#_M1012_g 0.00754412f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_258 N_A_27_74#_c_318_p N_A_208_368#_M1012_g 0.00406164f $X=3.57 $Y=0.665
+ $X2=0 $Y2=0
cc_259 N_A_27_74#_M1020_g N_A_208_368#_M1010_g 0.0112129f $X=5.64 $Y=0.94 $X2=0
+ $Y2=0
cc_260 N_A_27_74#_c_245_n N_A_208_368#_M1010_g 0.00712048f $X=5.64 $Y=1.3 $X2=0
+ $Y2=0
cc_261 N_A_27_74#_c_256_n N_A_208_368#_M1010_g 0.0154839f $X=5.55 $Y=0.455 $X2=0
+ $Y2=0
cc_262 N_A_27_74#_c_257_n N_A_208_368#_M1010_g 0.00486667f $X=5.55 $Y=0.455
+ $X2=0 $Y2=0
cc_263 N_A_27_74#_c_259_n N_A_208_368#_M1010_g 0.00342658f $X=4.65 $Y=0.52 $X2=0
+ $Y2=0
cc_264 N_A_27_74#_c_264_n N_A_208_368#_M1016_g 0.0197714f $X=5.18 $Y=2.045 $X2=0
+ $Y2=0
cc_265 N_A_27_74#_c_266_n N_A_208_368#_M1016_g 0.0132532f $X=5.34 $Y=1.97 $X2=0
+ $Y2=0
cc_266 N_A_27_74#_M1014_g N_A_208_368#_c_558_n 0.00684487f $X=0.95 $Y=2.4 $X2=0
+ $Y2=0
cc_267 N_A_27_74#_c_241_n N_A_208_368#_c_547_n 0.00422251f $X=1.135 $Y=1.22
+ $X2=0 $Y2=0
cc_268 N_A_27_74#_c_248_n N_A_208_368#_c_547_n 0.0309136f $X=0.88 $Y=1.34 $X2=0
+ $Y2=0
cc_269 N_A_27_74#_c_250_n N_A_208_368#_c_547_n 0.0266632f $X=2.375 $Y=0.815
+ $X2=0 $Y2=0
cc_270 N_A_27_74#_M1003_g N_A_208_368#_c_560_n 0.00558041f $X=3.175 $Y=2.75
+ $X2=0 $Y2=0
cc_271 N_A_27_74#_c_264_n N_A_208_368#_c_562_n 0.0194793f $X=5.18 $Y=2.045 $X2=0
+ $Y2=0
cc_272 N_A_27_74#_c_243_n N_A_208_368#_c_562_n 0.00426363f $X=5.34 $Y=1.895
+ $X2=0 $Y2=0
cc_273 N_A_27_74#_c_266_n N_A_208_368#_c_562_n 0.00559867f $X=5.34 $Y=1.97 $X2=0
+ $Y2=0
cc_274 N_A_27_74#_c_264_n N_A_208_368#_c_563_n 0.011237f $X=5.18 $Y=2.045 $X2=0
+ $Y2=0
cc_275 N_A_27_74#_M1014_g N_A_208_368#_c_548_n 0.00739547f $X=0.95 $Y=2.4 $X2=0
+ $Y2=0
cc_276 N_A_27_74#_c_268_n N_A_208_368#_c_548_n 0.00863354f $X=0.67 $Y=1.805
+ $X2=0 $Y2=0
cc_277 N_A_27_74#_c_249_n N_A_208_368#_c_548_n 0.00730627f $X=0.755 $Y=1.72
+ $X2=0 $Y2=0
cc_278 N_A_27_74#_c_250_n N_A_208_368#_c_548_n 0.00394693f $X=2.375 $Y=0.815
+ $X2=0 $Y2=0
cc_279 N_A_27_74#_c_258_n N_A_208_368#_c_548_n 0.0102005f $X=0.965 $Y=1.385
+ $X2=0 $Y2=0
cc_280 N_A_27_74#_c_260_n N_A_208_368#_c_548_n 0.00621043f $X=1.135 $Y=1.385
+ $X2=0 $Y2=0
cc_281 N_A_27_74#_M1014_g N_A_208_368#_c_549_n 0.00600128f $X=0.95 $Y=2.4 $X2=0
+ $Y2=0
cc_282 N_A_27_74#_c_250_n N_A_208_368#_c_549_n 6.67411e-19 $X=2.375 $Y=0.815
+ $X2=0 $Y2=0
cc_283 N_A_27_74#_c_260_n N_A_208_368#_c_549_n 0.00308767f $X=1.135 $Y=1.385
+ $X2=0 $Y2=0
cc_284 N_A_27_74#_M1014_g N_A_208_368#_c_567_n 0.0064732f $X=0.95 $Y=2.4 $X2=0
+ $Y2=0
cc_285 N_A_27_74#_M1003_g N_A_208_368#_c_618_n 0.0113296f $X=3.175 $Y=2.75 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_264_n N_A_208_368#_c_568_n 3.32479e-19 $X=5.18 $Y=2.045
+ $X2=0 $Y2=0
cc_287 N_A_27_74#_c_245_n N_A_208_368#_c_550_n 0.0194671f $X=5.64 $Y=1.3 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_c_266_n N_A_208_368#_c_551_n 2.48944e-19 $X=5.34 $Y=1.97 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_245_n N_A_208_368#_c_551_n 0.00191018f $X=5.64 $Y=1.3 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_c_264_n N_A_208_368#_c_571_n 0.00890066f $X=5.18 $Y=2.045
+ $X2=0 $Y2=0
cc_291 N_A_27_74#_c_243_n N_A_208_368#_c_552_n 3.37545e-19 $X=5.34 $Y=1.895
+ $X2=0 $Y2=0
cc_292 N_A_27_74#_c_243_n N_A_208_368#_c_553_n 0.0132532f $X=5.34 $Y=1.895 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_245_n N_A_208_368#_c_553_n 0.00503848f $X=5.64 $Y=1.3 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_c_248_n N_A_208_368#_c_554_n 8.50708e-19 $X=0.88 $Y=1.34 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_250_n N_A_208_368#_c_554_n 0.0174916f $X=2.375 $Y=0.815
+ $X2=0 $Y2=0
cc_296 N_A_27_74#_c_251_n N_A_208_368#_c_554_n 0.00268474f $X=2.46 $Y=0.73 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_260_n N_A_208_368#_c_554_n 0.0153188f $X=1.135 $Y=1.385
+ $X2=0 $Y2=0
cc_298 N_A_27_74#_c_256_n N_A_701_463#_M1008_d 0.00236045f $X=5.55 $Y=0.455
+ $X2=-0.19 $Y2=-0.245
cc_299 N_A_27_74#_c_259_n N_A_701_463#_M1008_d 0.00269557f $X=4.65 $Y=0.52
+ $X2=-0.19 $Y2=-0.245
cc_300 N_A_27_74#_M1003_g N_A_701_463#_c_771_n 0.00836419f $X=3.175 $Y=2.75
+ $X2=0 $Y2=0
cc_301 N_A_27_74#_c_271_n N_A_701_463#_c_771_n 0.00373919f $X=3.485 $Y=1.912
+ $X2=0 $Y2=0
cc_302 N_A_27_74#_c_272_n N_A_701_463#_c_771_n 0.0193084f $X=3.285 $Y=1.91 $X2=0
+ $Y2=0
cc_303 N_A_27_74#_c_252_n N_A_701_463#_c_772_n 6.92565e-19 $X=3.485 $Y=0.34
+ $X2=0 $Y2=0
cc_304 N_A_27_74#_c_254_n N_A_701_463#_c_772_n 0.00324162f $X=3.57 $Y=0.58 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_c_255_n N_A_701_463#_c_772_n 0.00835903f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_366_p N_A_701_463#_c_772_n 0.0131394f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_307 N_A_27_74#_c_259_n N_A_701_463#_c_772_n 7.80335e-19 $X=4.65 $Y=0.52 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_M1003_g N_A_701_463#_c_780_n 0.0428964f $X=3.175 $Y=2.75 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_271_n N_A_701_463#_c_780_n 9.77065e-19 $X=3.485 $Y=1.912
+ $X2=0 $Y2=0
cc_310 N_A_27_74#_c_255_n N_A_701_463#_c_773_n 0.0281658f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_366_p N_A_701_463#_c_773_n 0.0314351f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_c_243_n N_A_701_463#_c_774_n 3.19973e-19 $X=5.34 $Y=1.895
+ $X2=0 $Y2=0
cc_313 N_A_27_74#_c_256_n N_A_701_463#_c_775_n 0.0098544f $X=5.55 $Y=0.455 $X2=0
+ $Y2=0
cc_314 N_A_27_74#_c_259_n N_A_701_463#_c_775_n 0.0023898f $X=4.65 $Y=0.52 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_c_266_n N_A_701_463#_c_782_n 0.00175862f $X=5.34 $Y=1.97 $X2=0
+ $Y2=0
cc_316 N_A_27_74#_c_366_p N_A_701_463#_c_776_n 0.00546209f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_317 N_A_27_74#_c_259_n N_A_701_463#_c_776_n 0.00418601f $X=4.65 $Y=0.52 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_266_n N_A_701_463#_c_783_n 4.25482e-19 $X=5.34 $Y=1.97 $X2=0
+ $Y2=0
cc_319 N_A_27_74#_M1002_g N_A_701_463#_c_777_n 0.00849305f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_320 N_A_27_74#_c_255_n N_A_701_463#_c_777_n 0.0108304f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_366_p N_A_701_463#_c_777_n 0.00387233f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_c_264_n N_A_546_447#_M1011_g 0.00852739f $X=5.18 $Y=2.045
+ $X2=0 $Y2=0
cc_323 N_A_27_74#_c_366_p N_A_546_447#_M1008_g 0.00873882f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_324 N_A_27_74#_c_259_n N_A_546_447#_M1008_g 0.0142929f $X=4.65 $Y=0.52 $X2=0
+ $Y2=0
cc_325 N_A_27_74#_M1002_g N_A_546_447#_c_861_n 0.00503943f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_326 N_A_27_74#_M1003_g N_A_546_447#_c_861_n 0.00676836f $X=3.175 $Y=2.75
+ $X2=0 $Y2=0
cc_327 N_A_27_74#_c_271_n N_A_546_447#_c_861_n 0.024117f $X=3.485 $Y=1.912 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_272_n N_A_546_447#_c_861_n 0.00693674f $X=3.285 $Y=1.91
+ $X2=0 $Y2=0
cc_329 N_A_27_74#_c_255_n N_A_546_447#_c_861_n 0.00510602f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_M1003_g N_A_546_447#_c_868_n 0.012462f $X=3.175 $Y=2.75 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_271_n N_A_546_447#_c_868_n 0.0412232f $X=3.485 $Y=1.912
+ $X2=0 $Y2=0
cc_332 N_A_27_74#_c_272_n N_A_546_447#_c_868_n 0.00835874f $X=3.285 $Y=1.91
+ $X2=0 $Y2=0
cc_333 N_A_27_74#_M1002_g N_A_546_447#_c_862_n 0.0168077f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_334 N_A_27_74#_c_271_n N_A_546_447#_c_862_n 0.0146384f $X=3.485 $Y=1.912
+ $X2=0 $Y2=0
cc_335 N_A_27_74#_c_272_n N_A_546_447#_c_862_n 0.00591527f $X=3.285 $Y=1.91
+ $X2=0 $Y2=0
cc_336 N_A_27_74#_c_255_n N_A_546_447#_c_862_n 0.0139107f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_M1002_g N_A_546_447#_c_863_n 0.0161485f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_338 N_A_27_74#_c_252_n N_A_546_447#_c_863_n 0.0168505f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_255_n N_A_546_447#_c_863_n 0.0496115f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_318_p N_A_546_447#_c_863_n 0.0125189f $X=3.57 $Y=0.665 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_c_271_n N_A_546_447#_c_864_n 0.0154088f $X=3.485 $Y=1.912
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_c_255_n N_A_546_447#_c_864_n 0.00497917f $X=3.57 $Y=1.75 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_266_n N_A_546_447#_c_865_n 0.00852739f $X=5.34 $Y=1.97 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_257_n N_A_1191_120#_c_948_n 0.0201557f $X=5.55 $Y=0.455
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_M1020_g N_A_1191_120#_c_952_n 0.0201557f $X=5.64 $Y=0.94 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_256_n N_A_1005_120#_M1010_d 0.00339582f $X=5.55 $Y=0.455
+ $X2=-0.19 $Y2=-0.245
cc_347 N_A_27_74#_M1020_g N_A_1005_120#_c_1093_n 0.0146893f $X=5.64 $Y=0.94
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_245_n N_A_1005_120#_c_1093_n 0.0163607f $X=5.64 $Y=1.3 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_256_n N_A_1005_120#_c_1093_n 0.0346574f $X=5.55 $Y=0.455
+ $X2=0 $Y2=0
cc_350 N_A_27_74#_c_257_n N_A_1005_120#_c_1093_n 0.0017534f $X=5.55 $Y=0.455
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_c_264_n N_A_1005_120#_c_1094_n 0.00186114f $X=5.18 $Y=2.045
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_243_n N_A_1005_120#_c_1094_n 0.0123471f $X=5.34 $Y=1.895
+ $X2=0 $Y2=0
cc_353 N_A_27_74#_c_266_n N_A_1005_120#_c_1094_n 0.00613711f $X=5.34 $Y=1.97
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_M1020_g N_A_1005_120#_c_1096_n 0.00363885f $X=5.64 $Y=0.94
+ $X2=0 $Y2=0
cc_355 N_A_27_74#_c_245_n N_A_1005_120#_c_1096_n 0.00395369f $X=5.64 $Y=1.3
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_256_n N_A_1005_120#_c_1096_n 0.00318241f $X=5.55 $Y=0.455
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_268_n N_VPWR_M1015_d 0.001797f $X=0.67 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_358 N_A_27_74#_M1014_g N_VPWR_c_1227_n 0.0038373f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_267_n N_VPWR_c_1227_n 0.0297232f $X=0.275 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_268_n N_VPWR_c_1227_n 0.0159932f $X=0.67 $Y=1.805 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_M1014_g N_VPWR_c_1228_n 0.00304911f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_264_n N_VPWR_c_1232_n 0.00333867f $X=5.18 $Y=2.045 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_267_n N_VPWR_c_1234_n 0.011066f $X=0.275 $Y=1.985 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_M1014_g N_VPWR_c_1235_n 0.00519767f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_365 N_A_27_74#_M1003_g N_VPWR_c_1236_n 0.00365788f $X=3.175 $Y=2.75 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_M1014_g N_VPWR_c_1226_n 0.00983841f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_367 N_A_27_74#_M1003_g N_VPWR_c_1226_n 0.00449588f $X=3.175 $Y=2.75 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_264_n N_VPWR_c_1226_n 0.0043016f $X=5.18 $Y=2.045 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_267_n N_VPWR_c_1226_n 0.00915947f $X=0.275 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_M1002_g N_A_423_503#_c_1346_n 0.00273248f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_371 N_A_27_74#_M1002_g N_A_423_503#_c_1347_n 5.15818e-19 $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_c_252_n N_A_423_503#_c_1347_n 0.0125903f $X=3.485 $Y=0.34
+ $X2=0 $Y2=0
cc_373 N_A_27_74#_M1002_g N_A_423_503#_c_1348_n 0.0013209f $X=3.015 $Y=0.805
+ $X2=0 $Y2=0
cc_374 N_A_27_74#_c_250_n N_A_423_503#_c_1348_n 0.00580393f $X=2.375 $Y=0.815
+ $X2=0 $Y2=0
cc_375 N_A_27_74#_c_252_n N_A_423_503#_c_1348_n 0.00463789f $X=3.485 $Y=0.34
+ $X2=0 $Y2=0
cc_376 N_A_27_74#_c_283_n N_VGND_M1025_d 0.00203816f $X=0.67 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_377 N_A_27_74#_c_248_n N_VGND_M1025_d 0.00306381f $X=0.88 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_378 N_A_27_74#_c_438_p N_VGND_M1025_d 0.00481862f $X=0.88 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_379 N_A_27_74#_c_250_n N_VGND_M1009_s 0.0162449f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_c_251_n N_VGND_M1009_s 0.00220092f $X=2.46 $Y=0.73 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_366_p N_VGND_M1005_d 0.00784253f $X=4.48 $Y=0.52 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_241_n N_VGND_c_1447_n 0.00517914f $X=1.135 $Y=1.22 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_c_246_n N_VGND_c_1447_n 0.00830227f $X=0.28 $Y=0.73 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_283_n N_VGND_c_1447_n 0.00333414f $X=0.67 $Y=0.815 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_438_p N_VGND_c_1447_n 0.0288149f $X=0.88 $Y=0.815 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_c_260_n N_VGND_c_1447_n 6.03453e-19 $X=1.135 $Y=1.385 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_241_n N_VGND_c_1448_n 0.0018585f $X=1.135 $Y=1.22 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_c_250_n N_VGND_c_1448_n 0.0273135f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_389 N_A_27_74#_c_251_n N_VGND_c_1448_n 0.010507f $X=2.46 $Y=0.73 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_253_n N_VGND_c_1448_n 0.0149551f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_256_n N_VGND_c_1449_n 0.0154427f $X=5.55 $Y=0.455 $X2=0
+ $Y2=0
cc_392 N_A_27_74#_c_257_n N_VGND_c_1449_n 0.00357245f $X=5.55 $Y=0.455 $X2=0
+ $Y2=0
cc_393 N_A_27_74#_c_257_n N_VGND_c_1452_n 0.00761354f $X=5.55 $Y=0.455 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_c_366_p N_VGND_c_1452_n 0.00275846f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_259_n N_VGND_c_1452_n 0.0674522f $X=4.65 $Y=0.52 $X2=0 $Y2=0
cc_396 N_A_27_74#_c_246_n N_VGND_c_1456_n 0.0145323f $X=0.28 $Y=0.73 $X2=0 $Y2=0
cc_397 N_A_27_74#_c_283_n N_VGND_c_1456_n 0.00206038f $X=0.67 $Y=0.815 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_241_n N_VGND_c_1457_n 0.00336057f $X=1.135 $Y=1.22 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_250_n N_VGND_c_1457_n 0.0103557f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_438_p N_VGND_c_1457_n 8.51599e-19 $X=0.88 $Y=0.815 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_250_n N_VGND_c_1458_n 0.00241577f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_c_252_n N_VGND_c_1458_n 0.0721828f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_403 N_A_27_74#_c_253_n N_VGND_c_1458_n 0.0115448f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_404 N_A_27_74#_c_366_p N_VGND_c_1458_n 0.00530279f $X=4.48 $Y=0.52 $X2=0
+ $Y2=0
cc_405 N_A_27_74#_c_241_n N_VGND_c_1461_n 0.00439178f $X=1.135 $Y=1.22 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_246_n N_VGND_c_1461_n 0.0119861f $X=0.28 $Y=0.73 $X2=0 $Y2=0
cc_407 N_A_27_74#_c_283_n N_VGND_c_1461_n 0.00435273f $X=0.67 $Y=0.815 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_250_n N_VGND_c_1461_n 0.0239621f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_252_n N_VGND_c_1461_n 0.0377627f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_410 N_A_27_74#_c_253_n N_VGND_c_1461_n 0.00582224f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_411 N_A_27_74#_c_257_n N_VGND_c_1461_n 0.0109372f $X=5.55 $Y=0.455 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_c_438_p N_VGND_c_1461_n 0.00373489f $X=0.88 $Y=0.815 $X2=0
+ $Y2=0
cc_413 N_A_27_74#_c_366_p N_VGND_c_1461_n 0.0161936f $X=4.48 $Y=0.52 $X2=0 $Y2=0
cc_414 N_A_27_74#_c_259_n N_VGND_c_1461_n 0.0460173f $X=4.65 $Y=0.52 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_252_n N_VGND_c_1464_n 0.00873071f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_366_p N_VGND_c_1464_n 0.0244722f $X=4.48 $Y=0.52 $X2=0 $Y2=0
cc_417 N_A_27_74#_c_259_n N_VGND_c_1464_n 0.00868941f $X=4.65 $Y=0.52 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_254_n A_713_102# 7.77095e-19 $X=3.57 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_419 N_A_27_74#_c_255_n A_713_102# 0.00201594f $X=3.57 $Y=1.75 $X2=-0.19
+ $Y2=-0.245
cc_420 N_A_27_74#_c_366_p A_713_102# 0.0019187f $X=4.48 $Y=0.52 $X2=-0.19
+ $Y2=-0.245
cc_421 N_D_c_482_n N_A_208_368#_c_543_n 0.00903828f $X=2.585 $Y=1.125 $X2=0
+ $Y2=0
cc_422 N_D_c_481_n N_A_208_368#_c_555_n 0.0106711f $X=2.51 $Y=1.2 $X2=0 $Y2=0
cc_423 N_D_c_487_n N_A_208_368#_c_555_n 0.0032081f $X=1.995 $Y=2.025 $X2=0 $Y2=0
cc_424 N_D_c_484_n N_A_208_368#_c_555_n 0.0215245f $X=2.175 $Y=1.2 $X2=0 $Y2=0
cc_425 D N_A_208_368#_c_555_n 0.0181861f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_426 N_D_c_487_n N_A_208_368#_M1026_g 0.00103492f $X=1.995 $Y=2.025 $X2=0
+ $Y2=0
cc_427 N_D_c_488_n N_A_208_368#_M1026_g 2.67599e-19 $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_428 N_D_c_489_n N_A_208_368#_M1026_g 0.0188031f $X=2.025 $Y=2.19 $X2=0 $Y2=0
cc_429 N_D_M1021_g N_A_208_368#_c_558_n 0.00521764f $X=2.025 $Y=2.725 $X2=0
+ $Y2=0
cc_430 N_D_c_488_n N_A_208_368#_c_558_n 0.0192035f $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_431 N_D_c_489_n N_A_208_368#_c_558_n 0.00155202f $X=2.025 $Y=2.19 $X2=0 $Y2=0
cc_432 D N_A_208_368#_c_547_n 0.0196003f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_433 N_D_M1021_g N_A_208_368#_c_559_n 0.0106831f $X=2.025 $Y=2.725 $X2=0 $Y2=0
cc_434 N_D_c_488_n N_A_208_368#_c_559_n 0.0218569f $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_435 N_D_c_489_n N_A_208_368#_c_559_n 0.00506764f $X=2.025 $Y=2.19 $X2=0 $Y2=0
cc_436 N_D_M1021_g N_A_208_368#_c_560_n 7.62366e-19 $X=2.025 $Y=2.725 $X2=0
+ $Y2=0
cc_437 N_D_c_487_n N_A_208_368#_c_548_n 0.00836603f $X=1.995 $Y=2.025 $X2=0
+ $Y2=0
cc_438 N_D_c_488_n N_A_208_368#_c_548_n 0.00254579f $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_439 D N_A_208_368#_c_548_n 0.0262945f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_440 N_D_c_488_n N_A_208_368#_c_549_n 0.00124908f $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_441 N_D_c_489_n N_A_208_368#_c_549_n 0.02725f $X=2.025 $Y=2.19 $X2=0 $Y2=0
cc_442 N_D_M1021_g N_A_208_368#_c_567_n 0.00428146f $X=2.025 $Y=2.725 $X2=0
+ $Y2=0
cc_443 N_D_M1021_g N_A_208_368#_c_653_n 0.0155602f $X=2.025 $Y=2.725 $X2=0 $Y2=0
cc_444 N_D_c_488_n N_A_208_368#_c_653_n 0.00162457f $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_445 N_D_c_482_n N_A_208_368#_c_554_n 0.00840593f $X=2.585 $Y=1.125 $X2=0
+ $Y2=0
cc_446 D N_A_208_368#_c_554_n 0.00552936f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_447 N_D_c_484_n N_A_208_368#_c_554_n 0.0194048f $X=2.175 $Y=1.2 $X2=0 $Y2=0
cc_448 N_D_c_482_n N_A_546_447#_c_863_n 2.71831e-19 $X=2.585 $Y=1.125 $X2=0
+ $Y2=0
cc_449 N_D_M1021_g N_VPWR_c_1228_n 0.0065843f $X=2.025 $Y=2.725 $X2=0 $Y2=0
cc_450 N_D_M1021_g N_VPWR_c_1236_n 0.0050563f $X=2.025 $Y=2.725 $X2=0 $Y2=0
cc_451 N_D_M1021_g N_VPWR_c_1226_n 0.00645424f $X=2.025 $Y=2.725 $X2=0 $Y2=0
cc_452 N_D_c_481_n N_A_423_503#_c_1346_n 0.00450778f $X=2.51 $Y=1.2 $X2=0 $Y2=0
cc_453 N_D_c_487_n N_A_423_503#_c_1346_n 0.0106927f $X=1.995 $Y=2.025 $X2=0
+ $Y2=0
cc_454 N_D_c_488_n N_A_423_503#_c_1346_n 8.26298e-19 $X=1.995 $Y=2.19 $X2=0
+ $Y2=0
cc_455 D N_A_423_503#_c_1346_n 0.0411284f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_456 N_D_c_484_n N_A_423_503#_c_1346_n 0.00201648f $X=2.175 $Y=1.2 $X2=0 $Y2=0
cc_457 N_D_c_482_n N_A_423_503#_c_1347_n 0.0014192f $X=2.585 $Y=1.125 $X2=0
+ $Y2=0
cc_458 N_D_c_488_n N_A_423_503#_c_1350_n 0.024595f $X=1.995 $Y=2.19 $X2=0 $Y2=0
cc_459 N_D_c_489_n N_A_423_503#_c_1350_n 0.00342678f $X=2.025 $Y=2.19 $X2=0
+ $Y2=0
cc_460 D N_A_423_503#_c_1350_n 0.00113915f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_461 N_D_c_481_n N_A_423_503#_c_1348_n 0.00726186f $X=2.51 $Y=1.2 $X2=0 $Y2=0
cc_462 N_D_c_482_n N_A_423_503#_c_1348_n 0.00535172f $X=2.585 $Y=1.125 $X2=0
+ $Y2=0
cc_463 D N_A_423_503#_c_1348_n 0.00885757f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_464 N_D_c_482_n N_VGND_c_1448_n 3.16215e-19 $X=2.585 $Y=1.125 $X2=0 $Y2=0
cc_465 N_A_208_368#_c_561_n N_A_701_463#_M1011_d 0.0134358f $X=4.98 $Y=2.937
+ $X2=0 $Y2=0
cc_466 N_A_208_368#_c_562_n N_A_701_463#_M1011_d 0.00721113f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_467 N_A_208_368#_c_660_p N_A_701_463#_c_778_n 0.0134446f $X=4.3 $Y=2.67 $X2=0
+ $Y2=0
cc_468 N_A_208_368#_c_568_n N_A_701_463#_c_778_n 6.81363e-19 $X=4.385 $Y=2.67
+ $X2=0 $Y2=0
cc_469 N_A_208_368#_M1012_g N_A_701_463#_c_772_n 0.0408298f $X=3.49 $Y=0.72
+ $X2=0 $Y2=0
cc_470 N_A_208_368#_c_660_p N_A_701_463#_c_780_n 0.00335426f $X=4.3 $Y=2.67
+ $X2=0 $Y2=0
cc_471 N_A_208_368#_c_562_n N_A_701_463#_c_774_n 0.0076192f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_472 N_A_208_368#_c_550_n N_A_701_463#_c_774_n 0.0019033f $X=4.89 $Y=1.52
+ $X2=0 $Y2=0
cc_473 N_A_208_368#_c_551_n N_A_701_463#_c_774_n 0.0238337f $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_474 N_A_208_368#_M1010_g N_A_701_463#_c_775_n 0.00467243f $X=4.95 $Y=0.875
+ $X2=0 $Y2=0
cc_475 N_A_208_368#_c_550_n N_A_701_463#_c_775_n 0.00375305f $X=4.89 $Y=1.52
+ $X2=0 $Y2=0
cc_476 N_A_208_368#_c_551_n N_A_701_463#_c_775_n 0.00845643f $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_477 N_A_208_368#_c_561_n N_A_701_463#_c_782_n 0.0124498f $X=4.98 $Y=2.937
+ $X2=0 $Y2=0
cc_478 N_A_208_368#_c_562_n N_A_701_463#_c_782_n 0.0431061f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_479 N_A_208_368#_c_568_n N_A_701_463#_c_782_n 0.00210614f $X=4.385 $Y=2.67
+ $X2=0 $Y2=0
cc_480 N_A_208_368#_M1010_g N_A_701_463#_c_776_n 0.00435507f $X=4.95 $Y=0.875
+ $X2=0 $Y2=0
cc_481 N_A_208_368#_c_551_n N_A_701_463#_c_776_n 0.00119339f $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_482 N_A_208_368#_c_562_n N_A_701_463#_c_783_n 0.0134734f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_483 N_A_208_368#_c_568_n N_A_701_463#_c_783_n 5.26843e-19 $X=4.385 $Y=2.67
+ $X2=0 $Y2=0
cc_484 N_A_208_368#_c_550_n N_A_701_463#_c_783_n 0.00222583f $X=4.89 $Y=1.52
+ $X2=0 $Y2=0
cc_485 N_A_208_368#_c_551_n N_A_701_463#_c_783_n 0.00150313f $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_486 N_A_208_368#_c_560_n N_A_546_447#_M1026_d 0.00477186f $X=3.12 $Y=2.8
+ $X2=0 $Y2=0
cc_487 N_A_208_368#_c_561_n N_A_546_447#_M1011_g 0.00952701f $X=4.98 $Y=2.937
+ $X2=0 $Y2=0
cc_488 N_A_208_368#_c_562_n N_A_546_447#_M1011_g 0.00209938f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_489 N_A_208_368#_c_568_n N_A_546_447#_M1011_g 0.0216934f $X=4.385 $Y=2.67
+ $X2=0 $Y2=0
cc_490 N_A_208_368#_M1010_g N_A_546_447#_M1008_g 0.0221373f $X=4.95 $Y=0.875
+ $X2=0 $Y2=0
cc_491 N_A_208_368#_c_550_n N_A_546_447#_M1008_g 0.0203555f $X=4.89 $Y=1.52
+ $X2=0 $Y2=0
cc_492 N_A_208_368#_c_551_n N_A_546_447#_M1008_g 3.04229e-19 $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_493 N_A_208_368#_c_555_n N_A_546_447#_c_861_n 0.00407561f $X=2.55 $Y=1.74
+ $X2=0 $Y2=0
cc_494 N_A_208_368#_c_560_n N_A_546_447#_c_861_n 0.0131062f $X=3.12 $Y=2.8 $X2=0
+ $Y2=0
cc_495 N_A_208_368#_c_560_n N_A_546_447#_c_868_n 0.00668787f $X=3.12 $Y=2.8
+ $X2=0 $Y2=0
cc_496 N_A_208_368#_c_660_p N_A_546_447#_c_868_n 0.0681779f $X=4.3 $Y=2.67 $X2=0
+ $Y2=0
cc_497 N_A_208_368#_c_618_n N_A_546_447#_c_868_n 0.0111664f $X=3.205 $Y=2.67
+ $X2=0 $Y2=0
cc_498 N_A_208_368#_M1012_g N_A_546_447#_c_863_n 0.00185158f $X=3.49 $Y=0.72
+ $X2=0 $Y2=0
cc_499 N_A_208_368#_c_660_p N_A_546_447#_c_865_n 7.25328e-19 $X=4.3 $Y=2.67
+ $X2=0 $Y2=0
cc_500 N_A_208_368#_c_562_n N_A_546_447#_c_865_n 0.00123418f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_501 N_A_208_368#_c_563_n N_A_1191_120#_c_963_n 4.31611e-19 $X=5.82 $Y=2.99
+ $X2=0 $Y2=0
cc_502 N_A_208_368#_c_553_n N_A_1191_120#_c_952_n 0.00193829f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_503 N_A_208_368#_M1016_g N_A_1191_120#_c_967_n 0.0456348f $X=5.715 $Y=2.62
+ $X2=0 $Y2=0
cc_504 N_A_208_368#_c_564_n N_A_1191_120#_c_967_n 0.00717678f $X=5.905 $Y=2.905
+ $X2=0 $Y2=0
cc_505 N_A_208_368#_c_552_n N_A_1191_120#_c_958_n 0.0365678f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_506 N_A_208_368#_c_553_n N_A_1191_120#_c_958_n 0.00123628f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_507 N_A_208_368#_c_552_n N_A_1191_120#_c_959_n 4.21404e-19 $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_508 N_A_208_368#_c_553_n N_A_1191_120#_c_959_n 0.0177172f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_509 N_A_208_368#_c_563_n N_A_1005_120#_M1023_d 0.00205163f $X=5.82 $Y=2.99
+ $X2=0 $Y2=0
cc_510 N_A_208_368#_M1010_g N_A_1005_120#_c_1093_n 0.00837475f $X=4.95 $Y=0.875
+ $X2=0 $Y2=0
cc_511 N_A_208_368#_c_551_n N_A_1005_120#_c_1093_n 0.00362024f $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_512 N_A_208_368#_M1016_g N_A_1005_120#_c_1098_n 0.00460089f $X=5.715 $Y=2.62
+ $X2=0 $Y2=0
cc_513 N_A_208_368#_c_564_n N_A_1005_120#_c_1098_n 0.0173714f $X=5.905 $Y=2.905
+ $X2=0 $Y2=0
cc_514 N_A_208_368#_c_563_n N_A_1005_120#_c_1099_n 0.0184029f $X=5.82 $Y=2.99
+ $X2=0 $Y2=0
cc_515 N_A_208_368#_c_562_n N_A_1005_120#_c_1094_n 0.0512581f $X=5.065 $Y=2.8
+ $X2=0 $Y2=0
cc_516 N_A_208_368#_c_564_n N_A_1005_120#_c_1094_n 0.0080153f $X=5.905 $Y=2.905
+ $X2=0 $Y2=0
cc_517 N_A_208_368#_c_550_n N_A_1005_120#_c_1094_n 2.89229e-19 $X=4.89 $Y=1.52
+ $X2=0 $Y2=0
cc_518 N_A_208_368#_c_551_n N_A_1005_120#_c_1094_n 0.0231992f $X=5.065 $Y=1.52
+ $X2=0 $Y2=0
cc_519 N_A_208_368#_c_552_n N_A_1005_120#_c_1094_n 0.0248005f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_520 N_A_208_368#_c_553_n N_A_1005_120#_c_1094_n 0.00321912f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_521 N_A_208_368#_c_552_n N_A_1005_120#_c_1096_n 0.0199888f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_522 N_A_208_368#_c_553_n N_A_1005_120#_c_1096_n 0.00257163f $X=5.825 $Y=1.78
+ $X2=0 $Y2=0
cc_523 N_A_208_368#_c_559_n N_VPWR_M1021_s 0.0108037f $X=2.055 $Y=2.63 $X2=0
+ $Y2=0
cc_524 N_A_208_368#_c_660_p N_VPWR_M1019_d 0.0142515f $X=4.3 $Y=2.67 $X2=0 $Y2=0
cc_525 N_A_208_368#_c_567_n N_VPWR_c_1227_n 0.015735f $X=1.222 $Y=2.63 $X2=0
+ $Y2=0
cc_526 N_A_208_368#_c_559_n N_VPWR_c_1228_n 0.0244584f $X=2.055 $Y=2.63 $X2=0
+ $Y2=0
cc_527 N_A_208_368#_c_567_n N_VPWR_c_1228_n 0.00673603f $X=1.222 $Y=2.63 $X2=0
+ $Y2=0
cc_528 N_A_208_368#_M1016_g N_VPWR_c_1229_n 2.10745e-19 $X=5.715 $Y=2.62 $X2=0
+ $Y2=0
cc_529 N_A_208_368#_c_563_n N_VPWR_c_1229_n 0.0145031f $X=5.82 $Y=2.99 $X2=0
+ $Y2=0
cc_530 N_A_208_368#_c_564_n N_VPWR_c_1229_n 0.0222708f $X=5.905 $Y=2.905 $X2=0
+ $Y2=0
cc_531 N_A_208_368#_M1016_g N_VPWR_c_1232_n 8.50192e-19 $X=5.715 $Y=2.62 $X2=0
+ $Y2=0
cc_532 N_A_208_368#_c_660_p N_VPWR_c_1232_n 0.00321874f $X=4.3 $Y=2.67 $X2=0
+ $Y2=0
cc_533 N_A_208_368#_c_561_n N_VPWR_c_1232_n 0.0338079f $X=4.98 $Y=2.937 $X2=0
+ $Y2=0
cc_534 N_A_208_368#_c_563_n N_VPWR_c_1232_n 0.0549423f $X=5.82 $Y=2.99 $X2=0
+ $Y2=0
cc_535 N_A_208_368#_c_568_n N_VPWR_c_1232_n 0.0113002f $X=4.385 $Y=2.67 $X2=0
+ $Y2=0
cc_536 N_A_208_368#_c_571_n N_VPWR_c_1232_n 0.0119432f $X=5.065 $Y=2.937 $X2=0
+ $Y2=0
cc_537 N_A_208_368#_c_559_n N_VPWR_c_1235_n 0.00226527f $X=2.055 $Y=2.63 $X2=0
+ $Y2=0
cc_538 N_A_208_368#_c_567_n N_VPWR_c_1235_n 0.0166417f $X=1.222 $Y=2.63 $X2=0
+ $Y2=0
cc_539 N_A_208_368#_M1026_g N_VPWR_c_1236_n 7.25202e-19 $X=2.64 $Y=2.445 $X2=0
+ $Y2=0
cc_540 N_A_208_368#_c_559_n N_VPWR_c_1236_n 0.00255945f $X=2.055 $Y=2.63 $X2=0
+ $Y2=0
cc_541 N_A_208_368#_c_560_n N_VPWR_c_1236_n 0.02505f $X=3.12 $Y=2.8 $X2=0 $Y2=0
cc_542 N_A_208_368#_c_660_p N_VPWR_c_1236_n 0.00757438f $X=4.3 $Y=2.67 $X2=0
+ $Y2=0
cc_543 N_A_208_368#_c_653_n N_VPWR_c_1236_n 0.00416596f $X=2.14 $Y=2.63 $X2=0
+ $Y2=0
cc_544 N_A_208_368#_c_618_n N_VPWR_c_1236_n 0.00444253f $X=3.205 $Y=2.67 $X2=0
+ $Y2=0
cc_545 N_A_208_368#_c_559_n N_VPWR_c_1226_n 0.00989207f $X=2.055 $Y=2.63 $X2=0
+ $Y2=0
cc_546 N_A_208_368#_c_560_n N_VPWR_c_1226_n 0.0293925f $X=3.12 $Y=2.8 $X2=0
+ $Y2=0
cc_547 N_A_208_368#_c_660_p N_VPWR_c_1226_n 0.0196955f $X=4.3 $Y=2.67 $X2=0
+ $Y2=0
cc_548 N_A_208_368#_c_561_n N_VPWR_c_1226_n 0.019169f $X=4.98 $Y=2.937 $X2=0
+ $Y2=0
cc_549 N_A_208_368#_c_563_n N_VPWR_c_1226_n 0.0312462f $X=5.82 $Y=2.99 $X2=0
+ $Y2=0
cc_550 N_A_208_368#_c_567_n N_VPWR_c_1226_n 0.0149689f $X=1.222 $Y=2.63 $X2=0
+ $Y2=0
cc_551 N_A_208_368#_c_653_n N_VPWR_c_1226_n 0.00563155f $X=2.14 $Y=2.63 $X2=0
+ $Y2=0
cc_552 N_A_208_368#_c_618_n N_VPWR_c_1226_n 0.00495048f $X=3.205 $Y=2.67 $X2=0
+ $Y2=0
cc_553 N_A_208_368#_c_568_n N_VPWR_c_1226_n 0.005864f $X=4.385 $Y=2.67 $X2=0
+ $Y2=0
cc_554 N_A_208_368#_c_571_n N_VPWR_c_1226_n 0.00632998f $X=5.065 $Y=2.937 $X2=0
+ $Y2=0
cc_555 N_A_208_368#_c_660_p N_VPWR_c_1243_n 0.0289114f $X=4.3 $Y=2.67 $X2=0
+ $Y2=0
cc_556 N_A_208_368#_c_568_n N_VPWR_c_1243_n 0.01064f $X=4.385 $Y=2.67 $X2=0
+ $Y2=0
cc_557 N_A_208_368#_c_560_n N_A_423_503#_M1021_d 0.00557612f $X=3.12 $Y=2.8
+ $X2=0 $Y2=0
cc_558 N_A_208_368#_c_653_n N_A_423_503#_M1021_d 0.00558815f $X=2.14 $Y=2.63
+ $X2=0 $Y2=0
cc_559 N_A_208_368#_c_555_n N_A_423_503#_c_1346_n 0.0103878f $X=2.55 $Y=1.74
+ $X2=0 $Y2=0
cc_560 N_A_208_368#_M1026_g N_A_423_503#_c_1346_n 0.00683557f $X=2.64 $Y=2.445
+ $X2=0 $Y2=0
cc_561 N_A_208_368#_c_555_n N_A_423_503#_c_1350_n 0.00679505f $X=2.55 $Y=1.74
+ $X2=0 $Y2=0
cc_562 N_A_208_368#_M1026_g N_A_423_503#_c_1350_n 0.0102444f $X=2.64 $Y=2.445
+ $X2=0 $Y2=0
cc_563 N_A_208_368#_c_560_n N_A_423_503#_c_1350_n 0.015114f $X=3.12 $Y=2.8 $X2=0
+ $Y2=0
cc_564 N_A_208_368#_c_555_n N_A_423_503#_c_1348_n 0.00265578f $X=2.55 $Y=1.74
+ $X2=0 $Y2=0
cc_565 N_A_208_368#_c_554_n N_A_423_503#_c_1348_n 8.98793e-19 $X=1.635 $Y=1.485
+ $X2=0 $Y2=0
cc_566 N_A_208_368#_c_660_p A_653_508# 0.00323545f $X=4.3 $Y=2.67 $X2=-0.19
+ $Y2=-0.245
cc_567 N_A_208_368#_c_564_n A_1161_482# 0.00167911f $X=5.905 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_568 N_A_208_368#_c_544_n N_VGND_c_1447_n 0.002619f $X=1.8 $Y=0.18 $X2=0 $Y2=0
cc_569 N_A_208_368#_c_543_n N_VGND_c_1448_n 0.0244937f $X=3.415 $Y=0.18 $X2=0
+ $Y2=0
cc_570 N_A_208_368#_c_554_n N_VGND_c_1448_n 0.00813824f $X=1.635 $Y=1.485 $X2=0
+ $Y2=0
cc_571 N_A_208_368#_M1010_g N_VGND_c_1452_n 5.91945e-19 $X=4.95 $Y=0.875 $X2=0
+ $Y2=0
cc_572 N_A_208_368#_c_544_n N_VGND_c_1457_n 0.00596402f $X=1.8 $Y=0.18 $X2=0
+ $Y2=0
cc_573 N_A_208_368#_c_543_n N_VGND_c_1458_n 0.0291548f $X=3.415 $Y=0.18 $X2=0
+ $Y2=0
cc_574 N_A_208_368#_c_543_n N_VGND_c_1461_n 0.0363888f $X=3.415 $Y=0.18 $X2=0
+ $Y2=0
cc_575 N_A_208_368#_c_544_n N_VGND_c_1461_n 0.0067234f $X=1.8 $Y=0.18 $X2=0
+ $Y2=0
cc_576 N_A_208_368#_c_543_n N_VGND_c_1464_n 0.00317283f $X=3.415 $Y=0.18 $X2=0
+ $Y2=0
cc_577 N_A_208_368#_M1012_g N_VGND_c_1464_n 7.11128e-19 $X=3.49 $Y=0.72 $X2=0
+ $Y2=0
cc_578 N_A_701_463#_c_778_n N_A_546_447#_M1011_g 0.0087261f $X=3.595 $Y=2.465
+ $X2=0 $Y2=0
cc_579 N_A_701_463#_c_771_n N_A_546_447#_M1011_g 0.00815149f $X=3.735 $Y=2.315
+ $X2=0 $Y2=0
cc_580 N_A_701_463#_c_782_n N_A_546_447#_M1011_g 0.00910687f $X=4.725 $Y=2.42
+ $X2=0 $Y2=0
cc_581 N_A_701_463#_c_783_n N_A_546_447#_M1011_g 0.00439432f $X=4.725 $Y=1.94
+ $X2=0 $Y2=0
cc_582 N_A_701_463#_c_771_n N_A_546_447#_M1008_g 0.0046787f $X=3.735 $Y=2.315
+ $X2=0 $Y2=0
cc_583 N_A_701_463#_c_772_n N_A_546_447#_M1008_g 0.0185727f $X=3.85 $Y=1.04
+ $X2=0 $Y2=0
cc_584 N_A_701_463#_c_773_n N_A_546_447#_M1008_g 0.0116824f $X=4.45 $Y=1.192
+ $X2=0 $Y2=0
cc_585 N_A_701_463#_c_774_n N_A_546_447#_M1008_g 0.00710354f $X=4.535 $Y=1.855
+ $X2=0 $Y2=0
cc_586 N_A_701_463#_c_776_n N_A_546_447#_M1008_g 0.00962983f $X=4.45 $Y=1.015
+ $X2=0 $Y2=0
cc_587 N_A_701_463#_c_777_n N_A_546_447#_M1008_g 0.0246751f $X=3.85 $Y=1.23
+ $X2=0 $Y2=0
cc_588 N_A_701_463#_c_771_n N_A_546_447#_c_868_n 0.0097855f $X=3.735 $Y=2.315
+ $X2=0 $Y2=0
cc_589 N_A_701_463#_c_780_n N_A_546_447#_c_868_n 0.0112145f $X=3.735 $Y=2.39
+ $X2=0 $Y2=0
cc_590 N_A_701_463#_c_772_n N_A_546_447#_c_863_n 2.94886e-19 $X=3.85 $Y=1.04
+ $X2=0 $Y2=0
cc_591 N_A_701_463#_c_771_n N_A_546_447#_c_864_n 0.0062473f $X=3.735 $Y=2.315
+ $X2=0 $Y2=0
cc_592 N_A_701_463#_c_773_n N_A_546_447#_c_864_n 0.0152506f $X=4.45 $Y=1.192
+ $X2=0 $Y2=0
cc_593 N_A_701_463#_c_774_n N_A_546_447#_c_864_n 0.015765f $X=4.535 $Y=1.855
+ $X2=0 $Y2=0
cc_594 N_A_701_463#_c_782_n N_A_546_447#_c_864_n 0.00697091f $X=4.725 $Y=2.42
+ $X2=0 $Y2=0
cc_595 N_A_701_463#_c_783_n N_A_546_447#_c_864_n 0.0127452f $X=4.725 $Y=1.94
+ $X2=0 $Y2=0
cc_596 N_A_701_463#_c_777_n N_A_546_447#_c_864_n 4.9615e-19 $X=3.85 $Y=1.23
+ $X2=0 $Y2=0
cc_597 N_A_701_463#_c_771_n N_A_546_447#_c_865_n 0.0202334f $X=3.735 $Y=2.315
+ $X2=0 $Y2=0
cc_598 N_A_701_463#_c_773_n N_A_546_447#_c_865_n 0.00430875f $X=4.45 $Y=1.192
+ $X2=0 $Y2=0
cc_599 N_A_701_463#_c_774_n N_A_546_447#_c_865_n 0.0075693f $X=4.535 $Y=1.855
+ $X2=0 $Y2=0
cc_600 N_A_701_463#_c_783_n N_A_546_447#_c_865_n 0.00405068f $X=4.725 $Y=1.94
+ $X2=0 $Y2=0
cc_601 N_A_701_463#_c_777_n N_A_546_447#_c_865_n 0.00859211f $X=3.85 $Y=1.23
+ $X2=0 $Y2=0
cc_602 N_A_701_463#_c_775_n N_A_1005_120#_c_1093_n 0.0158988f $X=4.735 $Y=1.005
+ $X2=0 $Y2=0
cc_603 N_A_701_463#_c_778_n N_VPWR_c_1236_n 0.00383477f $X=3.595 $Y=2.465 $X2=0
+ $Y2=0
cc_604 N_A_701_463#_c_778_n N_VPWR_c_1226_n 0.00479598f $X=3.595 $Y=2.465 $X2=0
+ $Y2=0
cc_605 N_A_701_463#_c_778_n N_VPWR_c_1243_n 0.00447856f $X=3.595 $Y=2.465 $X2=0
+ $Y2=0
cc_606 N_A_701_463#_c_772_n N_VGND_c_1458_n 0.00365461f $X=3.85 $Y=1.04 $X2=0
+ $Y2=0
cc_607 N_A_701_463#_c_772_n N_VGND_c_1461_n 0.00502397f $X=3.85 $Y=1.04 $X2=0
+ $Y2=0
cc_608 N_A_701_463#_c_772_n N_VGND_c_1464_n 3.57863e-19 $X=3.85 $Y=1.04 $X2=0
+ $Y2=0
cc_609 N_A_546_447#_c_868_n N_VPWR_M1019_d 0.003889f $X=4.02 $Y=2.33 $X2=0 $Y2=0
cc_610 N_A_546_447#_c_864_n N_VPWR_M1019_d 0.00108265f $X=4.185 $Y=1.795 $X2=0
+ $Y2=0
cc_611 N_A_546_447#_M1011_g N_VPWR_c_1232_n 0.00335016f $X=4.425 $Y=2.54 $X2=0
+ $Y2=0
cc_612 N_A_546_447#_M1011_g N_VPWR_c_1226_n 0.0042684f $X=4.425 $Y=2.54 $X2=0
+ $Y2=0
cc_613 N_A_546_447#_M1011_g N_VPWR_c_1243_n 9.94773e-19 $X=4.425 $Y=2.54 $X2=0
+ $Y2=0
cc_614 N_A_546_447#_c_861_n N_A_423_503#_c_1346_n 0.0335416f $X=2.865 $Y=2.245
+ $X2=0 $Y2=0
cc_615 N_A_546_447#_c_862_n N_A_423_503#_c_1346_n 0.013911f $X=3.19 $Y=1.41
+ $X2=0 $Y2=0
cc_616 N_A_546_447#_c_863_n N_A_423_503#_c_1346_n 0.00585369f $X=3.23 $Y=0.77
+ $X2=0 $Y2=0
cc_617 N_A_546_447#_c_863_n N_A_423_503#_c_1347_n 0.0182668f $X=3.23 $Y=0.77
+ $X2=0 $Y2=0
cc_618 N_A_546_447#_c_861_n N_A_423_503#_c_1350_n 0.0147123f $X=2.865 $Y=2.245
+ $X2=0 $Y2=0
cc_619 N_A_546_447#_c_862_n N_A_423_503#_c_1348_n 0.0079066f $X=3.19 $Y=1.41
+ $X2=0 $Y2=0
cc_620 N_A_546_447#_c_863_n N_A_423_503#_c_1348_n 0.0128522f $X=3.23 $Y=0.77
+ $X2=0 $Y2=0
cc_621 N_A_546_447#_M1008_g N_VGND_c_1452_n 0.00423157f $X=4.44 $Y=0.655 $X2=0
+ $Y2=0
cc_622 N_A_546_447#_M1008_g N_VGND_c_1461_n 0.00542671f $X=4.44 $Y=0.655 $X2=0
+ $Y2=0
cc_623 N_A_546_447#_M1008_g N_VGND_c_1464_n 0.00389779f $X=4.44 $Y=0.655 $X2=0
+ $Y2=0
cc_624 N_A_1191_120#_M1006_g N_A_1005_120#_M1018_g 0.0197751f $X=7.59 $Y=0.74
+ $X2=0 $Y2=0
cc_625 N_A_1191_120#_c_955_n N_A_1005_120#_M1018_g 0.00663814f $X=6.805 $Y=0.645
+ $X2=0 $Y2=0
cc_626 N_A_1191_120#_c_956_n N_A_1005_120#_M1018_g 0.00896052f $X=7.3 $Y=0.935
+ $X2=0 $Y2=0
cc_627 N_A_1191_120#_c_957_n N_A_1005_120#_M1018_g 0.0041803f $X=6.97 $Y=0.935
+ $X2=0 $Y2=0
cc_628 N_A_1191_120#_c_962_n N_A_1005_120#_M1018_g 0.00357382f $X=7.515 $Y=1.35
+ $X2=0 $Y2=0
cc_629 N_A_1191_120#_c_948_n N_A_1005_120#_c_1091_n 3.87964e-19 $X=6.03 $Y=1.225
+ $X2=0 $Y2=0
cc_630 N_A_1191_120#_M1006_g N_A_1005_120#_c_1091_n 0.00426361f $X=7.59 $Y=0.74
+ $X2=0 $Y2=0
cc_631 N_A_1191_120#_c_952_n N_A_1005_120#_c_1091_n 0.00772793f $X=6.305 $Y=1.3
+ $X2=0 $Y2=0
cc_632 N_A_1191_120#_c_953_n N_A_1005_120#_c_1091_n 7.19653e-19 $X=6.395 $Y=1.55
+ $X2=0 $Y2=0
cc_633 N_A_1191_120#_c_956_n N_A_1005_120#_c_1091_n 0.00249534f $X=7.3 $Y=0.935
+ $X2=0 $Y2=0
cc_634 N_A_1191_120#_c_957_n N_A_1005_120#_c_1091_n 0.00335661f $X=6.97 $Y=0.935
+ $X2=0 $Y2=0
cc_635 N_A_1191_120#_c_958_n N_A_1005_120#_c_1091_n 0.00594113f $X=7.04 $Y=1.775
+ $X2=0 $Y2=0
cc_636 N_A_1191_120#_c_959_n N_A_1005_120#_c_1091_n 0.00611837f $X=6.395
+ $Y=1.715 $X2=0 $Y2=0
cc_637 N_A_1191_120#_c_960_n N_A_1005_120#_c_1091_n 0.00444742f $X=7.565
+ $Y=1.515 $X2=0 $Y2=0
cc_638 N_A_1191_120#_c_961_n N_A_1005_120#_c_1091_n 0.0185323f $X=7.565 $Y=1.515
+ $X2=0 $Y2=0
cc_639 N_A_1191_120#_c_962_n N_A_1005_120#_c_1091_n 0.00238376f $X=7.515 $Y=1.35
+ $X2=0 $Y2=0
cc_640 N_A_1191_120#_M1024_g N_A_1005_120#_M1001_g 0.0185f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_641 N_A_1191_120#_c_967_n N_A_1005_120#_M1001_g 0.00611837f $X=6.395 $Y=2.185
+ $X2=0 $Y2=0
cc_642 N_A_1191_120#_c_969_n N_A_1005_120#_M1001_g 0.00840951f $X=6.875 $Y=2.695
+ $X2=0 $Y2=0
cc_643 N_A_1191_120#_c_970_n N_A_1005_120#_M1001_g 0.0128186f $X=7.3 $Y=1.775
+ $X2=0 $Y2=0
cc_644 N_A_1191_120#_c_958_n N_A_1005_120#_M1001_g 0.0093215f $X=7.04 $Y=1.775
+ $X2=0 $Y2=0
cc_645 N_A_1191_120#_c_960_n N_A_1005_120#_M1001_g 2.5449e-19 $X=7.565 $Y=1.515
+ $X2=0 $Y2=0
cc_646 N_A_1191_120#_c_948_n N_A_1005_120#_c_1093_n 0.00155055f $X=6.03 $Y=1.225
+ $X2=0 $Y2=0
cc_647 N_A_1191_120#_c_953_n N_A_1005_120#_c_1095_n 8.9934e-19 $X=6.395 $Y=1.55
+ $X2=0 $Y2=0
cc_648 N_A_1191_120#_c_956_n N_A_1005_120#_c_1095_n 0.0115232f $X=7.3 $Y=0.935
+ $X2=0 $Y2=0
cc_649 N_A_1191_120#_c_957_n N_A_1005_120#_c_1095_n 0.01404f $X=6.97 $Y=0.935
+ $X2=0 $Y2=0
cc_650 N_A_1191_120#_c_970_n N_A_1005_120#_c_1095_n 0.00639324f $X=7.3 $Y=1.775
+ $X2=0 $Y2=0
cc_651 N_A_1191_120#_c_958_n N_A_1005_120#_c_1095_n 0.0201047f $X=7.04 $Y=1.775
+ $X2=0 $Y2=0
cc_652 N_A_1191_120#_c_962_n N_A_1005_120#_c_1095_n 0.0264444f $X=7.515 $Y=1.35
+ $X2=0 $Y2=0
cc_653 N_A_1191_120#_c_948_n N_A_1005_120#_c_1096_n 0.00626979f $X=6.03 $Y=1.225
+ $X2=0 $Y2=0
cc_654 N_A_1191_120#_c_952_n N_A_1005_120#_c_1096_n 0.0172282f $X=6.305 $Y=1.3
+ $X2=0 $Y2=0
cc_655 N_A_1191_120#_c_953_n N_A_1005_120#_c_1096_n 0.00208941f $X=6.395 $Y=1.55
+ $X2=0 $Y2=0
cc_656 N_A_1191_120#_c_957_n N_A_1005_120#_c_1096_n 0.0122939f $X=6.97 $Y=0.935
+ $X2=0 $Y2=0
cc_657 N_A_1191_120#_c_958_n N_A_1005_120#_c_1096_n 0.0389282f $X=7.04 $Y=1.775
+ $X2=0 $Y2=0
cc_658 N_A_1191_120#_c_959_n N_A_1005_120#_c_1096_n 0.00125196f $X=6.395
+ $Y=1.715 $X2=0 $Y2=0
cc_659 N_A_1191_120#_c_954_n N_A_1644_112#_M1000_g 0.0169957f $X=8.505 $Y=1.35
+ $X2=0 $Y2=0
cc_660 N_A_1191_120#_M1022_g N_A_1644_112#_M1027_g 0.0149415f $X=8.58 $Y=0.835
+ $X2=0 $Y2=0
cc_661 N_A_1191_120#_M1006_g N_A_1644_112#_c_1175_n 0.00156978f $X=7.59 $Y=0.74
+ $X2=0 $Y2=0
cc_662 N_A_1191_120#_M1022_g N_A_1644_112#_c_1175_n 0.0142937f $X=8.58 $Y=0.835
+ $X2=0 $Y2=0
cc_663 N_A_1191_120#_M1024_g N_A_1644_112#_c_1180_n 0.00175548f $X=7.605 $Y=2.4
+ $X2=0 $Y2=0
cc_664 N_A_1191_120#_c_950_n N_A_1644_112#_c_1180_n 0.00570762f $X=8.505
+ $Y=1.515 $X2=0 $Y2=0
cc_665 N_A_1191_120#_M1007_g N_A_1644_112#_c_1180_n 0.00971694f $X=8.595 $Y=2.26
+ $X2=0 $Y2=0
cc_666 N_A_1191_120#_M1022_g N_A_1644_112#_c_1176_n 0.00697058f $X=8.58 $Y=0.835
+ $X2=0 $Y2=0
cc_667 N_A_1191_120#_c_954_n N_A_1644_112#_c_1176_n 0.0132449f $X=8.505 $Y=1.35
+ $X2=0 $Y2=0
cc_668 N_A_1191_120#_M1022_g N_A_1644_112#_c_1177_n 0.0126574f $X=8.58 $Y=0.835
+ $X2=0 $Y2=0
cc_669 N_A_1191_120#_c_954_n N_A_1644_112#_c_1177_n 0.00652611f $X=8.505 $Y=1.35
+ $X2=0 $Y2=0
cc_670 N_A_1191_120#_c_950_n N_A_1644_112#_c_1178_n 0.0163108f $X=8.505 $Y=1.515
+ $X2=0 $Y2=0
cc_671 N_A_1191_120#_M1022_g N_A_1644_112#_c_1178_n 0.0010393f $X=8.58 $Y=0.835
+ $X2=0 $Y2=0
cc_672 N_A_1191_120#_c_954_n N_A_1644_112#_c_1178_n 0.00195703f $X=8.505 $Y=1.35
+ $X2=0 $Y2=0
cc_673 N_A_1191_120#_c_970_n N_VPWR_M1001_d 6.09984e-19 $X=7.3 $Y=1.775 $X2=0
+ $Y2=0
cc_674 N_A_1191_120#_c_960_n N_VPWR_M1001_d 0.0017826f $X=7.565 $Y=1.515 $X2=0
+ $Y2=0
cc_675 N_A_1191_120#_c_963_n N_VPWR_c_1229_n 0.0119707f $X=6.105 $Y=2.335 $X2=0
+ $Y2=0
cc_676 N_A_1191_120#_c_967_n N_VPWR_c_1229_n 0.00988509f $X=6.395 $Y=2.185 $X2=0
+ $Y2=0
cc_677 N_A_1191_120#_c_969_n N_VPWR_c_1229_n 0.0332024f $X=6.875 $Y=2.695 $X2=0
+ $Y2=0
cc_678 N_A_1191_120#_c_958_n N_VPWR_c_1229_n 0.0235084f $X=7.04 $Y=1.775 $X2=0
+ $Y2=0
cc_679 N_A_1191_120#_M1024_g N_VPWR_c_1230_n 0.00595969f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_680 N_A_1191_120#_c_969_n N_VPWR_c_1230_n 0.0217281f $X=6.875 $Y=2.695 $X2=0
+ $Y2=0
cc_681 N_A_1191_120#_c_970_n N_VPWR_c_1230_n 0.004312f $X=7.3 $Y=1.775 $X2=0
+ $Y2=0
cc_682 N_A_1191_120#_c_960_n N_VPWR_c_1230_n 0.0141554f $X=7.565 $Y=1.515 $X2=0
+ $Y2=0
cc_683 N_A_1191_120#_c_961_n N_VPWR_c_1230_n 3.95452e-19 $X=7.565 $Y=1.515 $X2=0
+ $Y2=0
cc_684 N_A_1191_120#_M1007_g N_VPWR_c_1231_n 0.0180689f $X=8.595 $Y=2.26 $X2=0
+ $Y2=0
cc_685 N_A_1191_120#_c_963_n N_VPWR_c_1232_n 0.0048655f $X=6.105 $Y=2.335 $X2=0
+ $Y2=0
cc_686 N_A_1191_120#_c_969_n N_VPWR_c_1237_n 0.00975961f $X=6.875 $Y=2.695 $X2=0
+ $Y2=0
cc_687 N_A_1191_120#_M1024_g N_VPWR_c_1238_n 0.005209f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_688 N_A_1191_120#_M1007_g N_VPWR_c_1238_n 0.00401533f $X=8.595 $Y=2.26 $X2=0
+ $Y2=0
cc_689 N_A_1191_120#_c_963_n N_VPWR_c_1226_n 0.00508748f $X=6.105 $Y=2.335 $X2=0
+ $Y2=0
cc_690 N_A_1191_120#_M1024_g N_VPWR_c_1226_n 0.00991972f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_691 N_A_1191_120#_M1007_g N_VPWR_c_1226_n 0.00465661f $X=8.595 $Y=2.26 $X2=0
+ $Y2=0
cc_692 N_A_1191_120#_c_969_n N_VPWR_c_1226_n 0.0111753f $X=6.875 $Y=2.695 $X2=0
+ $Y2=0
cc_693 N_A_1191_120#_M1006_g N_Q_c_1387_n 0.00946122f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_694 N_A_1191_120#_M1022_g N_Q_c_1387_n 0.00582178f $X=8.58 $Y=0.835 $X2=0
+ $Y2=0
cc_695 N_A_1191_120#_c_955_n N_Q_c_1387_n 0.00412382f $X=6.805 $Y=0.645 $X2=0
+ $Y2=0
cc_696 N_A_1191_120#_M1006_g N_Q_c_1388_n 0.00301591f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_697 N_A_1191_120#_c_950_n N_Q_c_1388_n 0.00621855f $X=8.505 $Y=1.515 $X2=0
+ $Y2=0
cc_698 N_A_1191_120#_c_960_n N_Q_c_1388_n 0.00618485f $X=7.565 $Y=1.515 $X2=0
+ $Y2=0
cc_699 N_A_1191_120#_c_962_n N_Q_c_1388_n 0.00501288f $X=7.515 $Y=1.35 $X2=0
+ $Y2=0
cc_700 N_A_1191_120#_M1024_g N_Q_c_1390_n 0.00270626f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_701 N_A_1191_120#_c_950_n N_Q_c_1390_n 0.00422012f $X=8.505 $Y=1.515 $X2=0
+ $Y2=0
cc_702 N_A_1191_120#_c_960_n N_Q_c_1390_n 0.00235997f $X=7.565 $Y=1.515 $X2=0
+ $Y2=0
cc_703 N_A_1191_120#_M1006_g N_Q_c_1389_n 0.00341467f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_704 N_A_1191_120#_M1024_g N_Q_c_1389_n 0.0051987f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_705 N_A_1191_120#_c_950_n N_Q_c_1389_n 0.0230273f $X=8.505 $Y=1.515 $X2=0
+ $Y2=0
cc_706 N_A_1191_120#_M1007_g N_Q_c_1389_n 0.00393262f $X=8.595 $Y=2.26 $X2=0
+ $Y2=0
cc_707 N_A_1191_120#_c_960_n N_Q_c_1389_n 0.0377164f $X=7.565 $Y=1.515 $X2=0
+ $Y2=0
cc_708 N_A_1191_120#_c_962_n N_Q_c_1389_n 0.00668697f $X=7.515 $Y=1.35 $X2=0
+ $Y2=0
cc_709 N_A_1191_120#_M1024_g Q 0.014097f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_710 N_A_1191_120#_M1007_g Q_N 3.73184e-19 $X=8.595 $Y=2.26 $X2=0 $Y2=0
cc_711 N_A_1191_120#_c_956_n N_VGND_M1018_d 0.00564413f $X=7.3 $Y=0.935 $X2=0
+ $Y2=0
cc_712 N_A_1191_120#_c_962_n N_VGND_M1018_d 0.00178719f $X=7.515 $Y=1.35 $X2=0
+ $Y2=0
cc_713 N_A_1191_120#_c_948_n N_VGND_c_1449_n 0.0109574f $X=6.03 $Y=1.225 $X2=0
+ $Y2=0
cc_714 N_A_1191_120#_c_952_n N_VGND_c_1449_n 0.00192045f $X=6.305 $Y=1.3 $X2=0
+ $Y2=0
cc_715 N_A_1191_120#_c_955_n N_VGND_c_1449_n 0.027608f $X=6.805 $Y=0.645 $X2=0
+ $Y2=0
cc_716 N_A_1191_120#_c_957_n N_VGND_c_1449_n 0.0121616f $X=6.97 $Y=0.935 $X2=0
+ $Y2=0
cc_717 N_A_1191_120#_M1006_g N_VGND_c_1450_n 0.00525427f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_718 N_A_1191_120#_c_956_n N_VGND_c_1450_n 0.0256676f $X=7.3 $Y=0.935 $X2=0
+ $Y2=0
cc_719 N_A_1191_120#_M1022_g N_VGND_c_1451_n 0.00492504f $X=8.58 $Y=0.835 $X2=0
+ $Y2=0
cc_720 N_A_1191_120#_c_948_n N_VGND_c_1452_n 0.00302627f $X=6.03 $Y=1.225 $X2=0
+ $Y2=0
cc_721 N_A_1191_120#_M1006_g N_VGND_c_1454_n 0.00434272f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_722 N_A_1191_120#_M1022_g N_VGND_c_1454_n 0.00434543f $X=8.58 $Y=0.835 $X2=0
+ $Y2=0
cc_723 N_A_1191_120#_c_955_n N_VGND_c_1459_n 0.00942501f $X=6.805 $Y=0.645 $X2=0
+ $Y2=0
cc_724 N_A_1191_120#_c_948_n N_VGND_c_1461_n 0.00370742f $X=6.03 $Y=1.225 $X2=0
+ $Y2=0
cc_725 N_A_1191_120#_M1006_g N_VGND_c_1461_n 0.00826311f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_726 N_A_1191_120#_M1022_g N_VGND_c_1461_n 0.00487769f $X=8.58 $Y=0.835 $X2=0
+ $Y2=0
cc_727 N_A_1191_120#_c_955_n N_VGND_c_1461_n 0.011246f $X=6.805 $Y=0.645 $X2=0
+ $Y2=0
cc_728 N_A_1191_120#_c_956_n N_VGND_c_1461_n 0.00605933f $X=7.3 $Y=0.935 $X2=0
+ $Y2=0
cc_729 N_A_1005_120#_M1001_g N_VPWR_c_1229_n 0.0037362f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_730 N_A_1005_120#_M1001_g N_VPWR_c_1230_n 0.00365529f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_731 N_A_1005_120#_M1001_g N_VPWR_c_1237_n 0.00567889f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_732 N_A_1005_120#_M1001_g N_VPWR_c_1226_n 0.00610055f $X=7.1 $Y=2.34 $X2=0
+ $Y2=0
cc_733 N_A_1005_120#_M1018_g N_Q_c_1387_n 7.09617e-19 $X=7.02 $Y=0.645 $X2=0
+ $Y2=0
cc_734 N_A_1005_120#_M1018_g N_VGND_c_1449_n 0.00695165f $X=7.02 $Y=0.645 $X2=0
+ $Y2=0
cc_735 N_A_1005_120#_c_1093_n N_VGND_c_1449_n 0.00815067f $X=5.405 $Y=1.38 $X2=0
+ $Y2=0
cc_736 N_A_1005_120#_c_1096_n N_VGND_c_1449_n 0.0243987f $X=6.8 $Y=1.355 $X2=0
+ $Y2=0
cc_737 N_A_1005_120#_M1018_g N_VGND_c_1450_n 0.00563133f $X=7.02 $Y=0.645 $X2=0
+ $Y2=0
cc_738 N_A_1005_120#_M1018_g N_VGND_c_1459_n 0.00436157f $X=7.02 $Y=0.645 $X2=0
+ $Y2=0
cc_739 N_A_1005_120#_M1018_g N_VGND_c_1461_n 0.00455189f $X=7.02 $Y=0.645 $X2=0
+ $Y2=0
cc_740 N_A_1644_112#_M1000_g N_VPWR_c_1231_n 0.00986253f $X=9.1 $Y=2.4 $X2=0
+ $Y2=0
cc_741 N_A_1644_112#_c_1180_n N_VPWR_c_1231_n 0.0302727f $X=8.37 $Y=1.985 $X2=0
+ $Y2=0
cc_742 N_A_1644_112#_c_1176_n N_VPWR_c_1231_n 0.0261911f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_743 N_A_1644_112#_c_1177_n N_VPWR_c_1231_n 0.00205259f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_744 N_A_1644_112#_c_1180_n N_VPWR_c_1238_n 0.0035402f $X=8.37 $Y=1.985 $X2=0
+ $Y2=0
cc_745 N_A_1644_112#_M1000_g N_VPWR_c_1239_n 0.005209f $X=9.1 $Y=2.4 $X2=0 $Y2=0
cc_746 N_A_1644_112#_M1000_g N_VPWR_c_1226_n 0.00990563f $X=9.1 $Y=2.4 $X2=0
+ $Y2=0
cc_747 N_A_1644_112#_c_1180_n N_VPWR_c_1226_n 0.00526929f $X=8.37 $Y=1.985 $X2=0
+ $Y2=0
cc_748 N_A_1644_112#_c_1175_n N_Q_c_1387_n 0.0471589f $X=8.365 $Y=0.835 $X2=0
+ $Y2=0
cc_749 N_A_1644_112#_c_1180_n N_Q_c_1389_n 0.0713906f $X=8.37 $Y=1.985 $X2=0
+ $Y2=0
cc_750 N_A_1644_112#_c_1178_n N_Q_c_1389_n 0.021634f $X=8.405 $Y=1.465 $X2=0
+ $Y2=0
cc_751 N_A_1644_112#_M1027_g N_Q_N_c_1422_n 0.00812323f $X=9.09 $Y=0.74 $X2=0
+ $Y2=0
cc_752 N_A_1644_112#_M1027_g N_Q_N_c_1423_n 0.00270338f $X=9.09 $Y=0.74 $X2=0
+ $Y2=0
cc_753 N_A_1644_112#_c_1176_n N_Q_N_c_1423_n 0.00275913f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_754 N_A_1644_112#_c_1177_n N_Q_N_c_1423_n 0.00255363f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_755 N_A_1644_112#_M1000_g Q_N 0.00329601f $X=9.1 $Y=2.4 $X2=0 $Y2=0
cc_756 N_A_1644_112#_c_1176_n Q_N 0.00102175f $X=9.06 $Y=1.465 $X2=0 $Y2=0
cc_757 N_A_1644_112#_c_1177_n Q_N 0.00152224f $X=9.06 $Y=1.465 $X2=0 $Y2=0
cc_758 N_A_1644_112#_M1000_g Q_N 0.0129762f $X=9.1 $Y=2.4 $X2=0 $Y2=0
cc_759 N_A_1644_112#_M1000_g N_Q_N_c_1424_n 0.00495575f $X=9.1 $Y=2.4 $X2=0
+ $Y2=0
cc_760 N_A_1644_112#_M1027_g N_Q_N_c_1424_n 0.00404757f $X=9.09 $Y=0.74 $X2=0
+ $Y2=0
cc_761 N_A_1644_112#_c_1176_n N_Q_N_c_1424_n 0.0262108f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_762 N_A_1644_112#_c_1177_n N_Q_N_c_1424_n 0.00787524f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_763 N_A_1644_112#_M1027_g N_VGND_c_1451_n 0.00536023f $X=9.09 $Y=0.74 $X2=0
+ $Y2=0
cc_764 N_A_1644_112#_c_1175_n N_VGND_c_1451_n 0.0180739f $X=8.365 $Y=0.835 $X2=0
+ $Y2=0
cc_765 N_A_1644_112#_c_1176_n N_VGND_c_1451_n 0.0216743f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_766 N_A_1644_112#_c_1177_n N_VGND_c_1451_n 0.00149092f $X=9.06 $Y=1.465 $X2=0
+ $Y2=0
cc_767 N_A_1644_112#_c_1175_n N_VGND_c_1454_n 0.00430431f $X=8.365 $Y=0.835
+ $X2=0 $Y2=0
cc_768 N_A_1644_112#_M1027_g N_VGND_c_1460_n 0.00434272f $X=9.09 $Y=0.74 $X2=0
+ $Y2=0
cc_769 N_A_1644_112#_M1027_g N_VGND_c_1461_n 0.00828991f $X=9.09 $Y=0.74 $X2=0
+ $Y2=0
cc_770 N_A_1644_112#_c_1175_n N_VGND_c_1461_n 0.00755262f $X=8.365 $Y=0.835
+ $X2=0 $Y2=0
cc_771 N_VPWR_c_1230_n N_Q_c_1390_n 0.0366401f $X=7.325 $Y=2.195 $X2=0 $Y2=0
cc_772 N_VPWR_c_1231_n Q 0.00957944f $X=8.82 $Y=1.985 $X2=0 $Y2=0
cc_773 N_VPWR_c_1238_n Q 0.0178955f $X=8.655 $Y=3.33 $X2=0 $Y2=0
cc_774 N_VPWR_c_1226_n Q 0.0147443f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_775 N_VPWR_c_1231_n Q_N 0.0445151f $X=8.82 $Y=1.985 $X2=0 $Y2=0
cc_776 N_VPWR_c_1239_n Q_N 0.0156645f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_777 N_VPWR_c_1226_n Q_N 0.0128976f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_778 N_Q_c_1387_n N_VGND_c_1450_n 0.0136846f $X=7.805 $Y=0.515 $X2=0 $Y2=0
cc_779 N_Q_c_1387_n N_VGND_c_1451_n 0.00798967f $X=7.805 $Y=0.515 $X2=0 $Y2=0
cc_780 N_Q_c_1387_n N_VGND_c_1454_n 0.019026f $X=7.805 $Y=0.515 $X2=0 $Y2=0
cc_781 N_Q_c_1387_n N_VGND_c_1461_n 0.0156917f $X=7.805 $Y=0.515 $X2=0 $Y2=0
cc_782 N_Q_N_c_1422_n N_VGND_c_1451_n 0.0299279f $X=9.305 $Y=0.515 $X2=0 $Y2=0
cc_783 N_Q_N_c_1422_n N_VGND_c_1460_n 0.0165719f $X=9.305 $Y=0.515 $X2=0 $Y2=0
cc_784 N_Q_N_c_1422_n N_VGND_c_1461_n 0.0136604f $X=9.305 $Y=0.515 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_231_132# CI VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.06802e+12p pd=6.52e+06u as=2.27012e+12p ps=1.57e+07u
M1001 a_410_58# a_811_379# a_879_55# VNB nlowvt w=640000u l=150000u
+  ad=2.6395e+11p pd=2.41e+06u as=4.9405e+11p ps=5.22e+06u
M1002 a_83_21# a_811_379# a_231_132# VNB nlowvt w=640000u l=150000u
+  ad=2.375e+11p pd=2.16e+06u as=3.808e+11p ps=3.75e+06u
M1003 a_644_104# a_231_132# VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.31125e+11p pd=3.21e+06u as=0p ps=0u
M1004 a_811_379# a_879_55# a_1852_374# VNB nlowvt w=640000u l=150000u
+  ad=6.528e+11p pd=3.32e+06u as=5.128e+11p ps=4.25e+06u
M1005 a_1023_379# a_879_55# a_1852_374# VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=1.57615e+12p ps=7.29e+06u
M1006 a_1023_379# a_879_55# a_1660_374# VNB nlowvt w=640000u l=150000u
+  ad=4.965e+11p pd=2.98e+06u as=5.157e+11p ps=4.37e+06u
M1007 VPWR a_410_58# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.5085e+11p ps=3.26e+06u
M1008 VGND a_410_58# COUT VNB nlowvt w=740000u l=150000u
+  ad=1.8144e+12p pd=1.292e+07u as=2.072e+11p ps=2.04e+06u
M1009 a_1660_374# B a_1023_379# VPB pshort w=840000u l=180000u
+  ad=5.782e+11p pd=5.13e+06u as=0p ps=0u
M1010 a_410_58# a_811_379# a_231_132# VPB pshort w=840000u l=180000u
+  ad=4.83e+11p pd=2.83e+06u as=0p ps=0u
M1011 a_1852_374# B a_811_379# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.688e+11p ps=2.32e+06u
M1012 a_231_132# CI VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_811_379# a_879_55# a_1660_374# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2342_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1015 VPWR a_83_21# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1016 a_231_132# a_1023_379# a_410_58# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_83_21# a_811_379# a_644_104# VPB pshort w=840000u l=180000u
+  ad=7.392e+11p pd=3.44e+06u as=0p ps=0u
M1018 VGND A a_1852_374# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_879_55# a_1023_379# a_410_58# VPB pshort w=840000u l=180000u
+  ad=3.742e+11p pd=2.95e+06u as=0p ps=0u
M1020 a_644_104# a_1023_379# a_83_21# VNB nlowvt w=640000u l=150000u
+  ad=4.1745e+11p pd=3.87e+06u as=0p ps=0u
M1021 VPWR B a_879_55# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_2342_48# a_1660_374# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND B a_879_55# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1660_374# B a_811_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_644_104# a_231_132# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_83_21# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1027 a_1852_374# B a_1023_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_231_132# a_1023_379# a_83_21# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2342_48# a_1660_374# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_1852_374# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2342_48# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

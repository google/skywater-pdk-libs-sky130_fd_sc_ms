# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__nand3_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__nand3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.847200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.535000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.847200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.130000 1.350000 3.715000 1.630000 ;
        RECT 2.560000 1.630000 3.715000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.847200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.140000 1.340000 6.115000 1.630000 ;
        RECT 4.495000 1.630000 6.115000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.904000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 1.725000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.950000 ;
        RECT 0.125000 1.950000 4.290000 2.120000 ;
        RECT 0.535000 0.595000 0.865000 1.010000 ;
        RECT 0.615000 2.120000 1.365000 2.980000 ;
        RECT 1.395000 0.595000 1.725000 1.010000 ;
        RECT 2.035000 1.820000 2.365000 1.950000 ;
        RECT 2.035000 2.120000 2.365000 2.980000 ;
        RECT 3.960000 1.820000 4.290000 1.950000 ;
        RECT 3.960000 2.120000 4.290000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.105000  0.255000 3.875000 0.425000 ;
      RECT 0.105000  0.425000 0.355000 0.840000 ;
      RECT 0.115000  2.290000 0.445000 3.245000 ;
      RECT 1.045000  0.425000 1.215000 0.840000 ;
      RECT 1.535000  2.290000 1.865000 3.245000 ;
      RECT 1.905000  0.425000 2.075000 1.170000 ;
      RECT 2.255000  0.595000 2.585000 0.920000 ;
      RECT 2.255000  0.920000 5.625000 1.170000 ;
      RECT 2.535000  2.290000 3.790000 3.245000 ;
      RECT 2.755000  0.425000 2.945000 0.750000 ;
      RECT 3.115000  0.595000 3.445000 0.920000 ;
      RECT 3.615000  0.425000 3.875000 0.750000 ;
      RECT 4.085000  0.085000 4.415000 0.750000 ;
      RECT 4.460000  1.950000 5.765000 3.245000 ;
      RECT 4.585000  0.390000 4.775000 0.920000 ;
      RECT 4.945000  0.085000 5.275000 0.750000 ;
      RECT 5.455000  0.390000 5.625000 0.920000 ;
      RECT 5.805000  0.085000 6.135000 1.170000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_ms__nand3_4

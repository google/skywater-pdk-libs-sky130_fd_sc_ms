* File: sky130_fd_sc_ms__and2_4.spice
* Created: Fri Aug 28 17:10:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and2_4.pex.spice"
.subckt sky130_fd_sc_ms__and2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_83_269#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_83_269#_M1001_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1001_d N_A_83_269#_M1003_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1591 PD=1.02 PS=1.17 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_83_269#_M1012_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13883 AS=0.1591 PD=1.17971 PS=1.17 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75001.6 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1004 N_A_504_119#_M1004_d N_B_M1004_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0976 AS=0.12007 PD=0.945 PS=1.02029 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75002.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_83_269#_M1002_d N_A_M1002_g N_A_504_119#_M1004_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.104 AS=0.0976 PD=0.965 PS=0.945 NRD=8.436 NRS=4.68 M=1 R=4.26667
+ SA=75002.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_83_269#_M1002_d N_A_M1005_g N_A_504_119#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.104 AS=0.096 PD=0.965 PS=0.94 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_504_119#_M1005_s N_B_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.096 AS=0.1824 PD=0.94 PS=1.85 NRD=3.744 NRS=0 M=1 R=4.26667 SA=75003.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_X_M1006_d N_A_83_269#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1006_d N_A_83_269#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1009_d N_A_83_269#_M1009_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.1512 PD=1.41 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1010 N_X_M1009_d N_A_83_269#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.211686 PD=1.41 PS=1.68571 NRD=2.6201 NRS=0 M=1 R=6.22222
+ SA=90001.6 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1013 N_A_83_269#_M1013_d N_B_M1013_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1239 AS=0.158764 PD=1.135 PS=1.26429 NRD=0 NRS=19.3454 M=1 R=4.66667
+ SA=90002.1 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_A_83_269#_M1013_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1239 AS=0.1239 PD=1.135 PS=1.135 NRD=4.6886 NRS=4.6886 M=1 R=4.66667
+ SA=90002.6 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1014 N_VPWR_M1011_d N_A_M1014_g N_A_83_269#_M1014_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1239 AS=0.1134 PD=1.135 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667 SA=90003
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1015 N_A_83_269#_M1014_s N_B_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90003.5
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_81 VPB 0 2.91098e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__and2_4.pxi.spice"
*
.ends
*
*

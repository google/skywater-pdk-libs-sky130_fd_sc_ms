* File: sky130_fd_sc_ms__decap_8.pxi.spice
* Created: Wed Sep  2 12:02:15 2020
* 
x_PM_SKY130_FD_SC_MS__DECAP_8%VGND N_VGND_M1001_s N_VGND_M1000_g N_VGND_M1002_g
+ N_VGND_c_30_n N_VGND_c_31_n N_VGND_c_32_n N_VGND_c_33_n N_VGND_c_34_n
+ N_VGND_c_35_n VGND N_VGND_c_36_n N_VGND_c_37_n N_VGND_c_38_n N_VGND_c_39_n
+ N_VGND_c_40_n N_VGND_c_41_n PM_SKY130_FD_SC_MS__DECAP_8%VGND
x_PM_SKY130_FD_SC_MS__DECAP_8%VPWR N_VPWR_M1000_s N_VPWR_c_74_n N_VPWR_c_75_n
+ N_VPWR_c_76_n N_VPWR_c_71_n N_VPWR_c_72_n N_VPWR_c_78_n N_VPWR_c_79_n
+ N_VPWR_c_80_n VPWR N_VPWR_M1001_g N_VPWR_M1003_g N_VPWR_c_81_n N_VPWR_c_73_n
+ N_VPWR_c_83_n PM_SKY130_FD_SC_MS__DECAP_8%VPWR
cc_1 VNB N_VGND_c_30_n 0.0180938f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.085
cc_2 VNB N_VGND_c_31_n 0.0675204f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.64
cc_3 VNB N_VGND_c_32_n 0.042044f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.42
cc_4 VNB N_VGND_c_33_n 0.00319093f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.64
cc_5 VNB N_VGND_c_34_n 0.0730389f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=0.64
cc_6 VNB N_VGND_c_35_n 0.0392248f $X=-0.19 $Y=-0.245 $X2=2.52 $Y2=1.42
cc_7 VNB N_VGND_c_36_n 0.0221481f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0
cc_8 VNB N_VGND_c_37_n 0.0178522f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0
cc_9 VNB N_VGND_c_38_n 0.0271236f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_10 VNB N_VGND_c_39_n 0.239022f $X=-0.19 $Y=-0.245 $X2=3.6 $Y2=0
cc_11 VNB N_VGND_c_40_n 0.0059813f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_12 VNB N_VGND_c_41_n 0.0128263f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0
cc_13 VNB N_VPWR_c_71_n 0.00208207f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.085
cc_14 VNB N_VPWR_c_72_n 0.32452f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.64
cc_15 VNB N_VPWR_c_73_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0
cc_16 VPB N_VGND_M1000_g 0.0989297f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=2.46
cc_17 VPB N_VGND_M1002_g 0.0927777f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.46
cc_18 VPB N_VGND_c_32_n 0.0193702f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.42
cc_19 VPB N_VGND_c_35_n 0.0189219f $X=-0.19 $Y=1.66 $X2=2.52 $Y2=1.42
cc_20 VPB N_VPWR_c_74_n 0.0113726f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.83
cc_21 VPB N_VPWR_c_75_n 0.056103f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=2.46
cc_22 VPB N_VPWR_c_76_n 0.0225322f $X=-0.19 $Y=1.66 $X2=2.185 $Y2=2.46
cc_23 VPB N_VPWR_c_71_n 0.00778682f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=0.085
cc_24 VPB N_VPWR_c_78_n 0.0519987f $X=-0.19 $Y=1.66 $X2=1.615 $Y2=0.64
cc_25 VPB N_VPWR_c_79_n 0.0180771f $X=-0.19 $Y=1.66 $X2=2.705 $Y2=1.42
cc_26 VPB N_VPWR_c_80_n 0.00613202f $X=-0.19 $Y=1.66 $X2=2.52 $Y2=1.42
cc_27 VPB N_VPWR_c_81_n 0.029192f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0
cc_28 VPB N_VPWR_c_73_n 0.0749347f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=0
cc_29 VPB N_VPWR_c_83_n 0.017094f $X=-0.19 $Y=1.66 $X2=3.6 $Y2=0
cc_30 N_VGND_M1000_g N_VPWR_c_75_n 0.0605103f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_31 N_VGND_c_31_n N_VPWR_c_75_n 0.0143348f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_32 N_VGND_M1000_g N_VPWR_c_76_n 0.0221223f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_33 N_VGND_M1000_g N_VPWR_c_71_n 0.107807f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_34 N_VGND_M1002_g N_VPWR_c_71_n 0.0975598f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_35 N_VGND_c_31_n N_VPWR_c_71_n 0.0138086f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_36 N_VGND_c_32_n N_VPWR_c_71_n 0.00993466f $X=0.575 $Y=1.42 $X2=0 $Y2=0
cc_37 N_VGND_c_33_n N_VPWR_c_71_n 0.0108665f $X=1.615 $Y=0.64 $X2=0 $Y2=0
cc_38 N_VGND_c_34_n N_VPWR_c_71_n 0.0189017f $X=2.89 $Y=0.64 $X2=0 $Y2=0
cc_39 N_VGND_c_35_n N_VPWR_c_71_n 0.0111522f $X=2.52 $Y=1.42 $X2=0 $Y2=0
cc_40 N_VGND_M1000_g N_VPWR_c_72_n 0.0139884f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_41 N_VGND_M1002_g N_VPWR_c_72_n 0.0208415f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_42 N_VGND_c_31_n N_VPWR_c_72_n 0.0861076f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_43 N_VGND_c_32_n N_VPWR_c_72_n 0.0267831f $X=0.575 $Y=1.42 $X2=0 $Y2=0
cc_44 N_VGND_c_33_n N_VPWR_c_72_n 0.0538668f $X=1.615 $Y=0.64 $X2=0 $Y2=0
cc_45 N_VGND_c_34_n N_VPWR_c_72_n 0.087653f $X=2.89 $Y=0.64 $X2=0 $Y2=0
cc_46 N_VGND_c_35_n N_VPWR_c_72_n 0.0367272f $X=2.52 $Y=1.42 $X2=0 $Y2=0
cc_47 N_VGND_c_36_n N_VPWR_c_72_n 0.0220076f $X=1.45 $Y=0 $X2=0 $Y2=0
cc_48 N_VGND_c_37_n N_VPWR_c_72_n 0.0178177f $X=2.355 $Y=0 $X2=0 $Y2=0
cc_49 N_VGND_c_39_n N_VPWR_c_72_n 0.0776326f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_50 N_VGND_M1002_g N_VPWR_c_78_n 0.0365849f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_51 N_VGND_c_34_n N_VPWR_c_78_n 0.0179872f $X=2.89 $Y=0.64 $X2=0 $Y2=0
cc_52 N_VGND_M1002_g N_VPWR_c_79_n 0.0178153f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_53 N_VGND_M1000_g N_VPWR_c_73_n 0.0434015f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_54 N_VGND_M1002_g N_VPWR_c_73_n 0.0349716f $X=2.185 $Y=2.46 $X2=0 $Y2=0

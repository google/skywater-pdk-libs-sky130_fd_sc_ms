* File: sky130_fd_sc_ms__and3b_1.spice
* Created: Fri Aug 28 17:12:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and3b_1.pex.spice"
.subckt sky130_fd_sc_ms__and3b_1  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_A_114_74#_M1006_d N_A_N_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.19525 AS=0.15675 PD=1.81 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1004 A_353_94# N_A_114_74#_M1004_g N_A_266_94#_M1004_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 A_431_94# N_B_M1005_g A_353_94# VNB NLOWVT L=0.15 W=0.64 AD=0.1248
+ AS=0.0768 PD=1.03 PS=0.88 NRD=26.244 NRS=12.18 M=1 R=4.26667 SA=75000.6
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g A_431_94# VNB NLOWVT L=0.15 W=0.64 AD=0.184162
+ AS=0.1248 PD=1.21043 PS=1.03 NRD=27.18 NRS=26.244 M=1 R=4.26667 SA=75001.1
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_266_94#_M1003_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.212938 PD=2.05 PS=1.39957 NRD=0 NRS=23.1 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_114_74#_M1002_d N_A_N_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.273 AS=0.2394 PD=2.33 PS=2.25 NRD=9.3772 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1009 N_VPWR_M1009_d N_A_114_74#_M1009_g N_A_266_94#_M1009_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1533 AS=0.2352 PD=1.205 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1000 N_A_266_94#_M1000_d N_B_M1000_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1155 AS=0.1533 PD=1.115 PS=1.205 NRD=0 NRS=9.3772 M=1 R=4.66667
+ SA=90000.7 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1008_d N_C_M1008_g N_A_266_94#_M1000_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1854 AS=0.1155 PD=1.30714 PS=1.115 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90001.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1001 N_X_M1001_d N_A_266_94#_M1001_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2472 PD=2.8 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__and3b_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand4_4.spice
* Created: Wed Sep  2 12:14:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4_4.pex.spice"
.subckt sky130_fd_sc_ms__nand4_4  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_M1006_g N_A_27_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1006_d N_D_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1295 PD=1.29 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1014_d N_D_M1019_g N_A_27_74#_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1295 PD=1.29 PS=1.09 NRD=32.424 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1001 N_A_554_74#_M1001_d N_C_M1001_g N_A_27_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.4 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1010 N_A_554_74#_M1001_d N_C_M1010_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75001 A=0.111 P=1.78 MULT=1
MM1011 N_A_554_74#_M1011_d N_C_M1011_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1020 N_A_554_74#_M1011_d N_C_M1020_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.19515 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_923_74#_M1003_d N_B_M1003_g N_A_554_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1969 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1004 N_A_923_74#_M1004_d N_B_M1004_g N_A_554_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1016 N_A_923_74#_M1004_d N_B_M1016_g N_A_554_74#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1021 N_A_923_74#_M1021_d N_B_M1021_g N_A_554_74#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_A_923_74#_M1021_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1002_d N_A_M1012_g N_A_923_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1015_d N_A_M1015_g N_A_923_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1628 AS=0.1036 PD=1.18 PS=1.02 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1023 N_Y_M1015_d N_A_M1023_g N_A_923_74#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1628 AS=0.1962 PD=1.18 PS=2.05 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_D_M1005_g N_Y_M1005_s VPB PSHORT L=0.18 W=1.12 AD=1.7192
+ AS=0.1792 PD=5.31 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.4 SB=90006.6
+ A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_D_M1007_g N_Y_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.9 SB=90006.1
+ A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_C_M1009_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1.12 AD=0.364
+ AS=0.1512 PD=1.77 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4 SB=90005.6
+ A=0.2016 P=2.6 MULT=1
MM1018 N_Y_M1009_d N_C_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12 AD=0.364
+ AS=0.4704 PD=1.77 PS=1.96 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2 SB=90004.8
+ A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1018_s N_B_M1000_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.4704
+ AS=0.364 PD=1.96 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2 SB=90003.8
+ A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1017_d N_B_M1017_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.9128
+ AS=0.364 PD=2.75 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.1 SB=90002.9
+ A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1017_d N_A_M1013_g N_Y_M1013_s VPB PSHORT L=0.18 W=1.12 AD=0.9128
+ AS=0.42 PD=2.75 PS=1.87 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.9 SB=90001.1
+ A=0.2016 P=2.6 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_Y_M1013_s VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.42 PD=2.8 PS=1.87 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.8 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__nand4_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor4bb_1.pxi.spice
* Created: Wed Sep  2 12:17:17 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4BB_1%C_N N_C_N_M1006_g N_C_N_c_77_n N_C_N_M1003_g C_N
+ N_C_N_c_79_n PM_SKY130_FD_SC_MS__NOR4BB_1%C_N
x_PM_SKY130_FD_SC_MS__NOR4BB_1%A N_A_M1010_g N_A_M1011_g A A N_A_c_103_n
+ N_A_c_104_n PM_SKY130_FD_SC_MS__NOR4BB_1%A
x_PM_SKY130_FD_SC_MS__NOR4BB_1%B N_B_M1009_g N_B_M1001_g B N_B_c_145_n
+ N_B_c_146_n PM_SKY130_FD_SC_MS__NOR4BB_1%B
x_PM_SKY130_FD_SC_MS__NOR4BB_1%A_27_112# N_A_27_112#_M1003_s N_A_27_112#_M1006_s
+ N_A_27_112#_M1002_g N_A_27_112#_M1008_g N_A_27_112#_c_181_n
+ N_A_27_112#_c_186_n N_A_27_112#_c_182_n N_A_27_112#_c_183_n
+ N_A_27_112#_c_189_n N_A_27_112#_c_190_n N_A_27_112#_c_191_n
+ N_A_27_112#_c_192_n N_A_27_112#_c_184_n PM_SKY130_FD_SC_MS__NOR4BB_1%A_27_112#
x_PM_SKY130_FD_SC_MS__NOR4BB_1%A_611_244# N_A_611_244#_M1004_d
+ N_A_611_244#_M1000_d N_A_611_244#_M1005_g N_A_611_244#_c_283_n
+ N_A_611_244#_M1007_g N_A_611_244#_c_292_n N_A_611_244#_c_293_n
+ N_A_611_244#_c_284_n N_A_611_244#_c_285_n N_A_611_244#_c_286_n
+ N_A_611_244#_c_295_n N_A_611_244#_c_309_n N_A_611_244#_c_287_n
+ N_A_611_244#_c_288_n N_A_611_244#_c_289_n N_A_611_244#_c_290_n
+ PM_SKY130_FD_SC_MS__NOR4BB_1%A_611_244#
x_PM_SKY130_FD_SC_MS__NOR4BB_1%D_N N_D_N_c_357_n N_D_N_M1000_g N_D_N_M1004_g D_N
+ N_D_N_c_359_n PM_SKY130_FD_SC_MS__NOR4BB_1%D_N
x_PM_SKY130_FD_SC_MS__NOR4BB_1%VPWR N_VPWR_M1006_d N_VPWR_M1000_s N_VPWR_c_391_n
+ VPWR N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_390_n N_VPWR_c_395_n
+ N_VPWR_c_396_n N_VPWR_c_397_n PM_SKY130_FD_SC_MS__NOR4BB_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR4BB_1%Y N_Y_M1010_d N_Y_M1008_d N_Y_M1005_d N_Y_c_440_n
+ N_Y_c_441_n N_Y_c_450_n N_Y_c_457_n N_Y_c_460_n N_Y_c_442_n Y N_Y_c_443_n
+ PM_SKY130_FD_SC_MS__NOR4BB_1%Y
x_PM_SKY130_FD_SC_MS__NOR4BB_1%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1007_d
+ N_VGND_c_501_n N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n VGND
+ N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n PM_SKY130_FD_SC_MS__NOR4BB_1%VGND
cc_1 VNB N_C_N_M1006_g 0.00451142f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_2 VNB N_C_N_c_77_n 0.0235244f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.22
cc_3 VNB C_N 0.00873016f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_C_N_c_79_n 0.0913571f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.415
cc_5 VNB N_A_M1010_g 0.0275783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_6 VNB N_A_c_103_n 0.00391014f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_7 VNB N_A_c_104_n 0.0360382f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_8 VNB N_B_M1009_g 0.0292581f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_9 VNB N_B_c_145_n 0.0309745f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_10 VNB N_B_c_146_n 0.00558343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_112#_M1008_g 0.0288172f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.415
cc_12 VNB N_A_27_112#_c_181_n 0.013952f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_A_27_112#_c_182_n 0.00208657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_112#_c_183_n 0.0270426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_112#_c_184_n 0.00361275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_611_244#_M1005_g 0.00446323f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.415
cc_17 VNB N_A_611_244#_c_283_n 0.0193467f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_18 VNB N_A_611_244#_c_284_n 0.0042639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_611_244#_c_285_n 0.00913271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_611_244#_c_286_n 0.0244614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_611_244#_c_287_n 0.00488535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_611_244#_c_288_n 0.0130414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_611_244#_c_289_n 0.0186936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_611_244#_c_290_n 0.057011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_D_N_c_357_n 0.0212192f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.61
cc_26 VNB N_D_N_M1004_g 0.0388469f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.835
cc_27 VNB N_D_N_c_359_n 0.00237576f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.415
cc_28 VNB N_VPWR_c_390_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_440_n 0.00280366f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_30 VNB N_Y_c_441_n 0.00582747f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_31 VNB N_Y_c_442_n 0.00264733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_443_n 0.00280529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_501_n 0.0233407f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_34 VNB N_VGND_c_502_n 0.0223553f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_35 VNB N_VGND_c_503_n 0.0295327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_504_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_505_n 0.0196163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_506_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_507_n 0.284156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_508_n 0.0185359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_509_n 0.0209009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_510_n 0.0148108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_C_N_M1006_g 0.0343084f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_44 VPB N_A_M1011_g 0.0231517f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.835
cc_45 VPB N_A_c_103_n 0.00139833f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_46 VPB N_A_c_104_n 0.0110892f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_47 VPB N_B_M1001_g 0.0235869f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.835
cc_48 VPB N_B_c_145_n 0.00849549f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_49 VPB N_B_c_146_n 0.00388201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_112#_M1002_g 0.024062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_27_112#_c_186_n 0.00394542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_112#_c_182_n 4.28226e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_112#_c_183_n 0.0056692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_112#_c_189_n 0.010553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_112#_c_190_n 0.00135146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_112#_c_191_n 0.00560699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_112#_c_192_n 0.0450155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_27_112#_c_184_n 0.00287517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_611_244#_M1005_g 0.0130714f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.415
cc_60 VPB N_A_611_244#_c_292_n 0.0339844f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.415
cc_61 VPB N_A_611_244#_c_293_n 0.0135162f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_62 VPB N_A_611_244#_c_284_n 0.0744494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_611_244#_c_295_n 0.0413842f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_611_244#_c_289_n 0.0209422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_D_N_c_357_n 0.0208485f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.61
cc_66 VPB N_D_N_M1000_g 0.0354979f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_67 VPB N_D_N_c_359_n 0.00161194f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.415
cc_68 VPB N_VPWR_c_391_n 0.0110663f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_69 VPB N_VPWR_c_392_n 0.0716443f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_70 VPB N_VPWR_c_393_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_390_n 0.0737493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_395_n 0.020284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_396_n 0.0297497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_397_n 0.00420575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_Y_c_441_n 0.00124557f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_76 N_C_N_c_77_n N_A_M1010_g 0.0167728f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_77 N_C_N_M1006_g N_A_c_103_n 0.00159301f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_78 N_C_N_c_79_n N_A_c_103_n 0.00112291f $X=0.505 $Y=1.415 $X2=0 $Y2=0
cc_79 N_C_N_M1006_g N_A_c_104_n 0.00127442f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_80 N_C_N_c_79_n N_A_c_104_n 0.0147979f $X=0.505 $Y=1.415 $X2=0 $Y2=0
cc_81 N_C_N_c_77_n N_A_27_112#_c_181_n 0.00666781f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_82 C_N N_A_27_112#_c_181_n 0.0264607f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_C_N_c_79_n N_A_27_112#_c_181_n 0.00933251f $X=0.505 $Y=1.415 $X2=0 $Y2=0
cc_84 N_C_N_M1006_g N_A_27_112#_c_186_n 8.08616e-19 $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_85 N_C_N_M1006_g N_A_27_112#_c_192_n 0.0473123f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_86 C_N N_A_27_112#_c_192_n 0.0191168f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_C_N_c_79_n N_A_27_112#_c_192_n 0.00267027f $X=0.505 $Y=1.415 $X2=0 $Y2=0
cc_88 N_C_N_M1006_g N_A_27_112#_c_184_n 0.00777797f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_89 N_C_N_c_77_n N_A_27_112#_c_184_n 0.00678818f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_90 C_N N_A_27_112#_c_184_n 0.0267372f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_91 N_C_N_c_79_n N_A_27_112#_c_184_n 0.0234888f $X=0.505 $Y=1.415 $X2=0 $Y2=0
cc_92 N_C_N_M1006_g N_VPWR_c_390_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_93 N_C_N_M1006_g N_VPWR_c_395_n 0.00371318f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_94 N_C_N_c_77_n N_VGND_c_501_n 0.0108888f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_95 N_C_N_c_77_n N_VGND_c_503_n 0.00390814f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_96 N_C_N_c_77_n N_VGND_c_507_n 0.00487769f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_97 N_A_M1010_g N_B_M1009_g 0.0212654f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A_M1011_g N_B_M1001_g 0.0473963f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_c_103_n N_B_M1001_g 2.55823e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_c_104_n N_B_c_145_n 0.0473963f $X=1.49 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A_c_104_n N_B_c_146_n 3.48537e-19 $X=1.49 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A_M1011_g N_A_27_112#_c_186_n 0.0195579f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_c_103_n N_A_27_112#_c_186_n 0.0114805f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A_M1011_g N_A_27_112#_c_192_n 0.0109123f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_M1010_g N_A_27_112#_c_184_n 0.00110337f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_M1011_g N_A_27_112#_c_184_n 0.00184987f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_c_103_n N_A_27_112#_c_184_n 0.0411461f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_c_104_n N_A_27_112#_c_184_n 0.00153543f $X=1.49 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A_c_103_n N_VPWR_M1006_d 0.0106395f $X=1.24 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_M1011_g N_VPWR_c_392_n 0.00386841f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_M1011_g N_VPWR_c_390_n 0.00488949f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_M1011_g N_VPWR_c_396_n 0.00723585f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_M1010_g N_Y_c_440_n 0.00670807f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_M1010_g N_Y_c_441_n 0.00508657f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_M1011_g N_Y_c_441_n 0.00787961f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A_c_103_n N_Y_c_441_n 0.0505976f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A_c_104_n N_Y_c_441_n 0.00687902f $X=1.49 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_M1011_g N_Y_c_450_n 0.0157443f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_c_103_n N_Y_c_450_n 0.00718422f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A_M1010_g N_Y_c_442_n 0.0041358f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_c_104_n N_Y_c_442_n 0.00481434f $X=1.49 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_M1010_g N_VGND_c_501_n 0.00970997f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_c_103_n N_VGND_c_501_n 0.0145292f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_c_104_n N_VGND_c_501_n 0.00151797f $X=1.49 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_M1010_g N_VGND_c_507_n 0.00825771f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_M1010_g N_VGND_c_508_n 0.00434272f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_M1010_g N_VGND_c_509_n 4.31196e-19 $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B_M1001_g N_A_27_112#_M1002_g 0.0365044f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B_c_146_n N_A_27_112#_M1002_g 2.55051e-19 $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_130 N_B_M1009_g N_A_27_112#_M1008_g 0.0132106f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B_M1001_g N_A_27_112#_c_186_n 0.0135959f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_132 N_B_c_145_n N_A_27_112#_c_182_n 3.9721e-19 $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_133 N_B_c_146_n N_A_27_112#_c_182_n 0.0251141f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_134 N_B_c_145_n N_A_27_112#_c_183_n 0.0175372f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B_c_146_n N_A_27_112#_c_183_n 0.00234681f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B_M1001_g N_A_27_112#_c_190_n 6.58171e-19 $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_137 N_B_c_146_n N_A_27_112#_c_190_n 0.0043213f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B_M1001_g N_VPWR_c_392_n 0.00386841f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_139 N_B_M1001_g N_VPWR_c_390_n 0.00486632f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B_M1009_g N_Y_c_440_n 0.00282538f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_141 N_B_M1009_g N_Y_c_441_n 0.0146597f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_142 N_B_c_146_n N_Y_c_441_n 0.0324918f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B_M1001_g N_Y_c_457_n 0.0232545f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_144 N_B_c_145_n N_Y_c_457_n 0.00120831f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_145 N_B_c_146_n N_Y_c_457_n 0.0187993f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_146 N_B_M1009_g N_Y_c_460_n 0.019134f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_147 N_B_c_145_n N_Y_c_460_n 0.00155436f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B_c_146_n N_Y_c_460_n 0.0161271f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_149 N_B_M1009_g N_Y_c_442_n 8.5887e-19 $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_150 N_B_M1009_g N_VGND_c_507_n 0.00753637f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B_M1009_g N_VGND_c_508_n 0.00383152f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_152 N_B_M1009_g N_VGND_c_509_n 0.00911669f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_27_112#_M1002_g N_A_611_244#_M1005_g 0.0480209f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_154 N_A_27_112#_c_186_n N_A_611_244#_M1005_g 0.0140727f $X=3.625 $Y=2.645
+ $X2=0 $Y2=0
cc_155 N_A_27_112#_c_182_n N_A_611_244#_M1005_g 8.93789e-19 $X=2.65 $Y=1.515
+ $X2=0 $Y2=0
cc_156 N_A_27_112#_c_183_n N_A_611_244#_M1005_g 0.0132769f $X=2.65 $Y=1.515
+ $X2=0 $Y2=0
cc_157 N_A_27_112#_c_189_n N_A_611_244#_M1005_g 0.0128629f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_158 N_A_27_112#_c_191_n N_A_611_244#_M1005_g 0.00176916f $X=3.71 $Y=2.56
+ $X2=0 $Y2=0
cc_159 N_A_27_112#_M1008_g N_A_611_244#_c_283_n 0.0198165f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_27_112#_c_186_n N_A_611_244#_c_292_n 0.00335276f $X=3.625 $Y=2.645
+ $X2=0 $Y2=0
cc_161 N_A_27_112#_c_186_n N_A_611_244#_c_284_n 0.010379f $X=3.625 $Y=2.645
+ $X2=0 $Y2=0
cc_162 N_A_27_112#_c_189_n N_A_611_244#_c_284_n 0.0090941f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_163 N_A_27_112#_c_191_n N_A_611_244#_c_284_n 0.0193753f $X=3.71 $Y=2.56 $X2=0
+ $Y2=0
cc_164 N_A_27_112#_c_189_n N_A_611_244#_c_285_n 0.00230969f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_165 N_A_27_112#_M1008_g N_A_611_244#_c_309_n 0.00151227f $X=2.74 $Y=0.74
+ $X2=0 $Y2=0
cc_166 N_A_27_112#_c_182_n N_A_611_244#_c_309_n 0.0114575f $X=2.65 $Y=1.515
+ $X2=0 $Y2=0
cc_167 N_A_27_112#_c_189_n N_A_611_244#_c_309_n 0.0410022f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_168 N_A_27_112#_c_189_n N_A_611_244#_c_287_n 0.0094058f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_169 N_A_27_112#_M1008_g N_A_611_244#_c_290_n 0.0132769f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_27_112#_c_182_n N_A_611_244#_c_290_n 0.00179414f $X=2.65 $Y=1.515
+ $X2=0 $Y2=0
cc_171 N_A_27_112#_c_189_n N_A_611_244#_c_290_n 0.0039236f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_172 N_A_27_112#_c_189_n N_D_N_c_357_n 0.00265493f $X=3.625 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_27_112#_c_191_n N_D_N_M1000_g 0.00418814f $X=3.71 $Y=2.56 $X2=0 $Y2=0
cc_174 N_A_27_112#_c_189_n N_D_N_c_359_n 0.00529505f $X=3.625 $Y=1.805 $X2=0
+ $Y2=0
cc_175 N_A_27_112#_c_186_n N_VPWR_M1006_d 0.0261396f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_27_112#_c_192_n N_VPWR_M1006_d 0.0139014f $X=0.28 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A_27_112#_c_186_n N_VPWR_c_391_n 0.0143757f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_178 N_A_27_112#_c_191_n N_VPWR_c_391_n 0.0346721f $X=3.71 $Y=2.56 $X2=0 $Y2=0
cc_179 N_A_27_112#_M1002_g N_VPWR_c_392_n 0.00386841f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_180 N_A_27_112#_c_186_n N_VPWR_c_392_n 0.0419797f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_181 N_A_27_112#_M1002_g N_VPWR_c_390_n 0.00487954f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_182 N_A_27_112#_c_186_n N_VPWR_c_390_n 0.0691461f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_183 N_A_27_112#_c_192_n N_VPWR_c_390_n 0.0170891f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_27_112#_c_192_n N_VPWR_c_395_n 0.0112128f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_27_112#_c_186_n N_VPWR_c_396_n 0.0425745f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_186 N_A_27_112#_c_192_n N_VPWR_c_396_n 0.0103275f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_27_112#_c_186_n A_316_368# 0.00343313f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_27_112#_c_186_n A_400_368# 0.0113106f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_27_112#_c_186_n A_533_368# 0.00782857f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_27_112#_c_189_n A_533_368# 0.00198757f $X=3.625 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_191 N_A_27_112#_c_190_n A_533_368# 0.00101345f $X=2.815 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_27_112#_c_186_n N_Y_M1005_d 0.00599241f $X=3.625 $Y=2.645 $X2=0 $Y2=0
cc_193 N_A_27_112#_c_189_n N_Y_M1005_d 0.00293923f $X=3.625 $Y=1.805 $X2=0 $Y2=0
cc_194 N_A_27_112#_c_186_n N_Y_c_450_n 0.00908059f $X=3.625 $Y=2.645 $X2=0 $Y2=0
cc_195 N_A_27_112#_M1002_g N_Y_c_457_n 0.0212232f $X=2.575 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_27_112#_c_186_n N_Y_c_457_n 0.101691f $X=3.625 $Y=2.645 $X2=0 $Y2=0
cc_197 N_A_27_112#_c_183_n N_Y_c_457_n 5.73996e-19 $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A_27_112#_c_189_n N_Y_c_457_n 0.0392224f $X=3.625 $Y=1.805 $X2=0 $Y2=0
cc_199 N_A_27_112#_c_190_n N_Y_c_457_n 0.0218101f $X=2.815 $Y=1.805 $X2=0 $Y2=0
cc_200 N_A_27_112#_c_191_n N_Y_c_457_n 0.0258892f $X=3.71 $Y=2.56 $X2=0 $Y2=0
cc_201 N_A_27_112#_M1008_g N_Y_c_460_n 0.0166532f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_27_112#_c_182_n N_Y_c_460_n 0.0145929f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A_27_112#_c_183_n N_Y_c_460_n 9.4439e-19 $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_204 N_A_27_112#_c_189_n N_Y_c_460_n 0.00614593f $X=3.625 $Y=1.805 $X2=0 $Y2=0
cc_205 N_A_27_112#_M1008_g N_Y_c_443_n 0.00282724f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_27_112#_c_181_n N_VGND_c_501_n 0.0271305f $X=0.605 $Y=0.845 $X2=0
+ $Y2=0
cc_207 N_A_27_112#_c_184_n N_VGND_c_501_n 0.00887541f $X=0.445 $Y=1.82 $X2=0
+ $Y2=0
cc_208 N_A_27_112#_c_181_n N_VGND_c_503_n 0.0104931f $X=0.605 $Y=0.845 $X2=0
+ $Y2=0
cc_209 N_A_27_112#_M1008_g N_VGND_c_505_n 0.00383152f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_27_112#_M1008_g N_VGND_c_507_n 0.00753637f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_211 N_A_27_112#_c_181_n N_VGND_c_507_n 0.0187574f $X=0.605 $Y=0.845 $X2=0
+ $Y2=0
cc_212 N_A_27_112#_M1008_g N_VGND_c_509_n 0.00923995f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_611_244#_c_284_n N_D_N_c_357_n 0.00982666f $X=3.665 $Y=3.035
+ $X2=-0.19 $Y2=-0.245
cc_214 N_A_611_244#_c_285_n N_D_N_c_357_n 0.00485457f $X=4.355 $Y=1.175
+ $X2=-0.19 $Y2=-0.245
cc_215 N_A_611_244#_c_289_n N_D_N_c_357_n 0.00983751f $X=4.52 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_611_244#_c_290_n N_D_N_c_357_n 0.0150445f $X=3.665 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_611_244#_c_292_n N_D_N_M1000_g 0.00982666f $X=3.59 $Y=3.11 $X2=0
+ $Y2=0
cc_218 N_A_611_244#_c_295_n N_D_N_M1000_g 0.0158442f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_219 N_A_611_244#_c_285_n N_D_N_M1004_g 0.0130612f $X=4.355 $Y=1.175 $X2=0
+ $Y2=0
cc_220 N_A_611_244#_c_286_n N_D_N_M1004_g 0.0150412f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_221 N_A_611_244#_c_287_n N_D_N_M1004_g 0.00101533f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_222 N_A_611_244#_c_288_n N_D_N_M1004_g 0.00508894f $X=4.52 $Y=1.175 $X2=0
+ $Y2=0
cc_223 N_A_611_244#_c_289_n N_D_N_M1004_g 0.0128589f $X=4.52 $Y=2.1 $X2=0 $Y2=0
cc_224 N_A_611_244#_c_290_n N_D_N_M1004_g 0.00455351f $X=3.665 $Y=1.385 $X2=0
+ $Y2=0
cc_225 N_A_611_244#_c_285_n N_D_N_c_359_n 0.0260399f $X=4.355 $Y=1.175 $X2=0
+ $Y2=0
cc_226 N_A_611_244#_c_287_n N_D_N_c_359_n 0.00674841f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_227 N_A_611_244#_c_289_n N_D_N_c_359_n 0.0250404f $X=4.52 $Y=2.1 $X2=0 $Y2=0
cc_228 N_A_611_244#_c_290_n N_D_N_c_359_n 0.00435647f $X=3.665 $Y=1.385 $X2=0
+ $Y2=0
cc_229 N_A_611_244#_c_284_n N_VPWR_c_391_n 0.0128698f $X=3.665 $Y=3.035 $X2=0
+ $Y2=0
cc_230 N_A_611_244#_c_295_n N_VPWR_c_391_n 0.0344689f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_231 N_A_611_244#_c_293_n N_VPWR_c_392_n 0.0170709f $X=3.235 $Y=3.11 $X2=0
+ $Y2=0
cc_232 N_A_611_244#_c_295_n N_VPWR_c_393_n 0.014549f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_233 N_A_611_244#_c_292_n N_VPWR_c_390_n 0.0156334f $X=3.59 $Y=3.11 $X2=0
+ $Y2=0
cc_234 N_A_611_244#_c_293_n N_VPWR_c_390_n 0.00675631f $X=3.235 $Y=3.11 $X2=0
+ $Y2=0
cc_235 N_A_611_244#_c_295_n N_VPWR_c_390_n 0.0119743f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_236 N_A_611_244#_M1005_g N_Y_c_457_n 0.0155199f $X=3.145 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_611_244#_c_284_n N_Y_c_457_n 0.00252041f $X=3.665 $Y=3.035 $X2=0
+ $Y2=0
cc_238 N_A_611_244#_c_283_n N_Y_c_460_n 0.00812308f $X=3.24 $Y=1.22 $X2=0 $Y2=0
cc_239 N_A_611_244#_c_309_n N_Y_c_460_n 0.0108526f $X=3.575 $Y=1.385 $X2=0 $Y2=0
cc_240 N_A_611_244#_c_290_n N_Y_c_460_n 0.00292421f $X=3.665 $Y=1.385 $X2=0
+ $Y2=0
cc_241 N_A_611_244#_c_283_n N_Y_c_443_n 0.00814444f $X=3.24 $Y=1.22 $X2=0 $Y2=0
cc_242 N_A_611_244#_c_285_n N_VGND_M1007_d 0.00472896f $X=4.355 $Y=1.175 $X2=0
+ $Y2=0
cc_243 N_A_611_244#_c_287_n N_VGND_M1007_d 0.00214094f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_244 N_A_611_244#_c_283_n N_VGND_c_502_n 0.0174322f $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_245 N_A_611_244#_c_286_n N_VGND_c_502_n 0.0144669f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_246 N_A_611_244#_c_309_n N_VGND_c_502_n 0.00873167f $X=3.575 $Y=1.385 $X2=0
+ $Y2=0
cc_247 N_A_611_244#_c_287_n N_VGND_c_502_n 0.0500172f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_248 N_A_611_244#_c_290_n N_VGND_c_502_n 0.00475493f $X=3.665 $Y=1.385 $X2=0
+ $Y2=0
cc_249 N_A_611_244#_c_283_n N_VGND_c_505_n 0.00383287f $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_250 N_A_611_244#_c_286_n N_VGND_c_506_n 0.00816527f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_251 N_A_611_244#_c_283_n N_VGND_c_507_n 0.00661688f $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_252 N_A_611_244#_c_286_n N_VGND_c_507_n 0.0106525f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_253 N_A_611_244#_c_283_n N_VGND_c_509_n 6.14575e-19 $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_254 N_D_N_c_357_n N_VPWR_c_391_n 0.0036051f $X=4.295 $Y=1.87 $X2=0 $Y2=0
cc_255 N_D_N_M1000_g N_VPWR_c_391_n 0.00472663f $X=4.295 $Y=2.54 $X2=0 $Y2=0
cc_256 N_D_N_c_359_n N_VPWR_c_391_n 0.0116968f $X=4.18 $Y=1.615 $X2=0 $Y2=0
cc_257 N_D_N_M1000_g N_VPWR_c_393_n 0.005209f $X=4.295 $Y=2.54 $X2=0 $Y2=0
cc_258 N_D_N_M1000_g N_VPWR_c_390_n 0.00987012f $X=4.295 $Y=2.54 $X2=0 $Y2=0
cc_259 N_D_N_M1004_g N_VGND_c_502_n 0.0124771f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_260 N_D_N_M1004_g N_VGND_c_506_n 0.0043356f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_261 N_D_N_M1004_g N_VGND_c_507_n 0.00487769f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_262 A_316_368# N_Y_c_441_n 0.00241994f $X=1.58 $Y=1.84 $X2=0.605 $Y2=0.845
cc_263 A_316_368# N_Y_c_450_n 0.001187f $X=1.58 $Y=1.84 $X2=0.545 $Y2=0.845
cc_264 A_316_368# N_Y_c_457_n 8.87649e-19 $X=1.58 $Y=1.84 $X2=0.69 $Y2=1.01
cc_265 A_400_368# N_Y_c_457_n 0.0152057f $X=2 $Y=1.84 $X2=0.69 $Y2=1.01
cc_266 A_533_368# N_Y_c_457_n 0.00638731f $X=2.665 $Y=1.84 $X2=0.69 $Y2=1.01
cc_267 N_Y_c_460_n N_VGND_M1009_d 0.0220163f $X=2.86 $Y=0.965 $X2=0 $Y2=0
cc_268 N_Y_c_440_n N_VGND_c_501_n 0.0206398f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_269 N_Y_c_442_n N_VGND_c_501_n 0.0109738f $X=1.61 $Y=0.965 $X2=0 $Y2=0
cc_270 N_Y_c_460_n N_VGND_c_502_n 0.00348012f $X=2.86 $Y=0.965 $X2=0 $Y2=0
cc_271 N_Y_c_443_n N_VGND_c_502_n 0.0439579f $X=3.025 $Y=0.515 $X2=0 $Y2=0
cc_272 N_Y_c_443_n N_VGND_c_505_n 0.0164719f $X=3.025 $Y=0.515 $X2=0 $Y2=0
cc_273 N_Y_c_440_n N_VGND_c_507_n 0.0119984f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_274 N_Y_c_443_n N_VGND_c_507_n 0.013457f $X=3.025 $Y=0.515 $X2=0 $Y2=0
cc_275 N_Y_c_440_n N_VGND_c_508_n 0.0145639f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_276 N_Y_c_440_n N_VGND_c_509_n 0.0146527f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_277 N_Y_c_460_n N_VGND_c_509_n 0.0449771f $X=2.86 $Y=0.965 $X2=0 $Y2=0
cc_278 N_Y_c_443_n N_VGND_c_509_n 0.0146682f $X=3.025 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__or3_4.pex.spice
* Created: Fri Aug 28 18:07:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR3_4%A 3 7 11 14 15 17 19 23 25 35 39 43
c89 43 0 1.22748e-19 $X=0.24 $Y=1.295
c90 19 0 1.25197e-19 $X=2.905 $Y=1.195
c91 7 0 6.61072e-20 $X=2.89 $Y=2.44
c92 3 0 8.47394e-20 $X=0.505 $Y=2.44
r93 41 43 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.27 $Y=1.28
+ $X2=0.27 $Y2=1.295
r94 35 37 40.5227 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.35 $Y=1.465
+ $X2=0.35 $Y2=1.63
r95 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r96 28 35 8.73518 $w=4.9e-07 $l=8e-08 $layer=POLY_cond $X=0.35 $Y=1.385 $X2=0.35
+ $Y2=1.465
r97 28 32 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=0.35 $Y=1.385
+ $X2=0.35 $Y2=1.125
r98 25 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.195
+ $X2=0.27 $Y2=1.28
r99 25 36 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.27 $Y=1.33
+ $X2=0.27 $Y2=1.465
r100 25 43 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.27 $Y=1.33
+ $X2=0.27 $Y2=1.295
r101 25 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.125 $X2=0.27 $Y2=1.125
r102 23 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.385
+ $X2=2.92 $Y2=1.55
r103 23 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.385
+ $X2=2.92 $Y2=1.22
r104 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.92
+ $Y=1.385 $X2=2.92 $Y2=1.385
r105 19 22 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=2.905 $Y=1.195
+ $X2=2.905 $Y2=1.385
r106 18 25 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=1.195
+ $X2=0.27 $Y2=1.195
r107 17 19 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.755 $Y=1.195
+ $X2=2.905 $Y2=1.195
r108 17 18 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=2.755 $Y=1.195
+ $X2=0.435 $Y2=1.195
r109 15 32 74.249 $w=4.9e-07 $l=6.8e-07 $layer=POLY_cond $X=0.35 $Y=0.445
+ $X2=0.35 $Y2=1.125
r110 14 15 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.445 $X2=0.27 $Y2=0.445
r111 12 25 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=1.195
r112 12 14 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=0.445
r113 11 39 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.93 $Y=0.74
+ $X2=2.93 $Y2=1.22
r114 7 40 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.89 $Y=2.44
+ $X2=2.89 $Y2=1.55
r115 3 37 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=0.505 $Y=2.44
+ $X2=0.505 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%B 3 7 11 13 14 15 16 22 27 28
c58 27 0 1.25197e-19 $X=2.38 $Y=1.615
c59 22 0 3.14127e-19 $X=0.97 $Y=1.615
c60 7 0 1.92271e-19 $X=2.39 $Y=2.44
c61 3 0 1.71217e-19 $X=0.955 $Y=2.44
r62 27 30 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.615
+ $X2=2.38 $Y2=1.78
r63 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.615
+ $X2=2.38 $Y2=1.45
r64 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.615 $X2=2.38 $Y2=1.615
r65 22 25 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.615
+ $X2=0.97 $Y2=1.78
r66 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.615 $X2=0.97 $Y2=1.615
r67 16 28 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=2.38 $Y2=1.615
r68 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=2.16 $Y2=1.615
r69 14 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.68 $Y2=1.615
r70 14 23 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=0.97 $Y2=1.615
r71 13 23 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.97 $Y2=1.615
r72 11 29 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.44 $Y=0.74
+ $X2=2.44 $Y2=1.45
r73 7 30 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.39 $Y=2.44 $X2=2.39
+ $Y2=1.78
r74 3 25 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=2.44
+ $X2=0.955 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%C 3 7 9 11 15 17 20 21
r53 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=0.435 $X2=1.215 $Y2=0.435
r54 17 21 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.215 $Y=0.555
+ $X2=1.215 $Y2=0.435
r55 15 16 9.34914 $w=2.32e-07 $l=4.5e-08 $layer=POLY_cond $X=1.885 $Y=1.345
+ $X2=1.93 $Y2=1.345
r56 14 15 93.4914 $w=2.32e-07 $l=4.5e-07 $layer=POLY_cond $X=1.435 $Y=1.345
+ $X2=1.885 $Y2=1.345
r57 13 20 93.7338 $w=4.45e-07 $l=7.5e-07 $layer=POLY_cond $X=1.272 $Y=1.185
+ $X2=1.272 $Y2=0.435
r58 13 14 33.8647 $w=2.32e-07 $l=2.29454e-07 $layer=POLY_cond $X=1.272 $Y=1.185
+ $X2=1.435 $Y2=1.345
r59 9 16 12.995 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.93 $Y=1.185 $X2=1.93
+ $Y2=1.345
r60 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.93 $Y=1.185
+ $X2=1.93 $Y2=0.74
r61 5 15 8.79421 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=1.885 $Y=1.505
+ $X2=1.885 $Y2=1.345
r62 5 7 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=1.885 $Y=1.505
+ $X2=1.885 $Y2=2.44
r63 1 14 8.79421 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=1.435 $Y=1.505
+ $X2=1.435 $Y2=1.345
r64 1 3 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=1.435 $Y=1.505
+ $X2=1.435 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%A_305_388# 1 2 3 12 16 20 24 28 32 36 40 44 46
+ 48 49 52 54 57 59 65 71 73 74 85
c163 85 0 1.56424e-19 $X=4.785 $Y=1.465
r164 84 85 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.775 $Y=1.465
+ $X2=4.785 $Y2=1.465
r165 81 82 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.325 $Y=1.465
+ $X2=4.355 $Y2=1.465
r166 80 81 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=3.875 $Y=1.465
+ $X2=4.325 $Y2=1.465
r167 79 80 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.865 $Y=1.465
+ $X2=3.875 $Y2=1.465
r168 75 77 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=3.425 $Y=1.465
+ $X2=3.43 $Y2=1.465
r169 69 71 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=2.075
+ $X2=1.825 $Y2=2.075
r170 66 84 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=4.52 $Y=1.465
+ $X2=4.775 $Y2=1.465
r171 66 82 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=1.465
+ $X2=4.355 $Y2=1.465
r172 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.465 $X2=4.52 $Y2=1.465
r173 63 79 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=3.5 $Y=1.465
+ $X2=3.865 $Y2=1.465
r174 63 77 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.5 $Y=1.465 $X2=3.43
+ $Y2=1.465
r175 62 65 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.5 $Y=1.465
+ $X2=4.52 $Y2=1.465
r176 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.5
+ $Y=1.465 $X2=3.5 $Y2=1.465
r177 60 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=1.465
+ $X2=3.31 $Y2=1.465
r178 60 62 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.395 $Y=1.465
+ $X2=3.5 $Y2=1.465
r179 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=1.63
+ $X2=3.31 $Y2=1.465
r180 58 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=1.63
+ $X2=3.31 $Y2=1.95
r181 57 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=1.3
+ $X2=3.31 $Y2=1.465
r182 56 57 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.31 $Y=0.94
+ $X2=3.31 $Y2=1.3
r183 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=0.855
+ $X2=2.715 $Y2=0.855
r184 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.225 $Y=0.855
+ $X2=3.31 $Y2=0.94
r185 54 55 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.225 $Y=0.855
+ $X2=2.88 $Y2=0.855
r186 50 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.77
+ $X2=2.715 $Y2=0.855
r187 50 52 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.715 $Y=0.77
+ $X2=2.715 $Y2=0.515
r188 48 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0.855
+ $X2=2.715 $Y2=0.855
r189 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.55 $Y=0.855
+ $X2=1.88 $Y2=0.855
r190 46 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.225 $Y=2.035
+ $X2=3.31 $Y2=1.95
r191 46 71 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.225 $Y=2.035
+ $X2=1.825 $Y2=2.035
r192 42 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.715 $Y=0.77
+ $X2=1.88 $Y2=0.855
r193 42 44 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.715 $Y=0.77
+ $X2=1.715 $Y2=0.515
r194 38 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=1.465
r195 38 40 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=0.74
r196 34 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.63
+ $X2=4.775 $Y2=1.465
r197 34 36 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.775 $Y=1.63
+ $X2=4.775 $Y2=2.4
r198 30 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=1.465
r199 30 32 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=0.74
r200 26 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.325 $Y=1.63
+ $X2=4.325 $Y2=1.465
r201 26 28 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.325 $Y=1.63
+ $X2=4.325 $Y2=2.4
r202 22 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=1.3
+ $X2=3.865 $Y2=1.465
r203 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.865 $Y=1.3
+ $X2=3.865 $Y2=0.74
r204 18 80 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=1.63
+ $X2=3.875 $Y2=1.465
r205 18 20 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.875 $Y=1.63
+ $X2=3.875 $Y2=2.4
r206 14 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.3
+ $X2=3.43 $Y2=1.465
r207 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.43 $Y=1.3
+ $X2=3.43 $Y2=0.74
r208 10 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.63
+ $X2=3.425 $Y2=1.465
r209 10 12 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.425 $Y=1.63
+ $X2=3.425 $Y2=2.4
r210 3 69 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.94 $X2=1.66 $Y2=2.1
r211 2 73 182 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.37 $X2=2.715 $Y2=0.855
r212 2 52 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.37 $X2=2.715 $Y2=0.515
r213 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.715 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%VPWR 1 2 3 4 13 15 21 25 27 29 31 33 41 46 55
+ 58 62
r67 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r69 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 50 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r72 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 47 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.06 $Y2=3.33
r75 47 49 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 46 61 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=5.097 $Y2=3.33
r77 46 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r79 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.2 $Y2=3.33
r82 42 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=4.06 $Y2=3.33
r84 41 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=3.6 $Y2=3.33
r85 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 34 52 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r89 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.2 $Y2=3.33
r91 33 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 31 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 31 37 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=0.72 $Y2=3.33
r94 31 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 27 61 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.097 $Y2=3.33
r96 27 29 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=2.305
r97 23 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=3.245
+ $X2=4.06 $Y2=3.33
r98 23 25 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.06 $Y=3.245
+ $X2=4.06 $Y2=2.305
r99 19 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=3.245 $X2=3.2
+ $Y2=3.33
r100 19 21 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.2 $Y=3.245
+ $X2=3.2 $Y2=2.455
r101 15 18 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.085
+ $X2=0.24 $Y2=2.795
r102 13 52 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r103 13 18 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.795
r104 4 29 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.84 $X2=5 $Y2=2.305
r105 3 25 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=3.965
+ $Y=1.84 $X2=4.1 $Y2=2.305
r106 2 21 300 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_PDIFF $count=2 $X=2.98
+ $Y=1.94 $X2=3.2 $Y2=2.455
r107 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.94 $X2=0.28 $Y2=2.795
r108 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.94 $X2=0.28 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%A_119_388# 1 2 9 13 15 17 19 22
c32 19 0 1.92271e-19 $X=2.665 $Y=2.795
c33 13 0 1.71217e-19 $X=0.73 $Y=2.795
c34 9 0 1.91378e-19 $X=0.73 $Y=2.115
r35 17 24 2.94173 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=2.665 $Y=2.54
+ $X2=2.665 $Y2=2.415
r36 17 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.665 $Y=2.54
+ $X2=2.665 $Y2=2.795
r37 16 22 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=2.455
+ $X2=0.69 $Y2=2.455
r38 15 24 4.82444 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.5 $Y=2.455
+ $X2=2.665 $Y2=2.415
r39 15 16 109.93 $w=1.68e-07 $l=1.685e-06 $layer=LI1_cond $X=2.5 $Y=2.455
+ $X2=0.815 $Y2=2.455
r40 11 22 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.54 $X2=0.69
+ $Y2=2.455
r41 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=2.54
+ $X2=0.69 $Y2=2.795
r42 7 22 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.37 $X2=0.69
+ $Y2=2.455
r43 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=2.37 $X2=0.69
+ $Y2=2.115
r44 2 24 600 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.94 $X2=2.665 $Y2=2.455
r45 2 19 600 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.94 $X2=2.665 $Y2=2.795
r46 1 22 600 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.94 $X2=0.73 $Y2=2.455
r47 1 13 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.94 $X2=0.73 $Y2=2.795
r48 1 9 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.94 $X2=0.73 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%A_209_388# 1 2 11
c14 11 0 1.50847e-19 $X=2.135 $Y=2.795
r15 8 11 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.195 $Y=2.835
+ $X2=2.135 $Y2=2.835
r16 2 11 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.94 $X2=2.135 $Y2=2.795
r17 1 8 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.94 $X2=1.195 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%X 1 2 3 4 15 19 23 24 25 26 29 35 37 39 41 42
+ 45 46
c79 37 0 1.56424e-19 $X=4.925 $Y=1.045
r80 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.665
r81 44 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=1.8
+ $X2=5.04 $Y2=1.665
r82 43 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=1.13
+ $X2=5.04 $Y2=1.295
r83 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=1.885
+ $X2=4.55 $Y2=1.885
r84 39 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.925 $Y=1.885
+ $X2=5.04 $Y2=1.8
r85 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.925 $Y=1.885
+ $X2=4.715 $Y2=1.885
r86 38 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.655 $Y=1.045
+ $X2=4.53 $Y2=1.045
r87 37 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.925 $Y=1.045
+ $X2=5.04 $Y2=1.13
r88 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.925 $Y=1.045
+ $X2=4.655 $Y2=1.045
r89 33 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.96
+ $X2=4.53 $Y2=1.045
r90 33 35 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.53 $Y=0.96
+ $X2=4.53 $Y2=0.515
r91 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.55 $Y=1.985
+ $X2=4.55 $Y2=2.815
r92 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=1.97 $X2=4.55
+ $Y2=1.885
r93 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.55 $Y=1.97
+ $X2=4.55 $Y2=1.985
r94 25 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=1.885
+ $X2=4.55 $Y2=1.885
r95 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.385 $Y=1.885
+ $X2=3.735 $Y2=1.885
r96 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.405 $Y=1.045
+ $X2=4.53 $Y2=1.045
r97 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.405 $Y=1.045
+ $X2=3.735 $Y2=1.045
r98 19 21 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.65 $Y=1.985
+ $X2=3.65 $Y2=2.815
r99 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.65 $Y=1.97
+ $X2=3.735 $Y2=1.885
r100 17 19 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.65 $Y=1.97
+ $X2=3.65 $Y2=1.985
r101 13 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.65 $Y=0.96
+ $X2=3.735 $Y2=1.045
r102 13 15 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.65 $Y=0.96
+ $X2=3.65 $Y2=0.515
r103 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.84 $X2=4.55 $Y2=2.815
r104 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.84 $X2=4.55 $Y2=1.985
r105 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.65 $Y2=2.815
r106 3 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.65 $Y2=1.985
r107 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.515
r108 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=0.37 $X2=3.65 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR3_4%VGND 1 2 3 4 15 17 21 25 27 29 31 33 41 46 52
+ 55 58 62
r74 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r75 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r76 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r77 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 50 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r79 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r80 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r81 47 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.04
+ $Y2=0
r82 47 49 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.56
+ $Y2=0
r83 46 61 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.057
+ $Y2=0
r84 46 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.56
+ $Y2=0
r85 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r86 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r87 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r88 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.215
+ $Y2=0
r89 42 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.6
+ $Y2=0
r90 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=4.04
+ $Y2=0
r91 41 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=3.6
+ $Y2=0
r92 40 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r93 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r94 36 40 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r95 35 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r96 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.215
+ $Y2=0
r98 33 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.68
+ $Y2=0
r99 31 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r100 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r101 27 61 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=0.085
+ $X2=5.057 $Y2=0
r102 27 29 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.61
r103 23 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r104 23 25 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.57
r105 19 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.085
+ $X2=3.215 $Y2=0
r106 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.215 $Y=0.085
+ $X2=3.215 $Y2=0.515
r107 18 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.215
+ $Y2=0
r108 17 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=3.215
+ $Y2=0
r109 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=2.38
+ $Y2=0
r110 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0
r111 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0.515
r112 4 29 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.61
r113 3 25 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=3.94
+ $Y=0.37 $X2=4.08 $Y2=0.57
r114 2 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.37 $X2=3.215 $Y2=0.515
r115 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.37 $X2=2.215 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__sdfxbp_1.spice
* Created: Wed Sep  2 12:31:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfxbp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfxbp_1  VNB VPB SCE D SCD CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_SCE_M1024_g N_A_31_74#_M1024_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1007 A_218_74# N_A_31_74#_M1007_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_296_74#_M1008_d N_D_M1008_g A_218_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1134 AS=0.0504 PD=0.96 PS=0.66 NRD=37.14 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 A_434_74# N_SCE_M1003_g N_A_296_74#_M1008_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1134 PD=0.66 PS=0.96 NRD=18.564 NRS=37.14 M=1 R=2.8 SA=75001.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_SCD_M1027_g A_434_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_A_612_74#_M1023_d N_CLK_M1023_g N_VGND_M1027_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=4.86 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_828_74#_M1015_d N_A_612_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.2805 PD=2.02 PS=2.25 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 N_A_1021_100#_M1030_d N_A_612_74#_M1030_g N_A_296_74#_M1030_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1155 PD=0.95 PS=1.39 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1006 A_1157_100# N_A_828_74#_M1006_g N_A_1021_100#_M1030_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0966 AS=0.1113 PD=0.88 PS=0.95 NRD=49.992 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1243_398#_M1016_g A_1157_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.172849 AS=0.0966 PD=1.19072 PS=0.88 NRD=101.868 NRS=49.992 M=1 R=2.8
+ SA=75001.5 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_1243_398#_M1011_d N_A_1021_100#_M1011_g N_VGND_M1016_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.078375 AS=0.226351 PD=0.835 PS=1.55928 NRD=1.08 NRS=72 M=1
+ R=3.66667 SA=75001.9 SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1010 N_A_1529_74#_M1010_d N_A_828_74#_M1010_g N_A_1243_398#_M1011_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.163696 AS=0.078375 PD=1.31546 PS=0.835 NRD=72 NRS=0 M=1
+ R=3.66667 SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1017 A_1681_74# N_A_612_74#_M1017_g N_A_1529_74#_M1010_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.125004 PD=0.63 PS=1.00454 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1723_48#_M1021_g A_1681_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.128793 AS=0.0441 PD=1.0132 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_A_1723_48#_M1001_d N_A_1529_74#_M1001_g N_VGND_M1021_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.168657 PD=1.67 PS=1.3268 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75003.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1012 N_Q_M1012_d N_A_1723_48#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_VGND_M1035_d N_A_1723_48#_M1035_g N_A_2216_112#_M1035_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.118548 AS=0.15675 PD=0.967829 PS=1.67 NRD=13.08 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1026 N_Q_N_M1026_d N_A_2216_112#_M1026_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.159502 PD=2.05 PS=1.30217 NRD=0 NRS=9.324 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_VPWR_M1022_d N_SCE_M1022_g N_A_31_74#_M1022_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.1792 PD=0.96 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.8 A=0.1152 P=1.64 MULT=1
MM1018 A_236_464# N_SCE_M1018_g N_VPWR_M1022_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90002.3 A=0.1152 P=1.64 MULT=1
MM1028 N_A_296_74#_M1028_d N_D_M1028_g A_236_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.1
+ SB=90001.9 A=0.1152 P=1.64 MULT=1
MM1032 A_410_464# N_A_31_74#_M1032_g N_A_296_74#_M1028_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1152 AS=0.0864 PD=1 PS=0.91 NRD=38.4741 NRS=0 M=1 R=3.55556
+ SA=90001.6 SB=90001.4 A=0.1152 P=1.64 MULT=1
MM1009 N_VPWR_M1009_d N_SCD_M1009_g A_410_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.166982 AS=0.1152 PD=1.2 PS=1 NRD=38.4741 NRS=38.4741 M=1 R=3.55556
+ SA=90002.1 SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1013 N_A_612_74#_M1013_d N_CLK_M1013_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.292218 PD=2.8 PS=2.1 NRD=0 NRS=21.9852 M=1 R=6.22222 SA=90001.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1025 N_A_828_74#_M1025_d N_A_612_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.5096 PD=2.77 PS=3.15 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1029 N_A_1021_100#_M1029_d N_A_828_74#_M1029_g N_A_296_74#_M1029_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1113 PD=0.69 PS=1.37 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90004.1 A=0.0756 P=1.2 MULT=1
MM1033 A_1183_496# N_A_612_74#_M1033_g N_A_1021_100#_M1029_d VPB PSHORT L=0.18
+ W=0.42 AD=0.063 AS=0.0567 PD=0.72 PS=0.69 NRD=44.5417 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90003.6 A=0.0756 P=1.2 MULT=1
MM1031 N_VPWR_M1031_d N_A_1243_398#_M1031_g A_1183_496# VPB PSHORT L=0.18 W=0.42
+ AD=0.1192 AS=0.063 PD=0.993333 PS=0.72 NRD=107.306 NRS=44.5417 M=1 R=2.33333
+ SA=90001.1 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1019 N_A_1243_398#_M1019_d N_A_1021_100#_M1019_g N_VPWR_M1031_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.3108 AS=0.2384 PD=1.58 PS=1.98667 NRD=0 NRS=53.6431 M=1
+ R=4.66667 SA=90001 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1000 N_A_1529_74#_M1000_d N_A_612_74#_M1000_g N_A_1243_398#_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1778 AS=0.3108 PD=1.59333 PS=1.58 NRD=0 NRS=99.6623 M=1
+ R=4.66667 SA=90001.9 SB=90001 A=0.1512 P=2.04 MULT=1
MM1020 A_1694_508# N_A_828_74#_M1020_g N_A_1529_74#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0889 PD=0.66 PS=0.796667 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90003 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_1723_48#_M1002_g A_1694_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.112454 AS=0.0504 PD=0.922817 PS=0.66 NRD=60.9715 NRS=30.4759 M=1
+ R=2.33333 SA=90003.4 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1014 N_A_1723_48#_M1014_d N_A_1529_74#_M1014_g N_VPWR_M1002_d VPB PSHORT
+ L=0.18 W=1 AD=0.26 AS=0.267746 PD=2.52 PS=2.19718 NRD=0 NRS=29.55 M=1
+ R=5.55556 SA=90001.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_Q_M1005_d N_A_1723_48#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_1723_48#_M1004_g N_A_2216_112#_M1004_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.2184 PD=1.23857 PS=2.2 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1034 N_Q_N_M1034_d N_A_2216_112#_M1034_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3024 AS=0.196 PD=2.78 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX36_noxref VNB VPB NWDIODE A=23.9196 P=29.44
c_142 VNB 0 1.65961e-19 $X=0 $Y=0
c_1886 A_434_74# 0 2.47416e-20 $X=2.17 $Y=0.37
*
.include "sky130_fd_sc_ms__sdfxbp_1.pxi.spice"
*
.ends
*
*

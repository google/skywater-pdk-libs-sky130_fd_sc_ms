* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_247_368# B2 a_84_48# VPB pshort w=1e+06u l=180000u
+  ad=8.2e+11p pd=7.64e+06u as=3.7e+11p ps=2.74e+06u
M1001 a_247_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.0496e+12p ps=6.26e+06u
M1002 a_84_48# B1 a_247_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_247_368# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A2 a_247_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_601_94# B1 a_84_48# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=4.032e+11p ps=2.54e+06u
M1006 a_259_94# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=6.004e+11p ps=4.48e+06u
M1007 a_337_94# A2 a_259_94# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1008 VPWR a_84_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1009 VGND B2 a_601_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_84_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_84_48# A1 a_337_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

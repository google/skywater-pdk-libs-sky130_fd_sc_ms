* File: sky130_fd_sc_ms__sdfrbp_2.pxi.spice
* Created: Fri Aug 28 18:11:50 2020
* 
x_PM_SKY130_FD_SC_MS__SDFRBP_2%SCE N_SCE_c_285_n N_SCE_M1009_g N_SCE_c_286_n
+ N_SCE_M1030_g N_SCE_c_295_n N_SCE_M1039_g N_SCE_M1031_g N_SCE_c_288_n
+ N_SCE_c_297_n N_SCE_c_289_n N_SCE_c_290_n N_SCE_c_291_n N_SCE_c_292_n SCE SCE
+ SCE N_SCE_c_299_n N_SCE_c_300_n PM_SKY130_FD_SC_MS__SDFRBP_2%SCE
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_27_79# N_A_27_79#_M1030_s N_A_27_79#_M1009_s
+ N_A_27_79#_M1012_g N_A_27_79#_M1027_g N_A_27_79#_c_374_n N_A_27_79#_c_375_n
+ N_A_27_79#_c_376_n N_A_27_79#_c_381_n N_A_27_79#_c_377_n N_A_27_79#_c_402_n
+ N_A_27_79#_c_382_n N_A_27_79#_c_378_n N_A_27_79#_c_383_n N_A_27_79#_c_384_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_27_79#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%D N_D_M1026_g N_D_M1006_g D N_D_c_459_n
+ N_D_c_460_n N_D_c_461_n PM_SKY130_FD_SC_MS__SDFRBP_2%D
x_PM_SKY130_FD_SC_MS__SDFRBP_2%SCD N_SCD_M1041_g N_SCD_M1013_g N_SCD_c_503_n
+ N_SCD_c_508_n SCD SCD N_SCD_c_505_n PM_SKY130_FD_SC_MS__SDFRBP_2%SCD
x_PM_SKY130_FD_SC_MS__SDFRBP_2%CLK N_CLK_c_547_n N_CLK_M1021_g N_CLK_M1019_g
+ N_CLK_c_548_n CLK N_CLK_c_550_n PM_SKY130_FD_SC_MS__SDFRBP_2%CLK
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_1025_119# N_A_1025_119#_M1033_d
+ N_A_1025_119#_M1036_d N_A_1025_119#_M1032_g N_A_1025_119#_c_599_n
+ N_A_1025_119#_M1015_g N_A_1025_119#_c_601_n N_A_1025_119#_M1017_g
+ N_A_1025_119#_c_602_n N_A_1025_119#_c_603_n N_A_1025_119#_M1042_g
+ N_A_1025_119#_c_604_n N_A_1025_119#_c_605_n N_A_1025_119#_c_606_n
+ N_A_1025_119#_c_607_n N_A_1025_119#_c_608_n N_A_1025_119#_c_609_n
+ N_A_1025_119#_c_779_p N_A_1025_119#_c_610_n N_A_1025_119#_c_611_n
+ N_A_1025_119#_c_612_n N_A_1025_119#_c_613_n N_A_1025_119#_c_614_n
+ N_A_1025_119#_c_615_n N_A_1025_119#_c_616_n N_A_1025_119#_c_617_n
+ N_A_1025_119#_c_624_n N_A_1025_119#_c_618_n N_A_1025_119#_c_619_n
+ N_A_1025_119#_c_627_n PM_SKY130_FD_SC_MS__SDFRBP_2%A_1025_119#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_1370_290# N_A_1370_290#_M1007_d
+ N_A_1370_290#_M1000_d N_A_1370_290#_M1020_g N_A_1370_290#_M1043_g
+ N_A_1370_290#_c_804_n N_A_1370_290#_c_805_n N_A_1370_290#_c_822_n
+ N_A_1370_290#_c_824_n N_A_1370_290#_c_812_n N_A_1370_290#_c_806_n
+ N_A_1370_290#_c_807_n N_A_1370_290#_c_808_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_1370_290#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%RESET_B N_RESET_B_M1003_g N_RESET_B_M1035_g
+ N_RESET_B_c_893_n N_RESET_B_c_894_n N_RESET_B_M1011_g N_RESET_B_c_896_n
+ N_RESET_B_c_897_n N_RESET_B_c_903_n N_RESET_B_M1034_g N_RESET_B_c_898_n
+ N_RESET_B_M1024_g N_RESET_B_M1023_g N_RESET_B_c_906_n N_RESET_B_c_900_n
+ N_RESET_B_c_908_n N_RESET_B_c_909_n N_RESET_B_c_910_n N_RESET_B_c_911_n
+ RESET_B N_RESET_B_c_913_n N_RESET_B_c_914_n N_RESET_B_c_915_n
+ N_RESET_B_c_916_n N_RESET_B_c_917_n N_RESET_B_c_918_n N_RESET_B_c_919_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%RESET_B
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_1223_119# N_A_1223_119#_M1014_d
+ N_A_1223_119#_M1032_d N_A_1223_119#_M1034_d N_A_1223_119#_M1007_g
+ N_A_1223_119#_M1000_g N_A_1223_119#_c_1121_n N_A_1223_119#_c_1108_n
+ N_A_1223_119#_c_1136_n N_A_1223_119#_c_1115_n N_A_1223_119#_c_1109_n
+ N_A_1223_119#_c_1110_n N_A_1223_119#_c_1111_n N_A_1223_119#_c_1112_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_1223_119#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_852_119# N_A_852_119#_M1021_s
+ N_A_852_119#_M1019_s N_A_852_119#_M1033_g N_A_852_119#_M1036_g
+ N_A_852_119#_c_1209_n N_A_852_119#_c_1210_n N_A_852_119#_c_1211_n
+ N_A_852_119#_c_1212_n N_A_852_119#_c_1213_n N_A_852_119#_c_1226_n
+ N_A_852_119#_c_1227_n N_A_852_119#_c_1214_n N_A_852_119#_M1014_g
+ N_A_852_119#_M1040_g N_A_852_119#_c_1229_n N_A_852_119#_M1004_g
+ N_A_852_119#_c_1215_n N_A_852_119#_c_1216_n N_A_852_119#_M1002_g
+ N_A_852_119#_c_1218_n N_A_852_119#_c_1233_n N_A_852_119#_c_1237_n
+ N_A_852_119#_c_1219_n N_A_852_119#_c_1220_n N_A_852_119#_c_1221_n
+ N_A_852_119#_c_1222_n N_A_852_119#_c_1223_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_852_119#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_2006_373# N_A_2006_373#_M1016_d
+ N_A_2006_373#_M1023_d N_A_2006_373#_M1022_g N_A_2006_373#_M1045_g
+ N_A_2006_373#_c_1391_n N_A_2006_373#_c_1392_n N_A_2006_373#_c_1383_n
+ N_A_2006_373#_c_1384_n N_A_2006_373#_c_1394_n N_A_2006_373#_c_1395_n
+ N_A_2006_373#_c_1385_n N_A_2006_373#_c_1386_n N_A_2006_373#_c_1387_n
+ N_A_2006_373#_c_1388_n N_A_2006_373#_c_1396_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_2006_373#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_1790_74# N_A_1790_74#_M1017_d
+ N_A_1790_74#_M1004_d N_A_1790_74#_M1016_g N_A_1790_74#_c_1497_n
+ N_A_1790_74#_M1028_g N_A_1790_74#_c_1498_n N_A_1790_74#_M1005_g
+ N_A_1790_74#_M1025_g N_A_1790_74#_M1008_g N_A_1790_74#_M1037_g
+ N_A_1790_74#_c_1502_n N_A_1790_74#_M1029_g N_A_1790_74#_M1010_g
+ N_A_1790_74#_c_1516_n N_A_1790_74#_c_1519_n N_A_1790_74#_c_1505_n
+ N_A_1790_74#_c_1506_n N_A_1790_74#_c_1507_n N_A_1790_74#_c_1529_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_1790_74#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_2607_392# N_A_2607_392#_M1010_d
+ N_A_2607_392#_M1029_d N_A_2607_392#_M1001_g N_A_2607_392#_M1018_g
+ N_A_2607_392#_M1044_g N_A_2607_392#_M1038_g N_A_2607_392#_c_1646_n
+ N_A_2607_392#_c_1647_n N_A_2607_392#_c_1648_n N_A_2607_392#_c_1649_n
+ N_A_2607_392#_c_1665_p N_A_2607_392#_c_1650_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%A_2607_392#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%VPWR N_VPWR_M1009_d N_VPWR_M1041_d N_VPWR_M1019_d
+ N_VPWR_M1020_d N_VPWR_M1000_s N_VPWR_M1022_d N_VPWR_M1028_d N_VPWR_M1008_s
+ N_VPWR_M1001_d N_VPWR_M1044_d N_VPWR_c_1693_n N_VPWR_c_1694_n N_VPWR_c_1695_n
+ N_VPWR_c_1696_n N_VPWR_c_1697_n N_VPWR_c_1698_n N_VPWR_c_1699_n
+ N_VPWR_c_1700_n N_VPWR_c_1701_n N_VPWR_c_1702_n N_VPWR_c_1703_n
+ N_VPWR_c_1704_n N_VPWR_c_1705_n N_VPWR_c_1706_n VPWR N_VPWR_c_1707_n
+ N_VPWR_c_1708_n N_VPWR_c_1709_n N_VPWR_c_1710_n N_VPWR_c_1711_n
+ N_VPWR_c_1712_n N_VPWR_c_1713_n N_VPWR_c_1714_n N_VPWR_c_1715_n
+ N_VPWR_c_1716_n N_VPWR_c_1717_n N_VPWR_c_1718_n N_VPWR_c_1719_n
+ N_VPWR_c_1720_n N_VPWR_c_1692_n PM_SKY130_FD_SC_MS__SDFRBP_2%VPWR
x_PM_SKY130_FD_SC_MS__SDFRBP_2%A_388_79# N_A_388_79#_M1026_d N_A_388_79#_M1014_s
+ N_A_388_79#_M1006_d N_A_388_79#_M1035_d N_A_388_79#_M1032_s
+ N_A_388_79#_c_1893_n N_A_388_79#_c_1874_n N_A_388_79#_c_1875_n
+ N_A_388_79#_c_1876_n N_A_388_79#_c_1904_n N_A_388_79#_c_1883_n
+ N_A_388_79#_c_1884_n N_A_388_79#_c_1877_n N_A_388_79#_c_1886_n
+ N_A_388_79#_c_1887_n N_A_388_79#_c_1888_n N_A_388_79#_c_1889_n
+ N_A_388_79#_c_1878_n N_A_388_79#_c_1890_n N_A_388_79#_c_1891_n
+ N_A_388_79#_c_1879_n N_A_388_79#_c_1880_n N_A_388_79#_c_1881_n
+ N_A_388_79#_c_1882_n PM_SKY130_FD_SC_MS__SDFRBP_2%A_388_79#
x_PM_SKY130_FD_SC_MS__SDFRBP_2%Q_N N_Q_N_M1025_d N_Q_N_M1005_d Q_N Q_N Q_N
+ N_Q_N_c_2045_n Q_N PM_SKY130_FD_SC_MS__SDFRBP_2%Q_N
x_PM_SKY130_FD_SC_MS__SDFRBP_2%Q N_Q_M1018_d N_Q_M1001_s Q N_Q_c_2072_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%Q
x_PM_SKY130_FD_SC_MS__SDFRBP_2%VGND N_VGND_M1030_d N_VGND_M1003_d N_VGND_M1021_d
+ N_VGND_M1011_d N_VGND_M1045_d N_VGND_M1025_s N_VGND_M1037_s N_VGND_M1018_s
+ N_VGND_M1038_s N_VGND_c_2088_n N_VGND_c_2089_n N_VGND_c_2090_n N_VGND_c_2091_n
+ N_VGND_c_2092_n N_VGND_c_2093_n N_VGND_c_2094_n N_VGND_c_2095_n
+ N_VGND_c_2096_n N_VGND_c_2097_n N_VGND_c_2098_n N_VGND_c_2099_n
+ N_VGND_c_2100_n N_VGND_c_2101_n N_VGND_c_2102_n N_VGND_c_2103_n VGND
+ N_VGND_c_2104_n N_VGND_c_2105_n N_VGND_c_2106_n N_VGND_c_2107_n
+ N_VGND_c_2108_n N_VGND_c_2109_n N_VGND_c_2110_n N_VGND_c_2111_n
+ N_VGND_c_2112_n N_VGND_c_2113_n N_VGND_c_2114_n
+ PM_SKY130_FD_SC_MS__SDFRBP_2%VGND
x_PM_SKY130_FD_SC_MS__SDFRBP_2%noxref_25 N_noxref_25_M1012_s N_noxref_25_M1013_d
+ N_noxref_25_c_2245_n N_noxref_25_c_2246_n N_noxref_25_c_2247_n
+ N_noxref_25_c_2248_n PM_SKY130_FD_SC_MS__SDFRBP_2%noxref_25
cc_1 VNB N_SCE_c_285_n 0.0443833f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.82
cc_2 VNB N_SCE_c_286_n 0.0211781f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.89
cc_3 VNB N_SCE_M1031_g 0.0363026f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_4 VNB N_SCE_c_288_n 0.0216296f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.965
cc_5 VNB N_SCE_c_289_n 0.00133979f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.82
cc_6 VNB N_SCE_c_290_n 0.00450757f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.49
cc_7 VNB N_SCE_c_291_n 0.0230028f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.455
cc_8 VNB N_SCE_c_292_n 0.0330707f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.455
cc_9 VNB N_A_27_79#_M1012_g 0.0455097f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.605
cc_10 VNB N_A_27_79#_c_374_n 0.0789787f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_11 VNB N_A_27_79#_c_375_n 0.0355558f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=0.965
cc_12 VNB N_A_27_79#_c_376_n 0.00354448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_79#_c_377_n 0.00484068f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.455
cc_14 VNB N_A_27_79#_c_378_n 0.0159647f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.985
cc_15 VNB N_D_M1006_g 0.0238331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_459_n 0.0310845f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_17 VNB N_D_c_460_n 0.00902418f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_18 VNB N_D_c_461_n 0.0162587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCD_M1013_g 0.042619f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.89
cc_20 VNB N_SCD_c_503_n 0.00499797f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_21 VNB SCD 0.00197778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_505_n 0.0164016f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=0.965
cc_23 VNB N_CLK_c_547_n 0.0164766f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.04
cc_24 VNB N_CLK_c_548_n 0.0436566f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.15
cc_25 VNB CLK 0.00857922f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_26 VNB N_CLK_c_550_n 0.0422129f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_27 VNB N_A_1025_119#_c_599_n 0.0264223f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_28 VNB N_A_1025_119#_M1015_g 0.0359456f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_29 VNB N_A_1025_119#_c_601_n 0.016501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_1025_119#_c_602_n 0.0226212f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.965
cc_31 VNB N_A_1025_119#_c_603_n 0.00721388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1025_119#_c_604_n 0.00630499f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.455
cc_33 VNB N_A_1025_119#_c_605_n 0.00151619f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_34 VNB N_A_1025_119#_c_606_n 0.0214463f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_35 VNB N_A_1025_119#_c_607_n 0.00390562f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.95
cc_36 VNB N_A_1025_119#_c_608_n 0.00204982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1025_119#_c_609_n 0.00174335f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=1.985
cc_38 VNB N_A_1025_119#_c_610_n 0.00706005f $X=-0.19 $Y=-0.245 $X2=1.385
+ $Y2=1.985
cc_39 VNB N_A_1025_119#_c_611_n 0.00245748f $X=-0.19 $Y=-0.245 $X2=1.385
+ $Y2=1.985
cc_40 VNB N_A_1025_119#_c_612_n 0.00157163f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.29
cc_41 VNB N_A_1025_119#_c_613_n 0.00388845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1025_119#_c_614_n 4.77558e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1025_119#_c_615_n 0.00358753f $X=-0.19 $Y=-0.245 $X2=1.71
+ $Y2=1.985
cc_44 VNB N_A_1025_119#_c_616_n 0.00460249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1025_119#_c_617_n 0.033082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1025_119#_c_618_n 0.0048475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1025_119#_c_619_n 0.0144077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1370_290#_M1043_g 0.0295995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1370_290#_c_804_n 0.00357226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1370_290#_c_805_n 0.0255382f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=0.965
cc_51 VNB N_A_1370_290#_c_806_n 0.00911531f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.95
cc_52 VNB N_A_1370_290#_c_807_n 0.00431592f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=1.95
cc_53 VNB N_A_1370_290#_c_808_n 0.00664491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_RESET_B_M1003_g 0.0519467f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_55 VNB N_RESET_B_c_893_n 0.267541f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.605
cc_56 VNB N_RESET_B_c_894_n 0.0126359f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.15
cc_57 VNB N_RESET_B_M1011_g 0.0292065f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=1.29
cc_58 VNB N_RESET_B_c_896_n 0.0258223f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_59 VNB N_RESET_B_c_897_n 0.0119677f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_60 VNB N_RESET_B_c_898_n 0.0223419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_M1024_g 0.0456332f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.62
cc_62 VNB N_RESET_B_c_900_n 0.0112292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1223_119#_M1007_g 0.0268435f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_64 VNB N_A_1223_119#_c_1108_n 0.0108902f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.82
cc_65 VNB N_A_1223_119#_c_1109_n 0.00155425f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.49
cc_66 VNB N_A_1223_119#_c_1110_n 0.00408417f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.455
cc_67 VNB N_A_1223_119#_c_1111_n 0.00984593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1223_119#_c_1112_n 0.0288317f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_69 VNB N_A_852_119#_c_1209_n 0.0120355f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=1.29
cc_70 VNB N_A_852_119#_c_1210_n 0.009011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_852_119#_c_1211_n 0.00287746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_852_119#_c_1212_n 0.0251275f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.965
cc_73 VNB N_A_852_119#_c_1213_n 0.00939473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_852_119#_c_1214_n 0.0162581f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.62
cc_75 VNB N_A_852_119#_c_1215_n 0.029955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_852_119#_c_1216_n 0.00540003f $X=-0.19 $Y=-0.245 $X2=1.37
+ $Y2=1.985
cc_77 VNB N_A_852_119#_M1002_g 0.0453681f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.985
cc_78 VNB N_A_852_119#_c_1218_n 0.00534438f $X=-0.19 $Y=-0.245 $X2=1.385
+ $Y2=1.985
cc_79 VNB N_A_852_119#_c_1219_n 6.69765e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_852_119#_c_1220_n 0.00560778f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.985
cc_81 VNB N_A_852_119#_c_1221_n 0.00619427f $X=-0.19 $Y=-0.245 $X2=1.71
+ $Y2=1.985
cc_82 VNB N_A_852_119#_c_1222_n 0.0141414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_852_119#_c_1223_n 0.0167287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2006_373#_M1045_g 0.0481405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2006_373#_c_1383_n 0.00410394f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.965
cc_86 VNB N_A_2006_373#_c_1384_n 0.00173724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2006_373#_c_1385_n 0.0070639f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.49
cc_88 VNB N_A_2006_373#_c_1386_n 0.00667447f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.455
cc_89 VNB N_A_2006_373#_c_1387_n 0.00230863f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.455
cc_90 VNB N_A_2006_373#_c_1388_n 0.00172407f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_91 VNB N_A_1790_74#_M1016_g 0.0262898f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.605
cc_92 VNB N_A_1790_74#_c_1497_n 0.0559917f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_93 VNB N_A_1790_74#_c_1498_n 0.0260795f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_94 VNB N_A_1790_74#_M1025_g 0.0197591f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.82
cc_95 VNB N_A_1790_74#_M1008_g 3.32386e-19 $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.49
cc_96 VNB N_A_1790_74#_M1037_g 0.0192815f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_97 VNB N_A_1790_74#_c_1502_n 0.0611909f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.95
cc_98 VNB N_A_1790_74#_M1029_g 0.00428291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1790_74#_M1010_g 0.027051f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.985
cc_100 VNB N_A_1790_74#_c_1505_n 0.00230536f $X=-0.19 $Y=-0.245 $X2=1.71
+ $Y2=1.985
cc_101 VNB N_A_1790_74#_c_1506_n 0.00223918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1790_74#_c_1507_n 0.021329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2607_392#_M1001_g 0.00188569f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.605
cc_104 VNB N_A_2607_392#_M1018_g 0.023917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2607_392#_M1044_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2607_392#_M1038_g 0.0268211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2607_392#_c_1646_n 0.0652038f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.82
cc_108 VNB N_A_2607_392#_c_1647_n 0.0484968f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.49
cc_109 VNB N_A_2607_392#_c_1648_n 0.0102396f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_110 VNB N_A_2607_392#_c_1649_n 7.2775e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2607_392#_c_1650_n 0.00109231f $X=-0.19 $Y=-0.245 $X2=1.385
+ $Y2=1.985
cc_112 VNB N_VPWR_c_1692_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_388_79#_c_1874_n 0.00214649f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.985
cc_114 VNB N_A_388_79#_c_1875_n 0.0235335f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.62
cc_115 VNB N_A_388_79#_c_1876_n 0.00417762f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.82
cc_116 VNB N_A_388_79#_c_1877_n 0.0041886f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_117 VNB N_A_388_79#_c_1878_n 7.44466e-19 $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=1.985
cc_118 VNB N_A_388_79#_c_1879_n 0.00627051f $X=-0.19 $Y=-0.245 $X2=1.385
+ $Y2=1.985
cc_119 VNB N_A_388_79#_c_1880_n 0.00155036f $X=-0.19 $Y=-0.245 $X2=2.57
+ $Y2=1.455
cc_120 VNB N_A_388_79#_c_1881_n 0.00308378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_388_79#_c_1882_n 0.00182366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB Q_N 0.00143966f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.605
cc_123 VNB N_Q_N_c_2045_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.605
cc_124 VNB N_Q_c_2072_n 0.0065793f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.15
cc_125 VNB N_VGND_c_2088_n 0.0153683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2089_n 0.0218542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2090_n 0.0139145f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.985
cc_128 VNB N_VGND_c_2091_n 0.00692506f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.985
cc_129 VNB N_VGND_c_2092_n 0.00869988f $X=-0.19 $Y=-0.245 $X2=2.57 $Y2=1.29
cc_130 VNB N_VGND_c_2093_n 0.0114612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2094_n 0.0225701f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.985
cc_132 VNB N_VGND_c_2095_n 0.00935384f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.985
cc_133 VNB N_VGND_c_2096_n 0.0108727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2097_n 0.0526431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2098_n 0.0649427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2099_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2100_n 0.0210202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2101_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2102_n 0.0583825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2103_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2104_n 0.0176416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2105_n 0.0276584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2106_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2107_n 0.0186734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2108_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2109_n 0.0605454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2110_n 0.0190049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2111_n 0.00478044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2112_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2113_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2114_n 0.772554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_noxref_25_c_2245_n 0.00622698f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.605
cc_153 VNB N_noxref_25_c_2246_n 0.017862f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_154 VNB N_noxref_25_c_2247_n 0.00386383f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.64
cc_155 VNB N_noxref_25_c_2248_n 0.00276768f $X=-0.19 $Y=-0.245 $X2=2.66
+ $Y2=0.605
cc_156 VPB N_SCE_c_285_n 0.013397f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.82
cc_157 VPB N_SCE_M1009_g 0.0322236f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_158 VPB N_SCE_c_295_n 0.013408f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.15
cc_159 VPB N_SCE_M1039_g 0.0286445f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.64
cc_160 VPB N_SCE_c_297_n 0.0213154f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.82
cc_161 VPB N_SCE_c_289_n 0.00700226f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.82
cc_162 VPB N_SCE_c_299_n 0.0564271f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.985
cc_163 VPB N_SCE_c_300_n 0.00222208f $X=-0.19 $Y=1.66 $X2=1.625 $Y2=1.985
cc_164 VPB N_A_27_79#_M1027_g 0.0292252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_27_79#_c_376_n 0.0311697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_27_79#_c_381_n 0.0211977f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.62
cc_167 VPB N_A_27_79#_c_382_n 0.00448364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_27_79#_c_383_n 0.00938146f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_169 VPB N_A_27_79#_c_384_n 0.0423597f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=1.985
cc_170 VPB N_D_M1006_g 0.057601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_SCD_M1041_g 0.0289341f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.15
cc_172 VPB N_SCD_c_503_n 0.0254895f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.64
cc_173 VPB N_SCD_c_508_n 0.0157901f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.64
cc_174 VPB SCD 0.00164304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_CLK_M1019_g 0.0233373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_CLK_c_548_n 0.0158596f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.15
cc_177 VPB N_A_1025_119#_M1032_g 0.038733f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.605
cc_178 VPB N_A_1025_119#_M1042_g 0.0241316f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.62
cc_179 VPB N_A_1025_119#_c_608_n 0.00192904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1025_119#_c_614_n 0.00266828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1025_119#_c_624_n 0.00660905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1025_119#_c_618_n 0.00417118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1025_119#_c_619_n 0.0160939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1025_119#_c_627_n 0.0316267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1370_290#_M1020_g 0.0455748f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.605
cc_186 VPB N_A_1370_290#_c_804_n 0.00212444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1370_290#_c_805_n 0.0186985f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=0.965
cc_188 VPB N_A_1370_290#_c_812_n 0.00229477f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.62
cc_189 VPB N_A_1370_290#_c_808_n 0.00165919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_M1003_g 0.00640222f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_191 VPB N_RESET_B_M1035_g 0.0339337f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.89
cc_192 VPB N_RESET_B_c_903_n 0.0206024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_RESET_B_c_898_n 0.00910493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_RESET_B_M1023_g 0.0270387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_RESET_B_c_906_n 0.0117122f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.95
cc_196 VPB N_RESET_B_c_900_n 0.00587573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_908_n 0.0214f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.985
cc_198 VPB N_RESET_B_c_909_n 0.00353357f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_199 VPB N_RESET_B_c_910_n 0.00850003f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_200 VPB N_RESET_B_c_911_n 0.00382672f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_201 VPB RESET_B 0.00298374f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_202 VPB N_RESET_B_c_913_n 0.047316f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.985
cc_203 VPB N_RESET_B_c_914_n 0.00208988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_915_n 0.052575f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.985
cc_205 VPB N_RESET_B_c_916_n 0.00231732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_917_n 0.0293981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_918_n 0.0120728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_RESET_B_c_919_n 0.0062794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1223_119#_M1000_g 0.0221395f $X=-0.19 $Y=1.66 $X2=2.66 $Y2=0.605
cc_210 VPB N_A_1223_119#_c_1108_n 0.0117f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.82
cc_211 VPB N_A_1223_119#_c_1115_n 0.00306967f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.82
cc_212 VPB N_A_1223_119#_c_1109_n 0.0151698f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.49
cc_213 VPB N_A_1223_119#_c_1111_n 0.00370269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1223_119#_c_1112_n 0.00500917f $X=-0.19 $Y=1.66 $X2=0.635
+ $Y2=1.95
cc_215 VPB N_A_852_119#_M1036_g 0.0212937f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.64
cc_216 VPB N_A_852_119#_c_1211_n 0.0740476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_852_119#_c_1226_n 0.053782f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.985
cc_218 VPB N_A_852_119#_c_1227_n 0.0106063f $X=-0.19 $Y=1.66 $X2=0.335 $Y2=1.82
cc_219 VPB N_A_852_119#_M1040_g 0.0413704f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.455
cc_220 VPB N_A_852_119#_c_1229_n 0.178706f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.95
cc_221 VPB N_A_852_119#_M1004_g 0.033537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_852_119#_c_1215_n 0.0303876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_852_119#_c_1216_n 0.00223926f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.985
cc_224 VPB N_A_852_119#_c_1233_n 0.00898883f $X=-0.19 $Y=1.66 $X2=1.385
+ $Y2=1.985
cc_225 VPB N_A_852_119#_c_1221_n 0.00511766f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.985
cc_226 VPB N_A_852_119#_c_1222_n 0.0100855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_2006_373#_M1022_g 0.0235027f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.605
cc_228 VPB N_A_2006_373#_M1045_g 0.0146783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_2006_373#_c_1391_n 0.00432037f $X=-0.19 $Y=1.66 $X2=0.41
+ $Y2=0.965
cc_230 VPB N_A_2006_373#_c_1392_n 0.0509674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2006_373#_c_1383_n 0.010942f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.965
cc_232 VPB N_A_2006_373#_c_1394_n 0.00269291f $X=-0.19 $Y=1.66 $X2=0.595
+ $Y2=1.985
cc_233 VPB N_A_2006_373#_c_1395_n 2.01178e-19 $X=-0.19 $Y=1.66 $X2=0.335
+ $Y2=1.82
cc_234 VPB N_A_2006_373#_c_1396_n 0.00556561f $X=-0.19 $Y=1.66 $X2=1.115
+ $Y2=1.95
cc_235 VPB N_A_1790_74#_M1028_g 0.0550921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1790_74#_M1005_g 0.0263295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1790_74#_M1008_g 0.0256608f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.49
cc_238 VPB N_A_1790_74#_M1029_g 0.0326348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1790_74#_c_1506_n 0.00736766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_2607_392#_M1001_g 0.025951f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.605
cc_241 VPB N_A_2607_392#_M1044_g 0.0274054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_2607_392#_c_1649_n 0.0194246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1693_n 0.00400995f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.95
cc_244 VPB N_VPWR_c_1694_n 0.00151893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1695_n 0.00801002f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_246 VPB N_VPWR_c_1696_n 0.0134255f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.455
cc_247 VPB N_VPWR_c_1697_n 0.0511217f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_248 VPB N_VPWR_c_1698_n 0.0223473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1699_n 0.0116888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1700_n 0.018127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1701_n 0.0109102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1702_n 0.0663346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1703_n 0.0330761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1704_n 0.00485379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1705_n 0.0565844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1706_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1707_n 0.0467369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1708_n 0.0237904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1709_n 0.0217361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1710_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1711_n 0.0206736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1712_n 0.0174144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1713_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1714_n 0.0261837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1715_n 0.00547828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1716_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1717_n 0.0389124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1718_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1719_n 0.00555219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1720_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1692_n 0.123152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_388_79#_c_1883_n 0.0069063f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.455
cc_273 VPB N_A_388_79#_c_1884_n 0.0073678f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.455
cc_274 VPB N_A_388_79#_c_1877_n 0.00479889f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.95
cc_275 VPB N_A_388_79#_c_1886_n 0.00507435f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.95
cc_276 VPB N_A_388_79#_c_1887_n 0.00868256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_388_79#_c_1888_n 0.0111306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_388_79#_c_1889_n 0.00619901f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.985
cc_279 VPB N_A_388_79#_c_1890_n 0.00574222f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.985
cc_280 VPB N_A_388_79#_c_1891_n 0.00191389f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=1.985
cc_281 VPB N_A_388_79#_c_1881_n 0.0054728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB Q_N 0.00231613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.605
cc_283 VPB N_Q_c_2072_n 0.00391262f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.15
cc_284 N_SCE_c_285_n N_A_27_79#_c_374_n 0.0181735f $X=0.41 $Y=1.82 $X2=0 $Y2=0
cc_285 N_SCE_c_290_n N_A_27_79#_c_374_n 0.00219996f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_286 N_SCE_c_299_n N_A_27_79#_c_374_n 0.0452379f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_287 N_SCE_c_300_n N_A_27_79#_c_374_n 0.00363355f $X=1.625 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_SCE_c_285_n N_A_27_79#_c_375_n 0.0127444f $X=0.41 $Y=1.82 $X2=0 $Y2=0
cc_289 N_SCE_c_286_n N_A_27_79#_c_375_n 0.00367837f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_290 N_SCE_c_288_n N_A_27_79#_c_375_n 0.0100023f $X=0.495 $Y=0.965 $X2=0 $Y2=0
cc_291 N_SCE_c_285_n N_A_27_79#_c_376_n 0.0140797f $X=0.41 $Y=1.82 $X2=0 $Y2=0
cc_292 N_SCE_c_297_n N_A_27_79#_c_376_n 0.0113427f $X=0.335 $Y=1.82 $X2=0 $Y2=0
cc_293 N_SCE_c_300_n N_A_27_79#_c_376_n 0.0192999f $X=1.625 $Y=1.985 $X2=0 $Y2=0
cc_294 N_SCE_M1009_g N_A_27_79#_c_381_n 0.0165225f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_295 N_SCE_c_285_n N_A_27_79#_c_377_n 0.0179853f $X=0.41 $Y=1.82 $X2=0 $Y2=0
cc_296 N_SCE_c_288_n N_A_27_79#_c_377_n 0.00327315f $X=0.495 $Y=0.965 $X2=0
+ $Y2=0
cc_297 N_SCE_c_297_n N_A_27_79#_c_377_n 0.00680735f $X=0.335 $Y=1.82 $X2=0 $Y2=0
cc_298 N_SCE_c_290_n N_A_27_79#_c_377_n 0.0155382f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_299 N_SCE_c_299_n N_A_27_79#_c_377_n 0.00253102f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_300 N_SCE_c_300_n N_A_27_79#_c_377_n 0.0494351f $X=1.625 $Y=1.985 $X2=0 $Y2=0
cc_301 N_SCE_M1009_g N_A_27_79#_c_402_n 0.0146414f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_302 N_SCE_M1039_g N_A_27_79#_c_402_n 0.0150497f $X=1.46 $Y=2.64 $X2=0 $Y2=0
cc_303 N_SCE_c_289_n N_A_27_79#_c_402_n 0.0119714f $X=1.71 $Y=1.82 $X2=0 $Y2=0
cc_304 N_SCE_c_299_n N_A_27_79#_c_402_n 0.0133402f $X=1.37 $Y=1.985 $X2=0 $Y2=0
cc_305 N_SCE_c_300_n N_A_27_79#_c_402_n 0.0735258f $X=1.625 $Y=1.985 $X2=0 $Y2=0
cc_306 N_SCE_c_289_n N_A_27_79#_c_382_n 0.0109466f $X=1.71 $Y=1.82 $X2=0 $Y2=0
cc_307 N_SCE_c_291_n N_A_27_79#_c_382_n 0.0221869f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_308 N_SCE_c_292_n N_A_27_79#_c_382_n 7.02495e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_309 N_SCE_c_285_n N_A_27_79#_c_378_n 0.00851213f $X=0.41 $Y=1.82 $X2=0 $Y2=0
cc_310 N_SCE_M1009_g N_A_27_79#_c_383_n 0.00469442f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_311 N_SCE_c_297_n N_A_27_79#_c_383_n 0.00204858f $X=0.335 $Y=1.82 $X2=0 $Y2=0
cc_312 N_SCE_c_289_n N_A_27_79#_c_384_n 0.00102331f $X=1.71 $Y=1.82 $X2=0 $Y2=0
cc_313 N_SCE_c_291_n N_A_27_79#_c_384_n 0.00193233f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_314 N_SCE_c_292_n N_A_27_79#_c_384_n 0.0202959f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_315 N_SCE_c_295_n N_D_M1006_g 0.0707626f $X=1.46 $Y=2.15 $X2=0 $Y2=0
cc_316 N_SCE_M1031_g N_D_M1006_g 8.48778e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_317 N_SCE_c_289_n N_D_M1006_g 0.0203296f $X=1.71 $Y=1.82 $X2=0 $Y2=0
cc_318 N_SCE_c_290_n N_D_M1006_g 0.00239218f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_319 N_SCE_c_291_n N_D_M1006_g 0.0189196f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_320 N_SCE_c_292_n N_D_M1006_g 0.00894005f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_321 N_SCE_M1031_g N_D_c_459_n 0.00730331f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_322 N_SCE_c_290_n N_D_c_459_n 7.56204e-19 $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_323 N_SCE_c_291_n N_D_c_459_n 0.002936f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_324 N_SCE_M1031_g N_D_c_460_n 5.42624e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_325 N_SCE_c_290_n N_D_c_460_n 0.0150217f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_326 N_SCE_c_291_n N_D_c_460_n 0.0224216f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_327 N_SCE_c_300_n N_D_c_460_n 0.0020111f $X=1.625 $Y=1.985 $X2=0 $Y2=0
cc_328 N_SCE_M1031_g N_D_c_461_n 0.00705002f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_329 N_SCE_M1031_g N_SCD_M1013_g 0.0628756f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_330 N_SCE_c_291_n N_SCD_M1013_g 5.04484e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_331 N_SCE_c_291_n SCD 0.0120234f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_332 N_SCE_c_292_n SCD 2.2546e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_333 N_SCE_c_291_n N_SCD_c_505_n 6.19299e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_334 N_SCE_c_292_n N_SCD_c_505_n 0.0113035f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_335 N_SCE_M1039_g N_VPWR_c_1707_n 0.00460063f $X=1.46 $Y=2.64 $X2=0 $Y2=0
cc_336 N_SCE_M1009_g N_VPWR_c_1713_n 0.005209f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_337 N_SCE_M1009_g N_VPWR_c_1714_n 0.00586566f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_338 N_SCE_M1039_g N_VPWR_c_1714_n 0.0112164f $X=1.46 $Y=2.64 $X2=0 $Y2=0
cc_339 N_SCE_M1009_g N_VPWR_c_1692_n 0.00541102f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_340 N_SCE_M1039_g N_VPWR_c_1692_n 0.00459004f $X=1.46 $Y=2.64 $X2=0 $Y2=0
cc_341 N_SCE_M1039_g N_A_388_79#_c_1893_n 8.35527e-19 $X=1.46 $Y=2.64 $X2=0
+ $Y2=0
cc_342 N_SCE_M1031_g N_A_388_79#_c_1874_n 0.0103246f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_343 N_SCE_M1031_g N_A_388_79#_c_1875_n 0.0087327f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_344 N_SCE_c_291_n N_A_388_79#_c_1875_n 0.00815275f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_345 N_SCE_M1031_g N_A_388_79#_c_1876_n 0.00327429f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_346 N_SCE_c_291_n N_A_388_79#_c_1876_n 0.0273677f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_347 N_SCE_c_292_n N_A_388_79#_c_1876_n 0.00449985f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_348 N_SCE_c_286_n N_VGND_c_2088_n 0.0143331f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_349 N_SCE_M1031_g N_VGND_c_2098_n 9.44495e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_350 N_SCE_c_286_n N_VGND_c_2104_n 0.00465077f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_351 N_SCE_c_286_n N_VGND_c_2114_n 0.00451796f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_352 N_SCE_c_286_n N_noxref_25_c_2245_n 7.27954e-19 $X=0.495 $Y=0.89 $X2=0
+ $Y2=0
cc_353 N_SCE_M1031_g N_noxref_25_c_2246_n 0.0128121f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_354 N_SCE_c_286_n N_noxref_25_c_2247_n 6.46792e-19 $X=0.495 $Y=0.89 $X2=0
+ $Y2=0
cc_355 N_SCE_M1031_g N_noxref_25_c_2248_n 0.00151906f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_356 N_A_27_79#_M1027_g N_D_M1006_g 0.0188494f $X=2.615 $Y=2.735 $X2=0 $Y2=0
cc_357 N_A_27_79#_c_374_n N_D_M1006_g 0.0185925f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_358 N_A_27_79#_c_377_n N_D_M1006_g 6.63701e-19 $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_359 N_A_27_79#_c_402_n N_D_M1006_g 0.0193772f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_360 N_A_27_79#_c_382_n N_D_M1006_g 0.00486063f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_361 N_A_27_79#_c_384_n N_D_M1006_g 0.0131037f $X=2.615 $Y=1.995 $X2=0 $Y2=0
cc_362 N_A_27_79#_M1012_g N_D_c_459_n 0.0200462f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_363 N_A_27_79#_M1012_g N_D_c_460_n 0.0109288f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_364 N_A_27_79#_M1012_g N_D_c_461_n 0.03521f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_365 N_A_27_79#_c_382_n N_SCD_c_503_n 0.0018886f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_366 N_A_27_79#_c_384_n N_SCD_c_503_n 0.035979f $X=2.615 $Y=1.995 $X2=0 $Y2=0
cc_367 N_A_27_79#_M1027_g N_SCD_c_508_n 0.035979f $X=2.615 $Y=2.735 $X2=0 $Y2=0
cc_368 N_A_27_79#_c_382_n SCD 0.0137339f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_369 N_A_27_79#_c_384_n SCD 0.00131174f $X=2.615 $Y=1.995 $X2=0 $Y2=0
cc_370 N_A_27_79#_c_402_n N_VPWR_M1009_d 0.0174232f $X=2.275 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_371 N_A_27_79#_M1027_g N_VPWR_c_1693_n 0.00170506f $X=2.615 $Y=2.735 $X2=0
+ $Y2=0
cc_372 N_A_27_79#_M1027_g N_VPWR_c_1707_n 0.00433125f $X=2.615 $Y=2.735 $X2=0
+ $Y2=0
cc_373 N_A_27_79#_c_381_n N_VPWR_c_1713_n 0.0145339f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_374 N_A_27_79#_c_381_n N_VPWR_c_1714_n 0.0102732f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_375 N_A_27_79#_c_402_n N_VPWR_c_1714_n 0.0409307f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_376 N_A_27_79#_M1027_g N_VPWR_c_1692_n 0.006833f $X=2.615 $Y=2.735 $X2=0
+ $Y2=0
cc_377 N_A_27_79#_c_381_n N_VPWR_c_1692_n 0.0119683f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_378 N_A_27_79#_c_402_n N_VPWR_c_1692_n 0.024692f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_379 N_A_27_79#_c_402_n A_310_464# 0.00387309f $X=2.275 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_79#_c_402_n N_A_388_79#_M1006_d 0.0157235f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_381 N_A_27_79#_M1027_g N_A_388_79#_c_1893_n 0.0197662f $X=2.615 $Y=2.735
+ $X2=0 $Y2=0
cc_382 N_A_27_79#_c_402_n N_A_388_79#_c_1893_n 0.0418114f $X=2.275 $Y=2.405
+ $X2=0 $Y2=0
cc_383 N_A_27_79#_c_384_n N_A_388_79#_c_1893_n 8.16359e-19 $X=2.615 $Y=1.995
+ $X2=0 $Y2=0
cc_384 N_A_27_79#_M1027_g N_A_388_79#_c_1904_n 0.00318734f $X=2.615 $Y=2.735
+ $X2=0 $Y2=0
cc_385 N_A_27_79#_M1027_g N_A_388_79#_c_1884_n 0.00218468f $X=2.615 $Y=2.735
+ $X2=0 $Y2=0
cc_386 N_A_27_79#_c_402_n N_A_388_79#_c_1884_n 0.0150238f $X=2.275 $Y=2.405
+ $X2=0 $Y2=0
cc_387 N_A_27_79#_M1012_g N_VGND_c_2088_n 5.90987e-19 $X=1.475 $Y=0.605 $X2=0
+ $Y2=0
cc_388 N_A_27_79#_c_374_n N_VGND_c_2088_n 0.00297438f $X=1.4 $Y=1.415 $X2=0
+ $Y2=0
cc_389 N_A_27_79#_c_375_n N_VGND_c_2088_n 0.0179429f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_390 N_A_27_79#_c_377_n N_VGND_c_2088_n 0.0148785f $X=1.23 $Y=1.415 $X2=0
+ $Y2=0
cc_391 N_A_27_79#_M1012_g N_VGND_c_2098_n 9.44495e-19 $X=1.475 $Y=0.605 $X2=0
+ $Y2=0
cc_392 N_A_27_79#_c_375_n N_VGND_c_2104_n 0.0100552f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_393 N_A_27_79#_c_375_n N_VGND_c_2114_n 0.00902019f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_394 N_A_27_79#_M1012_g N_noxref_25_c_2245_n 7.43016e-19 $X=1.475 $Y=0.605
+ $X2=0 $Y2=0
cc_395 N_A_27_79#_c_374_n N_noxref_25_c_2245_n 0.0048989f $X=1.4 $Y=1.415 $X2=0
+ $Y2=0
cc_396 N_A_27_79#_c_377_n N_noxref_25_c_2245_n 0.0106151f $X=1.23 $Y=1.415 $X2=0
+ $Y2=0
cc_397 N_A_27_79#_M1012_g N_noxref_25_c_2246_n 0.0154771f $X=1.475 $Y=0.605
+ $X2=0 $Y2=0
cc_398 N_D_M1006_g N_VPWR_c_1707_n 0.00521639f $X=1.88 $Y=2.64 $X2=0 $Y2=0
cc_399 N_D_M1006_g N_VPWR_c_1714_n 0.00138135f $X=1.88 $Y=2.64 $X2=0 $Y2=0
cc_400 N_D_M1006_g N_VPWR_c_1692_n 0.00538914f $X=1.88 $Y=2.64 $X2=0 $Y2=0
cc_401 N_D_c_460_n N_A_388_79#_M1026_d 0.00145733f $X=1.925 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_402 N_D_M1006_g N_A_388_79#_c_1893_n 0.0101718f $X=1.88 $Y=2.64 $X2=0 $Y2=0
cc_403 N_D_c_459_n N_A_388_79#_c_1874_n 3.29098e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_404 N_D_c_460_n N_A_388_79#_c_1874_n 0.0164816f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_405 N_D_c_461_n N_A_388_79#_c_1874_n 0.00523412f $X=1.925 $Y=0.925 $X2=0
+ $Y2=0
cc_406 N_D_c_459_n N_A_388_79#_c_1876_n 7.8315e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_407 N_D_c_460_n N_A_388_79#_c_1876_n 0.0148785f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_408 N_D_c_461_n N_VGND_c_2098_n 9.44495e-19 $X=1.925 $Y=0.925 $X2=0 $Y2=0
cc_409 N_D_c_460_n N_noxref_25_c_2245_n 0.00134475f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_410 N_D_c_459_n N_noxref_25_c_2246_n 5.75063e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_411 N_D_c_460_n N_noxref_25_c_2246_n 0.0127007f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_412 N_D_c_461_n N_noxref_25_c_2246_n 0.0123465f $X=1.925 $Y=0.925 $X2=0 $Y2=0
cc_413 N_D_c_460_n noxref_26 0.00197445f $X=1.925 $Y=1.09 $X2=-0.19 $Y2=-0.245
cc_414 N_SCD_M1013_g N_RESET_B_M1003_g 0.0292104f $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_415 SCD N_RESET_B_M1003_g 7.60177e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_416 N_SCD_c_505_n N_RESET_B_M1003_g 0.0196966f $X=3.11 $Y=1.605 $X2=0 $Y2=0
cc_417 N_SCD_M1041_g N_RESET_B_c_906_n 0.0257661f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_418 N_SCD_c_503_n N_RESET_B_c_906_n 0.0196966f $X=3.11 $Y=1.945 $X2=0 $Y2=0
cc_419 N_SCD_M1041_g N_VPWR_c_1693_n 0.0110718f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_420 N_SCD_M1041_g N_VPWR_c_1707_n 0.00616631f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_421 N_SCD_M1041_g N_VPWR_c_1692_n 0.00573258f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_422 N_SCD_M1041_g N_A_388_79#_c_1893_n 0.00244336f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_423 N_SCD_M1013_g N_A_388_79#_c_1874_n 0.00151803f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_424 N_SCD_M1013_g N_A_388_79#_c_1875_n 0.0127975f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_425 SCD N_A_388_79#_c_1875_n 0.0182456f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_426 N_SCD_c_505_n N_A_388_79#_c_1875_n 0.00113125f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_427 N_SCD_M1041_g N_A_388_79#_c_1883_n 0.0127324f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_428 N_SCD_c_508_n N_A_388_79#_c_1883_n 9.39545e-19 $X=3.11 $Y=2.11 $X2=0
+ $Y2=0
cc_429 SCD N_A_388_79#_c_1883_n 0.0266083f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_430 N_SCD_M1041_g N_A_388_79#_c_1884_n 0.00137019f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_431 N_SCD_M1041_g N_A_388_79#_c_1877_n 0.0031637f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_432 N_SCD_M1013_g N_A_388_79#_c_1877_n 0.00475298f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_433 SCD N_A_388_79#_c_1877_n 0.0534506f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_434 N_SCD_c_505_n N_A_388_79#_c_1877_n 0.00361663f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_435 N_SCD_M1041_g N_A_388_79#_c_1886_n 2.4222e-19 $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_436 N_SCD_M1013_g N_VGND_c_2089_n 2.27924e-19 $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_437 N_SCD_M1013_g N_VGND_c_2098_n 9.63557e-19 $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_438 N_SCD_M1013_g N_noxref_25_c_2246_n 0.0110567f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_439 N_SCD_M1013_g N_noxref_25_c_2248_n 0.00775324f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_440 N_CLK_M1019_g N_A_1025_119#_c_614_n 9.15039e-19 $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_441 N_CLK_c_548_n N_RESET_B_M1003_g 0.00289883f $X=4.62 $Y=1.61 $X2=0 $Y2=0
cc_442 CLK N_RESET_B_M1003_g 0.00168117f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_443 N_CLK_c_550_n N_RESET_B_M1003_g 0.0410462f $X=4.02 $Y=1.105 $X2=0 $Y2=0
cc_444 N_CLK_c_547_n N_RESET_B_c_893_n 0.0102747f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_445 N_CLK_c_550_n N_RESET_B_c_893_n 0.00658273f $X=4.02 $Y=1.105 $X2=0 $Y2=0
cc_446 N_CLK_M1019_g N_RESET_B_c_908_n 0.00239013f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_447 N_CLK_c_548_n N_RESET_B_c_908_n 0.00244269f $X=4.62 $Y=1.61 $X2=0 $Y2=0
cc_448 CLK N_RESET_B_c_908_n 3.47655e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_449 N_CLK_c_548_n N_RESET_B_c_909_n 0.00162803f $X=4.62 $Y=1.61 $X2=0 $Y2=0
cc_450 CLK N_RESET_B_c_909_n 0.00379332f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_451 N_CLK_M1019_g N_RESET_B_c_913_n 0.00538416f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_452 N_CLK_c_548_n N_RESET_B_c_913_n 0.0169131f $X=4.62 $Y=1.61 $X2=0 $Y2=0
cc_453 CLK N_RESET_B_c_913_n 8.25778e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_454 N_CLK_M1019_g N_RESET_B_c_914_n 4.97287e-19 $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_455 N_CLK_c_548_n N_RESET_B_c_914_n 0.00239604f $X=4.62 $Y=1.61 $X2=0 $Y2=0
cc_456 CLK N_RESET_B_c_914_n 0.0153258f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_M1019_g N_A_852_119#_M1036_g 0.0498506f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_458 N_CLK_M1019_g N_A_852_119#_c_1237_n 0.00532664f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_459 N_CLK_c_547_n N_A_852_119#_c_1219_n 0.012222f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_460 CLK N_A_852_119#_c_1219_n 0.0348825f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_461 N_CLK_c_550_n N_A_852_119#_c_1219_n 0.00268145f $X=4.02 $Y=1.105 $X2=0
+ $Y2=0
cc_462 N_CLK_c_547_n N_A_852_119#_c_1220_n 0.0032892f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_463 N_CLK_c_548_n N_A_852_119#_c_1220_n 0.00322677f $X=4.62 $Y=1.61 $X2=0
+ $Y2=0
cc_464 N_CLK_M1019_g N_A_852_119#_c_1221_n 0.0102555f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_465 N_CLK_c_548_n N_A_852_119#_c_1221_n 0.0400324f $X=4.62 $Y=1.61 $X2=0
+ $Y2=0
cc_466 CLK N_A_852_119#_c_1221_n 0.00843065f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_467 N_CLK_c_548_n N_A_852_119#_c_1222_n 0.0182297f $X=4.62 $Y=1.61 $X2=0
+ $Y2=0
cc_468 N_CLK_c_547_n N_A_852_119#_c_1223_n 0.0108777f $X=4.62 $Y=1.445 $X2=0
+ $Y2=0
cc_469 N_CLK_M1019_g N_VPWR_c_1694_n 0.017461f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_470 N_CLK_M1019_g N_VPWR_c_1703_n 0.00401239f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_471 N_CLK_M1019_g N_VPWR_c_1692_n 0.00589267f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_472 CLK N_A_388_79#_c_1875_n 0.0103709f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_473 N_CLK_c_550_n N_A_388_79#_c_1875_n 2.01872e-19 $X=4.02 $Y=1.105 $X2=0
+ $Y2=0
cc_474 N_CLK_c_548_n N_A_388_79#_c_1877_n 4.40341e-19 $X=4.62 $Y=1.61 $X2=0
+ $Y2=0
cc_475 CLK N_A_388_79#_c_1877_n 0.0205304f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_476 N_CLK_c_550_n N_A_388_79#_c_1877_n 4.5243e-19 $X=4.02 $Y=1.105 $X2=0
+ $Y2=0
cc_477 N_CLK_M1019_g N_A_388_79#_c_1886_n 0.00348169f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_478 N_CLK_M1019_g N_A_388_79#_c_1887_n 0.0110051f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_479 N_CLK_M1019_g N_A_388_79#_c_1888_n 0.0171874f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_480 N_CLK_c_548_n N_A_388_79#_c_1888_n 6.38984e-19 $X=4.62 $Y=1.61 $X2=0
+ $Y2=0
cc_481 N_CLK_c_547_n N_VGND_c_2089_n 0.00342867f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_482 CLK N_VGND_c_2089_n 0.00995577f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_483 N_CLK_c_550_n N_VGND_c_2089_n 0.00167099f $X=4.02 $Y=1.105 $X2=0 $Y2=0
cc_484 N_CLK_c_547_n N_VGND_c_2090_n 0.00294829f $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_485 N_CLK_c_547_n N_VGND_c_2114_n 9.39239e-19 $X=4.62 $Y=1.445 $X2=0 $Y2=0
cc_486 N_A_1025_119#_c_610_n N_A_1370_290#_M1007_d 0.00176891f $X=9.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_487 N_A_1025_119#_M1032_g N_A_1370_290#_M1020_g 0.00379368f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_488 N_A_1025_119#_M1015_g N_A_1370_290#_M1043_g 0.0462355f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_489 N_A_1025_119#_c_606_n N_A_1370_290#_M1043_g 0.00762221f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_490 N_A_1025_119#_c_615_n N_A_1370_290#_M1043_g 0.00542036f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_491 N_A_1025_119#_M1015_g N_A_1370_290#_c_805_n 0.0105382f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_492 N_A_1025_119#_c_615_n N_A_1370_290#_c_805_n 3.83611e-19 $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_493 N_A_1025_119#_c_619_n N_A_1370_290#_c_805_n 0.00192784f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_494 N_A_1025_119#_c_609_n N_A_1370_290#_c_822_n 0.00146445f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_495 N_A_1025_119#_c_615_n N_A_1370_290#_c_822_n 0.00967347f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_496 N_A_1025_119#_c_624_n N_A_1370_290#_c_824_n 0.0194909f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_497 N_A_1025_119#_c_627_n N_A_1370_290#_c_824_n 3.80268e-19 $X=9.7 $Y=2.03
+ $X2=0 $Y2=0
cc_498 N_A_1025_119#_M1042_g N_A_1370_290#_c_812_n 0.00121316f $X=9.7 $Y=2.565
+ $X2=0 $Y2=0
cc_499 N_A_1025_119#_c_609_n N_A_1370_290#_c_806_n 0.0737203f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_500 N_A_1025_119#_c_610_n N_A_1370_290#_c_806_n 0.00353238f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_501 N_A_1025_119#_c_601_n N_A_1370_290#_c_807_n 0.0114651f $X=8.875 $Y=1.085
+ $X2=0 $Y2=0
cc_502 N_A_1025_119#_c_603_n N_A_1370_290#_c_807_n 4.45722e-19 $X=8.95 $Y=1.16
+ $X2=0 $Y2=0
cc_503 N_A_1025_119#_c_610_n N_A_1370_290#_c_807_n 0.0229775f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_504 N_A_1025_119#_c_612_n N_A_1370_290#_c_807_n 0.0234316f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_505 N_A_1025_119#_c_616_n N_A_1370_290#_c_807_n 0.0157507f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_506 N_A_1025_119#_c_603_n N_A_1370_290#_c_808_n 0.006971f $X=8.95 $Y=1.16
+ $X2=0 $Y2=0
cc_507 N_A_1025_119#_c_616_n N_A_1370_290#_c_808_n 0.0107601f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_508 N_A_1025_119#_c_618_n N_A_1370_290#_c_808_n 0.0194909f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_509 N_A_1025_119#_M1015_g N_RESET_B_c_893_n 0.00880557f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_510 N_A_1025_119#_c_606_n N_RESET_B_c_893_n 0.0286159f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_511 N_A_1025_119#_c_607_n N_RESET_B_c_893_n 0.00755311f $X=5.43 $Y=0.395
+ $X2=0 $Y2=0
cc_512 N_A_1025_119#_c_615_n N_RESET_B_c_893_n 0.00357516f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_513 N_A_1025_119#_c_609_n N_RESET_B_M1011_g 0.0123884f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_514 N_A_1025_119#_c_615_n N_RESET_B_M1011_g 0.00727728f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_515 N_A_1025_119#_M1032_g N_RESET_B_c_908_n 0.00324919f $X=6.1 $Y=2.495 $X2=0
+ $Y2=0
cc_516 N_A_1025_119#_c_599_n N_RESET_B_c_908_n 0.00395271f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_517 N_A_1025_119#_c_608_n N_RESET_B_c_908_n 0.0134589f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_A_1025_119#_c_614_n N_RESET_B_c_908_n 0.0302208f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_519 N_A_1025_119#_c_619_n N_RESET_B_c_908_n 0.00369615f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_520 N_A_1025_119#_c_624_n N_RESET_B_c_910_n 0.0277328f $X=9.615 $Y=2.03 $X2=0
+ $Y2=0
cc_521 N_A_1025_119#_c_627_n N_RESET_B_c_910_n 0.00172094f $X=9.7 $Y=2.03 $X2=0
+ $Y2=0
cc_522 N_A_1025_119#_c_601_n N_A_1223_119#_M1007_g 0.0264029f $X=8.875 $Y=1.085
+ $X2=0 $Y2=0
cc_523 N_A_1025_119#_c_610_n N_A_1223_119#_M1007_g 0.0116384f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_524 N_A_1025_119#_c_599_n N_A_1223_119#_c_1121_n 6.10614e-19 $X=6.465
+ $Y=1.575 $X2=0 $Y2=0
cc_525 N_A_1025_119#_M1015_g N_A_1223_119#_c_1121_n 0.0146944f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_526 N_A_1025_119#_c_606_n N_A_1223_119#_c_1121_n 0.0431682f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_527 N_A_1025_119#_M1032_g N_A_1223_119#_c_1108_n 4.75534e-19 $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_528 N_A_1025_119#_M1015_g N_A_1223_119#_c_1108_n 0.00527914f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_529 N_A_1025_119#_M1032_g N_A_1223_119#_c_1115_n 0.00542781f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_530 N_A_1025_119#_c_599_n N_A_1223_119#_c_1115_n 0.00104855f $X=6.465
+ $Y=1.575 $X2=0 $Y2=0
cc_531 N_A_1025_119#_c_614_n N_A_852_119#_M1036_g 0.00764891f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_1025_119#_c_605_n N_A_852_119#_c_1209_n 0.00171313f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_533 N_A_1025_119#_c_614_n N_A_852_119#_c_1209_n 0.00704878f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_A_1025_119#_c_605_n N_A_852_119#_c_1210_n 0.00750167f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_535 N_A_1025_119#_c_613_n N_A_852_119#_c_1210_n 9.35297e-19 $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_536 N_A_1025_119#_M1032_g N_A_852_119#_c_1211_n 0.0271806f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_537 N_A_1025_119#_c_608_n N_A_852_119#_c_1211_n 0.00321388f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_1025_119#_c_614_n N_A_852_119#_c_1211_n 0.0189097f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_1025_119#_c_608_n N_A_852_119#_c_1212_n 0.00583367f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_1025_119#_c_619_n N_A_852_119#_c_1212_n 0.0127953f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_541 N_A_1025_119#_c_606_n N_A_852_119#_c_1213_n 0.00109326f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_542 N_A_1025_119#_c_613_n N_A_852_119#_c_1213_n 0.00835221f $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_543 N_A_1025_119#_M1032_g N_A_852_119#_c_1226_n 0.0107339f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_544 N_A_1025_119#_M1015_g N_A_852_119#_c_1214_n 0.0198517f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_545 N_A_1025_119#_c_604_n N_A_852_119#_c_1214_n 0.00427994f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_546 N_A_1025_119#_c_606_n N_A_852_119#_c_1214_n 0.00544855f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_547 N_A_1025_119#_c_613_n N_A_852_119#_c_1214_n 6.53033e-19 $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_548 N_A_1025_119#_M1032_g N_A_852_119#_M1040_g 0.0149938f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_549 N_A_1025_119#_c_599_n N_A_852_119#_M1040_g 0.00392883f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_550 N_A_1025_119#_M1042_g N_A_852_119#_M1004_g 0.0137144f $X=9.7 $Y=2.565
+ $X2=0 $Y2=0
cc_551 N_A_1025_119#_c_618_n N_A_852_119#_M1004_g 0.00731328f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_552 N_A_1025_119#_c_627_n N_A_852_119#_M1004_g 0.00884985f $X=9.7 $Y=2.03
+ $X2=0 $Y2=0
cc_553 N_A_1025_119#_c_602_n N_A_852_119#_c_1215_n 0.0219012f $X=9.31 $Y=1.16
+ $X2=0 $Y2=0
cc_554 N_A_1025_119#_c_616_n N_A_852_119#_c_1215_n 0.00157771f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_555 N_A_1025_119#_c_624_n N_A_852_119#_c_1215_n 7.40372e-19 $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_556 N_A_1025_119#_c_618_n N_A_852_119#_c_1215_n 0.0190498f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_557 N_A_1025_119#_c_627_n N_A_852_119#_c_1215_n 0.0185219f $X=9.7 $Y=2.03
+ $X2=0 $Y2=0
cc_558 N_A_1025_119#_c_603_n N_A_852_119#_c_1216_n 0.0219012f $X=8.95 $Y=1.16
+ $X2=0 $Y2=0
cc_559 N_A_1025_119#_c_610_n N_A_852_119#_M1002_g 0.00370958f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_560 N_A_1025_119#_c_612_n N_A_852_119#_M1002_g 0.00214927f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_561 N_A_1025_119#_c_616_n N_A_852_119#_M1002_g 0.00105258f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_562 N_A_1025_119#_c_617_n N_A_852_119#_M1002_g 0.0196932f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_563 N_A_1025_119#_c_618_n N_A_852_119#_M1002_g 0.00477388f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_564 N_A_1025_119#_c_605_n N_A_852_119#_c_1218_n 0.00158285f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_565 N_A_1025_119#_c_608_n N_A_852_119#_c_1218_n 0.00213243f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_566 N_A_1025_119#_c_614_n N_A_852_119#_c_1218_n 0.0011182f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_1025_119#_c_619_n N_A_852_119#_c_1218_n 0.0214031f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_568 N_A_1025_119#_c_614_n N_A_852_119#_c_1237_n 0.0060972f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_A_1025_119#_c_605_n N_A_852_119#_c_1221_n 0.00425568f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_570 N_A_1025_119#_c_613_n N_A_852_119#_c_1221_n 0.00806769f $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_571 N_A_1025_119#_c_614_n N_A_852_119#_c_1221_n 0.037353f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_572 N_A_1025_119#_c_613_n N_A_852_119#_c_1222_n 0.00463303f $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_573 N_A_1025_119#_c_614_n N_A_852_119#_c_1222_n 0.00322316f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_574 N_A_1025_119#_c_604_n N_A_852_119#_c_1223_n 0.00761662f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_575 N_A_1025_119#_c_605_n N_A_852_119#_c_1223_n 0.0033477f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_576 N_A_1025_119#_c_607_n N_A_852_119#_c_1223_n 6.62904e-19 $X=5.43 $Y=0.395
+ $X2=0 $Y2=0
cc_577 N_A_1025_119#_c_613_n N_A_852_119#_c_1223_n 0.00334503f $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_578 N_A_1025_119#_M1042_g N_A_2006_373#_M1022_g 0.0282074f $X=9.7 $Y=2.565
+ $X2=0 $Y2=0
cc_579 N_A_1025_119#_c_624_n N_A_2006_373#_c_1392_n 3.95315e-19 $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_580 N_A_1025_119#_c_627_n N_A_2006_373#_c_1392_n 0.0282074f $X=9.7 $Y=2.03
+ $X2=0 $Y2=0
cc_581 N_A_1025_119#_c_610_n N_A_1790_74#_M1017_d 0.00293623f $X=9.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_582 N_A_1025_119#_c_612_n N_A_1790_74#_M1017_d 0.0113447f $X=9.185 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_583 N_A_1025_119#_c_616_n N_A_1790_74#_M1017_d 0.00118465f $X=9.475 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_584 N_A_1025_119#_M1042_g N_A_1790_74#_c_1516_n 0.0207832f $X=9.7 $Y=2.565
+ $X2=0 $Y2=0
cc_585 N_A_1025_119#_c_624_n N_A_1790_74#_c_1516_n 0.0316643f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_586 N_A_1025_119#_c_627_n N_A_1790_74#_c_1516_n 0.0010406f $X=9.7 $Y=2.03
+ $X2=0 $Y2=0
cc_587 N_A_1025_119#_c_601_n N_A_1790_74#_c_1519_n 5.95394e-19 $X=8.875 $Y=1.085
+ $X2=0 $Y2=0
cc_588 N_A_1025_119#_c_610_n N_A_1790_74#_c_1519_n 0.00170833f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_589 N_A_1025_119#_c_612_n N_A_1790_74#_c_1519_n 0.0250265f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_590 N_A_1025_119#_c_616_n N_A_1790_74#_c_1519_n 0.0155252f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_591 N_A_1025_119#_c_617_n N_A_1790_74#_c_1519_n 0.00455646f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_592 N_A_1025_119#_c_612_n N_A_1790_74#_c_1505_n 0.00427034f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_593 N_A_1025_119#_c_616_n N_A_1790_74#_c_1505_n 0.00683662f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_594 N_A_1025_119#_c_624_n N_A_1790_74#_c_1506_n 0.0241297f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_595 N_A_1025_119#_c_618_n N_A_1790_74#_c_1506_n 0.0288004f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_596 N_A_1025_119#_c_627_n N_A_1790_74#_c_1506_n 0.00541216f $X=9.7 $Y=2.03
+ $X2=0 $Y2=0
cc_597 N_A_1025_119#_c_616_n N_A_1790_74#_c_1529_n 0.0103633f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_598 N_A_1025_119#_c_617_n N_A_1790_74#_c_1529_n 2.09861e-19 $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_599 N_A_1025_119#_c_618_n N_A_1790_74#_c_1529_n 0.00427046f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_600 N_A_1025_119#_M1042_g N_VPWR_c_1697_n 0.0041957f $X=9.7 $Y=2.565 $X2=0
+ $Y2=0
cc_601 N_A_1025_119#_M1032_g N_VPWR_c_1692_n 0.00113998f $X=6.1 $Y=2.495 $X2=0
+ $Y2=0
cc_602 N_A_1025_119#_M1042_g N_VPWR_c_1692_n 0.00587053f $X=9.7 $Y=2.565 $X2=0
+ $Y2=0
cc_603 N_A_1025_119#_M1036_d N_A_388_79#_c_1888_n 0.0058336f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_604 N_A_1025_119#_c_608_n N_A_388_79#_c_1888_n 7.56384e-19 $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_605 N_A_1025_119#_c_614_n N_A_388_79#_c_1888_n 0.0282747f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_606 N_A_1025_119#_M1032_g N_A_388_79#_c_1889_n 0.00219675f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_607 N_A_1025_119#_c_608_n N_A_388_79#_c_1889_n 6.01563e-19 $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_608 N_A_1025_119#_c_614_n N_A_388_79#_c_1889_n 0.00823921f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_609 N_A_1025_119#_M1015_g N_A_388_79#_c_1878_n 4.31453e-19 $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_610 N_A_1025_119#_c_604_n N_A_388_79#_c_1878_n 0.00733866f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_611 N_A_1025_119#_c_613_n N_A_388_79#_c_1878_n 0.0103323f $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_612 N_A_1025_119#_M1032_g N_A_388_79#_c_1890_n 0.0162038f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_613 N_A_1025_119#_c_599_n N_A_388_79#_c_1890_n 0.00260393f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_614 N_A_1025_119#_c_608_n N_A_388_79#_c_1890_n 0.0103323f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_615 N_A_1025_119#_c_619_n N_A_388_79#_c_1890_n 0.00122453f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_616 N_A_1025_119#_c_608_n N_A_388_79#_c_1891_n 0.0158752f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_617 N_A_1025_119#_c_614_n N_A_388_79#_c_1891_n 0.0130031f $X=5.405 $Y=1.665
+ $X2=0 $Y2=0
cc_618 N_A_1025_119#_c_619_n N_A_388_79#_c_1891_n 0.00234227f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_619 N_A_1025_119#_M1015_g N_A_388_79#_c_1879_n 0.00474699f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_620 N_A_1025_119#_c_606_n N_A_388_79#_c_1879_n 0.00414539f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_621 N_A_1025_119#_c_608_n N_A_388_79#_c_1879_n 0.0102296f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_622 N_A_1025_119#_c_619_n N_A_388_79#_c_1879_n 0.00755412f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_623 N_A_1025_119#_c_605_n N_A_388_79#_c_1880_n 0.00121012f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_624 N_A_1025_119#_c_608_n N_A_388_79#_c_1880_n 0.0121259f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_625 N_A_1025_119#_c_613_n N_A_388_79#_c_1880_n 0.0125313f $X=5.525 $Y=1.132
+ $X2=0 $Y2=0
cc_626 N_A_1025_119#_c_619_n N_A_388_79#_c_1880_n 6.96658e-19 $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_627 N_A_1025_119#_M1032_g N_A_388_79#_c_1881_n 0.00418686f $X=6.1 $Y=2.495
+ $X2=0 $Y2=0
cc_628 N_A_1025_119#_c_599_n N_A_388_79#_c_1881_n 0.0121437f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_629 N_A_1025_119#_M1015_g N_A_388_79#_c_1881_n 0.00569051f $X=6.54 $Y=0.805
+ $X2=0 $Y2=0
cc_630 N_A_1025_119#_c_605_n N_A_388_79#_c_1881_n 0.00534514f $X=5.525 $Y=1.5
+ $X2=0 $Y2=0
cc_631 N_A_1025_119#_c_608_n N_A_388_79#_c_1881_n 0.025654f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_632 N_A_1025_119#_c_619_n N_A_388_79#_c_1881_n 0.00206889f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_633 N_A_1025_119#_c_604_n N_A_388_79#_c_1882_n 0.0113657f $X=5.265 $Y=0.74
+ $X2=0 $Y2=0
cc_634 N_A_1025_119#_c_606_n N_A_388_79#_c_1882_n 0.0212057f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_635 N_A_1025_119#_c_609_n N_VGND_M1011_d 0.0231466f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_636 N_A_1025_119#_c_779_p N_VGND_M1011_d 0.00612573f $X=8.24 $Y=0.58 $X2=0
+ $Y2=0
cc_637 N_A_1025_119#_c_611_n N_VGND_M1011_d 0.0012599f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_638 N_A_1025_119#_c_604_n N_VGND_c_2090_n 0.0223626f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_639 N_A_1025_119#_c_607_n N_VGND_c_2090_n 0.0137189f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_640 N_A_1025_119#_c_601_n N_VGND_c_2102_n 0.00278271f $X=8.875 $Y=1.085 $X2=0
+ $Y2=0
cc_641 N_A_1025_119#_c_609_n N_VGND_c_2102_n 0.003347f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_642 N_A_1025_119#_c_610_n N_VGND_c_2102_n 0.0611382f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_643 N_A_1025_119#_c_611_n N_VGND_c_2102_n 0.0118998f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_644 N_A_1025_119#_c_606_n N_VGND_c_2109_n 0.0751677f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_645 N_A_1025_119#_c_607_n N_VGND_c_2109_n 0.0175158f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_646 N_A_1025_119#_c_609_n N_VGND_c_2109_n 0.00545957f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_647 N_A_1025_119#_c_615_n N_VGND_c_2109_n 0.00863901f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_648 N_A_1025_119#_c_609_n N_VGND_c_2110_n 0.0398776f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_649 N_A_1025_119#_c_611_n N_VGND_c_2110_n 0.014039f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_650 N_A_1025_119#_c_615_n N_VGND_c_2110_n 0.00577425f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_651 N_A_1025_119#_c_601_n N_VGND_c_2114_n 0.00358525f $X=8.875 $Y=1.085 $X2=0
+ $Y2=0
cc_652 N_A_1025_119#_c_606_n N_VGND_c_2114_n 0.0507418f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_653 N_A_1025_119#_c_607_n N_VGND_c_2114_n 0.0111521f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_654 N_A_1025_119#_c_609_n N_VGND_c_2114_n 0.015012f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_655 N_A_1025_119#_c_610_n N_VGND_c_2114_n 0.0343665f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_656 N_A_1025_119#_c_611_n N_VGND_c_2114_n 0.00655543f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_657 N_A_1025_119#_c_615_n N_VGND_c_2114_n 0.0055945f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_658 N_A_1025_119#_c_609_n A_1401_119# 5.60515e-19 $X=8.155 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_659 N_A_1025_119#_c_615_n A_1401_119# 0.00145656f $X=7.085 $Y=0.395 $X2=-0.19
+ $Y2=-0.245
cc_660 N_A_1370_290#_M1043_g N_RESET_B_c_893_n 0.00881802f $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_661 N_A_1370_290#_M1043_g N_RESET_B_M1011_g 0.0413828f $X=6.93 $Y=0.805 $X2=0
+ $Y2=0
cc_662 N_A_1370_290#_c_806_n N_RESET_B_M1011_g 0.0149052f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_663 N_A_1370_290#_c_806_n N_RESET_B_c_896_n 0.0110159f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_664 N_A_1370_290#_c_804_n N_RESET_B_c_897_n 0.00392043f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_665 N_A_1370_290#_c_805_n N_RESET_B_c_897_n 0.00184962f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_666 N_A_1370_290#_M1020_g N_RESET_B_c_898_n 0.00165672f $X=6.94 $Y=2.495
+ $X2=0 $Y2=0
cc_667 N_A_1370_290#_M1043_g N_RESET_B_c_898_n 0.00134145f $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_668 N_A_1370_290#_c_804_n N_RESET_B_c_898_n 4.1836e-19 $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_669 N_A_1370_290#_c_805_n N_RESET_B_c_898_n 0.00818789f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_670 N_A_1370_290#_M1020_g N_RESET_B_c_908_n 0.0119303f $X=6.94 $Y=2.495 $X2=0
+ $Y2=0
cc_671 N_A_1370_290#_c_804_n N_RESET_B_c_908_n 0.00636364f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_672 N_A_1370_290#_c_805_n N_RESET_B_c_908_n 0.00145933f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_673 N_A_1370_290#_M1000_d N_RESET_B_c_910_n 0.00365135f $X=8.59 $Y=1.735
+ $X2=0 $Y2=0
cc_674 N_A_1370_290#_c_812_n N_RESET_B_c_910_n 0.0384843f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_675 N_A_1370_290#_M1020_g N_RESET_B_c_915_n 0.0220571f $X=6.94 $Y=2.495 $X2=0
+ $Y2=0
cc_676 N_A_1370_290#_c_806_n N_A_1223_119#_M1007_g 0.01076f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_677 N_A_1370_290#_c_807_n N_A_1223_119#_M1007_g 0.0115167f $X=8.845 $Y=0.842
+ $X2=0 $Y2=0
cc_678 N_A_1370_290#_c_808_n N_A_1223_119#_M1007_g 0.00305733f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_679 N_A_1370_290#_c_812_n N_A_1223_119#_M1000_g 3.63477e-19 $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_680 N_A_1370_290#_M1043_g N_A_1223_119#_c_1108_n 0.00323506f $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_681 N_A_1370_290#_c_804_n N_A_1223_119#_c_1108_n 0.0500464f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_682 N_A_1370_290#_c_805_n N_A_1223_119#_c_1108_n 0.0114066f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_683 N_A_1370_290#_c_822_n N_A_1223_119#_c_1108_n 0.00869313f $X=7.21 $Y=1.005
+ $X2=0 $Y2=0
cc_684 N_A_1370_290#_M1020_g N_A_1223_119#_c_1136_n 0.0119163f $X=6.94 $Y=2.495
+ $X2=0 $Y2=0
cc_685 N_A_1370_290#_c_804_n N_A_1223_119#_c_1136_n 0.00226215f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_686 N_A_1370_290#_c_805_n N_A_1223_119#_c_1136_n 0.00227973f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_687 N_A_1370_290#_M1020_g N_A_1223_119#_c_1115_n 6.67944e-19 $X=6.94 $Y=2.495
+ $X2=0 $Y2=0
cc_688 N_A_1370_290#_M1020_g N_A_1223_119#_c_1109_n 0.00562338f $X=6.94 $Y=2.495
+ $X2=0 $Y2=0
cc_689 N_A_1370_290#_c_804_n N_A_1223_119#_c_1109_n 0.0148532f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_690 N_A_1370_290#_c_805_n N_A_1223_119#_c_1109_n 0.00180559f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_691 N_A_1370_290#_M1043_g N_A_1223_119#_c_1110_n 7.20903e-19 $X=6.93 $Y=0.805
+ $X2=0 $Y2=0
cc_692 N_A_1370_290#_c_804_n N_A_1223_119#_c_1110_n 0.0265063f $X=7.105 $Y=1.615
+ $X2=0 $Y2=0
cc_693 N_A_1370_290#_c_805_n N_A_1223_119#_c_1110_n 0.00122451f $X=7.105
+ $Y=1.615 $X2=0 $Y2=0
cc_694 N_A_1370_290#_c_806_n N_A_1223_119#_c_1110_n 0.0142918f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_695 N_A_1370_290#_c_806_n N_A_1223_119#_c_1111_n 0.080152f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_696 N_A_1370_290#_c_808_n N_A_1223_119#_c_1111_n 0.0250137f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_697 N_A_1370_290#_c_806_n N_A_1223_119#_c_1112_n 0.00251001f $X=8.495
+ $Y=0.842 $X2=0 $Y2=0
cc_698 N_A_1370_290#_c_807_n N_A_1223_119#_c_1112_n 0.00192164f $X=8.845
+ $Y=0.842 $X2=0 $Y2=0
cc_699 N_A_1370_290#_c_808_n N_A_1223_119#_c_1112_n 0.00590528f $X=8.785
+ $Y=1.745 $X2=0 $Y2=0
cc_700 N_A_1370_290#_M1020_g N_A_852_119#_M1040_g 0.0407278f $X=6.94 $Y=2.495
+ $X2=0 $Y2=0
cc_701 N_A_1370_290#_M1020_g N_A_852_119#_c_1229_n 0.0103216f $X=6.94 $Y=2.495
+ $X2=0 $Y2=0
cc_702 N_A_1370_290#_c_812_n N_A_852_119#_c_1229_n 0.00262042f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_703 N_A_1370_290#_c_824_n N_A_852_119#_M1004_g 0.00286004f $X=8.785 $Y=1.89
+ $X2=0 $Y2=0
cc_704 N_A_1370_290#_c_812_n N_A_852_119#_M1004_g 0.0174995f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_705 N_A_1370_290#_c_808_n N_A_852_119#_M1004_g 0.00298672f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_706 N_A_1370_290#_c_808_n N_A_852_119#_c_1216_n 0.00575991f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_707 N_A_1370_290#_c_812_n N_A_1790_74#_c_1516_n 0.0268436f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_708 N_A_1370_290#_M1020_g N_VPWR_c_1695_n 0.00349293f $X=6.94 $Y=2.495 $X2=0
+ $Y2=0
cc_709 N_A_1370_290#_c_812_n N_VPWR_c_1696_n 0.0341037f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_710 N_A_1370_290#_c_812_n N_VPWR_c_1697_n 0.00647129f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_711 N_A_1370_290#_M1020_g N_VPWR_c_1692_n 0.00113998f $X=6.94 $Y=2.495 $X2=0
+ $Y2=0
cc_712 N_A_1370_290#_c_812_n N_VPWR_c_1692_n 0.00789046f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_713 N_A_1370_290#_c_806_n N_VGND_M1011_d 0.0123333f $X=8.495 $Y=0.842 $X2=0
+ $Y2=0
cc_714 N_A_1370_290#_c_822_n A_1401_119# 0.00131009f $X=7.21 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_715 N_RESET_B_c_896_n N_A_1223_119#_M1007_g 0.00460948f $X=7.66 $Y=1.165
+ $X2=0 $Y2=0
cc_716 N_RESET_B_c_898_n N_A_1223_119#_M1000_g 0.00452045f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_910_n N_A_1223_119#_M1000_g 0.00792629f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_908_n N_A_1223_119#_c_1108_n 0.0243758f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_908_n N_A_1223_119#_c_1136_n 0.0191198f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_908_n N_A_1223_119#_c_1115_n 0.00956244f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_721 N_RESET_B_c_903_n N_A_1223_119#_c_1109_n 0.0200013f $X=7.525 $Y=2.165
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_898_n N_A_1223_119#_c_1109_n 0.00611723f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_723 N_RESET_B_c_908_n N_A_1223_119#_c_1109_n 0.0319179f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_724 N_RESET_B_c_911_n N_A_1223_119#_c_1109_n 0.00394987f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_915_n N_A_1223_119#_c_1109_n 0.0154752f $X=7.735 $Y=1.98
+ $X2=0 $Y2=0
cc_726 N_RESET_B_c_916_n N_A_1223_119#_c_1109_n 0.0379481f $X=7.825 $Y=1.96
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_897_n N_A_1223_119#_c_1110_n 0.00420432f $X=7.395 $Y=1.165
+ $X2=0 $Y2=0
cc_728 N_RESET_B_c_896_n N_A_1223_119#_c_1111_n 0.00254634f $X=7.66 $Y=1.165
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_898_n N_A_1223_119#_c_1111_n 0.0171699f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_730 N_RESET_B_c_908_n N_A_1223_119#_c_1111_n 0.00645679f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_910_n N_A_1223_119#_c_1111_n 0.0108447f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_RESET_B_c_911_n N_A_1223_119#_c_1111_n 0.00336108f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_915_n N_A_1223_119#_c_1111_n 0.00673793f $X=7.735 $Y=1.98
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_916_n N_A_1223_119#_c_1111_n 0.0174718f $X=7.825 $Y=1.96
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_898_n N_A_1223_119#_c_1112_n 0.00790704f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_908_n N_A_852_119#_M1019_s 0.00158238f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_908_n N_A_852_119#_M1036_g 0.00390692f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_908_n N_A_852_119#_c_1211_n 0.00269906f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_893_n N_A_852_119#_c_1214_n 0.00880557f $X=7.245 $Y=0.18
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_908_n N_A_852_119#_M1040_g 0.00299989f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_903_n N_A_852_119#_c_1229_n 0.0101913f $X=7.525 $Y=2.165
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_910_n N_A_852_119#_M1004_g 0.00995626f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_910_n N_A_852_119#_c_1215_n 0.00840564f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_744 N_RESET_B_M1035_g N_A_852_119#_c_1237_n 0.00274653f $X=3.585 $Y=2.735
+ $X2=0 $Y2=0
cc_745 N_RESET_B_c_908_n N_A_852_119#_c_1237_n 0.0101557f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_909_n N_A_852_119#_c_1237_n 0.00141079f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_913_n N_A_852_119#_c_1237_n 4.58098e-19 $X=3.95 $Y=1.985
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_914_n N_A_852_119#_c_1237_n 0.0111141f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_749 N_RESET_B_M1003_g N_A_852_119#_c_1220_n 5.20809e-19 $X=3.57 $Y=0.605
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_893_n N_A_852_119#_c_1220_n 0.00584017f $X=7.245 $Y=0.18
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_908_n N_A_852_119#_c_1221_n 0.0386239f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_909_n N_A_852_119#_c_1221_n 0.00142114f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_913_n N_A_852_119#_c_1221_n 6.26023e-19 $X=3.95 $Y=1.985
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_914_n N_A_852_119#_c_1221_n 0.0139322f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_893_n N_A_852_119#_c_1223_n 0.0101478f $X=7.245 $Y=0.18 $X2=0
+ $Y2=0
cc_756 N_RESET_B_M1023_g N_A_2006_373#_M1022_g 0.00842708f $X=11.005 $Y=2.565
+ $X2=0 $Y2=0
cc_757 N_RESET_B_M1024_g N_A_2006_373#_M1045_g 0.0455699f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_918_n N_A_2006_373#_M1045_g 0.00569933f $X=10.945 $Y=1.82
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1023_g N_A_2006_373#_c_1391_n 0.00287022f $X=11.005 $Y=2.565
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_910_n N_A_2006_373#_c_1391_n 0.0257703f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_761 RESET_B N_A_2006_373#_c_1391_n 0.00275621f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_762 N_RESET_B_c_917_n N_A_2006_373#_c_1391_n 5.14527e-19 $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_918_n N_A_2006_373#_c_1391_n 0.00379957f $X=10.945 $Y=1.82
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_919_n N_A_2006_373#_c_1391_n 0.0241058f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_765 N_RESET_B_M1023_g N_A_2006_373#_c_1392_n 0.00182434f $X=11.005 $Y=2.565
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_910_n N_A_2006_373#_c_1392_n 0.0143374f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_767 RESET_B N_A_2006_373#_c_1392_n 0.00149024f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_768 N_RESET_B_c_917_n N_A_2006_373#_c_1392_n 0.0189581f $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_919_n N_A_2006_373#_c_1392_n 0.00155699f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_900_n N_A_2006_373#_c_1383_n 0.012737f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_910_n N_A_2006_373#_c_1383_n 0.00282721f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_772 RESET_B N_A_2006_373#_c_1383_n 0.00310808f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_773 N_RESET_B_c_917_n N_A_2006_373#_c_1383_n 0.00313906f $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_918_n N_A_2006_373#_c_1383_n 0.00306368f $X=10.945 $Y=1.82
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_919_n N_A_2006_373#_c_1383_n 0.0505438f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_M1023_g N_A_2006_373#_c_1394_n 0.0116913f $X=11.005 $Y=2.565
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_900_n N_A_2006_373#_c_1394_n 4.02079e-19 $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_778 N_RESET_B_c_910_n N_A_2006_373#_c_1394_n 0.00318931f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_779 RESET_B N_A_2006_373#_c_1394_n 0.00772021f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_780 N_RESET_B_c_917_n N_A_2006_373#_c_1394_n 0.00248288f $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_919_n N_A_2006_373#_c_1394_n 0.0232211f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_782 N_RESET_B_M1024_g N_A_2006_373#_c_1385_n 9.65407e-19 $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_783 N_RESET_B_M1024_g N_A_2006_373#_c_1387_n 6.07222e-19 $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_784 N_RESET_B_M1023_g N_A_2006_373#_c_1396_n 0.01203f $X=11.005 $Y=2.565
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_917_n N_A_2006_373#_c_1396_n 3.45297e-19 $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_919_n N_A_2006_373#_c_1396_n 0.0276612f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_910_n N_A_1790_74#_M1004_d 0.00808489f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_788 N_RESET_B_M1024_g N_A_1790_74#_M1016_g 0.0556926f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_789 N_RESET_B_M1024_g N_A_1790_74#_c_1497_n 0.0094439f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_900_n N_A_1790_74#_c_1497_n 0.00511143f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_917_n N_A_1790_74#_c_1497_n 0.00126375f $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_792 N_RESET_B_M1023_g N_A_1790_74#_M1028_g 0.017447f $X=11.005 $Y=2.565 $X2=0
+ $Y2=0
cc_793 N_RESET_B_c_917_n N_A_1790_74#_M1028_g 0.0168019f $X=10.945 $Y=1.985
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_918_n N_A_1790_74#_M1028_g 0.00511143f $X=10.945 $Y=1.82
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_919_n N_A_1790_74#_M1028_g 0.00839981f $X=10.8 $Y=2.035 $X2=0
+ $Y2=0
cc_796 N_RESET_B_c_910_n N_A_1790_74#_c_1516_n 0.0195034f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_910_n N_A_1790_74#_c_1506_n 0.0213448f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_M1024_g N_A_1790_74#_c_1507_n 0.0184362f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_799 N_RESET_B_c_900_n N_A_1790_74#_c_1507_n 0.00370089f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_908_n N_VPWR_M1019_d 0.00277212f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_801 N_RESET_B_c_910_n N_VPWR_M1000_s 0.00198285f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_802 N_RESET_B_M1035_g N_VPWR_c_1693_n 0.00520262f $X=3.585 $Y=2.735 $X2=0
+ $Y2=0
cc_803 N_RESET_B_c_903_n N_VPWR_c_1695_n 0.0031993f $X=7.525 $Y=2.165 $X2=0
+ $Y2=0
cc_804 N_RESET_B_c_903_n N_VPWR_c_1696_n 0.0057797f $X=7.525 $Y=2.165 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_898_n N_VPWR_c_1696_n 4.74228e-19 $X=7.735 $Y=1.795 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_910_n N_VPWR_c_1696_n 0.0236795f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_911_n N_VPWR_c_1696_n 0.0027362f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_915_n N_VPWR_c_1696_n 0.00134605f $X=7.735 $Y=1.98 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_916_n N_VPWR_c_1696_n 0.0258087f $X=7.825 $Y=1.96 $X2=0 $Y2=0
cc_810 N_RESET_B_c_919_n N_VPWR_c_1698_n 0.0233946f $X=10.8 $Y=2.035 $X2=0 $Y2=0
cc_811 N_RESET_B_M1035_g N_VPWR_c_1703_n 0.00572074f $X=3.585 $Y=2.735 $X2=0
+ $Y2=0
cc_812 N_RESET_B_M1023_g N_VPWR_c_1709_n 0.00523383f $X=11.005 $Y=2.565 $X2=0
+ $Y2=0
cc_813 N_RESET_B_M1023_g N_VPWR_c_1717_n 0.00523928f $X=11.005 $Y=2.565 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_910_n N_VPWR_c_1717_n 0.00135184f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_815 N_RESET_B_M1035_g N_VPWR_c_1692_n 0.00760006f $X=3.585 $Y=2.735 $X2=0
+ $Y2=0
cc_816 N_RESET_B_c_903_n N_VPWR_c_1692_n 0.00113998f $X=7.525 $Y=2.165 $X2=0
+ $Y2=0
cc_817 N_RESET_B_M1023_g N_VPWR_c_1692_n 0.00587053f $X=11.005 $Y=2.565 $X2=0
+ $Y2=0
cc_818 N_RESET_B_M1003_g N_A_388_79#_c_1875_n 0.011739f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_819 N_RESET_B_M1003_g N_A_388_79#_c_1877_n 0.0216891f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_820 N_RESET_B_M1035_g N_A_388_79#_c_1877_n 0.00922847f $X=3.585 $Y=2.735
+ $X2=0 $Y2=0
cc_821 N_RESET_B_c_906_n N_A_388_79#_c_1877_n 0.0092617f $X=3.585 $Y=1.985 $X2=0
+ $Y2=0
cc_822 N_RESET_B_c_909_n N_A_388_79#_c_1877_n 0.00108246f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_823 N_RESET_B_c_914_n N_A_388_79#_c_1877_n 0.0228178f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_824 N_RESET_B_M1035_g N_A_388_79#_c_1886_n 0.0218371f $X=3.585 $Y=2.735 $X2=0
+ $Y2=0
cc_825 N_RESET_B_c_909_n N_A_388_79#_c_1886_n 0.0014753f $X=4.225 $Y=2.035 $X2=0
+ $Y2=0
cc_826 N_RESET_B_c_913_n N_A_388_79#_c_1886_n 0.00943655f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_827 N_RESET_B_c_914_n N_A_388_79#_c_1886_n 0.016893f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_828 N_RESET_B_M1035_g N_A_388_79#_c_1887_n 0.00809035f $X=3.585 $Y=2.735
+ $X2=0 $Y2=0
cc_829 N_RESET_B_c_908_n N_A_388_79#_c_1888_n 0.0232417f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_909_n N_A_388_79#_c_1888_n 0.00643846f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_831 N_RESET_B_c_913_n N_A_388_79#_c_1888_n 0.00177112f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_832 N_RESET_B_c_914_n N_A_388_79#_c_1888_n 0.00610606f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_833 N_RESET_B_c_908_n N_A_388_79#_c_1889_n 0.0011812f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_834 N_RESET_B_c_908_n N_A_388_79#_c_1890_n 0.0218219f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_835 N_RESET_B_c_908_n N_A_388_79#_c_1891_n 0.01661f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_836 N_RESET_B_c_908_n N_A_388_79#_c_1881_n 0.00666387f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_837 N_RESET_B_M1003_g N_VGND_c_2089_n 0.00773148f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_838 N_RESET_B_c_893_n N_VGND_c_2089_n 0.0192978f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_839 N_RESET_B_c_894_n N_VGND_c_2089_n 0.00321798f $X=3.645 $Y=0.18 $X2=0
+ $Y2=0
cc_840 N_RESET_B_c_893_n N_VGND_c_2090_n 0.0170937f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_841 N_RESET_B_M1024_g N_VGND_c_2091_n 0.0122664f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_842 N_RESET_B_c_894_n N_VGND_c_2098_n 0.00564095f $X=3.645 $Y=0.18 $X2=0
+ $Y2=0
cc_843 N_RESET_B_c_893_n N_VGND_c_2100_n 0.0237488f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_844 N_RESET_B_M1024_g N_VGND_c_2105_n 0.00383152f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_845 N_RESET_B_c_893_n N_VGND_c_2109_n 0.0558684f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_846 N_RESET_B_c_893_n N_VGND_c_2110_n 0.0109384f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_847 N_RESET_B_c_893_n N_VGND_c_2114_n 0.0936844f $X=7.245 $Y=0.18 $X2=0 $Y2=0
cc_848 N_RESET_B_c_894_n N_VGND_c_2114_n 0.0110707f $X=3.645 $Y=0.18 $X2=0 $Y2=0
cc_849 N_RESET_B_M1024_g N_VGND_c_2114_n 0.0075694f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_850 N_RESET_B_M1003_g N_noxref_25_c_2246_n 0.00204561f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_851 N_RESET_B_M1003_g N_noxref_25_c_2248_n 0.0037218f $X=3.57 $Y=0.605 $X2=0
+ $Y2=0
cc_852 N_A_1223_119#_c_1115_n N_A_852_119#_c_1226_n 0.00352096f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_853 N_A_1223_119#_c_1108_n N_A_852_119#_M1040_g 0.00180133f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_854 N_A_1223_119#_c_1115_n N_A_852_119#_M1040_g 0.0143382f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_855 N_A_1223_119#_M1000_g N_A_852_119#_c_1229_n 0.0123711f $X=8.5 $Y=2.235
+ $X2=0 $Y2=0
cc_856 N_A_1223_119#_c_1136_n N_A_852_119#_c_1229_n 0.00275389f $X=7.38 $Y=2.425
+ $X2=0 $Y2=0
cc_857 N_A_1223_119#_c_1115_n N_A_852_119#_c_1229_n 0.00213073f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_858 N_A_1223_119#_c_1109_n N_A_852_119#_c_1229_n 0.00632319f $X=7.465 $Y=2.32
+ $X2=0 $Y2=0
cc_859 N_A_1223_119#_M1000_g N_A_852_119#_M1004_g 0.00893939f $X=8.5 $Y=2.235
+ $X2=0 $Y2=0
cc_860 N_A_1223_119#_c_1112_n N_A_852_119#_c_1216_n 0.00893939f $X=8.425 $Y=1.41
+ $X2=0 $Y2=0
cc_861 N_A_1223_119#_c_1136_n N_VPWR_M1020_d 0.00669455f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_862 N_A_1223_119#_c_1136_n N_VPWR_c_1695_n 0.0178778f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_863 N_A_1223_119#_c_1115_n N_VPWR_c_1695_n 8.68772e-19 $X=6.83 $Y=2.425 $X2=0
+ $Y2=0
cc_864 N_A_1223_119#_c_1109_n N_VPWR_c_1695_n 0.00274181f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_865 N_A_1223_119#_M1000_g N_VPWR_c_1696_n 0.0166824f $X=8.5 $Y=2.235 $X2=0
+ $Y2=0
cc_866 N_A_1223_119#_c_1109_n N_VPWR_c_1696_n 0.0295996f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_867 N_A_1223_119#_c_1111_n N_VPWR_c_1696_n 0.0170364f $X=8.425 $Y=1.41 $X2=0
+ $Y2=0
cc_868 N_A_1223_119#_c_1112_n N_VPWR_c_1696_n 0.00347843f $X=8.425 $Y=1.41 $X2=0
+ $Y2=0
cc_869 N_A_1223_119#_c_1115_n N_VPWR_c_1705_n 0.00987805f $X=6.83 $Y=2.425 $X2=0
+ $Y2=0
cc_870 N_A_1223_119#_c_1109_n N_VPWR_c_1708_n 0.00742407f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_871 N_A_1223_119#_M1000_g N_VPWR_c_1692_n 9.455e-19 $X=8.5 $Y=2.235 $X2=0
+ $Y2=0
cc_872 N_A_1223_119#_c_1136_n N_VPWR_c_1692_n 0.00963217f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_873 N_A_1223_119#_c_1115_n N_VPWR_c_1692_n 0.019007f $X=6.83 $Y=2.425 $X2=0
+ $Y2=0
cc_874 N_A_1223_119#_c_1109_n N_VPWR_c_1692_n 0.0152355f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_875 N_A_1223_119#_c_1108_n N_A_388_79#_c_1889_n 0.00326197f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_876 N_A_1223_119#_c_1115_n N_A_388_79#_c_1889_n 0.0119294f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_877 N_A_1223_119#_c_1108_n N_A_388_79#_c_1878_n 0.00327725f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_878 N_A_1223_119#_c_1108_n N_A_388_79#_c_1890_n 0.0130386f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_879 N_A_1223_119#_c_1115_n N_A_388_79#_c_1890_n 0.0209731f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_880 N_A_1223_119#_c_1121_n N_A_388_79#_c_1879_n 0.0240423f $X=6.66 $Y=0.8
+ $X2=0 $Y2=0
cc_881 N_A_1223_119#_c_1108_n N_A_388_79#_c_1879_n 0.0135678f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_882 N_A_1223_119#_c_1108_n N_A_388_79#_c_1881_n 0.0518294f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_883 N_A_1223_119#_c_1115_n A_1328_457# 0.00139756f $X=6.83 $Y=2.425 $X2=-0.19
+ $Y2=-0.245
cc_884 N_A_1223_119#_M1007_g N_VGND_c_2102_n 0.00278271f $X=8.445 $Y=0.69 $X2=0
+ $Y2=0
cc_885 N_A_1223_119#_M1007_g N_VGND_c_2110_n 0.00116012f $X=8.445 $Y=0.69 $X2=0
+ $Y2=0
cc_886 N_A_1223_119#_M1007_g N_VGND_c_2114_n 0.00358525f $X=8.445 $Y=0.69 $X2=0
+ $Y2=0
cc_887 N_A_1223_119#_c_1121_n A_1323_119# 0.0012023f $X=6.66 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_888 N_A_852_119#_M1002_g N_A_2006_373#_M1045_g 0.0830829f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_889 N_A_852_119#_M1004_g N_A_1790_74#_c_1516_n 0.0038297f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_890 N_A_852_119#_M1002_g N_A_1790_74#_c_1519_n 0.0113037f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_891 N_A_852_119#_M1002_g N_A_1790_74#_c_1505_n 0.00782202f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_892 N_A_852_119#_c_1215_n N_A_1790_74#_c_1506_n 0.00624492f $X=9.85 $Y=1.55
+ $X2=0 $Y2=0
cc_893 N_A_852_119#_M1002_g N_A_1790_74#_c_1506_n 0.0034675f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_894 N_A_852_119#_M1002_g N_A_1790_74#_c_1529_n 0.00668941f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_895 N_A_852_119#_c_1221_n N_VPWR_M1019_d 0.00173132f $X=4.49 $Y=1.717 $X2=0
+ $Y2=0
cc_896 N_A_852_119#_M1036_g N_VPWR_c_1694_n 0.0104793f $X=5.095 $Y=2.495 $X2=0
+ $Y2=0
cc_897 N_A_852_119#_c_1211_n N_VPWR_c_1694_n 0.00212623f $X=5.595 $Y=3.075 $X2=0
+ $Y2=0
cc_898 N_A_852_119#_c_1227_n N_VPWR_c_1694_n 7.14853e-19 $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_899 N_A_852_119#_M1040_g N_VPWR_c_1695_n 0.00683756f $X=6.55 $Y=2.495 $X2=0
+ $Y2=0
cc_900 N_A_852_119#_c_1229_n N_VPWR_c_1695_n 0.0209699f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_901 N_A_852_119#_c_1229_n N_VPWR_c_1696_n 0.0210786f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_902 N_A_852_119#_M1004_g N_VPWR_c_1696_n 0.00679318f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_903 N_A_852_119#_c_1229_n N_VPWR_c_1697_n 0.0188909f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_904 N_A_852_119#_M1036_g N_VPWR_c_1705_n 0.00401239f $X=5.095 $Y=2.495 $X2=0
+ $Y2=0
cc_905 N_A_852_119#_c_1227_n N_VPWR_c_1705_n 0.0464425f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_906 N_A_852_119#_c_1229_n N_VPWR_c_1708_n 0.0266609f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_907 N_A_852_119#_M1036_g N_VPWR_c_1692_n 0.00499124f $X=5.095 $Y=2.495 $X2=0
+ $Y2=0
cc_908 N_A_852_119#_c_1226_n N_VPWR_c_1692_n 0.0228136f $X=6.46 $Y=3.15 $X2=0
+ $Y2=0
cc_909 N_A_852_119#_c_1227_n N_VPWR_c_1692_n 0.00586733f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_910 N_A_852_119#_c_1229_n N_VPWR_c_1692_n 0.0676591f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_911 N_A_852_119#_c_1233_n N_VPWR_c_1692_n 0.00508464f $X=6.55 $Y=3.15 $X2=0
+ $Y2=0
cc_912 N_A_852_119#_M1019_s N_A_388_79#_c_1888_n 0.00756732f $X=4.275 $Y=1.935
+ $X2=0 $Y2=0
cc_913 N_A_852_119#_M1036_g N_A_388_79#_c_1888_n 0.0160071f $X=5.095 $Y=2.495
+ $X2=0 $Y2=0
cc_914 N_A_852_119#_c_1211_n N_A_388_79#_c_1888_n 0.013906f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_915 N_A_852_119#_c_1237_n N_A_388_79#_c_1888_n 0.0143912f $X=4.42 $Y=2.11
+ $X2=0 $Y2=0
cc_916 N_A_852_119#_c_1221_n N_A_388_79#_c_1888_n 0.00799706f $X=4.49 $Y=1.717
+ $X2=0 $Y2=0
cc_917 N_A_852_119#_c_1211_n N_A_388_79#_c_1889_n 0.0077784f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_918 N_A_852_119#_c_1226_n N_A_388_79#_c_1889_n 0.0044661f $X=6.46 $Y=3.15
+ $X2=0 $Y2=0
cc_919 N_A_852_119#_c_1212_n N_A_388_79#_c_1878_n 0.00325896f $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_920 N_A_852_119#_c_1214_n N_A_388_79#_c_1878_n 0.00764854f $X=6.04 $Y=1.11
+ $X2=0 $Y2=0
cc_921 N_A_852_119#_M1040_g N_A_388_79#_c_1890_n 0.00131556f $X=6.55 $Y=2.495
+ $X2=0 $Y2=0
cc_922 N_A_852_119#_c_1211_n N_A_388_79#_c_1891_n 0.00122663f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_923 N_A_852_119#_c_1212_n N_A_388_79#_c_1879_n 0.00745866f $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_924 N_A_852_119#_c_1212_n N_A_388_79#_c_1880_n 0.00542357f $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_925 N_A_852_119#_c_1210_n N_A_388_79#_c_1881_n 0.00225242f $X=5.595 $Y=1.445
+ $X2=0 $Y2=0
cc_926 N_A_852_119#_c_1212_n N_A_388_79#_c_1882_n 5.07577e-19 $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_927 N_A_852_119#_c_1213_n N_A_388_79#_c_1882_n 0.00489735f $X=5.67 $Y=1.185
+ $X2=0 $Y2=0
cc_928 N_A_852_119#_c_1214_n N_A_388_79#_c_1882_n 0.00209515f $X=6.04 $Y=1.11
+ $X2=0 $Y2=0
cc_929 N_A_852_119#_c_1220_n N_VGND_c_2089_n 0.0150337f $X=4.405 $Y=0.75 $X2=0
+ $Y2=0
cc_930 N_A_852_119#_c_1220_n N_VGND_c_2090_n 0.00945897f $X=4.405 $Y=0.75 $X2=0
+ $Y2=0
cc_931 N_A_852_119#_c_1221_n N_VGND_c_2090_n 0.0150964f $X=4.49 $Y=1.717 $X2=0
+ $Y2=0
cc_932 N_A_852_119#_c_1223_n N_VGND_c_2090_n 9.24546e-19 $X=5.14 $Y=1.445 $X2=0
+ $Y2=0
cc_933 N_A_852_119#_M1002_g N_VGND_c_2091_n 0.00120934f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_934 N_A_852_119#_c_1220_n N_VGND_c_2100_n 0.00693131f $X=4.405 $Y=0.75 $X2=0
+ $Y2=0
cc_935 N_A_852_119#_M1002_g N_VGND_c_2102_n 0.00298877f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_936 N_A_852_119#_M1002_g N_VGND_c_2114_n 0.00370514f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_937 N_A_852_119#_c_1220_n N_VGND_c_2114_n 0.00873938f $X=4.405 $Y=0.75 $X2=0
+ $Y2=0
cc_938 N_A_852_119#_c_1223_n N_VGND_c_2114_n 7.82699e-19 $X=5.14 $Y=1.445 $X2=0
+ $Y2=0
cc_939 N_A_2006_373#_c_1385_n N_A_1790_74#_M1016_g 0.00658176f $X=11.29 $Y=0.58
+ $X2=0 $Y2=0
cc_940 N_A_2006_373#_c_1387_n N_A_1790_74#_M1016_g 0.00562994f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_941 N_A_2006_373#_c_1388_n N_A_1790_74#_M1016_g 0.00311727f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_942 N_A_2006_373#_c_1383_n N_A_1790_74#_c_1497_n 0.0111503f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_943 N_A_2006_373#_c_1386_n N_A_1790_74#_c_1497_n 0.00258531f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_944 N_A_2006_373#_c_1387_n N_A_1790_74#_c_1497_n 0.0075729f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_945 N_A_2006_373#_c_1388_n N_A_1790_74#_c_1497_n 0.00284108f $X=11.775
+ $Y=1.48 $X2=0 $Y2=0
cc_946 N_A_2006_373#_c_1383_n N_A_1790_74#_M1028_g 0.00955274f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_947 N_A_2006_373#_c_1396_n N_A_1790_74#_M1028_g 0.00756118f $X=11.23 $Y=2.405
+ $X2=0 $Y2=0
cc_948 N_A_2006_373#_c_1383_n N_A_1790_74#_c_1498_n 0.0109994f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_949 N_A_2006_373#_c_1386_n N_A_1790_74#_c_1498_n 0.00113849f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_950 N_A_2006_373#_c_1388_n N_A_1790_74#_c_1498_n 0.0180935f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_951 N_A_2006_373#_c_1383_n N_A_1790_74#_M1005_g 5.67655e-19 $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_952 N_A_2006_373#_c_1385_n N_A_1790_74#_M1025_g 0.00446735f $X=11.29 $Y=0.58
+ $X2=0 $Y2=0
cc_953 N_A_2006_373#_c_1386_n N_A_1790_74#_M1025_g 0.00377396f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_954 N_A_2006_373#_c_1388_n N_A_1790_74#_M1025_g 0.00455681f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_955 N_A_2006_373#_M1022_g N_A_1790_74#_c_1516_n 0.0154851f $X=10.12 $Y=2.565
+ $X2=0 $Y2=0
cc_956 N_A_2006_373#_M1045_g N_A_1790_74#_c_1519_n 0.00245703f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_957 N_A_2006_373#_M1045_g N_A_1790_74#_c_1505_n 0.00544577f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_958 N_A_2006_373#_M1022_g N_A_1790_74#_c_1506_n 0.00327425f $X=10.12 $Y=2.565
+ $X2=0 $Y2=0
cc_959 N_A_2006_373#_M1045_g N_A_1790_74#_c_1506_n 0.0092441f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_960 N_A_2006_373#_c_1391_n N_A_1790_74#_c_1506_n 0.0474407f $X=10.405 $Y=2.03
+ $X2=0 $Y2=0
cc_961 N_A_2006_373#_c_1392_n N_A_1790_74#_c_1506_n 0.00892164f $X=10.405
+ $Y=2.03 $X2=0 $Y2=0
cc_962 N_A_2006_373#_c_1384_n N_A_1790_74#_c_1506_n 0.0135848f $X=10.545
+ $Y=1.565 $X2=0 $Y2=0
cc_963 N_A_2006_373#_c_1395_n N_A_1790_74#_c_1506_n 0.00308334f $X=10.545
+ $Y=2.405 $X2=0 $Y2=0
cc_964 N_A_2006_373#_M1045_g N_A_1790_74#_c_1507_n 0.0192761f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_965 N_A_2006_373#_c_1392_n N_A_1790_74#_c_1507_n 0.00397248f $X=10.405
+ $Y=2.03 $X2=0 $Y2=0
cc_966 N_A_2006_373#_c_1383_n N_A_1790_74#_c_1507_n 0.0718198f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_967 N_A_2006_373#_c_1384_n N_A_1790_74#_c_1507_n 0.0235777f $X=10.545
+ $Y=1.565 $X2=0 $Y2=0
cc_968 N_A_2006_373#_c_1386_n N_A_1790_74#_c_1507_n 0.00476671f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_969 N_A_2006_373#_c_1387_n N_A_1790_74#_c_1507_n 0.026725f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_970 N_A_2006_373#_c_1388_n N_A_1790_74#_c_1507_n 0.0207312f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_971 N_A_2006_373#_c_1394_n N_VPWR_M1022_d 0.00447642f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_972 N_A_2006_373#_c_1395_n N_VPWR_M1022_d 0.00475326f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_973 N_A_2006_373#_M1022_g N_VPWR_c_1697_n 0.00499688f $X=10.12 $Y=2.565 $X2=0
+ $Y2=0
cc_974 N_A_2006_373#_c_1383_n N_VPWR_c_1698_n 0.0223748f $X=11.69 $Y=1.565 $X2=0
+ $Y2=0
cc_975 N_A_2006_373#_c_1396_n N_VPWR_c_1698_n 0.0171971f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_976 N_A_2006_373#_c_1396_n N_VPWR_c_1709_n 0.00795735f $X=11.23 $Y=2.405
+ $X2=0 $Y2=0
cc_977 N_A_2006_373#_M1022_g N_VPWR_c_1717_n 0.00565381f $X=10.12 $Y=2.565 $X2=0
+ $Y2=0
cc_978 N_A_2006_373#_c_1392_n N_VPWR_c_1717_n 0.00121634f $X=10.405 $Y=2.03
+ $X2=0 $Y2=0
cc_979 N_A_2006_373#_c_1394_n N_VPWR_c_1717_n 0.0239763f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_980 N_A_2006_373#_c_1395_n N_VPWR_c_1717_n 0.0237576f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_981 N_A_2006_373#_c_1396_n N_VPWR_c_1717_n 0.00511833f $X=11.23 $Y=2.405
+ $X2=0 $Y2=0
cc_982 N_A_2006_373#_M1022_g N_VPWR_c_1692_n 0.00587053f $X=10.12 $Y=2.565 $X2=0
+ $Y2=0
cc_983 N_A_2006_373#_c_1394_n N_VPWR_c_1692_n 0.00761719f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_984 N_A_2006_373#_c_1395_n N_VPWR_c_1692_n 0.0010136f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_985 N_A_2006_373#_c_1396_n N_VPWR_c_1692_n 0.0104796f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_986 N_A_2006_373#_c_1383_n Q_N 0.0138022f $X=11.69 $Y=1.565 $X2=0 $Y2=0
cc_987 N_A_2006_373#_c_1386_n N_Q_N_c_2045_n 0.00970057f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_988 N_A_2006_373#_c_1388_n N_Q_N_c_2045_n 0.00199024f $X=11.775 $Y=1.48 $X2=0
+ $Y2=0
cc_989 N_A_2006_373#_c_1388_n Q_N 0.0415299f $X=11.775 $Y=1.48 $X2=0 $Y2=0
cc_990 N_A_2006_373#_c_1386_n N_VGND_M1025_s 0.00517852f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_991 N_A_2006_373#_c_1388_n N_VGND_M1025_s 0.00675628f $X=11.775 $Y=1.48 $X2=0
+ $Y2=0
cc_992 N_A_2006_373#_M1045_g N_VGND_c_2091_n 0.0105628f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_993 N_A_2006_373#_c_1385_n N_VGND_c_2091_n 0.0118606f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_994 N_A_2006_373#_c_1387_n N_VGND_c_2091_n 0.00372607f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_995 N_A_2006_373#_c_1385_n N_VGND_c_2092_n 0.0139523f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_996 N_A_2006_373#_c_1386_n N_VGND_c_2092_n 0.0181192f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_997 N_A_2006_373#_M1045_g N_VGND_c_2102_n 0.00383152f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_998 N_A_2006_373#_c_1385_n N_VGND_c_2105_n 0.0142949f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_999 N_A_2006_373#_c_1386_n N_VGND_c_2105_n 0.00298753f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_1000 N_A_2006_373#_M1045_g N_VGND_c_2114_n 0.0075694f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_1001 N_A_2006_373#_c_1385_n N_VGND_c_2114_n 0.011894f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_1002 N_A_2006_373#_c_1386_n N_VGND_c_2114_n 0.00611276f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_1003 N_A_1790_74#_c_1502_n N_A_2607_392#_c_1646_n 0.0166552f $X=12.945
+ $Y=1.585 $X2=0 $Y2=0
cc_1004 N_A_1790_74#_M1029_g N_A_2607_392#_c_1646_n 0.00200517f $X=12.945
+ $Y=2.46 $X2=0 $Y2=0
cc_1005 N_A_1790_74#_M1010_g N_A_2607_392#_c_1648_n 0.0121223f $X=12.99 $Y=0.69
+ $X2=0 $Y2=0
cc_1006 N_A_1790_74#_M1029_g N_A_2607_392#_c_1649_n 0.0138753f $X=12.945 $Y=2.46
+ $X2=0 $Y2=0
cc_1007 N_A_1790_74#_c_1502_n N_A_2607_392#_c_1650_n 0.0099279f $X=12.945
+ $Y=1.585 $X2=0 $Y2=0
cc_1008 N_A_1790_74#_M1029_g N_A_2607_392#_c_1650_n 0.00145958f $X=12.945
+ $Y=2.46 $X2=0 $Y2=0
cc_1009 N_A_1790_74#_c_1516_n N_VPWR_c_1697_n 0.016504f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_1010 N_A_1790_74#_M1028_g N_VPWR_c_1698_n 0.0132718f $X=11.455 $Y=2.565 $X2=0
+ $Y2=0
cc_1011 N_A_1790_74#_c_1498_n N_VPWR_c_1698_n 0.00119756f $X=11.9 $Y=1.422 $X2=0
+ $Y2=0
cc_1012 N_A_1790_74#_M1005_g N_VPWR_c_1698_n 0.00545542f $X=11.99 $Y=2.4 $X2=0
+ $Y2=0
cc_1013 N_A_1790_74#_M1008_g N_VPWR_c_1699_n 0.00332832f $X=12.44 $Y=2.4 $X2=0
+ $Y2=0
cc_1014 N_A_1790_74#_c_1502_n N_VPWR_c_1699_n 0.00560381f $X=12.945 $Y=1.585
+ $X2=0 $Y2=0
cc_1015 N_A_1790_74#_M1029_g N_VPWR_c_1699_n 0.00366678f $X=12.945 $Y=2.46 $X2=0
+ $Y2=0
cc_1016 N_A_1790_74#_M1029_g N_VPWR_c_1700_n 0.00487483f $X=12.945 $Y=2.46 $X2=0
+ $Y2=0
cc_1017 N_A_1790_74#_M1028_g N_VPWR_c_1709_n 0.00523383f $X=11.455 $Y=2.565
+ $X2=0 $Y2=0
cc_1018 N_A_1790_74#_M1005_g N_VPWR_c_1710_n 0.0049824f $X=11.99 $Y=2.4 $X2=0
+ $Y2=0
cc_1019 N_A_1790_74#_M1008_g N_VPWR_c_1710_n 0.0054356f $X=12.44 $Y=2.4 $X2=0
+ $Y2=0
cc_1020 N_A_1790_74#_M1029_g N_VPWR_c_1711_n 0.00553757f $X=12.945 $Y=2.46 $X2=0
+ $Y2=0
cc_1021 N_A_1790_74#_M1028_g N_VPWR_c_1692_n 0.00587053f $X=11.455 $Y=2.565
+ $X2=0 $Y2=0
cc_1022 N_A_1790_74#_M1005_g N_VPWR_c_1692_n 0.00914025f $X=11.99 $Y=2.4 $X2=0
+ $Y2=0
cc_1023 N_A_1790_74#_M1008_g N_VPWR_c_1692_n 0.0105528f $X=12.44 $Y=2.4 $X2=0
+ $Y2=0
cc_1024 N_A_1790_74#_M1029_g N_VPWR_c_1692_n 0.0109377f $X=12.945 $Y=2.46 $X2=0
+ $Y2=0
cc_1025 N_A_1790_74#_c_1516_n N_VPWR_c_1692_n 0.0290699f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_1026 N_A_1790_74#_c_1516_n A_1958_471# 0.00341864f $X=9.925 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_1027 N_A_1790_74#_M1028_g Q_N 0.00111704f $X=11.455 $Y=2.565 $X2=0 $Y2=0
cc_1028 N_A_1790_74#_M1005_g Q_N 0.0236261f $X=11.99 $Y=2.4 $X2=0 $Y2=0
cc_1029 N_A_1790_74#_M1025_g Q_N 0.00434424f $X=12.085 $Y=0.74 $X2=0 $Y2=0
cc_1030 N_A_1790_74#_M1008_g Q_N 0.020668f $X=12.44 $Y=2.4 $X2=0 $Y2=0
cc_1031 N_A_1790_74#_M1037_g Q_N 0.00444052f $X=12.515 $Y=0.74 $X2=0 $Y2=0
cc_1032 N_A_1790_74#_c_1502_n Q_N 0.0354989f $X=12.945 $Y=1.585 $X2=0 $Y2=0
cc_1033 N_A_1790_74#_M1029_g Q_N 0.0017566f $X=12.945 $Y=2.46 $X2=0 $Y2=0
cc_1034 N_A_1790_74#_M1025_g N_Q_N_c_2045_n 0.0129348f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1035 N_A_1790_74#_M1037_g N_Q_N_c_2045_n 0.0062067f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1036 N_A_1790_74#_M1010_g N_Q_N_c_2045_n 2.82358e-19 $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1037 N_A_1790_74#_M1025_g Q_N 0.00845569f $X=12.085 $Y=0.74 $X2=0 $Y2=0
cc_1038 N_A_1790_74#_M1037_g Q_N 0.00357919f $X=12.515 $Y=0.74 $X2=0 $Y2=0
cc_1039 N_A_1790_74#_M1016_g N_VGND_c_2091_n 0.00182072f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1040 N_A_1790_74#_c_1519_n N_VGND_c_2091_n 0.0208351f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1041 N_A_1790_74#_c_1505_n N_VGND_c_2091_n 0.00424796f $X=10.01 $Y=1.045
+ $X2=0 $Y2=0
cc_1042 N_A_1790_74#_c_1507_n N_VGND_c_2091_n 0.0223381f $X=11.355 $Y=1.175
+ $X2=0 $Y2=0
cc_1043 N_A_1790_74#_M1016_g N_VGND_c_2092_n 0.00310691f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1044 N_A_1790_74#_M1025_g N_VGND_c_2092_n 0.00814486f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1045 N_A_1790_74#_M1037_g N_VGND_c_2093_n 0.0030832f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1046 N_A_1790_74#_c_1502_n N_VGND_c_2093_n 0.00643338f $X=12.945 $Y=1.585
+ $X2=0 $Y2=0
cc_1047 N_A_1790_74#_M1010_g N_VGND_c_2093_n 0.00352391f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1048 N_A_1790_74#_M1010_g N_VGND_c_2094_n 0.00461464f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1049 N_A_1790_74#_M1010_g N_VGND_c_2095_n 0.00385314f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1050 N_A_1790_74#_c_1519_n N_VGND_c_2102_n 0.0202724f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1051 N_A_1790_74#_M1016_g N_VGND_c_2105_n 0.00434272f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1052 N_A_1790_74#_M1025_g N_VGND_c_2106_n 0.00434272f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1053 N_A_1790_74#_M1037_g N_VGND_c_2106_n 0.00434272f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1054 N_A_1790_74#_M1016_g N_VGND_c_2114_n 0.00825669f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1055 N_A_1790_74#_M1025_g N_VGND_c_2114_n 0.00826269f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1056 N_A_1790_74#_M1037_g N_VGND_c_2114_n 0.00820493f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1057 N_A_1790_74#_M1010_g N_VGND_c_2114_n 0.00912981f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1058 N_A_1790_74#_c_1519_n N_VGND_c_2114_n 0.0221648f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1059 N_A_1790_74#_c_1519_n A_2000_74# 0.00371855f $X=9.925 $Y=0.57 $X2=-0.19
+ $Y2=-0.245
cc_1060 N_A_1790_74#_c_1505_n A_2000_74# 5.09211e-19 $X=10.01 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_1061 N_A_2607_392#_c_1649_n N_VPWR_c_1699_n 0.0037413f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1062 N_A_2607_392#_M1001_g N_VPWR_c_1700_n 0.0204468f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1063 N_A_2607_392#_M1044_g N_VPWR_c_1700_n 7.00033e-19 $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1064 N_A_2607_392#_c_1646_n N_VPWR_c_1700_n 0.00687596f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1065 N_A_2607_392#_c_1649_n N_VPWR_c_1700_n 0.07922f $X=13.17 $Y=2.105 $X2=0
+ $Y2=0
cc_1066 N_A_2607_392#_c_1665_p N_VPWR_c_1700_n 0.0252753f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1067 N_A_2607_392#_M1044_g N_VPWR_c_1702_n 0.0053556f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1068 N_A_2607_392#_c_1649_n N_VPWR_c_1711_n 0.0115122f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1069 N_A_2607_392#_M1001_g N_VPWR_c_1712_n 0.00460063f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1070 N_A_2607_392#_M1044_g N_VPWR_c_1712_n 0.005209f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1071 N_A_2607_392#_M1001_g N_VPWR_c_1692_n 0.00908554f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1072 N_A_2607_392#_M1044_g N_VPWR_c_1692_n 0.009853f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1073 N_A_2607_392#_c_1649_n N_VPWR_c_1692_n 0.0095288f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1074 N_A_2607_392#_c_1648_n Q_N 0.00105746f $X=13.205 $Y=0.515 $X2=0 $Y2=0
cc_1075 N_A_2607_392#_M1001_g N_Q_c_2072_n 0.00565021f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1076 N_A_2607_392#_M1018_g N_Q_c_2072_n 0.00531072f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1077 N_A_2607_392#_M1044_g N_Q_c_2072_n 0.0246155f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1078 N_A_2607_392#_M1038_g N_Q_c_2072_n 0.00534388f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1079 N_A_2607_392#_c_1647_n N_Q_c_2072_n 0.0309742f $X=14.4 $Y=1.465 $X2=0
+ $Y2=0
cc_1080 N_A_2607_392#_c_1665_p N_Q_c_2072_n 0.0258081f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1081 N_A_2607_392#_c_1648_n N_VGND_c_2093_n 0.0303376f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1082 N_A_2607_392#_c_1648_n N_VGND_c_2094_n 0.0115122f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1083 N_A_2607_392#_M1018_g N_VGND_c_2095_n 0.00508752f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1084 N_A_2607_392#_c_1646_n N_VGND_c_2095_n 0.00391367f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1085 N_A_2607_392#_c_1648_n N_VGND_c_2095_n 0.0350664f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1086 N_A_2607_392#_c_1665_p N_VGND_c_2095_n 0.014168f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1087 N_A_2607_392#_M1038_g N_VGND_c_2097_n 0.00543765f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1088 N_A_2607_392#_M1018_g N_VGND_c_2107_n 0.00461464f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1089 N_A_2607_392#_M1038_g N_VGND_c_2107_n 0.00461464f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1090 N_A_2607_392#_M1018_g N_VGND_c_2114_n 0.00913331f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1091 N_A_2607_392#_M1038_g N_VGND_c_2114_n 0.00911154f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1092 N_A_2607_392#_c_1648_n N_VGND_c_2114_n 0.0095288f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1093 N_VPWR_c_1693_n N_A_388_79#_c_1893_n 0.0175614f $X=3.28 $Y=2.78 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1707_n N_A_388_79#_c_1893_n 0.0284119f $X=3.115 $Y=3.33 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1714_n N_A_388_79#_c_1893_n 0.00580252f $X=1.4 $Y=3.072 $X2=0
+ $Y2=0
cc_1096 N_VPWR_c_1692_n N_A_388_79#_c_1893_n 0.0333838f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1097 N_VPWR_M1041_d N_A_388_79#_c_1883_n 0.00274897f $X=3.125 $Y=2.415 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1693_n N_A_388_79#_c_1883_n 0.0211681f $X=3.28 $Y=2.78 $X2=0
+ $Y2=0
cc_1099 N_VPWR_c_1692_n N_A_388_79#_c_1883_n 0.00600976f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1692_n N_A_388_79#_c_1886_n 0.00593542f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1703_n N_A_388_79#_c_1887_n 0.0216794f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1692_n N_A_388_79#_c_1887_n 0.01427f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1103 N_VPWR_M1019_d N_A_388_79#_c_1888_n 0.00406554f $X=4.735 $Y=1.935 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1694_n N_A_388_79#_c_1888_n 0.016342f $X=4.87 $Y=2.88 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1703_n N_A_388_79#_c_1888_n 0.0103633f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1106 N_VPWR_c_1705_n N_A_388_79#_c_1888_n 0.00954247f $X=7.07 $Y=3.33 $X2=0
+ $Y2=0
cc_1107 N_VPWR_c_1692_n N_A_388_79#_c_1888_n 0.0364796f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1108 N_VPWR_c_1705_n N_A_388_79#_c_1889_n 0.00586463f $X=7.07 $Y=3.33 $X2=0
+ $Y2=0
cc_1109 N_VPWR_c_1692_n N_A_388_79#_c_1889_n 0.00739256f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1110 N_VPWR_c_1698_n Q_N 0.0430319f $X=11.765 $Y=1.985 $X2=0 $Y2=0
cc_1111 N_VPWR_c_1699_n Q_N 0.0387363f $X=12.665 $Y=2.085 $X2=0 $Y2=0
cc_1112 N_VPWR_c_1710_n Q_N 0.0144623f $X=12.54 $Y=3.33 $X2=0 $Y2=0
cc_1113 N_VPWR_c_1692_n Q_N 0.0118344f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1700_n N_Q_c_2072_n 0.0430489f $X=13.71 $Y=1.985 $X2=0 $Y2=0
cc_1115 N_VPWR_c_1702_n N_Q_c_2072_n 0.0437503f $X=14.61 $Y=1.985 $X2=0 $Y2=0
cc_1116 N_VPWR_c_1712_n N_Q_c_2072_n 0.0118717f $X=14.495 $Y=3.33 $X2=0 $Y2=0
cc_1117 N_VPWR_c_1692_n N_Q_c_2072_n 0.00975826f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1118 N_A_388_79#_c_1893_n A_541_483# 0.00218234f $X=2.775 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1119 N_A_388_79#_c_1904_n A_541_483# 0.00152243f $X=2.86 $Y=2.66 $X2=-0.19
+ $Y2=-0.245
cc_1120 N_A_388_79#_c_1884_n A_541_483# 0.00102652f $X=2.945 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_1121 N_A_388_79#_M1026_d N_noxref_25_c_2246_n 0.011077f $X=1.94 $Y=0.395
+ $X2=0 $Y2=0
cc_1122 N_A_388_79#_c_1874_n N_noxref_25_c_2246_n 0.0217278f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1123 N_A_388_79#_c_1875_n N_noxref_25_c_2246_n 0.0118204f $X=3.445 $Y=1.09
+ $X2=0 $Y2=0
cc_1124 N_A_388_79#_c_1874_n N_noxref_25_c_2248_n 0.00763776f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1125 N_A_388_79#_c_1875_n N_noxref_25_c_2248_n 0.0271448f $X=3.445 $Y=1.09
+ $X2=0 $Y2=0
cc_1126 N_Q_N_c_2045_n N_VGND_c_2092_n 0.010788f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1127 N_Q_N_c_2045_n N_VGND_c_2093_n 0.0272093f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1128 N_Q_N_c_2045_n N_VGND_c_2106_n 0.0144922f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1129 N_Q_N_c_2045_n N_VGND_c_2114_n 0.0118826f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1130 N_Q_c_2072_n N_VGND_c_2095_n 0.00251281f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1131 N_Q_c_2072_n N_VGND_c_2097_n 0.0305242f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1132 N_Q_c_2072_n N_VGND_c_2107_n 0.0119584f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1133 N_Q_c_2072_n N_VGND_c_2114_n 0.00989813f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1134 N_VGND_c_2088_n N_noxref_25_c_2245_n 0.0278855f $X=0.71 $Y=0.605 $X2=0
+ $Y2=0
cc_1135 N_VGND_c_2089_n N_noxref_25_c_2246_n 0.0121474f $X=3.805 $Y=0.605 $X2=0
+ $Y2=0
cc_1136 N_VGND_c_2098_n N_noxref_25_c_2246_n 0.136372f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1137 N_VGND_c_2114_n N_noxref_25_c_2246_n 0.078753f $X=14.64 $Y=0 $X2=0 $Y2=0
cc_1138 N_VGND_c_2088_n N_noxref_25_c_2247_n 0.0125436f $X=0.71 $Y=0.605 $X2=0
+ $Y2=0
cc_1139 N_VGND_c_2098_n N_noxref_25_c_2247_n 0.0177095f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1140 N_VGND_c_2114_n N_noxref_25_c_2247_n 0.00967952f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1141 N_VGND_c_2089_n N_noxref_25_c_2248_n 0.0270493f $X=3.805 $Y=0.605 $X2=0
+ $Y2=0
cc_1142 N_noxref_25_c_2246_n noxref_26 0.00198134f $X=3.1 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1143 N_noxref_25_c_2246_n noxref_27 0.00246354f $X=3.1 $Y=0.34 $X2=-0.19
+ $Y2=-0.245

* File: sky130_fd_sc_ms__a32oi_4.spice
* Created: Wed Sep  2 11:56:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a32oi_4.pex.spice"
.subckt sky130_fd_sc_ms__a32oi_4  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_74#_M1008_d N_B2_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1015 N_A_27_74#_M1015_d N_B2_M1015_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1032 N_A_27_74#_M1015_d N_B2_M1032_g N_VGND_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12765 PD=1.02 PS=1.085 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1035 N_A_27_74#_M1035_d N_B2_M1035_g N_VGND_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12765 PD=1.02 PS=1.085 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75001.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1035_d N_B1_M1018_g N_Y_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1028 N_A_27_74#_M1028_d N_B1_M1028_g N_Y_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1028_d N_B1_M1033_g N_Y_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1038 N_A_27_74#_M1038_d N_B1_M1038_g N_Y_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_868_74#_M1005_d N_A1_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1029 N_A_868_74#_M1029_d N_A1_M1029_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1034 N_A_868_74#_M1029_d N_A1_M1034_g N_Y_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1036 N_A_868_74#_M1036_d N_A1_M1036_g N_Y_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1001 N_A_868_74#_M1036_d N_A2_M1001_g N_A_1313_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1006 N_A_868_74#_M1006_d N_A2_M1006_g N_A_1313_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1022 N_A_868_74#_M1006_d N_A2_M1022_g N_A_1313_74#_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_A_868_74#_M1023_d N_A2_M1023_g N_A_1313_74#_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A3_M1004_g N_A_1313_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A3_M1024_g N_A_1313_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1037 N_VGND_M1024_d N_A3_M1037_g N_A_1313_74#_M1037_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1039 N_VGND_M1039_d N_A3_M1039_g N_A_1313_74#_M1037_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g N_A_27_368#_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.3192 PD=1.435 PS=2.81 NRD=7.0329 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90009.7 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1000_d N_B2_M1007_g N_A_27_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.1512 PD=1.435 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90009.2 A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1010_d N_B2_M1010_g N_A_27_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90008.8 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1010_d N_B2_M1014_g N_A_27_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.6
+ SB=90008.3 A=0.2016 P=2.6 MULT=1
MM1009 N_A_27_368#_M1014_s N_B1_M1009_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.1
+ SB=90007.8 A=0.2016 P=2.6 MULT=1
MM1011 N_A_27_368#_M1011_d N_B1_M1011_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.6
+ SB=90007.3 A=0.2016 P=2.6 MULT=1
MM1012 N_A_27_368#_M1011_d N_B1_M1012_g N_Y_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.1
+ SB=90006.8 A=0.2016 P=2.6 MULT=1
MM1013 N_A_27_368#_M1013_d N_B1_M1013_g N_Y_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2576 AS=0.1792 PD=1.58 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.6
+ SB=90006.3 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_A1_M1016_g N_A_27_368#_M1013_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2576 PD=1.44 PS=1.58 NRD=0 NRS=23.7385 M=1 R=6.22222 SA=90004.2
+ SB=90005.7 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1016_d N_A1_M1017_g N_A_27_368#_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90004.7
+ SB=90005.2 A=0.2016 P=2.6 MULT=1
MM1025 N_VPWR_M1025_d N_A1_M1025_g N_A_27_368#_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90005.2
+ SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1031 N_VPWR_M1025_d N_A1_M1031_g N_A_27_368#_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1568 PD=1.49 PS=1.4 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90005.7
+ SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_27_368#_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.1568 PD=1.48 PS=1.4 NRD=6.1464 NRS=0.8668 M=1 R=6.22222
+ SA=90006.2 SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1002_d N_A2_M1020_g N_A_27_368#_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.1512 PD=1.48 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90006.7
+ SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1026 N_VPWR_M1026_d N_A2_M1026_g N_A_27_368#_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90007.2
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1030 N_VPWR_M1026_d N_A2_M1030_g N_A_27_368#_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90007.7
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1003 N_A_27_368#_M1030_s N_A3_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90008.2
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1019 N_A_27_368#_M1019_d N_A3_M1019_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90008.7
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1021 N_A_27_368#_M1019_d N_A3_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.21 PD=1.44 PS=1.495 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90009.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1027 N_A_27_368#_M1027_d N_A3_M1027_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.21 PD=2.8 PS=1.495 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90009.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.3484 P=25.6
*
.include "sky130_fd_sc_ms__a32oi_4.pxi.spice"
*
.ends
*
*

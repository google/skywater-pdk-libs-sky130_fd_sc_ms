# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__bufinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.250600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.350000 1.390000 0.880000 ;
        RECT 1.060000 0.880000 3.250000 0.960000 ;
        RECT 1.060000 0.960000 4.250000 1.130000 ;
        RECT 1.060000 1.130000 1.390000 1.800000 ;
        RECT 1.060000 1.800000 4.225000 2.070000 ;
        RECT 2.060000 0.350000 2.250000 0.880000 ;
        RECT 2.920000 0.350000 3.250000 0.880000 ;
        RECT 3.920000 0.350000 4.250000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  1.950000 0.445000 2.240000 ;
      RECT 0.115000  2.240000 4.565000 2.410000 ;
      RECT 0.115000  2.410000 0.445000 2.980000 ;
      RECT 0.130000  0.350000 0.380000 1.010000 ;
      RECT 0.130000  1.010000 0.890000 1.180000 ;
      RECT 0.560000  0.085000 0.890000 0.840000 ;
      RECT 0.615000  2.580000 0.945000 3.245000 ;
      RECT 0.720000  1.180000 0.890000 2.240000 ;
      RECT 1.515000  2.580000 1.845000 3.245000 ;
      RECT 1.560000  0.085000 1.890000 0.710000 ;
      RECT 1.665000  1.300000 4.820000 1.630000 ;
      RECT 2.415000  2.580000 2.745000 3.245000 ;
      RECT 2.420000  0.085000 2.750000 0.710000 ;
      RECT 3.315000  2.580000 3.645000 3.245000 ;
      RECT 3.420000  0.085000 3.750000 0.790000 ;
      RECT 4.345000  2.580000 4.675000 3.245000 ;
      RECT 4.395000  1.800000 5.605000 1.970000 ;
      RECT 4.395000  1.970000 4.565000 2.240000 ;
      RECT 4.420000  0.085000 4.750000 0.710000 ;
      RECT 4.650000  0.880000 6.125000 1.130000 ;
      RECT 4.650000  1.130000 4.820000 1.300000 ;
      RECT 4.845000  2.140000 6.125000 2.310000 ;
      RECT 4.845000  2.310000 5.175000 2.980000 ;
      RECT 4.920000  0.350000 5.125000 0.880000 ;
      RECT 4.990000  1.320000 5.605000 1.800000 ;
      RECT 5.295000  0.085000 5.625000 0.710000 ;
      RECT 5.345000  2.480000 5.675000 3.245000 ;
      RECT 5.795000  0.350000 6.125000 0.880000 ;
      RECT 5.795000  1.130000 6.125000 2.140000 ;
      RECT 5.845000  2.310000 6.125000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_ms__bufinv_8
END LIBRARY

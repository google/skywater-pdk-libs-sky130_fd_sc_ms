* NGSPICE file created from sky130_fd_sc_ms__clkinv_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__clkinv_2 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=6.16e+11p ps=5.58e+06u
M1001 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=2.394e+11p pd=2.82e+06u as=3.276e+11p ps=2.4e+06u
M1003 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


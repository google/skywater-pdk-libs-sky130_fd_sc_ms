* File: sky130_fd_sc_ms__and4_4.spice
* Created: Fri Aug 28 17:13:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4_4.pex.spice"
.subckt sky130_fd_sc_ms__and4_4  VNB VPB A B D C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* D	D
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_A_119_119#_M1005_d N_B_M1005_g N_A_32_119#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_119_392#_M1003_d N_A_M1003_g N_A_119_119#_M1005_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1006 N_A_119_392#_M1003_d N_A_M1006_g N_A_119_119#_M1006_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1018 N_A_119_119#_M1006_s N_B_M1018_g N_A_32_119#_M1018_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_463_119#_M1019_d N_C_M1019_g N_A_32_119#_M1018_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1016 N_VGND_M1016_d N_D_M1016_g N_A_463_119#_M1019_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.170525 AS=0.0896 PD=1.285 PS=0.92 NRD=39.636 NRS=0 M=1 R=4.26667
+ SA=75002.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1016_d N_D_M1020_g N_A_463_119#_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.170525 AS=0.0896 PD=1.285 PS=0.92 NRD=39.636 NRS=0 M=1 R=4.26667
+ SA=75002.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_463_119#_M1020_s N_C_M1021_g N_A_32_119#_M1021_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1705 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_A_119_392#_M1008_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2405 AS=0.1147 PD=2.13 PS=1.05 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_119_392#_M1017_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1147 PD=1.09 PS=1.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1017_d N_A_119_392#_M1022_g N_X_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_119_392#_M1023_g N_X_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.1036 PD=2.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_119_392#_M1001_d N_B_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_119_392#_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90005.4 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1002_d N_A_M1004_g N_A_119_392#_M1004_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.1425 PD=1.27 PS=1.285 NRD=0 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1014 N_A_119_392#_M1004_s N_B_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1
+ AD=0.1425 AS=0.16 PD=1.285 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1014_s N_C_M1011_g N_A_119_392#_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.135 PD=1.32 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90002.1
+ SB=90004 A=0.18 P=2.36 MULT=1
MM1012 N_A_119_392#_M1011_s N_D_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.3525 PD=1.27 PS=1.705 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.5
+ SB=90003.6 A=0.18 P=2.36 MULT=1
MM1015 N_A_119_392#_M1015_d N_D_M1015_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.3525 PD=1.32 PS=1.705 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90003.4
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_C_M1013_g N_A_119_392#_M1015_d VPB PSHORT L=0.18 W=1
+ AD=0.193396 AS=0.16 PD=1.41509 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90003.9 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_119_392#_M1000_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.216604 PD=1.44 PS=1.58491 NRD=7.8997 NRS=9.6727 M=1 R=6.22222
+ SA=90004 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1000_d N_A_119_392#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1009_d N_A_119_392#_M1009_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.9
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1010 N_X_M1009_d N_A_119_392#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90005.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_73 VNB 0 4.03451e-19 $X=0 $Y=0
c_135 VPB 0 7.60421e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__and4_4.pxi.spice"
*
.ends
*
*

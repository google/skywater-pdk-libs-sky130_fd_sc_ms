* File: sky130_fd_sc_ms__and4_2.pex.spice
* Created: Wed Sep  2 11:58:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4_2%A 3 7 9 10 11 15
c29 10 0 1.05466e-19 $X=0.505 $Y=1.3
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.465 $X2=0.28 $Y2=1.465
r31 11 15 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.28 $Y=1.665 $X2=0.28
+ $Y2=1.465
r32 9 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.28 $Y2=1.465
r33 9 10 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=1.3
r34 5 10 34.7346 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=0.64 $Y=1.3
+ $X2=0.505 $Y2=1.3
r35 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.64 $Y=1.3 $X2=0.64
+ $Y2=0.74
r36 1 10 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=0.595 $Y=1.63
+ $X2=0.505 $Y2=1.3
r37 1 3 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=0.595 $Y=1.63
+ $X2=0.595 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%B 3 6 8 9 10 15 17
c37 8 0 1.05466e-19 $X=1.2 $Y=0.555
r38 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.385
+ $X2=1.12 $Y2=1.55
r39 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.385
+ $X2=1.12 $Y2=1.22
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.385 $X2=1.12 $Y2=1.385
r41 10 16 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.385
r42 9 10 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.925
+ $X2=1.135 $Y2=1.295
r43 8 9 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.555
+ $X2=1.135 $Y2=0.925
r44 6 18 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=1.045 $Y=2.46
+ $X2=1.045 $Y2=1.55
r45 3 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.03 $Y=0.74 $X2=1.03
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%C 3 6 8 9 10 15 17
c35 17 0 1.05261e-19 $X=1.69 $Y=1.22
r36 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.55
r37 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=1.69 $Y2=1.22
r38 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.385 $X2=1.69 $Y2=1.385
r39 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.385
r40 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.295
r41 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.555 $X2=1.69
+ $Y2=0.925
r42 6 18 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=1.705 $Y=2.46
+ $X2=1.705 $Y2=1.55
r43 3 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.6 $Y=0.74 $X2=1.6
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%D 1 3 6 9 10 13 14 15
c38 14 0 1.05261e-19 $X=2.26 $Y=1.385
r39 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.385
+ $X2=2.26 $Y2=1.55
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.385
+ $X2=2.26 $Y2=1.22
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.385 $X2=2.26 $Y2=1.385
r42 10 14 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.365 $X2=2.26
+ $Y2=1.365
r43 9 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.17 $Y=1.79 $X2=2.17
+ $Y2=1.55
r44 6 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.17 $Y=0.74 $X2=2.17
+ $Y2=1.22
r45 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.155 $Y=1.88 $X2=2.155
+ $Y2=1.79
r46 1 3 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.155 $Y=1.88
+ $X2=2.155 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%A_56_74# 1 2 3 12 16 20 24 26 33 36 39 43 48
+ 51 53 57 58 62 64 65
r110 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.465 $X2=3.57 $Y2=1.465
r111 55 57 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.57 $Y=2.32
+ $X2=3.57 $Y2=1.465
r112 54 65 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=2.405
+ $X2=1.93 $Y2=2.405
r113 53 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.405 $Y=2.405
+ $X2=3.57 $Y2=2.32
r114 53 54 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.405 $Y=2.405
+ $X2=2.095 $Y2=2.405
r115 49 65 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.49
+ $X2=1.93 $Y2=2.405
r116 49 51 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.93 $Y=2.49
+ $X2=1.93 $Y2=2.815
r117 46 65 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=2.32
+ $X2=1.93 $Y2=2.405
r118 46 48 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.93 $Y=2.32
+ $X2=1.93 $Y2=2.105
r119 45 48 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.93 $Y=1.89
+ $X2=1.93 $Y2=2.105
r120 44 64 3.05049 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.985 $Y=1.805
+ $X2=0.8 $Y2=1.805
r121 43 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.765 $Y=1.805
+ $X2=1.93 $Y2=1.89
r122 43 44 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.765 $Y=1.805
+ $X2=0.985 $Y2=1.805
r123 39 41 22.1144 $w=3.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.8 $Y=2.105
+ $X2=0.8 $Y2=2.815
r124 37 64 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.89 $X2=0.8
+ $Y2=1.805
r125 37 39 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.8 $Y=1.89
+ $X2=0.8 $Y2=2.105
r126 36 64 3.46198 $w=2.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.7 $Y=1.72
+ $X2=0.8 $Y2=1.805
r127 35 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.13 $X2=0.7
+ $Y2=1.045
r128 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.7 $Y=1.13 $X2=0.7
+ $Y2=1.72
r129 31 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.425 $Y=1.045
+ $X2=0.7 $Y2=1.045
r130 31 33 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.425 $Y=0.96
+ $X2=0.425 $Y2=0.515
r131 29 30 8.60714 $w=3.08e-07 $l=5.5e-08 $layer=POLY_cond $X=3.17 $Y=1.465
+ $X2=3.225 $Y2=1.465
r132 26 58 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.315 $Y=1.465
+ $X2=3.57 $Y2=1.465
r133 26 30 13.428 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.315 $Y=1.465
+ $X2=3.225 $Y2=1.465
r134 22 30 15.3289 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=1.63
+ $X2=3.225 $Y2=1.465
r135 22 24 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.225 $Y=1.63
+ $X2=3.225 $Y2=2.4
r136 18 29 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.3
+ $X2=3.17 $Y2=1.465
r137 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.17 $Y=1.3
+ $X2=3.17 $Y2=0.74
r138 14 29 61.8149 $w=3.08e-07 $l=3.95e-07 $layer=POLY_cond $X=2.775 $Y=1.465
+ $X2=3.17 $Y2=1.465
r139 14 27 5.47727 $w=3.08e-07 $l=3.5e-08 $layer=POLY_cond $X=2.775 $Y=1.465
+ $X2=2.74 $Y2=1.465
r140 14 16 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=2.775 $Y=1.6
+ $X2=2.775 $Y2=2.4
r141 10 27 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.3
+ $X2=2.74 $Y2=1.465
r142 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.74 $Y=1.3
+ $X2=2.74 $Y2=0.74
r143 3 51 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.96 $X2=1.93 $Y2=2.815
r144 3 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.96 $X2=1.93 $Y2=2.105
r145 2 41 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=1.96 $X2=0.82 $Y2=2.815
r146 2 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=1.96 $X2=0.82 $Y2=2.105
r147 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.28
+ $Y=0.37 $X2=0.425 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%VPWR 1 2 3 4 13 15 21 25 27 29 32 33 35 36 37
+ 46 55
r50 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 49 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 46 54 4.96106 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.605 $Y2=3.33
r55 46 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 45 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 39 51 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r61 39 41 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 37 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 37 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 35 44 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33 $X2=2.16
+ $Y2=3.33
r65 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.465 $Y2=3.33
r66 34 48 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=2.465 $Y2=3.33
r68 32 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.215 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=3.33
+ $X2=1.38 $Y2=3.33
r70 31 44 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.38 $Y2=3.33
r72 27 54 3.01886 $w=3.55e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.547 $Y=3.245
+ $X2=3.605 $Y2=3.33
r73 27 29 14.6084 $w=3.53e-07 $l=4.5e-07 $layer=LI1_cond $X=3.547 $Y=3.245
+ $X2=3.547 $Y2=2.795
r74 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=3.33
r75 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=2.795
r76 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=3.245
+ $X2=1.38 $Y2=3.33
r77 19 21 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=1.38 $Y=3.245
+ $X2=1.38 $Y2=2.195
r78 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r79 13 51 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r80 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r81 4 29 600 $w=1.7e-07 $l=1.0638e-06 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.84 $X2=3.545 $Y2=2.795
r82 3 25 600 $w=1.7e-07 $l=9.38576e-07 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.96 $X2=2.465 $Y2=2.795
r83 2 21 300 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.96 $X2=1.38 $Y2=2.195
r84 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r85 1 15 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%X 1 2 7 8 9 10 26
r20 10 21 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=3.035 $Y=2.035
+ $X2=3.035 $Y2=1.985
r21 9 21 9.21954 $w=3.98e-07 $l=3.2e-07 $layer=LI1_cond $X=3.035 $Y=1.665
+ $X2=3.035 $Y2=1.985
r22 8 9 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.665
r23 8 30 4.75383 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=1.295
+ $X2=3.035 $Y2=1.13
r24 7 30 5.45223 $w=4.43e-07 $l=2.05e-07 $layer=LI1_cond $X=3.012 $Y=0.925
+ $X2=3.012 $Y2=1.13
r25 7 26 0.388464 $w=4.43e-07 $l=1.5e-08 $layer=LI1_cond $X=3.012 $Y=0.925
+ $X2=3.012 $Y2=0.91
r26 2 21 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.84 $X2=3 $Y2=1.985
r27 1 26 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_2%VGND 1 2 9 11 12 15 18 19 21 23 32 38
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r43 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 32 37 5.51088 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.53
+ $Y2=0
r46 32 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.12
+ $Y2=0
r47 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r48 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 26 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r50 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r52 23 27 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r53 21 22 4.31883 $w=4.33e-07 $l=8.5e-08 $layer=LI1_cond $X=3.437 $Y=0.515
+ $X2=3.437 $Y2=0.6
r54 18 30 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.16
+ $Y2=0
r55 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.43
+ $Y2=0
r56 17 34 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=3.12
+ $Y2=0
r57 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.43
+ $Y2=0
r58 15 22 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.53 $Y=0.915
+ $X2=3.53 $Y2=0.6
r59 12 21 3.49707 $w=4.33e-07 $l=1.32e-07 $layer=LI1_cond $X=3.437 $Y=0.383
+ $X2=3.437 $Y2=0.515
r60 11 37 3.16431 $w=4.35e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.53 $Y2=0
r61 11 12 7.8949 $w=4.33e-07 $l=2.98e-07 $layer=LI1_cond $X=3.437 $Y=0.085
+ $X2=3.437 $Y2=0.383
r62 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.085 $X2=2.43
+ $Y2=0
r63 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.43 $Y=0.085 $X2=2.43
+ $Y2=0.495
r64 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.37 $X2=3.385 $Y2=0.515
r65 2 15 182 $w=1.7e-07 $l=6.56163e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.37 $X2=3.49 $Y2=0.915
r66 1 9 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.37 $X2=2.43 $Y2=0.495
.ends


* NGSPICE file created from sky130_fd_sc_ms__sedfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1377_368# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=3.44925e+12p ps=2.926e+07u
M1001 a_141_74# D a_32_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.835e+11p ps=3.03e+06u
M1002 VPWR a_575_87# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1003 VPWR a_183_290# a_135_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1004 a_1586_74# a_1377_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.61097e+12p ps=2.285e+07u
M1005 a_32_74# a_575_87# a_527_113# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_575_87# a_2675_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 a_2417_74# a_2013_71# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 a_1586_74# a_1377_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1009 a_691_113# a_661_87# a_32_74# VNB nlowvt w=420000u l=150000u
+  ad=3.885e+11p pd=4.37e+06u as=0p ps=0u
M1010 a_2489_74# a_1586_74# a_2417_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1011 a_2591_74# a_1377_368# a_2489_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_575_87# a_2489_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 VPWR DE a_183_290# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1014 VPWR SCE a_661_87# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1015 a_1784_97# a_1586_74# a_691_113# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.76e+11p ps=5.08e+06u
M1016 VPWR a_2013_71# a_1947_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1017 a_1091_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_2013_71# a_1784_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1019 a_1947_508# a_1377_368# a_1784_97# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND DE a_183_290# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1021 a_527_113# a_183_290# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_575_87# a_2591_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_575_87# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1024 a_32_74# a_575_87# a_581_462# VPB pshort w=640000u l=180000u
+  ad=3.52e+11p pd=3.66e+06u as=1.344e+11p ps=1.7e+06u
M1025 VGND a_2013_71# a_1920_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.953e+11p ps=1.77e+06u
M1026 Q a_2489_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1027 a_135_464# D a_32_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_691_113# SCE a_32_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1377_368# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1030 a_2675_508# a_1586_74# a_2489_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.115e+11p ps=2.71e+06u
M1031 a_1091_453# SCD VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1032 a_2013_71# a_1784_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1033 a_691_113# SCE a_1091_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2489_74# a_1377_368# a_2377_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.75e+11p ps=3.55e+06u
M1035 a_1784_97# a_1377_368# a_691_113# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1036 Q a_2489_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1037 VGND SCE a_661_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1038 a_1920_97# a_1586_74# a_1784_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_2489_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_691_113# a_661_87# a_1091_453# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_575_87# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND DE a_141_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_2377_392# a_2013_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_575_87# a_2489_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1045 a_581_462# DE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Q_N a_575_87# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_2489_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


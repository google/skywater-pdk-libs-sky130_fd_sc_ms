# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ms__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__a22o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.450000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 0.255000 5.320000 0.505000 ;
        RECT 4.955000 0.505000 5.125000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.495000 1.435000 3.825000 1.765000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.435000 3.325000 1.765000 ;
        RECT 3.155000 1.765000 3.325000 1.935000 ;
        RECT 3.155000 1.935000 4.195000 2.150000 ;
        RECT 4.025000 1.440000 4.655000 1.770000 ;
        RECT 4.025000 1.770000 4.195000 1.935000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 2.515000 1.180000 ;
        RECT 0.125000 1.180000 1.855000 1.410000 ;
        RECT 0.705000 1.410000 1.855000 1.650000 ;
        RECT 0.705000 1.650000 0.875000 2.980000 ;
        RECT 1.405000 0.480000 1.655000 1.010000 ;
        RECT 1.405000 1.010000 2.515000 1.140000 ;
        RECT 1.525000 1.650000 1.855000 2.980000 ;
        RECT 2.265000 0.480000 2.515000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 7.200000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 7.390000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.175000  1.900000 0.505000 3.245000 ;
      RECT 0.975000  0.085000 1.225000 0.970000 ;
      RECT 1.075000  1.820000 1.325000 3.245000 ;
      RECT 1.835000  0.085000 2.085000 0.840000 ;
      RECT 2.025000  1.350000 2.855000 1.680000 ;
      RECT 2.055000  1.850000 2.305000 3.245000 ;
      RECT 2.475000  1.680000 2.645000 2.905000 ;
      RECT 2.475000  2.905000 4.415000 2.980000 ;
      RECT 2.475000  2.980000 3.515000 3.075000 ;
      RECT 2.685000  1.095000 6.055000 1.265000 ;
      RECT 2.685000  1.265000 2.855000 1.350000 ;
      RECT 2.695000  0.085000 3.025000 0.925000 ;
      RECT 2.815000  1.940000 2.985000 2.320000 ;
      RECT 2.815000  2.320000 4.865000 2.490000 ;
      RECT 2.815000  2.490000 2.985000 2.735000 ;
      RECT 3.185000  2.660000 4.415000 2.905000 ;
      RECT 3.200000  0.580000 4.355000 0.830000 ;
      RECT 3.630000  1.000000 3.960000 1.095000 ;
      RECT 4.140000  0.830000 4.355000 0.925000 ;
      RECT 4.535000  0.085000 4.785000 0.925000 ;
      RECT 4.615000  1.940000 4.865000 1.950000 ;
      RECT 4.615000  1.950000 6.910000 2.120000 ;
      RECT 4.615000  2.120000 4.865000 2.320000 ;
      RECT 4.615000  2.490000 4.865000 2.980000 ;
      RECT 5.035000  2.290000 5.510000 3.245000 ;
      RECT 5.295000  0.675000 6.405000 0.845000 ;
      RECT 5.680000  2.120000 5.930000 2.980000 ;
      RECT 5.725000  1.015000 6.055000 1.095000 ;
      RECT 5.725000  1.265000 6.055000 1.275000 ;
      RECT 6.130000  2.290000 6.460000 3.245000 ;
      RECT 6.235000  0.595000 6.405000 0.675000 ;
      RECT 6.235000  0.845000 6.405000 1.275000 ;
      RECT 6.585000  0.085000 6.915000 1.275000 ;
      RECT 6.660000  1.940000 6.910000 1.950000 ;
      RECT 6.660000  2.120000 6.910000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_ms__a22o_4
END LIBRARY

* NGSPICE file created from sky130_fd_sc_ms__clkdlyinv5sd2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__clkdlyinv5sd2_1 A VGND VNB VPB VPWR Y
M1000 a_549_74# a_288_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=7.371e+11p ps=6.03e+06u
M1001 VGND a_549_74# a_682_74# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.457e+11p ps=2.01e+06u
M1002 Y a_682_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 a_549_74# a_288_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=1.6512e+12p ps=9.66e+06u
M1004 VPWR a_549_74# a_682_74# VPB pshort w=1e+06u l=250000u
+  ad=0p pd=0u as=5.1e+11p ps=3.02e+06u
M1005 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1007 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 Y a_682_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1009 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__nor4bb_1.spice
* Created: Wed Sep  2 12:17:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4bb_1.pex.spice"
.subckt sky130_fd_sc_ms__nor4bb_1  VNB VPB C_N A B D_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D_N	D_N
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_C_N_M1003_g N_A_27_112#_M1003_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.142488 AS=0.3025 PD=1.04457 PS=2.2 NRD=30 NRS=0 M=1 R=3.66667 SA=75000.5
+ SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.191712 PD=1.09 PS=1.40543 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.9
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_Y_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.25715 AS=0.1295 PD=1.435 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_A_27_112#_M1008_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.25715 PD=1.09 PS=1.435 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_611_244#_M1007_g N_Y_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.38024 AS=0.1295 PD=1.89876 PS=1.09 NRD=18.648 NRS=0 M=1 R=4.93333
+ SA=75002.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_611_244#_M1004_d N_D_N_M1004_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.15675 AS=0.28261 PD=1.67 PS=1.41124 NRD=0 NRS=18 M=1 R=3.66667
+ SA=75004 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1006 N_VPWR_M1006_d N_C_N_M1006_g N_A_27_112#_M1006_s VPB PSHORT L=0.18 W=0.84
+ AD=0.425121 AS=0.2352 PD=1.79571 PS=2.24 NRD=105.789 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.8 A=0.1512 P=2.04 MULT=1
MM1011 A_316_368# N_A_M1011_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.566829 PD=1.36 PS=2.39429 NRD=11.426 NRS=14.9326 M=1 R=6.22222 SA=90001
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1001 A_400_368# N_B_M1001_g A_316_368# VPB PSHORT L=0.18 W=1.12 AD=0.2716
+ AS=0.1344 PD=1.605 PS=1.36 NRD=32.9778 NRS=11.426 M=1 R=6.22222 SA=90001.5
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1002 A_533_368# N_A_27_112#_M1002_g A_400_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.2184 AS=0.2716 PD=1.51 PS=1.605 NRD=24.6053 NRS=32.9778 M=1 R=6.22222
+ SA=90002.1 SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_A_611_244#_M1005_g A_533_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90002.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_611_244#_M1000_d N_D_N_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2184 PD=2.24 PS=2.2 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
DX12_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__nor4bb_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfrtp_4.pxi.spice
* Created: Fri Aug 28 17:23:10 2020
* 
x_PM_SKY130_FD_SC_MS__DFRTP_4%D N_D_c_276_n N_D_c_281_n N_D_M1034_g N_D_M1017_g
+ N_D_c_283_n D D D N_D_c_278_n N_D_c_279_n N_D_c_285_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%D
x_PM_SKY130_FD_SC_MS__DFRTP_4%CLK N_CLK_M1010_g N_CLK_M1001_g CLK N_CLK_c_313_n
+ N_CLK_c_314_n N_CLK_c_317_n PM_SKY130_FD_SC_MS__DFRTP_4%CLK
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_497_395# N_A_497_395#_M1002_d
+ N_A_497_395#_M1013_d N_A_497_395#_c_359_n N_A_497_395#_M1014_g
+ N_A_497_395#_c_360_n N_A_497_395#_c_361_n N_A_497_395#_M1036_g
+ N_A_497_395#_c_363_n N_A_497_395#_M1004_g N_A_497_395#_c_364_n
+ N_A_497_395#_c_365_n N_A_497_395#_M1007_g N_A_497_395#_c_383_n
+ N_A_497_395#_c_366_n N_A_497_395#_c_367_n N_A_497_395#_c_368_n
+ N_A_497_395#_c_369_n N_A_497_395#_c_370_n N_A_497_395#_c_371_n
+ N_A_497_395#_c_372_n N_A_497_395#_c_373_n N_A_497_395#_c_374_n
+ N_A_497_395#_c_375_n N_A_497_395#_c_376_n N_A_497_395#_c_377_n
+ N_A_497_395#_c_386_n PM_SKY130_FD_SC_MS__DFRTP_4%A_497_395#
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_834_355# N_A_834_355#_M1011_d
+ N_A_834_355#_M1015_d N_A_834_355#_M1006_g N_A_834_355#_M1024_g
+ N_A_834_355#_c_558_n N_A_834_355#_c_563_n N_A_834_355#_c_574_n
+ N_A_834_355#_c_559_n N_A_834_355#_c_576_n N_A_834_355#_c_602_p
+ N_A_834_355#_c_577_n N_A_834_355#_c_565_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%A_834_355#
x_PM_SKY130_FD_SC_MS__DFRTP_4%RESET_B N_RESET_B_M1005_g N_RESET_B_c_648_n
+ N_RESET_B_M1035_g N_RESET_B_c_649_n N_RESET_B_c_650_n N_RESET_B_M1033_g
+ N_RESET_B_M1016_g N_RESET_B_c_652_n N_RESET_B_M1026_g N_RESET_B_M1030_g
+ N_RESET_B_c_654_n N_RESET_B_c_663_n N_RESET_B_c_664_n N_RESET_B_c_665_n
+ N_RESET_B_c_666_n N_RESET_B_c_667_n N_RESET_B_c_668_n N_RESET_B_c_669_n
+ N_RESET_B_c_670_n RESET_B N_RESET_B_c_671_n N_RESET_B_c_655_n
+ N_RESET_B_c_656_n N_RESET_B_c_673_n N_RESET_B_c_674_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%RESET_B
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_303_395# N_A_303_395#_M1001_s
+ N_A_303_395#_M1010_s N_A_303_395#_c_889_n N_A_303_395#_M1013_g
+ N_A_303_395#_c_877_n N_A_303_395#_M1002_g N_A_303_395#_c_890_n
+ N_A_303_395#_c_891_n N_A_303_395#_c_892_n N_A_303_395#_c_878_n
+ N_A_303_395#_c_879_n N_A_303_395#_c_880_n N_A_303_395#_M1000_g
+ N_A_303_395#_M1019_g N_A_303_395#_c_895_n N_A_303_395#_c_896_n
+ N_A_303_395#_c_881_n N_A_303_395#_M1020_g N_A_303_395#_c_882_n
+ N_A_303_395#_M1037_g N_A_303_395#_c_900_n N_A_303_395#_c_884_n
+ N_A_303_395#_c_914_n N_A_303_395#_c_885_n N_A_303_395#_c_901_n
+ N_A_303_395#_c_902_n N_A_303_395#_c_886_n N_A_303_395#_c_903_n
+ N_A_303_395#_c_887_n N_A_303_395#_c_905_n N_A_303_395#_c_906_n
+ N_A_303_395#_c_888_n PM_SKY130_FD_SC_MS__DFRTP_4%A_303_395#
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_702_463# N_A_702_463#_M1000_d
+ N_A_702_463#_M1014_d N_A_702_463#_M1016_d N_A_702_463#_c_1103_n
+ N_A_702_463#_M1011_g N_A_702_463#_c_1112_n N_A_702_463#_M1015_g
+ N_A_702_463#_c_1104_n N_A_702_463#_c_1105_n N_A_702_463#_c_1106_n
+ N_A_702_463#_c_1107_n N_A_702_463#_c_1143_n N_A_702_463#_c_1108_n
+ N_A_702_463#_c_1109_n N_A_702_463#_c_1110_n N_A_702_463#_c_1111_n
+ N_A_702_463#_c_1117_n N_A_702_463#_c_1118_n N_A_702_463#_c_1119_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%A_702_463#
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_1678_395# N_A_1678_395#_M1031_d
+ N_A_1678_395#_M1026_d N_A_1678_395#_M1012_g N_A_1678_395#_M1022_g
+ N_A_1678_395#_c_1242_n N_A_1678_395#_c_1251_n N_A_1678_395#_c_1243_n
+ N_A_1678_395#_c_1252_n N_A_1678_395#_c_1253_n N_A_1678_395#_c_1254_n
+ N_A_1678_395#_c_1244_n N_A_1678_395#_c_1245_n N_A_1678_395#_c_1246_n
+ N_A_1678_395#_c_1247_n N_A_1678_395#_c_1256_n N_A_1678_395#_c_1248_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%A_1678_395#
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_1353_392# N_A_1353_392#_M1004_d
+ N_A_1353_392#_M1020_d N_A_1353_392#_M1031_g N_A_1353_392#_M1027_g
+ N_A_1353_392#_c_1364_n N_A_1353_392#_M1008_g N_A_1353_392#_c_1365_n
+ N_A_1353_392#_M1025_g N_A_1353_392#_c_1366_n N_A_1353_392#_M1018_g
+ N_A_1353_392#_c_1367_n N_A_1353_392#_c_1368_n N_A_1353_392#_c_1369_n
+ N_A_1353_392#_c_1370_n N_A_1353_392#_c_1391_n N_A_1353_392#_c_1371_n
+ N_A_1353_392#_c_1372_n N_A_1353_392#_c_1406_n N_A_1353_392#_c_1385_n
+ N_A_1353_392#_c_1373_n N_A_1353_392#_c_1374_n N_A_1353_392#_c_1375_n
+ N_A_1353_392#_c_1376_n PM_SKY130_FD_SC_MS__DFRTP_4%A_1353_392#
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_2013_409# N_A_2013_409#_M1018_d
+ N_A_2013_409#_M1008_s N_A_2013_409#_M1009_g N_A_2013_409#_c_1527_n
+ N_A_2013_409#_M1021_g N_A_2013_409#_M1003_g N_A_2013_409#_c_1530_n
+ N_A_2013_409#_c_1531_n N_A_2013_409#_M1023_g N_A_2013_409#_M1028_g
+ N_A_2013_409#_M1032_g N_A_2013_409#_M1029_g N_A_2013_409#_M1038_g
+ N_A_2013_409#_c_1548_n N_A_2013_409#_c_1537_n N_A_2013_409#_c_1538_n
+ N_A_2013_409#_c_1539_n N_A_2013_409#_c_1540_n N_A_2013_409#_c_1541_n
+ N_A_2013_409#_c_1542_n N_A_2013_409#_c_1543_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%A_2013_409#
x_PM_SKY130_FD_SC_MS__DFRTP_4%VPWR N_VPWR_M1034_s N_VPWR_M1035_d N_VPWR_M1010_d
+ N_VPWR_M1006_d N_VPWR_M1015_s N_VPWR_M1012_d N_VPWR_M1027_d N_VPWR_M1025_d
+ N_VPWR_M1021_s N_VPWR_M1029_s N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n
+ N_VPWR_c_1656_n N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n
+ N_VPWR_c_1660_n N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n
+ N_VPWR_c_1664_n N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1667_n
+ N_VPWR_c_1668_n N_VPWR_c_1669_n N_VPWR_c_1670_n VPWR N_VPWR_c_1671_n
+ N_VPWR_c_1672_n N_VPWR_c_1673_n N_VPWR_c_1674_n N_VPWR_c_1675_n
+ N_VPWR_c_1676_n N_VPWR_c_1677_n N_VPWR_c_1678_n N_VPWR_c_1679_n
+ N_VPWR_c_1680_n N_VPWR_c_1681_n N_VPWR_c_1652_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%VPWR
x_PM_SKY130_FD_SC_MS__DFRTP_4%A_37_78# N_A_37_78#_M1017_s N_A_37_78#_M1000_s
+ N_A_37_78#_M1034_d N_A_37_78#_M1014_s N_A_37_78#_c_1822_n N_A_37_78#_c_1829_n
+ N_A_37_78#_c_1823_n N_A_37_78#_c_1831_n N_A_37_78#_c_1824_n
+ N_A_37_78#_c_1832_n N_A_37_78#_c_1825_n N_A_37_78#_c_1826_n
+ N_A_37_78#_c_1827_n N_A_37_78#_c_1828_n N_A_37_78#_c_1834_n
+ N_A_37_78#_c_1835_n PM_SKY130_FD_SC_MS__DFRTP_4%A_37_78#
x_PM_SKY130_FD_SC_MS__DFRTP_4%Q N_Q_M1003_s N_Q_M1032_s N_Q_M1009_d N_Q_M1028_d
+ N_Q_c_1950_n N_Q_c_1951_n N_Q_c_1952_n N_Q_c_1943_n N_Q_c_1944_n N_Q_c_1945_n
+ N_Q_c_1953_n N_Q_c_1946_n N_Q_c_1947_n N_Q_c_1948_n Q
+ PM_SKY130_FD_SC_MS__DFRTP_4%Q
x_PM_SKY130_FD_SC_MS__DFRTP_4%VGND N_VGND_M1005_d N_VGND_M1001_d N_VGND_M1033_d
+ N_VGND_M1022_d N_VGND_M1018_s N_VGND_M1003_d N_VGND_M1023_d N_VGND_M1038_d
+ N_VGND_c_2015_n N_VGND_c_2016_n N_VGND_c_2017_n N_VGND_c_2018_n
+ N_VGND_c_2019_n N_VGND_c_2020_n N_VGND_c_2021_n N_VGND_c_2022_n
+ N_VGND_c_2023_n N_VGND_c_2024_n N_VGND_c_2025_n N_VGND_c_2026_n VGND
+ N_VGND_c_2027_n N_VGND_c_2028_n N_VGND_c_2029_n N_VGND_c_2030_n
+ N_VGND_c_2031_n N_VGND_c_2032_n N_VGND_c_2033_n N_VGND_c_2034_n
+ N_VGND_c_2035_n N_VGND_c_2036_n N_VGND_c_2037_n N_VGND_c_2038_n
+ PM_SKY130_FD_SC_MS__DFRTP_4%VGND
cc_1 VNB N_D_c_276_n 0.0407866f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.81
cc_2 VNB N_D_M1017_g 0.0286444f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_3 VNB N_D_c_278_n 0.0249067f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_279_n 0.0295836f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB CLK 0.00319184f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_6 VNB N_CLK_c_313_n 0.0309384f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_7 VNB N_CLK_c_314_n 0.0141294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_497_395#_c_359_n 0.00905176f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_9 VNB N_A_497_395#_c_360_n 0.00919935f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_10 VNB N_A_497_395#_c_361_n 0.021231f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.35
cc_11 VNB N_A_497_395#_M1036_g 0.0235332f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A_497_395#_c_363_n 0.0216455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_497_395#_c_364_n 0.0206494f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.165
cc_14 VNB N_A_497_395#_c_365_n 0.00999606f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_15 VNB N_A_497_395#_c_366_n 0.00701139f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_16 VNB N_A_497_395#_c_367_n 0.0319818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_497_395#_c_368_n 0.0030128f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_18 VNB N_A_497_395#_c_369_n 0.0255302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_497_395#_c_370_n 0.00585827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_497_395#_c_371_n 0.00192671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_497_395#_c_372_n 0.0152924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_497_395#_c_373_n 0.00355484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_497_395#_c_374_n 0.00607047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_497_395#_c_375_n 0.00241598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_497_395#_c_376_n 0.030848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_497_395#_c_377_n 0.00738738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_834_355#_M1024_g 0.034709f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.35
cc_28 VNB N_A_834_355#_c_558_n 0.00382242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_834_355#_c_559_n 0.00906432f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1
cc_30 VNB N_RESET_B_M1005_g 0.0222451f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.245
cc_31 VNB N_RESET_B_c_648_n 0.0275322f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_32 VNB N_RESET_B_c_649_n 0.275673f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_33 VNB N_RESET_B_c_650_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_RESET_B_M1033_g 0.03486f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_35 VNB N_RESET_B_c_652_n 0.021059f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_36 VNB N_RESET_B_M1030_g 0.0519609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_RESET_B_c_654_n 0.0175891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_RESET_B_c_655_n 0.0319596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_c_656_n 0.00562946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_303_395#_c_877_n 0.0140494f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_41 VNB N_A_303_395#_c_878_n 0.0308361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_303_395#_c_879_n 0.0668917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_303_395#_c_880_n 0.0162572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_303_395#_c_881_n 0.0368611f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_45 VNB N_A_303_395#_c_882_n 0.0331371f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_46 VNB N_A_303_395#_M1037_g 0.0499146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_303_395#_c_884_n 0.0142811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_303_395#_c_885_n 4.56294e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_303_395#_c_886_n 0.00285158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_303_395#_c_887_n 0.00952752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_303_395#_c_888_n 0.00625184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_702_463#_c_1103_n 0.0239206f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.6
cc_53 VNB N_A_702_463#_c_1104_n 0.0175129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_702_463#_c_1105_n 0.0496729f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.165
cc_55 VNB N_A_702_463#_c_1106_n 0.00824647f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_56 VNB N_A_702_463#_c_1107_n 0.00401724f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.01
cc_57 VNB N_A_702_463#_c_1108_n 0.00102843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_702_463#_c_1109_n 0.00109066f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.665
cc_59 VNB N_A_702_463#_c_1110_n 0.0134696f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_60 VNB N_A_702_463#_c_1111_n 0.00211834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1678_395#_M1022_g 0.0226108f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_62 VNB N_A_1678_395#_c_1242_n 0.0147871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1678_395#_c_1243_n 0.0161902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1678_395#_c_1244_n 0.0100185f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.01
cc_65 VNB N_A_1678_395#_c_1245_n 0.00724983f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.295
cc_66 VNB N_A_1678_395#_c_1246_n 0.00408177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1678_395#_c_1247_n 0.0315912f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=2.035
cc_68 VNB N_A_1678_395#_c_1248_n 0.00985953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1353_392#_M1031_g 0.0443312f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1
cc_70 VNB N_A_1353_392#_c_1364_n 0.00790233f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_71 VNB N_A_1353_392#_c_1365_n 0.0119253f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_72 VNB N_A_1353_392#_c_1366_n 0.0144823f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.165
cc_73 VNB N_A_1353_392#_c_1367_n 0.0103775f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.665
cc_74 VNB N_A_1353_392#_c_1368_n 0.00465131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1353_392#_c_1369_n 0.0189463f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.845
cc_76 VNB N_A_1353_392#_c_1370_n 0.0167302f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=2.035
cc_77 VNB N_A_1353_392#_c_1371_n 0.00538628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1353_392#_c_1372_n 0.0041539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1353_392#_c_1373_n 0.00737056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1353_392#_c_1374_n 0.00664015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1353_392#_c_1375_n 0.00100027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1353_392#_c_1376_n 0.0239677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2013_409#_M1009_g 0.00170702f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1
cc_84 VNB N_A_2013_409#_c_1527_n 0.0102302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2013_409#_M1021_g 0.00249279f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_86 VNB N_A_2013_409#_M1003_g 0.0250105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2013_409#_c_1530_n 0.0263854f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_88 VNB N_A_2013_409#_c_1531_n 0.0222317f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_89 VNB N_A_2013_409#_M1023_g 0.0223949f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_90 VNB N_A_2013_409#_M1028_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2013_409#_M1032_g 0.02888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2013_409#_M1029_g 0.0017572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2013_409#_M1038_g 0.0378399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2013_409#_c_1537_n 0.00142943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2013_409#_c_1538_n 0.00371217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2013_409#_c_1539_n 0.0128657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2013_409#_c_1540_n 0.0109985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2013_409#_c_1541_n 0.0048999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2013_409#_c_1542_n 0.011911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2013_409#_c_1543_n 0.0536028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VPWR_c_1652_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_37_78#_c_1822_n 0.00234939f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.35
cc_103 VNB N_A_37_78#_c_1823_n 0.0151278f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.165
cc_104 VNB N_A_37_78#_c_1824_n 0.00218843f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_105 VNB N_A_37_78#_c_1825_n 0.00552249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_37_78#_c_1826_n 0.00175492f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_107 VNB N_A_37_78#_c_1827_n 0.00344986f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_108 VNB N_A_37_78#_c_1828_n 0.0222792f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_109 VNB N_Q_c_1943_n 0.00250883f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_110 VNB N_Q_c_1944_n 0.00280896f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1
cc_111 VNB N_Q_c_1945_n 0.00323677f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_112 VNB N_Q_c_1946_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_113 VNB N_Q_c_1947_n 0.00131414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_Q_c_1948_n 2.04518e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB Q 0.0222191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2015_n 0.00749944f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.01
cc_117 VNB N_VGND_c_2016_n 0.0125405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2017_n 0.0151521f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_119 VNB N_VGND_c_2018_n 0.0133586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2019_n 0.0179738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2020_n 0.00503034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2021_n 0.0117082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2022_n 0.0382127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2023_n 0.0309871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2024_n 0.00226387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2025_n 0.0344576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2026_n 0.00528956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2027_n 0.0203404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2028_n 0.0611822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2029_n 0.0798951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2030_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2031_n 0.0187248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2032_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2033_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2034_n 0.0136561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2035_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2036_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2037_n 0.00606636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2038_n 0.706765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VPB N_D_c_276_n 0.0132401f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.81
cc_141 VPB N_D_c_281_n 0.0172277f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.245
cc_142 VPB N_D_M1034_g 0.0293003f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_143 VPB N_D_c_283_n 0.0100802f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.35
cc_144 VPB N_D_c_279_n 0.0247385f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_145 VPB N_D_c_285_n 0.0231943f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_146 VPB CLK 0.00219035f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_147 VPB N_CLK_c_313_n 0.0124972f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.6
cc_148 VPB N_CLK_c_317_n 0.0201585f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.35
cc_149 VPB N_A_497_395#_c_359_n 0.0188377f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_150 VPB N_A_497_395#_M1014_g 0.0351244f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_151 VPB N_A_497_395#_c_360_n 0.00981759f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.6
cc_152 VPB N_A_497_395#_c_361_n 0.00689031f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.35
cc_153 VPB N_A_497_395#_M1007_g 0.0267279f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.845
cc_154 VPB N_A_497_395#_c_383_n 0.00601711f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=2.01
cc_155 VPB N_A_497_395#_c_370_n 0.00688356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_497_395#_c_373_n 0.00541034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_497_395#_c_386_n 0.041097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_834_355#_M1006_g 0.0239659f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_159 VPB N_A_834_355#_M1024_g 0.00601276f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.35
cc_160 VPB N_A_834_355#_c_558_n 0.00190944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_834_355#_c_563_n 0.0445642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_834_355#_c_559_n 0.00253652f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1
cc_163 VPB N_A_834_355#_c_565_n 0.00708598f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.035
cc_164 VPB N_RESET_B_c_648_n 0.0228693f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_165 VPB N_RESET_B_M1035_g 0.0430097f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_166 VPB N_RESET_B_M1016_g 0.0321763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_RESET_B_c_652_n 7.13987e-19 $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_168 VPB N_RESET_B_M1026_g 0.0236708f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_169 VPB N_RESET_B_M1030_g 0.0152075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_RESET_B_c_663_n 0.0106508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_RESET_B_c_664_n 0.0278436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_RESET_B_c_665_n 0.00389604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_RESET_B_c_666_n 0.0267148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_RESET_B_c_667_n 0.00376976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_RESET_B_c_668_n 0.0151376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_RESET_B_c_669_n 0.00293589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_RESET_B_c_670_n 0.00604009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_c_671_n 0.0464745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_RESET_B_c_656_n 0.00125931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_RESET_B_c_673_n 0.0286073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_RESET_B_c_674_n 0.0283585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_303_395#_c_889_n 0.0170113f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_183 VPB N_A_303_395#_c_890_n 0.0687783f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_184 VPB N_A_303_395#_c_891_n 0.0539077f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_185 VPB N_A_303_395#_c_892_n 0.00992448f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_186 VPB N_A_303_395#_c_879_n 0.0143337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_303_395#_M1019_g 0.0374349f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.845
cc_188 VPB N_A_303_395#_c_895_n 0.106212f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_189 VPB N_A_303_395#_c_896_n 0.0375897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_303_395#_c_881_n 0.00527407f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_191 VPB N_A_303_395#_M1020_g 0.0303468f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_192 VPB N_A_303_395#_c_882_n 0.0503144f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_193 VPB N_A_303_395#_c_900_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_303_395#_c_901_n 0.00410718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_303_395#_c_902_n 0.00425266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_303_395#_c_903_n 0.008639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_303_395#_c_887_n 0.00295293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_303_395#_c_905_n 0.00400792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_303_395#_c_906_n 0.0464113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_702_463#_c_1112_n 0.00658077f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_201 VPB N_A_702_463#_M1015_g 0.02266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_702_463#_c_1106_n 0.00436657f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_203 VPB N_A_702_463#_c_1107_n 0.0107882f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=2.01
cc_204 VPB N_A_702_463#_c_1108_n 0.00423545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_702_463#_c_1117_n 0.00269421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_702_463#_c_1118_n 0.00191819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_702_463#_c_1119_n 0.00334423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1678_395#_M1012_g 0.0296597f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_209 VPB N_A_1678_395#_c_1242_n 0.017829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1678_395#_c_1251_n 0.00952112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1678_395#_c_1252_n 0.0031426f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_212 VPB N_A_1678_395#_c_1253_n 0.00693697f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1
cc_213 VPB N_A_1678_395#_c_1254_n 0.00169772f $X=-0.19 $Y=1.66 $X2=0.42
+ $Y2=1.845
cc_214 VPB N_A_1678_395#_c_1245_n 0.00167634f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.295
cc_215 VPB N_A_1678_395#_c_1256_n 0.00962782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1353_392#_M1027_g 0.0505453f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.35
cc_217 VPB N_A_1353_392#_c_1364_n 0.00374484f $X=-0.19 $Y=1.66 $X2=0.155
+ $Y2=1.58
cc_218 VPB N_A_1353_392#_M1008_g 0.028763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1353_392#_c_1365_n 0.00385745f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_220 VPB N_A_1353_392#_M1025_g 0.0300483f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_221 VPB N_A_1353_392#_c_1367_n 8.59645e-19 $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.665
cc_222 VPB N_A_1353_392#_c_1368_n 0.00184123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1353_392#_c_1371_n 0.0164109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1353_392#_c_1385_n 0.00772124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1353_392#_c_1373_n 0.00974213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1353_392#_c_1374_n 2.91644e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1353_392#_c_1375_n 3.14732e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1353_392#_c_1376_n 0.00359861f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_2013_409#_M1009_g 0.0244008f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1
cc_230 VPB N_A_2013_409#_M1021_g 0.0282845f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_231 VPB N_A_2013_409#_M1028_g 0.0271366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_2013_409#_M1029_g 0.0256142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_2013_409#_c_1548_n 0.004415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1653_n 0.0104926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1654_n 0.0312148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1655_n 0.0085187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1656_n 4.20494e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1657_n 0.00927888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1658_n 0.0068774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1659_n 0.0199781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1660_n 0.00921168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1661_n 0.00705994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1662_n 0.0122424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1663_n 0.0149023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1664_n 0.0511073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1665_n 0.0667644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1666_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1667_n 0.020793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1668_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1669_n 0.0184712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1670_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1671_n 0.0181107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1672_n 0.0200512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1673_n 0.0576704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1674_n 0.0303917f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1675_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1676_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1677_n 0.00612764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1678_n 0.00436893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1679_n 0.00436844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1680_n 0.00622306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1681_n 0.0135346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1652_n 0.121277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_37_78#_c_1829_n 0.00227613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_37_78#_c_1823_n 0.0127824f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.165
cc_266 VPB N_A_37_78#_c_1831_n 0.0135562f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_267 VPB N_A_37_78#_c_1832_n 0.00392603f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=2.01
cc_268 VPB N_A_37_78#_c_1827_n 0.00498525f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_269 VPB N_A_37_78#_c_1834_n 0.00444479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_37_78#_c_1835_n 0.00708249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_Q_c_1950_n 0.00275653f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_272 VPB N_Q_c_1951_n 0.00560979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_Q_c_1952_n 0.00289401f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.165
cc_274 VPB N_Q_c_1953_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB Q 0.0122269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 N_D_M1017_g N_RESET_B_M1005_g 0.0206939f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_277 N_D_c_276_n N_RESET_B_c_648_n 0.0206939f $X=0.42 $Y=1.81 $X2=0 $Y2=0
cc_278 N_D_c_281_n N_RESET_B_M1035_g 0.0206939f $X=0.515 $Y=2.245 $X2=0 $Y2=0
cc_279 N_D_M1034_g N_RESET_B_M1035_g 0.0174986f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_280 N_D_c_278_n N_RESET_B_c_655_n 0.0206939f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_281 N_D_c_285_n N_RESET_B_c_673_n 0.0206939f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_282 N_D_M1034_g N_VPWR_c_1654_n 0.00477201f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_283 N_D_c_279_n N_VPWR_c_1654_n 0.0134569f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_284 N_D_c_285_n N_VPWR_c_1654_n 7.3436e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_285 N_D_M1034_g N_VPWR_c_1655_n 4.09929e-19 $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_286 N_D_M1034_g N_VPWR_c_1671_n 0.005209f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_287 N_D_M1034_g N_VPWR_c_1652_n 0.00986101f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_288 N_D_M1017_g N_A_37_78#_c_1822_n 0.0116103f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_289 N_D_c_279_n N_A_37_78#_c_1822_n 0.00144733f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_290 N_D_M1034_g N_A_37_78#_c_1829_n 0.00527901f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_291 N_D_M1034_g N_A_37_78#_c_1823_n 8.86329e-19 $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_292 N_D_M1017_g N_A_37_78#_c_1823_n 0.0162507f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_293 N_D_c_279_n N_A_37_78#_c_1823_n 0.0891656f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_294 N_D_M1017_g N_A_37_78#_c_1828_n 0.00807807f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_295 N_D_c_278_n N_A_37_78#_c_1828_n 0.00188146f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_296 N_D_c_279_n N_A_37_78#_c_1828_n 0.0285087f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_297 N_D_M1034_g N_A_37_78#_c_1834_n 0.00740192f $X=0.5 $Y=2.75 $X2=0 $Y2=0
cc_298 N_D_c_283_n N_A_37_78#_c_1834_n 0.00138105f $X=0.515 $Y=2.35 $X2=0 $Y2=0
cc_299 N_D_M1017_g N_VGND_c_2015_n 0.00180389f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_300 N_D_M1017_g N_VGND_c_2023_n 0.00429844f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_301 N_D_M1017_g N_VGND_c_2038_n 0.00539454f $X=0.545 $Y=0.6 $X2=0 $Y2=0
cc_302 N_CLK_c_317_n N_A_497_395#_c_383_n 8.9774e-19 $X=1.93 $Y=1.885 $X2=0
+ $Y2=0
cc_303 N_CLK_c_313_n N_RESET_B_c_648_n 0.00977857f $X=1.93 $Y=1.61 $X2=0 $Y2=0
cc_304 N_CLK_c_317_n N_RESET_B_c_648_n 0.0053618f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_305 N_CLK_c_314_n N_RESET_B_c_649_n 0.0104164f $X=1.93 $Y=1.41 $X2=0 $Y2=0
cc_306 CLK N_RESET_B_c_664_n 0.0142361f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_307 N_CLK_c_313_n N_RESET_B_c_664_n 0.00301605f $X=1.93 $Y=1.61 $X2=0 $Y2=0
cc_308 N_CLK_c_317_n N_RESET_B_c_664_n 0.00656313f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_309 N_CLK_c_314_n N_RESET_B_c_655_n 0.00323598f $X=1.93 $Y=1.41 $X2=0 $Y2=0
cc_310 N_CLK_c_317_n N_RESET_B_c_656_n 2.51239e-19 $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_311 CLK N_A_303_395#_M1001_s 4.93455e-19 $X=2.075 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_312 N_CLK_c_317_n N_A_303_395#_c_889_n 0.0471711f $X=1.93 $Y=1.885 $X2=0
+ $Y2=0
cc_313 CLK N_A_303_395#_c_877_n 7.73725e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_314 N_CLK_c_314_n N_A_303_395#_c_877_n 0.0187765f $X=1.93 $Y=1.41 $X2=0 $Y2=0
cc_315 CLK N_A_303_395#_c_879_n 0.00323328f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_316 N_CLK_c_313_n N_A_303_395#_c_879_n 0.0320746f $X=1.93 $Y=1.61 $X2=0 $Y2=0
cc_317 N_CLK_c_314_n N_A_303_395#_c_884_n 0.00312263f $X=1.93 $Y=1.41 $X2=0
+ $Y2=0
cc_318 CLK N_A_303_395#_c_914_n 0.0262776f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_319 N_CLK_c_313_n N_A_303_395#_c_914_n 2.75938e-19 $X=1.93 $Y=1.61 $X2=0
+ $Y2=0
cc_320 N_CLK_c_314_n N_A_303_395#_c_914_n 0.0129975f $X=1.93 $Y=1.41 $X2=0 $Y2=0
cc_321 CLK N_A_303_395#_c_885_n 0.0363665f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_322 N_CLK_c_313_n N_A_303_395#_c_885_n 2.65287e-19 $X=1.93 $Y=1.61 $X2=0
+ $Y2=0
cc_323 N_CLK_c_314_n N_A_303_395#_c_885_n 9.92384e-19 $X=1.93 $Y=1.41 $X2=0
+ $Y2=0
cc_324 CLK N_A_303_395#_c_886_n 0.00201688f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_325 N_CLK_c_313_n N_A_303_395#_c_886_n 0.0015915f $X=1.93 $Y=1.61 $X2=0 $Y2=0
cc_326 CLK N_A_303_395#_c_903_n 6.63104e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_327 N_CLK_c_313_n N_A_303_395#_c_903_n 0.00165188f $X=1.93 $Y=1.61 $X2=0
+ $Y2=0
cc_328 N_CLK_c_317_n N_A_303_395#_c_903_n 0.00375038f $X=1.93 $Y=1.885 $X2=0
+ $Y2=0
cc_329 CLK N_A_303_395#_c_887_n 0.0366934f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_330 N_CLK_c_313_n N_A_303_395#_c_887_n 0.00575696f $X=1.93 $Y=1.61 $X2=0
+ $Y2=0
cc_331 N_CLK_c_314_n N_A_303_395#_c_887_n 0.00253494f $X=1.93 $Y=1.41 $X2=0
+ $Y2=0
cc_332 N_CLK_c_317_n N_A_303_395#_c_887_n 2.11312e-19 $X=1.93 $Y=1.885 $X2=0
+ $Y2=0
cc_333 N_CLK_c_317_n N_VPWR_c_1655_n 0.00739434f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_334 N_CLK_c_317_n N_VPWR_c_1656_n 0.0138887f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_335 N_CLK_c_317_n N_VPWR_c_1672_n 0.00583607f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_336 N_CLK_c_317_n N_VPWR_c_1652_n 0.0066554f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_337 CLK N_A_37_78#_c_1831_n 0.00454075f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_338 N_CLK_c_313_n N_A_37_78#_c_1831_n 0.00176727f $X=1.93 $Y=1.61 $X2=0 $Y2=0
cc_339 N_CLK_c_317_n N_A_37_78#_c_1831_n 0.0171077f $X=1.93 $Y=1.885 $X2=0 $Y2=0
cc_340 CLK N_VGND_M1001_d 0.00232932f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_341 N_CLK_c_314_n N_VGND_c_2016_n 0.00119784f $X=1.93 $Y=1.41 $X2=0 $Y2=0
cc_342 N_CLK_c_314_n N_VGND_c_2038_n 9.39239e-19 $X=1.93 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_497_395#_c_369_n N_A_834_355#_M1011_d 0.0186644f $X=8.105 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_344 N_A_497_395#_c_361_n N_A_834_355#_M1024_g 0.00574617f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_345 N_A_497_395#_M1036_g N_A_834_355#_M1024_g 0.0491928f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_346 N_A_497_395#_c_368_n N_A_834_355#_M1024_g 3.87813e-19 $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_347 N_A_497_395#_c_374_n N_A_834_355#_M1024_g 0.00758607f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_348 N_A_497_395#_M1036_g N_A_834_355#_c_558_n 5.34274e-19 $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_349 N_A_497_395#_c_359_n N_A_834_355#_c_563_n 0.00121772f $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_350 N_A_497_395#_M1014_g N_A_834_355#_c_563_n 0.00389351f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_351 N_A_497_395#_c_368_n N_A_834_355#_c_574_n 0.00512559f $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_352 N_A_497_395#_c_374_n N_A_834_355#_c_574_n 0.0116732f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_353 N_A_497_395#_c_369_n N_A_834_355#_c_576_n 0.0530777f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_354 N_A_497_395#_c_368_n N_A_834_355#_c_577_n 0.050878f $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_355 N_A_497_395#_c_369_n N_A_834_355#_c_577_n 0.00379885f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_356 N_A_497_395#_c_375_n N_A_834_355#_c_577_n 0.0123656f $X=5.48 $Y=0.34
+ $X2=0 $Y2=0
cc_357 N_A_497_395#_M1036_g N_RESET_B_c_649_n 0.00526413f $X=3.985 $Y=0.9 $X2=0
+ $Y2=0
cc_358 N_A_497_395#_c_367_n N_RESET_B_c_649_n 0.0245672f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_359 N_A_497_395#_c_368_n N_RESET_B_c_649_n 0.00239679f $X=5.395 $Y=0.625
+ $X2=0 $Y2=0
cc_360 N_A_497_395#_c_372_n N_RESET_B_c_649_n 0.0110537f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_361 N_A_497_395#_c_374_n N_RESET_B_c_649_n 0.00182747f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_362 N_A_497_395#_c_368_n N_RESET_B_M1033_g 0.0127957f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_363 N_A_497_395#_c_374_n N_RESET_B_M1033_g 0.00659147f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_364 N_A_497_395#_c_375_n N_RESET_B_M1033_g 0.00440016f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_A_497_395#_c_359_n N_RESET_B_c_664_n 2.55325e-19 $X=3.42 $Y=1.89 $X2=0
+ $Y2=0
cc_366 N_A_497_395#_M1014_g N_RESET_B_c_664_n 0.00663018f $X=3.42 $Y=2.525 $X2=0
+ $Y2=0
cc_367 N_A_497_395#_c_360_n N_RESET_B_c_664_n 0.00437182f $X=3.8 $Y=1.665 $X2=0
+ $Y2=0
cc_368 N_A_497_395#_c_361_n N_RESET_B_c_664_n 2.83397e-19 $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_369 N_A_497_395#_c_383_n N_RESET_B_c_664_n 0.0223775f $X=2.845 $Y=2.082 $X2=0
+ $Y2=0
cc_370 N_A_497_395#_c_373_n N_RESET_B_c_664_n 0.0304395f $X=3.355 $Y=1.725 $X2=0
+ $Y2=0
cc_371 N_A_497_395#_c_370_n N_RESET_B_c_666_n 0.0224618f $X=7.905 $Y=2.14 $X2=0
+ $Y2=0
cc_372 N_A_497_395#_c_386_n N_RESET_B_c_666_n 0.00379291f $X=8.06 $Y=2.14 $X2=0
+ $Y2=0
cc_373 N_A_497_395#_c_383_n N_A_303_395#_c_889_n 0.00613446f $X=2.845 $Y=2.082
+ $X2=0 $Y2=0
cc_374 N_A_497_395#_c_373_n N_A_303_395#_c_889_n 3.48066e-19 $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_375 N_A_497_395#_c_366_n N_A_303_395#_c_877_n 0.00498881f $X=2.93 $Y=1.56
+ $X2=0 $Y2=0
cc_376 N_A_497_395#_c_372_n N_A_303_395#_c_877_n 0.0031356f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_377 N_A_497_395#_M1014_g N_A_303_395#_c_890_n 0.0262877f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_378 N_A_497_395#_c_383_n N_A_303_395#_c_890_n 0.00485691f $X=2.845 $Y=2.082
+ $X2=0 $Y2=0
cc_379 N_A_497_395#_c_373_n N_A_303_395#_c_890_n 0.00939366f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_380 N_A_497_395#_M1014_g N_A_303_395#_c_891_n 0.0123546f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_381 N_A_497_395#_c_359_n N_A_303_395#_c_878_n 0.0195256f $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_382 N_A_497_395#_c_360_n N_A_303_395#_c_878_n 0.00184099f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_383 N_A_497_395#_c_367_n N_A_303_395#_c_878_n 5.79793e-19 $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_384 N_A_497_395#_c_373_n N_A_303_395#_c_878_n 0.00623128f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_385 N_A_497_395#_c_359_n N_A_303_395#_c_879_n 0.0213222f $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_386 N_A_497_395#_c_383_n N_A_303_395#_c_879_n 0.00581358f $X=2.845 $Y=2.082
+ $X2=0 $Y2=0
cc_387 N_A_497_395#_c_366_n N_A_303_395#_c_879_n 0.0180555f $X=2.93 $Y=1.56
+ $X2=0 $Y2=0
cc_388 N_A_497_395#_c_367_n N_A_303_395#_c_879_n 0.00344397f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_389 N_A_497_395#_c_372_n N_A_303_395#_c_879_n 0.00526006f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_390 N_A_497_395#_c_373_n N_A_303_395#_c_879_n 0.0156744f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_391 N_A_497_395#_M1036_g N_A_303_395#_c_880_n 0.0183299f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_392 N_A_497_395#_c_367_n N_A_303_395#_c_880_n 0.00349197f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_393 N_A_497_395#_c_372_n N_A_303_395#_c_880_n 0.00450148f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_394 N_A_497_395#_M1014_g N_A_303_395#_M1019_g 0.0170083f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_395 N_A_497_395#_c_360_n N_A_303_395#_M1019_g 0.0052298f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_396 N_A_497_395#_c_365_n N_A_303_395#_c_881_n 0.00558264f $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_397 N_A_497_395#_c_365_n N_A_303_395#_c_882_n 0.0477631f $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_398 N_A_497_395#_c_370_n N_A_303_395#_c_882_n 0.0163868f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_399 N_A_497_395#_c_377_n N_A_303_395#_c_882_n 0.0018416f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_400 N_A_497_395#_c_386_n N_A_303_395#_c_882_n 0.023403f $X=8.06 $Y=2.14 $X2=0
+ $Y2=0
cc_401 N_A_497_395#_c_369_n N_A_303_395#_M1037_g 0.0088085f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_402 N_A_497_395#_c_370_n N_A_303_395#_M1037_g 0.00916962f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_403 N_A_497_395#_c_371_n N_A_303_395#_M1037_g 0.0233298f $X=8.19 $Y=1.015
+ $X2=0 $Y2=0
cc_404 N_A_497_395#_c_376_n N_A_303_395#_M1037_g 0.0213806f $X=7.71 $Y=1.18
+ $X2=0 $Y2=0
cc_405 N_A_497_395#_c_377_n N_A_303_395#_M1037_g 0.0144366f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_406 N_A_497_395#_M1002_d N_A_303_395#_c_914_n 0.00263826f $X=2.545 $Y=0.595
+ $X2=0 $Y2=0
cc_407 N_A_497_395#_c_366_n N_A_303_395#_c_914_n 0.0136886f $X=2.93 $Y=1.56
+ $X2=0 $Y2=0
cc_408 N_A_497_395#_c_372_n N_A_303_395#_c_914_n 0.00641127f $X=2.78 $Y=0.415
+ $X2=0 $Y2=0
cc_409 N_A_497_395#_M1002_d N_A_303_395#_c_885_n 0.0017515f $X=2.545 $Y=0.595
+ $X2=0 $Y2=0
cc_410 N_A_497_395#_c_383_n N_A_303_395#_c_885_n 0.016387f $X=2.845 $Y=2.082
+ $X2=0 $Y2=0
cc_411 N_A_497_395#_c_366_n N_A_303_395#_c_885_n 0.0308188f $X=2.93 $Y=1.56
+ $X2=0 $Y2=0
cc_412 N_A_497_395#_c_373_n N_A_303_395#_c_885_n 0.0166149f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_413 N_A_497_395#_c_383_n N_A_303_395#_c_903_n 0.00329212f $X=2.845 $Y=2.082
+ $X2=0 $Y2=0
cc_414 N_A_497_395#_c_365_n N_A_303_395#_c_888_n 7.01297e-19 $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_415 N_A_497_395#_c_369_n N_A_702_463#_c_1103_n 0.013057f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_416 N_A_497_395#_c_375_n N_A_702_463#_c_1103_n 0.00165256f $X=5.48 $Y=0.34
+ $X2=0 $Y2=0
cc_417 N_A_497_395#_M1014_g N_A_702_463#_c_1107_n 4.20006e-19 $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_418 N_A_497_395#_c_361_n N_A_702_463#_c_1107_n 0.00787964f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_419 N_A_497_395#_M1036_g N_A_702_463#_c_1107_n 0.00772225f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_420 N_A_497_395#_c_360_n N_A_702_463#_c_1111_n 7.41936e-19 $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_421 N_A_497_395#_c_361_n N_A_702_463#_c_1111_n 0.00282934f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_422 N_A_497_395#_M1036_g N_A_702_463#_c_1111_n 0.0116997f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_423 N_A_497_395#_c_367_n N_A_702_463#_c_1111_n 0.0325837f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_424 N_A_497_395#_c_374_n N_A_702_463#_c_1111_n 0.00153321f $X=4.39 $Y=0.415
+ $X2=0 $Y2=0
cc_425 N_A_497_395#_M1014_g N_A_702_463#_c_1117_n 7.94952e-19 $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_426 N_A_497_395#_M1007_g N_A_1678_395#_M1012_g 0.0281156f $X=8.06 $Y=2.675
+ $X2=0 $Y2=0
cc_427 N_A_497_395#_c_369_n N_A_1678_395#_M1022_g 0.00112332f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_428 N_A_497_395#_c_371_n N_A_1678_395#_M1022_g 0.00454635f $X=8.19 $Y=1.015
+ $X2=0 $Y2=0
cc_429 N_A_497_395#_c_377_n N_A_1678_395#_M1022_g 4.94468e-19 $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_430 N_A_497_395#_c_370_n N_A_1678_395#_c_1251_n 3.41992e-19 $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_431 N_A_497_395#_c_386_n N_A_1678_395#_c_1251_n 0.0281156f $X=8.06 $Y=2.14
+ $X2=0 $Y2=0
cc_432 N_A_497_395#_c_370_n N_A_1678_395#_c_1246_n 8.76782e-19 $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_433 N_A_497_395#_c_377_n N_A_1678_395#_c_1246_n 0.026059f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_434 N_A_497_395#_c_377_n N_A_1678_395#_c_1247_n 0.00189496f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_435 N_A_497_395#_c_369_n N_A_1353_392#_M1004_d 0.00949814f $X=8.105 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_436 N_A_497_395#_c_363_n N_A_1353_392#_c_1391_n 0.00759713f $X=7.11 $Y=1.195
+ $X2=0 $Y2=0
cc_437 N_A_497_395#_c_369_n N_A_1353_392#_c_1391_n 0.00844204f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_438 N_A_497_395#_c_363_n N_A_1353_392#_c_1371_n 0.0120402f $X=7.11 $Y=1.195
+ $X2=0 $Y2=0
cc_439 N_A_497_395#_c_364_n N_A_1353_392#_c_1371_n 0.00910494f $X=7.545 $Y=1.27
+ $X2=0 $Y2=0
cc_440 N_A_497_395#_c_365_n N_A_1353_392#_c_1371_n 0.00382426f $X=7.185 $Y=1.27
+ $X2=0 $Y2=0
cc_441 N_A_497_395#_M1007_g N_A_1353_392#_c_1371_n 0.00352564f $X=8.06 $Y=2.675
+ $X2=0 $Y2=0
cc_442 N_A_497_395#_c_370_n N_A_1353_392#_c_1371_n 0.036911f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_443 N_A_497_395#_c_376_n N_A_1353_392#_c_1371_n 6.23735e-19 $X=7.71 $Y=1.18
+ $X2=0 $Y2=0
cc_444 N_A_497_395#_c_377_n N_A_1353_392#_c_1371_n 0.0212415f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_445 N_A_497_395#_c_386_n N_A_1353_392#_c_1371_n 0.00548394f $X=8.06 $Y=2.14
+ $X2=0 $Y2=0
cc_446 N_A_497_395#_c_364_n N_A_1353_392#_c_1372_n 0.00633476f $X=7.545 $Y=1.27
+ $X2=0 $Y2=0
cc_447 N_A_497_395#_c_369_n N_A_1353_392#_c_1372_n 0.0424696f $X=8.105 $Y=0.34
+ $X2=0 $Y2=0
cc_448 N_A_497_395#_c_371_n N_A_1353_392#_c_1372_n 0.0196081f $X=8.19 $Y=1.015
+ $X2=0 $Y2=0
cc_449 N_A_497_395#_c_376_n N_A_1353_392#_c_1372_n 0.00746605f $X=7.71 $Y=1.18
+ $X2=0 $Y2=0
cc_450 N_A_497_395#_c_377_n N_A_1353_392#_c_1372_n 0.030444f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_451 N_A_497_395#_M1007_g N_A_1353_392#_c_1406_n 0.0147394f $X=8.06 $Y=2.675
+ $X2=0 $Y2=0
cc_452 N_A_497_395#_c_370_n N_A_1353_392#_c_1406_n 0.0232787f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_453 N_A_497_395#_c_386_n N_A_1353_392#_c_1406_n 0.00155184f $X=8.06 $Y=2.14
+ $X2=0 $Y2=0
cc_454 N_A_497_395#_c_370_n N_A_1353_392#_c_1385_n 0.045021f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_455 N_A_497_395#_c_386_n N_A_1353_392#_c_1385_n 0.00587378f $X=8.06 $Y=2.14
+ $X2=0 $Y2=0
cc_456 N_A_497_395#_c_370_n N_A_1353_392#_c_1374_n 0.0145381f $X=7.905 $Y=2.14
+ $X2=0 $Y2=0
cc_457 N_A_497_395#_c_377_n N_A_1353_392#_c_1374_n 0.00286183f $X=8.19 $Y=1.18
+ $X2=0 $Y2=0
cc_458 N_A_497_395#_M1007_g N_VPWR_c_1665_n 0.00469675f $X=8.06 $Y=2.675 $X2=0
+ $Y2=0
cc_459 N_A_497_395#_M1013_d N_VPWR_c_1652_n 0.00367888f $X=2.485 $Y=1.975 $X2=0
+ $Y2=0
cc_460 N_A_497_395#_M1014_g N_VPWR_c_1652_n 0.00112709f $X=3.42 $Y=2.525 $X2=0
+ $Y2=0
cc_461 N_A_497_395#_M1007_g N_VPWR_c_1652_n 0.00626544f $X=8.06 $Y=2.675 $X2=0
+ $Y2=0
cc_462 N_A_497_395#_M1013_d N_A_37_78#_c_1831_n 0.00597109f $X=2.485 $Y=1.975
+ $X2=0 $Y2=0
cc_463 N_A_497_395#_c_383_n N_A_37_78#_c_1831_n 0.0232729f $X=2.845 $Y=2.082
+ $X2=0 $Y2=0
cc_464 N_A_497_395#_c_373_n N_A_37_78#_c_1831_n 0.0129779f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_465 N_A_497_395#_M1036_g N_A_37_78#_c_1824_n 5.96704e-19 $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_466 N_A_497_395#_c_367_n N_A_37_78#_c_1824_n 0.0198808f $X=4.305 $Y=0.415
+ $X2=0 $Y2=0
cc_467 N_A_497_395#_c_372_n N_A_37_78#_c_1824_n 0.042559f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_468 N_A_497_395#_c_359_n N_A_37_78#_c_1832_n 3.579e-19 $X=3.42 $Y=1.89 $X2=0
+ $Y2=0
cc_469 N_A_497_395#_M1014_g N_A_37_78#_c_1832_n 0.0129286f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_470 N_A_497_395#_c_360_n N_A_37_78#_c_1832_n 0.00289451f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_471 N_A_497_395#_c_373_n N_A_37_78#_c_1832_n 0.00532454f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_472 N_A_497_395#_c_359_n N_A_37_78#_c_1825_n 0.00143239f $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_473 N_A_497_395#_c_360_n N_A_37_78#_c_1825_n 0.00292226f $X=3.8 $Y=1.665
+ $X2=0 $Y2=0
cc_474 N_A_497_395#_M1036_g N_A_37_78#_c_1825_n 0.00194262f $X=3.985 $Y=0.9
+ $X2=0 $Y2=0
cc_475 N_A_497_395#_c_373_n N_A_37_78#_c_1825_n 0.00144971f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_476 N_A_497_395#_c_359_n N_A_37_78#_c_1826_n 9.32078e-19 $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_477 N_A_497_395#_c_366_n N_A_37_78#_c_1826_n 0.0130768f $X=2.93 $Y=1.56 $X2=0
+ $Y2=0
cc_478 N_A_497_395#_c_373_n N_A_37_78#_c_1826_n 0.0209626f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_479 N_A_497_395#_c_359_n N_A_37_78#_c_1827_n 0.00239275f $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_480 N_A_497_395#_M1014_g N_A_37_78#_c_1827_n 0.00263548f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_481 N_A_497_395#_c_360_n N_A_37_78#_c_1827_n 0.0129748f $X=3.8 $Y=1.665 $X2=0
+ $Y2=0
cc_482 N_A_497_395#_c_361_n N_A_37_78#_c_1827_n 0.00458963f $X=3.985 $Y=1.385
+ $X2=0 $Y2=0
cc_483 N_A_497_395#_c_366_n N_A_37_78#_c_1827_n 0.00496978f $X=2.93 $Y=1.56
+ $X2=0 $Y2=0
cc_484 N_A_497_395#_c_373_n N_A_37_78#_c_1827_n 0.0325128f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_485 N_A_497_395#_c_359_n N_A_37_78#_c_1835_n 8.44622e-19 $X=3.42 $Y=1.89
+ $X2=0 $Y2=0
cc_486 N_A_497_395#_M1014_g N_A_37_78#_c_1835_n 0.0103984f $X=3.42 $Y=2.525
+ $X2=0 $Y2=0
cc_487 N_A_497_395#_c_373_n N_A_37_78#_c_1835_n 0.0254745f $X=3.355 $Y=1.725
+ $X2=0 $Y2=0
cc_488 N_A_497_395#_c_368_n N_VGND_M1033_d 0.0148411f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_489 N_A_497_395#_c_375_n N_VGND_M1033_d 0.00624194f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_490 N_A_497_395#_c_372_n N_VGND_c_2016_n 0.0315755f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_491 N_A_497_395#_c_369_n N_VGND_c_2017_n 0.00808546f $X=8.105 $Y=0.34 $X2=0
+ $Y2=0
cc_492 N_A_497_395#_c_371_n N_VGND_c_2017_n 0.0105982f $X=8.19 $Y=1.015 $X2=0
+ $Y2=0
cc_493 N_A_497_395#_c_367_n N_VGND_c_2028_n 0.0564819f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_494 N_A_497_395#_c_368_n N_VGND_c_2028_n 0.0091991f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_495 N_A_497_395#_c_372_n N_VGND_c_2028_n 0.0223109f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_496 N_A_497_395#_c_374_n N_VGND_c_2028_n 0.007809f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_497 N_A_497_395#_c_363_n N_VGND_c_2029_n 0.00278271f $X=7.11 $Y=1.195 $X2=0
+ $Y2=0
cc_498 N_A_497_395#_c_368_n N_VGND_c_2029_n 0.00371184f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_499 N_A_497_395#_c_369_n N_VGND_c_2029_n 0.174907f $X=8.105 $Y=0.34 $X2=0
+ $Y2=0
cc_500 N_A_497_395#_c_375_n N_VGND_c_2029_n 0.0116868f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_501 N_A_497_395#_c_368_n N_VGND_c_2034_n 0.0242401f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_502 N_A_497_395#_c_374_n N_VGND_c_2034_n 0.00168902f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_503 N_A_497_395#_c_375_n N_VGND_c_2034_n 0.00911749f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_504 N_A_497_395#_c_363_n N_VGND_c_2038_n 0.00363426f $X=7.11 $Y=1.195 $X2=0
+ $Y2=0
cc_505 N_A_497_395#_c_367_n N_VGND_c_2038_n 0.0410726f $X=4.305 $Y=0.415 $X2=0
+ $Y2=0
cc_506 N_A_497_395#_c_368_n N_VGND_c_2038_n 0.0183804f $X=5.395 $Y=0.625 $X2=0
+ $Y2=0
cc_507 N_A_497_395#_c_369_n N_VGND_c_2038_n 0.100739f $X=8.105 $Y=0.34 $X2=0
+ $Y2=0
cc_508 N_A_497_395#_c_372_n N_VGND_c_2038_n 0.0154876f $X=2.78 $Y=0.415 $X2=0
+ $Y2=0
cc_509 N_A_497_395#_c_374_n N_VGND_c_2038_n 0.0054919f $X=4.39 $Y=0.415 $X2=0
+ $Y2=0
cc_510 N_A_497_395#_c_375_n N_VGND_c_2038_n 0.00646475f $X=5.48 $Y=0.34 $X2=0
+ $Y2=0
cc_511 N_A_497_395#_c_368_n A_890_138# 0.00133041f $X=5.395 $Y=0.625 $X2=-0.19
+ $Y2=-0.245
cc_512 N_A_834_355#_M1024_g N_RESET_B_c_649_n 0.00540258f $X=4.375 $Y=0.9 $X2=0
+ $Y2=0
cc_513 N_A_834_355#_M1024_g N_RESET_B_M1033_g 0.0417267f $X=4.375 $Y=0.9 $X2=0
+ $Y2=0
cc_514 N_A_834_355#_c_558_n N_RESET_B_M1033_g 0.00472366f $X=4.405 $Y=1.94 $X2=0
+ $Y2=0
cc_515 N_A_834_355#_c_577_n N_RESET_B_M1033_g 0.0136619f $X=5.735 $Y=0.885 $X2=0
+ $Y2=0
cc_516 N_A_834_355#_M1006_g N_RESET_B_M1016_g 0.0178212f $X=4.26 $Y=2.525 $X2=0
+ $Y2=0
cc_517 N_A_834_355#_M1024_g N_RESET_B_c_652_n 0.0107658f $X=4.375 $Y=0.9 $X2=0
+ $Y2=0
cc_518 N_A_834_355#_c_558_n N_RESET_B_c_652_n 0.00104148f $X=4.405 $Y=1.94 $X2=0
+ $Y2=0
cc_519 N_A_834_355#_c_577_n N_RESET_B_c_654_n 0.00316016f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_520 N_A_834_355#_M1024_g N_RESET_B_c_663_n 0.00382675f $X=4.375 $Y=0.9 $X2=0
+ $Y2=0
cc_521 N_A_834_355#_c_558_n N_RESET_B_c_663_n 8.0459e-19 $X=4.405 $Y=1.94 $X2=0
+ $Y2=0
cc_522 N_A_834_355#_c_563_n N_RESET_B_c_663_n 0.0215869f $X=4.405 $Y=1.94 $X2=0
+ $Y2=0
cc_523 N_A_834_355#_c_558_n N_RESET_B_c_664_n 0.0222661f $X=4.405 $Y=1.94 $X2=0
+ $Y2=0
cc_524 N_A_834_355#_c_563_n N_RESET_B_c_664_n 0.00911976f $X=4.405 $Y=1.94 $X2=0
+ $Y2=0
cc_525 N_A_834_355#_c_559_n N_RESET_B_c_666_n 0.00270434f $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_526 N_A_834_355#_c_565_n N_RESET_B_c_666_n 0.0278833f $X=6.45 $Y=2.125 $X2=0
+ $Y2=0
cc_527 N_A_834_355#_c_559_n N_RESET_B_c_667_n 4.50751e-19 $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_528 N_A_834_355#_c_565_n N_RESET_B_c_667_n 0.0020002f $X=6.45 $Y=2.125 $X2=0
+ $Y2=0
cc_529 N_A_834_355#_c_559_n N_RESET_B_c_668_n 0.00890742f $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_530 N_A_834_355#_c_565_n N_RESET_B_c_668_n 0.00333678f $X=6.45 $Y=2.125 $X2=0
+ $Y2=0
cc_531 N_A_834_355#_M1006_g N_A_303_395#_M1019_g 0.0411652f $X=4.26 $Y=2.525
+ $X2=0 $Y2=0
cc_532 N_A_834_355#_M1006_g N_A_303_395#_c_895_n 0.0118309f $X=4.26 $Y=2.525
+ $X2=0 $Y2=0
cc_533 N_A_834_355#_c_559_n N_A_303_395#_c_881_n 0.00372027f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_534 N_A_834_355#_c_602_p N_A_303_395#_c_881_n 0.00811989f $X=6.825 $Y=0.885
+ $X2=0 $Y2=0
cc_535 N_A_834_355#_c_565_n N_A_303_395#_c_881_n 0.00181011f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_536 N_A_834_355#_c_565_n N_A_303_395#_M1020_g 0.00418835f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_537 N_A_834_355#_c_602_p N_A_303_395#_c_882_n 8.72478e-19 $X=6.825 $Y=0.885
+ $X2=0 $Y2=0
cc_538 N_A_834_355#_M1015_d N_A_303_395#_c_901_n 0.00464376f $X=6.315 $Y=1.96
+ $X2=0 $Y2=0
cc_539 N_A_834_355#_c_565_n N_A_303_395#_c_901_n 0.0234932f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_540 N_A_834_355#_c_559_n N_A_303_395#_c_902_n 0.012635f $X=6.24 $Y=1.94 $X2=0
+ $Y2=0
cc_541 N_A_834_355#_c_565_n N_A_303_395#_c_902_n 0.0138472f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_542 N_A_834_355#_c_559_n N_A_303_395#_c_888_n 0.0254145f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_543 N_A_834_355#_c_602_p N_A_303_395#_c_888_n 0.0309014f $X=6.825 $Y=0.885
+ $X2=0 $Y2=0
cc_544 N_A_834_355#_c_565_n N_A_303_395#_c_888_n 0.00452315f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_545 N_A_834_355#_c_559_n N_A_702_463#_c_1103_n 0.00417334f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_546 N_A_834_355#_c_576_n N_A_702_463#_c_1103_n 0.00865527f $X=6.325 $Y=0.885
+ $X2=0 $Y2=0
cc_547 N_A_834_355#_c_577_n N_A_702_463#_c_1103_n 0.010622f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_548 N_A_834_355#_c_559_n N_A_702_463#_c_1112_n 0.00359669f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_549 N_A_834_355#_c_559_n N_A_702_463#_M1015_g 0.00429581f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_550 N_A_834_355#_c_565_n N_A_702_463#_M1015_g 0.0124484f $X=6.45 $Y=2.125
+ $X2=0 $Y2=0
cc_551 N_A_834_355#_c_559_n N_A_702_463#_c_1105_n 0.0135266f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_552 N_A_834_355#_c_576_n N_A_702_463#_c_1105_n 0.0125532f $X=6.325 $Y=0.885
+ $X2=0 $Y2=0
cc_553 N_A_834_355#_c_559_n N_A_702_463#_c_1106_n 0.00813214f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_554 N_A_834_355#_M1024_g N_A_702_463#_c_1107_n 0.00444711f $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_555 N_A_834_355#_c_558_n N_A_702_463#_c_1107_n 0.0769404f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_556 N_A_834_355#_c_563_n N_A_702_463#_c_1107_n 0.00746781f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_557 N_A_834_355#_M1006_g N_A_702_463#_c_1143_n 0.00907016f $X=4.26 $Y=2.525
+ $X2=0 $Y2=0
cc_558 N_A_834_355#_c_558_n N_A_702_463#_c_1143_n 0.00794189f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_559 N_A_834_355#_c_563_n N_A_702_463#_c_1143_n 0.00120561f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_560 N_A_834_355#_M1006_g N_A_702_463#_c_1108_n 0.00147703f $X=4.26 $Y=2.525
+ $X2=0 $Y2=0
cc_561 N_A_834_355#_M1024_g N_A_702_463#_c_1108_n 6.92887e-19 $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_562 N_A_834_355#_c_558_n N_A_702_463#_c_1108_n 0.0439058f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_563 N_A_834_355#_c_563_n N_A_702_463#_c_1108_n 0.00159342f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_564 N_A_834_355#_M1024_g N_A_702_463#_c_1109_n 6.42461e-19 $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_565 N_A_834_355#_c_558_n N_A_702_463#_c_1109_n 0.0233608f $X=4.405 $Y=1.94
+ $X2=0 $Y2=0
cc_566 N_A_834_355#_c_577_n N_A_702_463#_c_1109_n 0.0110525f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_567 N_A_834_355#_c_559_n N_A_702_463#_c_1110_n 0.0211767f $X=6.24 $Y=1.94
+ $X2=0 $Y2=0
cc_568 N_A_834_355#_c_577_n N_A_702_463#_c_1110_n 0.0767028f $X=5.735 $Y=0.885
+ $X2=0 $Y2=0
cc_569 N_A_834_355#_M1024_g N_A_702_463#_c_1111_n 0.00193581f $X=4.375 $Y=0.9
+ $X2=0 $Y2=0
cc_570 N_A_834_355#_c_574_n N_A_702_463#_c_1111_n 0.0145807f $X=4.57 $Y=0.965
+ $X2=0 $Y2=0
cc_571 N_A_834_355#_M1006_g N_A_702_463#_c_1118_n 0.010875f $X=4.26 $Y=2.525
+ $X2=0 $Y2=0
cc_572 N_A_834_355#_M1006_g N_A_702_463#_c_1119_n 0.0012415f $X=4.26 $Y=2.525
+ $X2=0 $Y2=0
cc_573 N_A_834_355#_M1006_g N_VPWR_c_1657_n 0.00300462f $X=4.26 $Y=2.525 $X2=0
+ $Y2=0
cc_574 N_A_834_355#_M1006_g N_VPWR_c_1652_n 0.00112709f $X=4.26 $Y=2.525 $X2=0
+ $Y2=0
cc_575 N_A_834_355#_c_577_n N_VGND_M1033_d 0.017178f $X=5.735 $Y=0.885 $X2=0
+ $Y2=0
cc_576 N_A_834_355#_c_558_n A_890_138# 7.01113e-19 $X=4.405 $Y=1.94 $X2=-0.19
+ $Y2=-0.245
cc_577 N_A_834_355#_c_574_n A_890_138# 6.42914e-19 $X=4.57 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_578 N_A_834_355#_c_577_n A_890_138# 0.00300161f $X=5.735 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_579 N_RESET_B_c_664_n N_A_303_395#_M1010_s 4.43317e-19 $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_664_n N_A_303_395#_c_889_n 0.00825897f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_649_n N_A_303_395#_c_877_n 0.0104164f $X=4.69 $Y=0.18 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_649_n N_A_303_395#_c_880_n 0.00526413f $X=4.69 $Y=0.18 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_664_n N_A_303_395#_M1019_g 0.00280858f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_RESET_B_M1016_g N_A_303_395#_c_895_n 0.0118683f $X=4.87 $Y=2.525 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_666_n N_A_303_395#_c_881_n 0.0164749f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_666_n N_A_303_395#_M1020_g 0.00554859f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_587 N_RESET_B_M1005_g N_A_303_395#_c_884_n 0.00344772f $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_649_n N_A_303_395#_c_884_n 0.00989069f $X=4.69 $Y=0.18 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_664_n N_A_303_395#_c_885_n 0.00201936f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_RESET_B_c_666_n N_A_303_395#_c_901_n 0.0252115f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_591 N_RESET_B_c_666_n N_A_303_395#_c_902_n 0.0163819f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_592 N_RESET_B_M1005_g N_A_303_395#_c_886_n 0.00128044f $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_656_n N_A_303_395#_c_886_n 8.29766e-19 $X=1.155 $Y=1.295
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_648_n N_A_303_395#_c_903_n 0.0047307f $X=1.09 $Y=1.91 $X2=0
+ $Y2=0
cc_595 N_RESET_B_M1035_g N_A_303_395#_c_903_n 0.00147539f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_664_n N_A_303_395#_c_903_n 0.0305196f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_665_n N_A_303_395#_c_903_n 0.00147353f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_RESET_B_c_665_n N_A_303_395#_c_887_n 0.00140842f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_599 N_RESET_B_c_655_n N_A_303_395#_c_887_n 0.0047307f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_600 N_RESET_B_c_656_n N_A_303_395#_c_887_n 0.0730334f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_601 N_RESET_B_c_666_n N_A_303_395#_c_905_n 0.00253684f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_667_n N_A_303_395#_c_905_n 0.00819203f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_668_n N_A_303_395#_c_905_n 0.0158138f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_604 N_RESET_B_M1016_g N_A_303_395#_c_906_n 0.015006f $X=4.87 $Y=2.525 $X2=0
+ $Y2=0
cc_605 N_RESET_B_c_666_n N_A_303_395#_c_906_n 0.00100516f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_606 N_RESET_B_c_667_n N_A_303_395#_c_906_n 0.00764771f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_RESET_B_c_668_n N_A_303_395#_c_906_n 0.00798692f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_608 N_RESET_B_c_671_n N_A_303_395#_c_906_n 0.00688662f $X=5.25 $Y=1.835 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_666_n N_A_303_395#_c_888_n 0.00684899f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_RESET_B_c_654_n N_A_702_463#_c_1103_n 0.00129161f $X=4.885 $Y=1.26
+ $X2=0 $Y2=0
cc_611 N_RESET_B_c_666_n N_A_702_463#_M1015_g 0.00314953f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_612 N_RESET_B_c_667_n N_A_702_463#_M1015_g 0.00156943f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_652_n N_A_702_463#_c_1104_n 0.00381437f $X=4.885 $Y=1.67
+ $X2=0 $Y2=0
cc_614 N_RESET_B_c_666_n N_A_702_463#_c_1104_n 0.0095029f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_RESET_B_c_668_n N_A_702_463#_c_1106_n 0.00388048f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_616 N_RESET_B_c_671_n N_A_702_463#_c_1106_n 0.00334448f $X=5.25 $Y=1.835
+ $X2=0 $Y2=0
cc_617 N_RESET_B_c_664_n N_A_702_463#_c_1107_n 0.0143029f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_618 N_RESET_B_c_664_n N_A_702_463#_c_1143_n 0.0088891f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_619 N_RESET_B_M1016_g N_A_702_463#_c_1108_n 0.00948975f $X=4.87 $Y=2.525
+ $X2=0 $Y2=0
cc_620 N_RESET_B_c_652_n N_A_702_463#_c_1108_n 0.0090051f $X=4.885 $Y=1.67 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_663_n N_A_702_463#_c_1108_n 0.00990343f $X=4.87 $Y=1.835
+ $X2=0 $Y2=0
cc_622 N_RESET_B_c_664_n N_A_702_463#_c_1108_n 0.0210119f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_623 N_RESET_B_c_667_n N_A_702_463#_c_1108_n 0.00125371f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_624 N_RESET_B_c_668_n N_A_702_463#_c_1108_n 0.0325452f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_652_n N_A_702_463#_c_1109_n 0.00273309f $X=4.885 $Y=1.67
+ $X2=0 $Y2=0
cc_626 N_RESET_B_c_654_n N_A_702_463#_c_1109_n 0.0056443f $X=4.885 $Y=1.26 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_652_n N_A_702_463#_c_1110_n 0.00501004f $X=4.885 $Y=1.67
+ $X2=0 $Y2=0
cc_628 N_RESET_B_c_654_n N_A_702_463#_c_1110_n 0.00303885f $X=4.885 $Y=1.26
+ $X2=0 $Y2=0
cc_629 N_RESET_B_c_664_n N_A_702_463#_c_1110_n 0.0065884f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_630 N_RESET_B_c_666_n N_A_702_463#_c_1110_n 0.0103027f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_631 N_RESET_B_c_667_n N_A_702_463#_c_1110_n 0.0023311f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_632 N_RESET_B_c_668_n N_A_702_463#_c_1110_n 0.0429796f $X=5.52 $Y=2.035 $X2=0
+ $Y2=0
cc_633 N_RESET_B_c_671_n N_A_702_463#_c_1110_n 0.0124264f $X=5.25 $Y=1.835 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_664_n N_A_702_463#_c_1117_n 0.00725122f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_635 N_RESET_B_M1016_g N_A_702_463#_c_1118_n 7.97141e-19 $X=4.87 $Y=2.525
+ $X2=0 $Y2=0
cc_636 N_RESET_B_c_664_n N_A_702_463#_c_1118_n 0.00673934f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_637 N_RESET_B_M1016_g N_A_702_463#_c_1119_n 0.0169316f $X=4.87 $Y=2.525 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_664_n N_A_702_463#_c_1119_n 0.00883222f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_639 N_RESET_B_c_668_n N_A_702_463#_c_1119_n 0.00739632f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_640 N_RESET_B_c_671_n N_A_702_463#_c_1119_n 0.00440403f $X=5.25 $Y=1.835
+ $X2=0 $Y2=0
cc_641 N_RESET_B_M1026_g N_A_1678_395#_M1012_g 0.0106369f $X=9.02 $Y=2.675 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_669_n N_A_1678_395#_M1012_g 3.76177e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_643 N_RESET_B_c_670_n N_A_1678_395#_M1012_g 0.0011165f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_674_n N_A_1678_395#_M1012_g 0.00759212f $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_645 N_RESET_B_M1030_g N_A_1678_395#_M1022_g 0.0119923f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_646 N_RESET_B_M1030_g N_A_1678_395#_c_1242_n 0.0189876f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_647 N_RESET_B_c_666_n N_A_1678_395#_c_1242_n 0.00170338f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_648 N_RESET_B_c_669_n N_A_1678_395#_c_1242_n 7.09824e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_649 N_RESET_B_c_670_n N_A_1678_395#_c_1242_n 0.00127122f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_650 N_RESET_B_c_674_n N_A_1678_395#_c_1242_n 0.0114583f $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_651 N_RESET_B_c_666_n N_A_1678_395#_c_1251_n 0.00856922f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_652 N_RESET_B_c_669_n N_A_1678_395#_c_1251_n 3.05552e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_653 N_RESET_B_M1030_g N_A_1678_395#_c_1243_n 0.0151687f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_654 N_RESET_B_M1026_g N_A_1678_395#_c_1252_n 0.00339122f $X=9.02 $Y=2.675
+ $X2=0 $Y2=0
cc_655 N_RESET_B_c_669_n N_A_1678_395#_c_1252_n 5.78327e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_656 N_RESET_B_c_670_n N_A_1678_395#_c_1252_n 0.016871f $X=8.88 $Y=2.035 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_674_n N_A_1678_395#_c_1252_n 6.89219e-19 $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_658 N_RESET_B_M1030_g N_A_1678_395#_c_1254_n 0.00130041f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_659 N_RESET_B_c_669_n N_A_1678_395#_c_1254_n 7.6951e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_660 N_RESET_B_c_670_n N_A_1678_395#_c_1254_n 0.0098343f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_661 N_RESET_B_c_674_n N_A_1678_395#_c_1254_n 3.78573e-19 $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_662 N_RESET_B_M1030_g N_A_1678_395#_c_1244_n 0.00227582f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_663 N_RESET_B_M1030_g N_A_1678_395#_c_1246_n 0.00118187f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_664 N_RESET_B_M1030_g N_A_1678_395#_c_1247_n 0.021263f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_665 N_RESET_B_M1026_g N_A_1678_395#_c_1256_n 0.00676827f $X=9.02 $Y=2.675
+ $X2=0 $Y2=0
cc_666 N_RESET_B_c_670_n N_A_1678_395#_c_1256_n 0.00477377f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_667 N_RESET_B_c_674_n N_A_1678_395#_c_1256_n 7.88034e-19 $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_668 N_RESET_B_c_666_n N_A_1353_392#_M1020_d 0.00366961f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_669 N_RESET_B_M1030_g N_A_1353_392#_M1031_g 0.0569104f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_670 N_RESET_B_M1026_g N_A_1353_392#_M1027_g 0.01567f $X=9.02 $Y=2.675 $X2=0
+ $Y2=0
cc_671 N_RESET_B_M1030_g N_A_1353_392#_M1027_g 0.0128751f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_670_n N_A_1353_392#_M1027_g 4.39619e-19 $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_673 N_RESET_B_c_674_n N_A_1353_392#_M1027_g 0.0180965f $X=8.975 $Y=2.11 $X2=0
+ $Y2=0
cc_674 N_RESET_B_c_666_n N_A_1353_392#_c_1371_n 0.0218301f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_675 N_RESET_B_c_666_n N_A_1353_392#_c_1406_n 0.0242722f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_676 N_RESET_B_M1026_g N_A_1353_392#_c_1385_n 7.7939e-19 $X=9.02 $Y=2.675
+ $X2=0 $Y2=0
cc_677 N_RESET_B_c_666_n N_A_1353_392#_c_1385_n 0.023506f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_678 N_RESET_B_c_669_n N_A_1353_392#_c_1385_n 0.00234791f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_679 N_RESET_B_c_670_n N_A_1353_392#_c_1385_n 0.0125499f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_680 N_RESET_B_c_674_n N_A_1353_392#_c_1385_n 3.65035e-19 $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_681 N_RESET_B_M1030_g N_A_1353_392#_c_1373_n 0.0116508f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_682 N_RESET_B_c_666_n N_A_1353_392#_c_1373_n 0.0123609f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_683 N_RESET_B_c_669_n N_A_1353_392#_c_1373_n 0.00816472f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_684 N_RESET_B_c_670_n N_A_1353_392#_c_1373_n 0.0203289f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_685 N_RESET_B_c_674_n N_A_1353_392#_c_1373_n 0.00113257f $X=8.975 $Y=2.11
+ $X2=0 $Y2=0
cc_686 N_RESET_B_M1030_g N_A_1353_392#_c_1375_n 0.00118604f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_687 N_RESET_B_M1030_g N_A_1353_392#_c_1376_n 0.0213066f $X=9.06 $Y=0.615
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_664_n N_VPWR_M1010_d 0.00244277f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_689 N_RESET_B_c_666_n N_VPWR_M1015_s 0.00677602f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_690 N_RESET_B_M1035_g N_VPWR_c_1655_n 0.00861602f $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_691 N_RESET_B_M1016_g N_VPWR_c_1657_n 0.0033842f $X=4.87 $Y=2.525 $X2=0 $Y2=0
cc_692 N_RESET_B_M1026_g N_VPWR_c_1659_n 0.00384525f $X=9.02 $Y=2.675 $X2=0
+ $Y2=0
cc_693 N_RESET_B_c_666_n N_VPWR_c_1659_n 0.00679776f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_694 N_RESET_B_c_669_n N_VPWR_c_1659_n 0.0023649f $X=8.88 $Y=2.035 $X2=0 $Y2=0
cc_695 N_RESET_B_c_670_n N_VPWR_c_1659_n 0.0114656f $X=8.88 $Y=2.035 $X2=0 $Y2=0
cc_696 N_RESET_B_c_674_n N_VPWR_c_1659_n 0.00230627f $X=8.975 $Y=2.11 $X2=0
+ $Y2=0
cc_697 N_RESET_B_M1026_g N_VPWR_c_1667_n 0.00600227f $X=9.02 $Y=2.675 $X2=0
+ $Y2=0
cc_698 N_RESET_B_M1035_g N_VPWR_c_1671_n 0.00439065f $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_699 N_RESET_B_M1035_g N_VPWR_c_1652_n 0.00441441f $X=0.95 $Y=2.75 $X2=0 $Y2=0
cc_700 N_RESET_B_M1016_g N_VPWR_c_1652_n 0.00112709f $X=4.87 $Y=2.525 $X2=0
+ $Y2=0
cc_701 N_RESET_B_M1026_g N_VPWR_c_1652_n 0.00626544f $X=9.02 $Y=2.675 $X2=0
+ $Y2=0
cc_702 N_RESET_B_M1005_g N_A_37_78#_c_1822_n 7.80212e-19 $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_703 N_RESET_B_M1035_g N_A_37_78#_c_1829_n 2.23847e-19 $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_704 N_RESET_B_M1005_g N_A_37_78#_c_1823_n 0.0177928f $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_705 N_RESET_B_c_665_n N_A_37_78#_c_1823_n 0.0018287f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_706 N_RESET_B_c_656_n N_A_37_78#_c_1823_n 0.0729934f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_707 N_RESET_B_M1035_g N_A_37_78#_c_1831_n 0.01601f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_664_n N_A_37_78#_c_1831_n 0.0280435f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_709 N_RESET_B_c_665_n N_A_37_78#_c_1831_n 0.00879083f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_656_n N_A_37_78#_c_1831_n 0.0112881f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_711 N_RESET_B_c_673_n N_A_37_78#_c_1831_n 0.00265097f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_664_n N_A_37_78#_c_1832_n 0.0135548f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_664_n N_A_37_78#_c_1825_n 0.00509385f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_714 N_RESET_B_c_664_n N_A_37_78#_c_1827_n 0.0118532f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_715 N_RESET_B_M1005_g N_A_37_78#_c_1828_n 8.54775e-19 $X=0.935 $Y=0.6 $X2=0
+ $Y2=0
cc_716 N_RESET_B_M1035_g N_A_37_78#_c_1834_n 0.00609315f $X=0.95 $Y=2.75 $X2=0
+ $Y2=0
cc_717 N_RESET_B_c_664_n N_A_37_78#_c_1835_n 0.00965531f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_718 N_RESET_B_M1005_g N_VGND_c_2015_n 0.00252332f $X=0.935 $Y=0.6 $X2=0 $Y2=0
cc_719 N_RESET_B_c_649_n N_VGND_c_2015_n 0.0155925f $X=4.69 $Y=0.18 $X2=0 $Y2=0
cc_720 N_RESET_B_c_655_n N_VGND_c_2015_n 0.00122895f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_721 N_RESET_B_c_656_n N_VGND_c_2015_n 0.00978084f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_722 N_RESET_B_c_649_n N_VGND_c_2016_n 0.0257653f $X=4.69 $Y=0.18 $X2=0 $Y2=0
cc_723 N_RESET_B_M1030_g N_VGND_c_2017_n 0.00393134f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_724 N_RESET_B_c_650_n N_VGND_c_2023_n 0.00796123f $X=1.01 $Y=0.18 $X2=0 $Y2=0
cc_725 N_RESET_B_M1030_g N_VGND_c_2025_n 0.00552345f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_726 N_RESET_B_c_649_n N_VGND_c_2027_n 0.0227427f $X=4.69 $Y=0.18 $X2=0 $Y2=0
cc_727 N_RESET_B_c_649_n N_VGND_c_2028_n 0.0563402f $X=4.69 $Y=0.18 $X2=0 $Y2=0
cc_728 N_RESET_B_c_649_n N_VGND_c_2034_n 0.010027f $X=4.69 $Y=0.18 $X2=0 $Y2=0
cc_729 N_RESET_B_c_649_n N_VGND_c_2038_n 0.0937549f $X=4.69 $Y=0.18 $X2=0 $Y2=0
cc_730 N_RESET_B_c_650_n N_VGND_c_2038_n 0.0114838f $X=1.01 $Y=0.18 $X2=0 $Y2=0
cc_731 N_RESET_B_M1030_g N_VGND_c_2038_n 0.00534666f $X=9.06 $Y=0.615 $X2=0
+ $Y2=0
cc_732 N_A_303_395#_c_881_n N_A_702_463#_c_1112_n 0.0242353f $X=6.675 $Y=1.735
+ $X2=0 $Y2=0
cc_733 N_A_303_395#_c_896_n N_A_702_463#_M1015_g 0.00549932f $X=5.385 $Y=3.075
+ $X2=0 $Y2=0
cc_734 N_A_303_395#_M1020_g N_A_702_463#_M1015_g 0.0242353f $X=6.675 $Y=2.46
+ $X2=0 $Y2=0
cc_735 N_A_303_395#_c_901_n N_A_702_463#_M1015_g 0.0141165f $X=6.785 $Y=2.49
+ $X2=0 $Y2=0
cc_736 N_A_303_395#_c_905_n N_A_702_463#_M1015_g 7.93468e-19 $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_737 N_A_303_395#_c_906_n N_A_702_463#_M1015_g 0.0104403f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_738 N_A_303_395#_c_906_n N_A_702_463#_c_1104_n 0.00125125f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_739 N_A_303_395#_c_881_n N_A_702_463#_c_1105_n 0.0214503f $X=6.675 $Y=1.735
+ $X2=0 $Y2=0
cc_740 N_A_303_395#_c_888_n N_A_702_463#_c_1105_n 3.74234e-19 $X=6.87 $Y=1.425
+ $X2=0 $Y2=0
cc_741 N_A_303_395#_c_881_n N_A_702_463#_c_1106_n 0.00590001f $X=6.675 $Y=1.735
+ $X2=0 $Y2=0
cc_742 N_A_303_395#_c_880_n N_A_702_463#_c_1107_n 6.23807e-19 $X=3.485 $Y=1.185
+ $X2=0 $Y2=0
cc_743 N_A_303_395#_M1019_g N_A_702_463#_c_1107_n 0.00143908f $X=3.87 $Y=2.525
+ $X2=0 $Y2=0
cc_744 N_A_303_395#_c_895_n N_A_702_463#_c_1143_n 0.00138474f $X=5.31 $Y=3.15
+ $X2=0 $Y2=0
cc_745 N_A_303_395#_c_906_n N_A_702_463#_c_1108_n 5.16665e-19 $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_746 N_A_303_395#_c_880_n N_A_702_463#_c_1111_n 0.00204771f $X=3.485 $Y=1.185
+ $X2=0 $Y2=0
cc_747 N_A_303_395#_c_891_n N_A_702_463#_c_1117_n 0.00314225f $X=3.78 $Y=3.15
+ $X2=0 $Y2=0
cc_748 N_A_303_395#_M1019_g N_A_702_463#_c_1117_n 0.0156337f $X=3.87 $Y=2.525
+ $X2=0 $Y2=0
cc_749 N_A_303_395#_c_895_n N_A_702_463#_c_1118_n 0.00255153f $X=5.31 $Y=3.15
+ $X2=0 $Y2=0
cc_750 N_A_303_395#_c_895_n N_A_702_463#_c_1119_n 0.00475781f $X=5.31 $Y=3.15
+ $X2=0 $Y2=0
cc_751 N_A_303_395#_c_905_n N_A_702_463#_c_1119_n 0.0190155f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_752 N_A_303_395#_c_906_n N_A_702_463#_c_1119_n 0.0069024f $X=5.56 $Y=2.375
+ $X2=0 $Y2=0
cc_753 N_A_303_395#_M1037_g N_A_1678_395#_M1022_g 0.0378955f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_754 N_A_303_395#_c_882_n N_A_1678_395#_c_1242_n 0.0216911f $X=8.085 $Y=1.66
+ $X2=0 $Y2=0
cc_755 N_A_303_395#_M1037_g N_A_1678_395#_c_1246_n 4.34985e-19 $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_756 N_A_303_395#_M1037_g N_A_1678_395#_c_1247_n 0.0216911f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_757 N_A_303_395#_c_901_n N_A_1353_392#_M1020_d 0.00477838f $X=6.785 $Y=2.49
+ $X2=0 $Y2=0
cc_758 N_A_303_395#_c_902_n N_A_1353_392#_M1020_d 0.00633951f $X=6.87 $Y=2.405
+ $X2=0 $Y2=0
cc_759 N_A_303_395#_c_881_n N_A_1353_392#_c_1371_n 0.00127705f $X=6.675 $Y=1.735
+ $X2=0 $Y2=0
cc_760 N_A_303_395#_M1020_g N_A_1353_392#_c_1371_n 0.00977626f $X=6.675 $Y=2.46
+ $X2=0 $Y2=0
cc_761 N_A_303_395#_c_882_n N_A_1353_392#_c_1371_n 0.013648f $X=8.085 $Y=1.66
+ $X2=0 $Y2=0
cc_762 N_A_303_395#_c_901_n N_A_1353_392#_c_1371_n 0.0140222f $X=6.785 $Y=2.49
+ $X2=0 $Y2=0
cc_763 N_A_303_395#_c_902_n N_A_1353_392#_c_1371_n 0.051078f $X=6.87 $Y=2.405
+ $X2=0 $Y2=0
cc_764 N_A_303_395#_c_888_n N_A_1353_392#_c_1371_n 0.0231503f $X=6.87 $Y=1.425
+ $X2=0 $Y2=0
cc_765 N_A_303_395#_M1037_g N_A_1353_392#_c_1372_n 0.00507341f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_766 N_A_303_395#_c_882_n N_A_1353_392#_c_1385_n 2.44969e-19 $X=8.085 $Y=1.66
+ $X2=0 $Y2=0
cc_767 N_A_303_395#_M1037_g N_A_1353_392#_c_1374_n 0.00153073f $X=8.16 $Y=0.615
+ $X2=0 $Y2=0
cc_768 N_A_303_395#_c_901_n N_VPWR_M1015_s 0.00535876f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_769 N_A_303_395#_c_889_n N_VPWR_c_1656_n 0.0136934f $X=2.395 $Y=1.885 $X2=0
+ $Y2=0
cc_770 N_A_303_395#_c_890_n N_VPWR_c_1656_n 0.00260315f $X=2.905 $Y=3.075 $X2=0
+ $Y2=0
cc_771 N_A_303_395#_M1019_g N_VPWR_c_1657_n 0.00610747f $X=3.87 $Y=2.525 $X2=0
+ $Y2=0
cc_772 N_A_303_395#_c_895_n N_VPWR_c_1657_n 0.0250293f $X=5.31 $Y=3.15 $X2=0
+ $Y2=0
cc_773 N_A_303_395#_c_896_n N_VPWR_c_1657_n 0.00529092f $X=5.385 $Y=3.075 $X2=0
+ $Y2=0
cc_774 N_A_303_395#_c_896_n N_VPWR_c_1658_n 0.0101782f $X=5.385 $Y=3.075 $X2=0
+ $Y2=0
cc_775 N_A_303_395#_M1020_g N_VPWR_c_1658_n 0.00165549f $X=6.675 $Y=2.46 $X2=0
+ $Y2=0
cc_776 N_A_303_395#_c_901_n N_VPWR_c_1658_n 0.0216308f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_777 N_A_303_395#_M1020_g N_VPWR_c_1665_n 0.00406265f $X=6.675 $Y=2.46 $X2=0
+ $Y2=0
cc_778 N_A_303_395#_c_901_n N_VPWR_c_1665_n 0.0094867f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_779 N_A_303_395#_c_889_n N_VPWR_c_1673_n 0.00583607f $X=2.395 $Y=1.885 $X2=0
+ $Y2=0
cc_780 N_A_303_395#_c_892_n N_VPWR_c_1673_n 0.0441814f $X=2.98 $Y=3.15 $X2=0
+ $Y2=0
cc_781 N_A_303_395#_c_895_n N_VPWR_c_1674_n 0.0212613f $X=5.31 $Y=3.15 $X2=0
+ $Y2=0
cc_782 N_A_303_395#_c_901_n N_VPWR_c_1674_n 0.00150121f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_783 N_A_303_395#_c_905_n N_VPWR_c_1674_n 0.00478946f $X=5.56 $Y=2.375 $X2=0
+ $Y2=0
cc_784 N_A_303_395#_M1010_s N_VPWR_c_1652_n 0.00377894f $X=1.515 $Y=1.975 $X2=0
+ $Y2=0
cc_785 N_A_303_395#_c_889_n N_VPWR_c_1652_n 0.00541847f $X=2.395 $Y=1.885 $X2=0
+ $Y2=0
cc_786 N_A_303_395#_c_891_n N_VPWR_c_1652_n 0.022687f $X=3.78 $Y=3.15 $X2=0
+ $Y2=0
cc_787 N_A_303_395#_c_892_n N_VPWR_c_1652_n 0.00567376f $X=2.98 $Y=3.15 $X2=0
+ $Y2=0
cc_788 N_A_303_395#_c_895_n N_VPWR_c_1652_n 0.0407681f $X=5.31 $Y=3.15 $X2=0
+ $Y2=0
cc_789 N_A_303_395#_M1020_g N_VPWR_c_1652_n 0.00535823f $X=6.675 $Y=2.46 $X2=0
+ $Y2=0
cc_790 N_A_303_395#_c_900_n N_VPWR_c_1652_n 0.00494927f $X=3.87 $Y=3.15 $X2=0
+ $Y2=0
cc_791 N_A_303_395#_c_901_n N_VPWR_c_1652_n 0.0232028f $X=6.785 $Y=2.49 $X2=0
+ $Y2=0
cc_792 N_A_303_395#_c_905_n N_VPWR_c_1652_n 0.00841698f $X=5.56 $Y=2.375 $X2=0
+ $Y2=0
cc_793 N_A_303_395#_c_884_n N_A_37_78#_c_1823_n 0.00463142f $X=1.69 $Y=0.715
+ $X2=0 $Y2=0
cc_794 N_A_303_395#_c_886_n N_A_37_78#_c_1823_n 0.00556056f $X=1.665 $Y=1.055
+ $X2=0 $Y2=0
cc_795 N_A_303_395#_c_903_n N_A_37_78#_c_1823_n 0.00242029f $X=1.64 $Y=2.135
+ $X2=0 $Y2=0
cc_796 N_A_303_395#_M1010_s N_A_37_78#_c_1831_n 0.00711239f $X=1.515 $Y=1.975
+ $X2=0 $Y2=0
cc_797 N_A_303_395#_c_889_n N_A_37_78#_c_1831_n 0.0138781f $X=2.395 $Y=1.885
+ $X2=0 $Y2=0
cc_798 N_A_303_395#_c_890_n N_A_37_78#_c_1831_n 0.0123779f $X=2.905 $Y=3.075
+ $X2=0 $Y2=0
cc_799 N_A_303_395#_c_903_n N_A_37_78#_c_1831_n 0.0253284f $X=1.64 $Y=2.135
+ $X2=0 $Y2=0
cc_800 N_A_303_395#_c_878_n N_A_37_78#_c_1824_n 0.00683285f $X=3.41 $Y=1.26
+ $X2=0 $Y2=0
cc_801 N_A_303_395#_c_880_n N_A_37_78#_c_1824_n 0.00878411f $X=3.485 $Y=1.185
+ $X2=0 $Y2=0
cc_802 N_A_303_395#_M1019_g N_A_37_78#_c_1832_n 0.00240447f $X=3.87 $Y=2.525
+ $X2=0 $Y2=0
cc_803 N_A_303_395#_c_878_n N_A_37_78#_c_1825_n 0.00831879f $X=3.41 $Y=1.26
+ $X2=0 $Y2=0
cc_804 N_A_303_395#_c_878_n N_A_37_78#_c_1826_n 0.00522272f $X=3.41 $Y=1.26
+ $X2=0 $Y2=0
cc_805 N_A_303_395#_c_879_n N_A_37_78#_c_1826_n 0.00110212f $X=3.02 $Y=1.26
+ $X2=0 $Y2=0
cc_806 N_A_303_395#_c_879_n N_A_37_78#_c_1827_n 0.00176032f $X=3.02 $Y=1.26
+ $X2=0 $Y2=0
cc_807 N_A_303_395#_c_890_n N_A_37_78#_c_1835_n 0.00971976f $X=2.905 $Y=3.075
+ $X2=0 $Y2=0
cc_808 N_A_303_395#_c_891_n N_A_37_78#_c_1835_n 0.00524628f $X=3.78 $Y=3.15
+ $X2=0 $Y2=0
cc_809 N_A_303_395#_M1019_g N_A_37_78#_c_1835_n 5.36766e-19 $X=3.87 $Y=2.525
+ $X2=0 $Y2=0
cc_810 N_A_303_395#_c_914_n N_VGND_M1001_d 0.00639859f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_811 N_A_303_395#_c_884_n N_VGND_c_2015_n 0.0317977f $X=1.69 $Y=0.715 $X2=0
+ $Y2=0
cc_812 N_A_303_395#_c_877_n N_VGND_c_2016_n 0.00119784f $X=2.47 $Y=1.41 $X2=0
+ $Y2=0
cc_813 N_A_303_395#_c_884_n N_VGND_c_2016_n 0.0295324f $X=1.69 $Y=0.715 $X2=0
+ $Y2=0
cc_814 N_A_303_395#_c_914_n N_VGND_c_2016_n 0.0208278f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_815 N_A_303_395#_c_884_n N_VGND_c_2027_n 0.0186352f $X=1.69 $Y=0.715 $X2=0
+ $Y2=0
cc_816 N_A_303_395#_M1037_g N_VGND_c_2029_n 9.33926e-19 $X=8.16 $Y=0.615 $X2=0
+ $Y2=0
cc_817 N_A_303_395#_c_877_n N_VGND_c_2038_n 9.39239e-19 $X=2.47 $Y=1.41 $X2=0
+ $Y2=0
cc_818 N_A_303_395#_c_884_n N_VGND_c_2038_n 0.0137621f $X=1.69 $Y=0.715 $X2=0
+ $Y2=0
cc_819 N_A_702_463#_c_1143_n N_VPWR_M1006_d 0.00750623f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_820 N_A_702_463#_c_1143_n N_VPWR_c_1657_n 0.0255562f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_821 N_A_702_463#_c_1118_n N_VPWR_c_1657_n 0.00285906f $X=4.23 $Y=2.587 $X2=0
+ $Y2=0
cc_822 N_A_702_463#_c_1119_n N_VPWR_c_1657_n 0.00110155f $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_823 N_A_702_463#_M1015_g N_VPWR_c_1658_n 0.00976492f $X=6.225 $Y=2.46 $X2=0
+ $Y2=0
cc_824 N_A_702_463#_c_1119_n N_VPWR_c_1658_n 3.02124e-19 $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_825 N_A_702_463#_M1015_g N_VPWR_c_1665_n 0.00337973f $X=6.225 $Y=2.46 $X2=0
+ $Y2=0
cc_826 N_A_702_463#_c_1143_n N_VPWR_c_1673_n 0.00183105f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_827 N_A_702_463#_c_1117_n N_VPWR_c_1673_n 0.0154923f $X=3.965 $Y=2.587 $X2=0
+ $Y2=0
cc_828 N_A_702_463#_c_1119_n N_VPWR_c_1674_n 0.00791714f $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_829 N_A_702_463#_M1015_g N_VPWR_c_1652_n 0.00439578f $X=6.225 $Y=2.46 $X2=0
+ $Y2=0
cc_830 N_A_702_463#_c_1143_n N_VPWR_c_1652_n 0.00519397f $X=4.745 $Y=2.485 $X2=0
+ $Y2=0
cc_831 N_A_702_463#_c_1117_n N_VPWR_c_1652_n 0.0187716f $X=3.965 $Y=2.587 $X2=0
+ $Y2=0
cc_832 N_A_702_463#_c_1119_n N_VPWR_c_1652_n 0.0110248f $X=4.83 $Y=2.525 $X2=0
+ $Y2=0
cc_833 N_A_702_463#_c_1107_n N_A_37_78#_c_1824_n 0.0046376f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_834 N_A_702_463#_c_1111_n N_A_37_78#_c_1824_n 0.014524f $X=3.77 $Y=0.86 $X2=0
+ $Y2=0
cc_835 N_A_702_463#_c_1107_n N_A_37_78#_c_1832_n 0.013816f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_836 N_A_702_463#_c_1117_n N_A_37_78#_c_1832_n 0.0173919f $X=3.965 $Y=2.587
+ $X2=0 $Y2=0
cc_837 N_A_702_463#_c_1107_n N_A_37_78#_c_1825_n 0.0135526f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_838 N_A_702_463#_c_1111_n N_A_37_78#_c_1825_n 0.0160421f $X=3.77 $Y=0.86
+ $X2=0 $Y2=0
cc_839 N_A_702_463#_c_1107_n N_A_37_78#_c_1827_n 0.0519798f $X=4.05 $Y=2.4 $X2=0
+ $Y2=0
cc_840 N_A_702_463#_c_1107_n N_A_37_78#_c_1835_n 0.00211076f $X=4.05 $Y=2.4
+ $X2=0 $Y2=0
cc_841 N_A_702_463#_c_1117_n N_A_37_78#_c_1835_n 0.013112f $X=3.965 $Y=2.587
+ $X2=0 $Y2=0
cc_842 N_A_702_463#_c_1107_n A_792_463# 2.74036e-19 $X=4.05 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_843 N_A_702_463#_c_1118_n A_792_463# 2.73178e-19 $X=4.23 $Y=2.587 $X2=-0.19
+ $Y2=-0.245
cc_844 N_A_702_463#_c_1103_n N_VGND_c_2029_n 0.00278271f $X=5.685 $Y=1.22 $X2=0
+ $Y2=0
cc_845 N_A_702_463#_c_1103_n N_VGND_c_2034_n 4.07279e-19 $X=5.685 $Y=1.22 $X2=0
+ $Y2=0
cc_846 N_A_702_463#_c_1103_n N_VGND_c_2038_n 0.00363426f $X=5.685 $Y=1.22 $X2=0
+ $Y2=0
cc_847 N_A_702_463#_c_1107_n A_812_138# 4.92957e-19 $X=4.05 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_848 N_A_702_463#_c_1111_n A_812_138# 0.00171007f $X=3.77 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_849 N_A_1678_395#_c_1243_n N_A_1353_392#_M1031_g 0.0108485f $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_850 N_A_1678_395#_c_1244_n N_A_1353_392#_M1031_g 0.0168963f $X=9.665 $Y=0.615
+ $X2=0 $Y2=0
cc_851 N_A_1678_395#_c_1245_n N_A_1353_392#_M1031_g 0.00530998f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_852 N_A_1678_395#_c_1248_n N_A_1353_392#_M1031_g 0.00445436f $X=9.722 $Y=1.12
+ $X2=0 $Y2=0
cc_853 N_A_1678_395#_c_1252_n N_A_1353_392#_M1027_g 0.0124793f $X=9.395 $Y=2.445
+ $X2=0 $Y2=0
cc_854 N_A_1678_395#_c_1253_n N_A_1353_392#_M1027_g 0.00808979f $X=9.775 $Y=1.96
+ $X2=0 $Y2=0
cc_855 N_A_1678_395#_c_1254_n N_A_1353_392#_M1027_g 0.00374598f $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_856 N_A_1678_395#_c_1245_n N_A_1353_392#_M1027_g 0.00340775f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_857 N_A_1678_395#_c_1256_n N_A_1353_392#_M1027_g 0.00962273f $X=9.395
+ $Y=2.675 $X2=0 $Y2=0
cc_858 N_A_1678_395#_c_1245_n N_A_1353_392#_c_1364_n 0.00646442f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_859 N_A_1678_395#_c_1248_n N_A_1353_392#_c_1364_n 0.00210562f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_860 N_A_1678_395#_c_1252_n N_A_1353_392#_M1008_g 0.00139999f $X=9.395
+ $Y=2.445 $X2=0 $Y2=0
cc_861 N_A_1678_395#_c_1253_n N_A_1353_392#_M1008_g 0.00718285f $X=9.775 $Y=1.96
+ $X2=0 $Y2=0
cc_862 N_A_1678_395#_c_1245_n N_A_1353_392#_M1008_g 0.00347834f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_863 N_A_1678_395#_c_1245_n N_A_1353_392#_c_1366_n 2.16647e-19 $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_864 N_A_1678_395#_c_1245_n N_A_1353_392#_c_1367_n 0.00420863f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_865 N_A_1678_395#_c_1248_n N_A_1353_392#_c_1369_n 0.00110652f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_866 N_A_1678_395#_c_1245_n N_A_1353_392#_c_1370_n 0.00382761f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_867 N_A_1678_395#_c_1248_n N_A_1353_392#_c_1370_n 4.03357e-19 $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_868 N_A_1678_395#_M1012_g N_A_1353_392#_c_1406_n 0.00723124f $X=8.48 $Y=2.675
+ $X2=0 $Y2=0
cc_869 N_A_1678_395#_M1012_g N_A_1353_392#_c_1385_n 0.00781998f $X=8.48 $Y=2.675
+ $X2=0 $Y2=0
cc_870 N_A_1678_395#_c_1242_n N_A_1353_392#_c_1385_n 0.00937113f $X=8.492
+ $Y=1.975 $X2=0 $Y2=0
cc_871 N_A_1678_395#_c_1251_n N_A_1353_392#_c_1385_n 0.00314765f $X=8.492
+ $Y=2.125 $X2=0 $Y2=0
cc_872 N_A_1678_395#_c_1242_n N_A_1353_392#_c_1373_n 0.0106324f $X=8.492
+ $Y=1.975 $X2=0 $Y2=0
cc_873 N_A_1678_395#_c_1251_n N_A_1353_392#_c_1373_n 0.0010085f $X=8.492
+ $Y=2.125 $X2=0 $Y2=0
cc_874 N_A_1678_395#_c_1243_n N_A_1353_392#_c_1373_n 0.0259611f $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_875 N_A_1678_395#_c_1254_n N_A_1353_392#_c_1373_n 0.00291458f $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_876 N_A_1678_395#_c_1246_n N_A_1353_392#_c_1373_n 0.0236067f $X=8.61 $Y=1.12
+ $X2=0 $Y2=0
cc_877 N_A_1678_395#_c_1247_n N_A_1353_392#_c_1373_n 0.00125903f $X=8.61 $Y=1.2
+ $X2=0 $Y2=0
cc_878 N_A_1678_395#_c_1243_n N_A_1353_392#_c_1375_n 0.0111296f $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_879 N_A_1678_395#_c_1253_n N_A_1353_392#_c_1375_n 0.00903277f $X=9.775
+ $Y=1.96 $X2=0 $Y2=0
cc_880 N_A_1678_395#_c_1254_n N_A_1353_392#_c_1375_n 0.0107527f $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_881 N_A_1678_395#_c_1245_n N_A_1353_392#_c_1375_n 0.0237947f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_882 N_A_1678_395#_c_1248_n N_A_1353_392#_c_1375_n 0.00870087f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_883 N_A_1678_395#_c_1243_n N_A_1353_392#_c_1376_n 2.04435e-19 $X=9.5 $Y=1.12
+ $X2=0 $Y2=0
cc_884 N_A_1678_395#_c_1253_n N_A_1353_392#_c_1376_n 0.00306014f $X=9.775
+ $Y=1.96 $X2=0 $Y2=0
cc_885 N_A_1678_395#_c_1254_n N_A_1353_392#_c_1376_n 2.63281e-19 $X=9.48 $Y=1.96
+ $X2=0 $Y2=0
cc_886 N_A_1678_395#_c_1245_n N_A_1353_392#_c_1376_n 0.00218969f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_887 N_A_1678_395#_c_1248_n N_A_1353_392#_c_1376_n 0.00294175f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_888 N_A_1678_395#_c_1253_n N_A_2013_409#_c_1548_n 0.013857f $X=9.775 $Y=1.96
+ $X2=0 $Y2=0
cc_889 N_A_1678_395#_c_1245_n N_A_2013_409#_c_1548_n 0.0176781f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_890 N_A_1678_395#_c_1245_n N_A_2013_409#_c_1538_n 0.0137366f $X=9.86 $Y=1.875
+ $X2=0 $Y2=0
cc_891 N_A_1678_395#_c_1245_n N_A_2013_409#_c_1539_n 0.00265607f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_892 N_A_1678_395#_c_1248_n N_A_2013_409#_c_1539_n 0.00237986f $X=9.722
+ $Y=1.12 $X2=0 $Y2=0
cc_893 N_A_1678_395#_c_1245_n N_A_2013_409#_c_1541_n 0.00529677f $X=9.86
+ $Y=1.875 $X2=0 $Y2=0
cc_894 N_A_1678_395#_c_1253_n N_VPWR_M1027_d 0.00184301f $X=9.775 $Y=1.96 $X2=0
+ $Y2=0
cc_895 N_A_1678_395#_M1012_g N_VPWR_c_1659_n 0.00424898f $X=8.48 $Y=2.675 $X2=0
+ $Y2=0
cc_896 N_A_1678_395#_c_1251_n N_VPWR_c_1659_n 5.77237e-19 $X=8.492 $Y=2.125
+ $X2=0 $Y2=0
cc_897 N_A_1678_395#_c_1256_n N_VPWR_c_1659_n 0.0193003f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_898 N_A_1678_395#_c_1253_n N_VPWR_c_1660_n 0.0100122f $X=9.775 $Y=1.96 $X2=0
+ $Y2=0
cc_899 N_A_1678_395#_c_1256_n N_VPWR_c_1660_n 0.0355217f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_900 N_A_1678_395#_M1012_g N_VPWR_c_1665_n 0.00611098f $X=8.48 $Y=2.675 $X2=0
+ $Y2=0
cc_901 N_A_1678_395#_c_1256_n N_VPWR_c_1667_n 0.0129427f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_902 N_A_1678_395#_M1012_g N_VPWR_c_1652_n 0.00626544f $X=8.48 $Y=2.675 $X2=0
+ $Y2=0
cc_903 N_A_1678_395#_c_1256_n N_VPWR_c_1652_n 0.0137485f $X=9.395 $Y=2.675 $X2=0
+ $Y2=0
cc_904 N_A_1678_395#_M1022_g N_VGND_c_2017_n 0.00207012f $X=8.55 $Y=0.615 $X2=0
+ $Y2=0
cc_905 N_A_1678_395#_c_1243_n N_VGND_c_2017_n 0.0139742f $X=9.5 $Y=1.12 $X2=0
+ $Y2=0
cc_906 N_A_1678_395#_c_1244_n N_VGND_c_2017_n 0.00732847f $X=9.665 $Y=0.615
+ $X2=0 $Y2=0
cc_907 N_A_1678_395#_c_1246_n N_VGND_c_2017_n 0.0115305f $X=8.61 $Y=1.12 $X2=0
+ $Y2=0
cc_908 N_A_1678_395#_c_1247_n N_VGND_c_2017_n 0.00115479f $X=8.61 $Y=1.2 $X2=0
+ $Y2=0
cc_909 N_A_1678_395#_c_1244_n N_VGND_c_2018_n 0.0362241f $X=9.665 $Y=0.615 $X2=0
+ $Y2=0
cc_910 N_A_1678_395#_c_1248_n N_VGND_c_2018_n 0.00818535f $X=9.722 $Y=1.12 $X2=0
+ $Y2=0
cc_911 N_A_1678_395#_c_1244_n N_VGND_c_2025_n 0.0127604f $X=9.665 $Y=0.615 $X2=0
+ $Y2=0
cc_912 N_A_1678_395#_M1022_g N_VGND_c_2029_n 0.00551028f $X=8.55 $Y=0.615 $X2=0
+ $Y2=0
cc_913 N_A_1678_395#_M1022_g N_VGND_c_2038_n 0.00534666f $X=8.55 $Y=0.615 $X2=0
+ $Y2=0
cc_914 N_A_1678_395#_c_1244_n N_VGND_c_2038_n 0.011834f $X=9.665 $Y=0.615 $X2=0
+ $Y2=0
cc_915 N_A_1353_392#_c_1368_n N_A_2013_409#_M1009_g 0.0146425f $X=10.425 $Y=1.63
+ $X2=0 $Y2=0
cc_916 N_A_1353_392#_c_1366_n N_A_2013_409#_c_1527_n 0.0146425f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_917 N_A_1353_392#_c_1366_n N_A_2013_409#_c_1531_n 0.00125363f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_918 N_A_1353_392#_c_1370_n N_A_2013_409#_c_1531_n 4.19636e-19 $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_919 N_A_1353_392#_M1008_g N_A_2013_409#_c_1548_n 0.00333791f $X=9.975
+ $Y=2.465 $X2=0 $Y2=0
cc_920 N_A_1353_392#_c_1365_n N_A_2013_409#_c_1548_n 0.00471727f $X=10.335
+ $Y=1.63 $X2=0 $Y2=0
cc_921 N_A_1353_392#_M1025_g N_A_2013_409#_c_1548_n 0.0213472f $X=10.425
+ $Y=2.465 $X2=0 $Y2=0
cc_922 N_A_1353_392#_c_1368_n N_A_2013_409#_c_1548_n 0.00143923f $X=10.425
+ $Y=1.63 $X2=0 $Y2=0
cc_923 N_A_1353_392#_c_1366_n N_A_2013_409#_c_1537_n 0.00840659f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_924 N_A_1353_392#_c_1368_n N_A_2013_409#_c_1537_n 0.00862712f $X=10.425
+ $Y=1.63 $X2=0 $Y2=0
cc_925 N_A_1353_392#_c_1370_n N_A_2013_409#_c_1537_n 0.00194299f $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_926 N_A_1353_392#_c_1365_n N_A_2013_409#_c_1538_n 0.00614927f $X=10.335
+ $Y=1.63 $X2=0 $Y2=0
cc_927 N_A_1353_392#_c_1366_n N_A_2013_409#_c_1538_n 0.00148617f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_928 N_A_1353_392#_c_1368_n N_A_2013_409#_c_1538_n 6.95643e-19 $X=10.425
+ $Y=1.63 $X2=0 $Y2=0
cc_929 N_A_1353_392#_c_1369_n N_A_2013_409#_c_1539_n 0.0127757f $X=10.475
+ $Y=1.185 $X2=0 $Y2=0
cc_930 N_A_1353_392#_c_1370_n N_A_2013_409#_c_1539_n 0.00490997f $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_931 N_A_1353_392#_c_1366_n N_A_2013_409#_c_1541_n 0.0026095f $X=10.44
+ $Y=1.555 $X2=0 $Y2=0
cc_932 N_A_1353_392#_c_1370_n N_A_2013_409#_c_1541_n 0.00200729f $X=10.475
+ $Y=1.335 $X2=0 $Y2=0
cc_933 N_A_1353_392#_c_1385_n N_VPWR_c_1659_n 0.00177329f $X=8.325 $Y=2.475
+ $X2=0 $Y2=0
cc_934 N_A_1353_392#_M1027_g N_VPWR_c_1660_n 0.00443836f $X=9.47 $Y=2.675 $X2=0
+ $Y2=0
cc_935 N_A_1353_392#_M1008_g N_VPWR_c_1660_n 0.00971757f $X=9.975 $Y=2.465 $X2=0
+ $Y2=0
cc_936 N_A_1353_392#_M1025_g N_VPWR_c_1660_n 5.19678e-19 $X=10.425 $Y=2.465
+ $X2=0 $Y2=0
cc_937 N_A_1353_392#_M1025_g N_VPWR_c_1661_n 0.00296024f $X=10.425 $Y=2.465
+ $X2=0 $Y2=0
cc_938 N_A_1353_392#_c_1371_n N_VPWR_c_1665_n 0.00505902f $X=7.245 $Y=2.475
+ $X2=0 $Y2=0
cc_939 N_A_1353_392#_c_1406_n N_VPWR_c_1665_n 0.0235999f $X=8.24 $Y=2.64 $X2=0
+ $Y2=0
cc_940 N_A_1353_392#_M1027_g N_VPWR_c_1667_n 0.00533576f $X=9.47 $Y=2.675 $X2=0
+ $Y2=0
cc_941 N_A_1353_392#_M1008_g N_VPWR_c_1669_n 0.00575164f $X=9.975 $Y=2.465 $X2=0
+ $Y2=0
cc_942 N_A_1353_392#_M1025_g N_VPWR_c_1669_n 0.00601158f $X=10.425 $Y=2.465
+ $X2=0 $Y2=0
cc_943 N_A_1353_392#_M1027_g N_VPWR_c_1652_n 0.00626544f $X=9.47 $Y=2.675 $X2=0
+ $Y2=0
cc_944 N_A_1353_392#_M1008_g N_VPWR_c_1652_n 0.00577812f $X=9.975 $Y=2.465 $X2=0
+ $Y2=0
cc_945 N_A_1353_392#_M1025_g N_VPWR_c_1652_n 0.00626544f $X=10.425 $Y=2.465
+ $X2=0 $Y2=0
cc_946 N_A_1353_392#_c_1371_n N_VPWR_c_1652_n 0.00669727f $X=7.245 $Y=2.475
+ $X2=0 $Y2=0
cc_947 N_A_1353_392#_c_1406_n N_VPWR_c_1652_n 0.0343488f $X=8.24 $Y=2.64 $X2=0
+ $Y2=0
cc_948 N_A_1353_392#_c_1406_n A_1630_493# 0.00250904f $X=8.24 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_949 N_A_1353_392#_M1031_g N_VGND_c_2018_n 0.00460851f $X=9.45 $Y=0.615 $X2=0
+ $Y2=0
cc_950 N_A_1353_392#_c_1365_n N_VGND_c_2018_n 0.0015097f $X=10.335 $Y=1.63 $X2=0
+ $Y2=0
cc_951 N_A_1353_392#_c_1369_n N_VGND_c_2018_n 0.0197658f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_952 N_A_1353_392#_c_1370_n N_VGND_c_2018_n 8.25701e-19 $X=10.475 $Y=1.335
+ $X2=0 $Y2=0
cc_953 N_A_1353_392#_c_1369_n N_VGND_c_2019_n 0.00422452f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_954 N_A_1353_392#_M1031_g N_VGND_c_2025_n 0.00527282f $X=9.45 $Y=0.615 $X2=0
+ $Y2=0
cc_955 N_A_1353_392#_c_1369_n N_VGND_c_2030_n 0.00434272f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_956 N_A_1353_392#_M1031_g N_VGND_c_2038_n 0.00534666f $X=9.45 $Y=0.615 $X2=0
+ $Y2=0
cc_957 N_A_1353_392#_c_1369_n N_VGND_c_2038_n 0.00830058f $X=10.475 $Y=1.185
+ $X2=0 $Y2=0
cc_958 N_A_2013_409#_c_1548_n N_VPWR_c_1660_n 0.0143519f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_959 N_A_2013_409#_M1009_g N_VPWR_c_1661_n 0.017977f $X=10.93 $Y=2.4 $X2=0
+ $Y2=0
cc_960 N_A_2013_409#_M1021_g N_VPWR_c_1661_n 5.94112e-19 $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_961 N_A_2013_409#_c_1548_n N_VPWR_c_1661_n 0.0332253f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_962 N_A_2013_409#_c_1537_n N_VPWR_c_1661_n 0.00110837f $X=10.56 $Y=1.545
+ $X2=0 $Y2=0
cc_963 N_A_2013_409#_c_1541_n N_VPWR_c_1661_n 0.0137311f $X=10.725 $Y=1.465
+ $X2=0 $Y2=0
cc_964 N_A_2013_409#_M1021_g N_VPWR_c_1662_n 0.00667517f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_965 N_A_2013_409#_M1028_g N_VPWR_c_1662_n 0.00667517f $X=12.35 $Y=2.4 $X2=0
+ $Y2=0
cc_966 N_A_2013_409#_M1029_g N_VPWR_c_1664_n 0.00394849f $X=12.8 $Y=2.4 $X2=0
+ $Y2=0
cc_967 N_A_2013_409#_c_1543_n N_VPWR_c_1664_n 5.6762e-19 $X=12.8 $Y=1.48 $X2=0
+ $Y2=0
cc_968 N_A_2013_409#_c_1548_n N_VPWR_c_1669_n 0.00841313f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_969 N_A_2013_409#_M1009_g N_VPWR_c_1675_n 0.00475445f $X=10.93 $Y=2.4 $X2=0
+ $Y2=0
cc_970 N_A_2013_409#_M1021_g N_VPWR_c_1675_n 0.005209f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_971 N_A_2013_409#_M1028_g N_VPWR_c_1676_n 0.005209f $X=12.35 $Y=2.4 $X2=0
+ $Y2=0
cc_972 N_A_2013_409#_M1029_g N_VPWR_c_1676_n 0.005209f $X=12.8 $Y=2.4 $X2=0
+ $Y2=0
cc_973 N_A_2013_409#_M1009_g N_VPWR_c_1652_n 0.00939102f $X=10.93 $Y=2.4 $X2=0
+ $Y2=0
cc_974 N_A_2013_409#_M1021_g N_VPWR_c_1652_n 0.00987168f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_975 N_A_2013_409#_M1028_g N_VPWR_c_1652_n 0.00986727f $X=12.35 $Y=2.4 $X2=0
+ $Y2=0
cc_976 N_A_2013_409#_M1029_g N_VPWR_c_1652_n 0.00985721f $X=12.8 $Y=2.4 $X2=0
+ $Y2=0
cc_977 N_A_2013_409#_c_1548_n N_VPWR_c_1652_n 0.00870638f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_978 N_A_2013_409#_M1009_g N_Q_c_1950_n 4.36913e-19 $X=10.93 $Y=2.4 $X2=0
+ $Y2=0
cc_979 N_A_2013_409#_M1021_g N_Q_c_1950_n 0.0183863f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_980 N_A_2013_409#_M1021_g N_Q_c_1951_n 0.0150541f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_981 N_A_2013_409#_c_1530_n N_Q_c_1951_n 0.0138254f $X=11.95 $Y=1.465 $X2=0
+ $Y2=0
cc_982 N_A_2013_409#_M1028_g N_Q_c_1951_n 0.0165635f $X=12.35 $Y=2.4 $X2=0 $Y2=0
cc_983 N_A_2013_409#_c_1540_n N_Q_c_1951_n 0.0650941f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_984 N_A_2013_409#_M1009_g N_Q_c_1952_n 7.29949e-19 $X=10.93 $Y=2.4 $X2=0
+ $Y2=0
cc_985 N_A_2013_409#_M1021_g N_Q_c_1952_n 0.00133968f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_986 N_A_2013_409#_c_1548_n N_Q_c_1952_n 0.0026242f $X=10.2 $Y=2.19 $X2=0
+ $Y2=0
cc_987 N_A_2013_409#_c_1540_n N_Q_c_1952_n 0.0276603f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_988 N_A_2013_409#_c_1542_n N_Q_c_1952_n 0.00272801f $X=11.23 $Y=1.465 $X2=0
+ $Y2=0
cc_989 N_A_2013_409#_M1003_g N_Q_c_1943_n 2.01997e-19 $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_990 N_A_2013_409#_c_1530_n N_Q_c_1943_n 0.00454265f $X=11.95 $Y=1.465 $X2=0
+ $Y2=0
cc_991 N_A_2013_409#_c_1540_n N_Q_c_1943_n 0.0265674f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_992 N_A_2013_409#_M1003_g N_Q_c_1944_n 3.0578e-19 $X=11.5 $Y=0.74 $X2=0 $Y2=0
cc_993 N_A_2013_409#_M1023_g N_Q_c_1944_n 2.92386e-19 $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_994 N_A_2013_409#_M1023_g N_Q_c_1945_n 0.0154071f $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_995 N_A_2013_409#_M1032_g N_Q_c_1945_n 0.0148564f $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_996 N_A_2013_409#_c_1540_n N_Q_c_1945_n 0.0248822f $X=12.075 $Y=1.465 $X2=0
+ $Y2=0
cc_997 N_A_2013_409#_c_1543_n N_Q_c_1945_n 0.00876922f $X=12.8 $Y=1.48 $X2=0
+ $Y2=0
cc_998 N_A_2013_409#_M1028_g N_Q_c_1953_n 0.0184131f $X=12.35 $Y=2.4 $X2=0 $Y2=0
cc_999 N_A_2013_409#_M1029_g N_Q_c_1953_n 0.0129396f $X=12.8 $Y=2.4 $X2=0 $Y2=0
cc_1000 N_A_2013_409#_M1023_g N_Q_c_1946_n 5.92753e-19 $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_1001 N_A_2013_409#_M1032_g N_Q_c_1946_n 0.00800161f $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1002 N_A_2013_409#_M1038_g N_Q_c_1946_n 3.97481e-19 $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1003 N_A_2013_409#_M1023_g N_Q_c_1947_n 6.59139e-19 $X=12.025 $Y=0.74 $X2=0
+ $Y2=0
cc_1004 N_A_2013_409#_M1032_g N_Q_c_1947_n 0.00385048f $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1005 N_A_2013_409#_M1038_g N_Q_c_1947_n 0.00355386f $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1006 N_A_2013_409#_M1032_g N_Q_c_1948_n 7.39274e-19 $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1007 N_A_2013_409#_M1038_g N_Q_c_1948_n 6.05444e-19 $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1008 N_A_2013_409#_M1028_g Q 0.0109106f $X=12.35 $Y=2.4 $X2=0 $Y2=0
cc_1009 N_A_2013_409#_M1032_g Q 0.0055056f $X=12.525 $Y=0.74 $X2=0 $Y2=0
cc_1010 N_A_2013_409#_M1029_g Q 0.0241643f $X=12.8 $Y=2.4 $X2=0 $Y2=0
cc_1011 N_A_2013_409#_M1038_g Q 0.0162652f $X=12.955 $Y=0.74 $X2=0 $Y2=0
cc_1012 N_A_2013_409#_c_1540_n Q 0.0167026f $X=12.075 $Y=1.465 $X2=0 $Y2=0
cc_1013 N_A_2013_409#_c_1543_n Q 0.0236847f $X=12.8 $Y=1.48 $X2=0 $Y2=0
cc_1014 N_A_2013_409#_c_1537_n N_VGND_c_2018_n 0.00116291f $X=10.56 $Y=1.545
+ $X2=0 $Y2=0
cc_1015 N_A_2013_409#_c_1538_n N_VGND_c_2018_n 0.0146779f $X=10.365 $Y=1.545
+ $X2=0 $Y2=0
cc_1016 N_A_2013_409#_c_1539_n N_VGND_c_2018_n 0.0308054f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1017 N_A_2013_409#_M1003_g N_VGND_c_2019_n 0.00531367f $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1018 N_A_2013_409#_c_1531_n N_VGND_c_2019_n 0.00481677f $X=11.575 $Y=1.465
+ $X2=0 $Y2=0
cc_1019 N_A_2013_409#_c_1539_n N_VGND_c_2019_n 0.0520772f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1020 N_A_2013_409#_c_1540_n N_VGND_c_2019_n 0.0247375f $X=12.075 $Y=1.465
+ $X2=0 $Y2=0
cc_1021 N_A_2013_409#_c_1542_n N_VGND_c_2019_n 5.70705e-19 $X=11.23 $Y=1.465
+ $X2=0 $Y2=0
cc_1022 N_A_2013_409#_M1003_g N_VGND_c_2020_n 4.65028e-19 $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1023 N_A_2013_409#_M1023_g N_VGND_c_2020_n 0.00807752f $X=12.025 $Y=0.74
+ $X2=0 $Y2=0
cc_1024 N_A_2013_409#_M1032_g N_VGND_c_2020_n 0.00355746f $X=12.525 $Y=0.74
+ $X2=0 $Y2=0
cc_1025 N_A_2013_409#_M1032_g N_VGND_c_2022_n 5.9507e-19 $X=12.525 $Y=0.74 $X2=0
+ $Y2=0
cc_1026 N_A_2013_409#_M1038_g N_VGND_c_2022_n 0.0138049f $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1027 N_A_2013_409#_c_1539_n N_VGND_c_2030_n 0.0145639f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1028 N_A_2013_409#_M1003_g N_VGND_c_2031_n 0.00461464f $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1029 N_A_2013_409#_M1023_g N_VGND_c_2031_n 0.00398535f $X=12.025 $Y=0.74
+ $X2=0 $Y2=0
cc_1030 N_A_2013_409#_M1032_g N_VGND_c_2032_n 0.00434272f $X=12.525 $Y=0.74
+ $X2=0 $Y2=0
cc_1031 N_A_2013_409#_M1038_g N_VGND_c_2032_n 0.00383152f $X=12.955 $Y=0.74
+ $X2=0 $Y2=0
cc_1032 N_A_2013_409#_M1003_g N_VGND_c_2038_n 0.00913308f $X=11.5 $Y=0.74 $X2=0
+ $Y2=0
cc_1033 N_A_2013_409#_M1023_g N_VGND_c_2038_n 0.00788407f $X=12.025 $Y=0.74
+ $X2=0 $Y2=0
cc_1034 N_A_2013_409#_M1032_g N_VGND_c_2038_n 0.00820718f $X=12.525 $Y=0.74
+ $X2=0 $Y2=0
cc_1035 N_A_2013_409#_M1038_g N_VGND_c_2038_n 0.0075754f $X=12.955 $Y=0.74 $X2=0
+ $Y2=0
cc_1036 N_A_2013_409#_c_1539_n N_VGND_c_2038_n 0.0119984f $X=10.725 $Y=0.515
+ $X2=0 $Y2=0
cc_1037 N_VPWR_c_1654_n N_A_37_78#_c_1829_n 0.0126913f $X=0.275 $Y=2.75 $X2=0
+ $Y2=0
cc_1038 N_VPWR_c_1655_n N_A_37_78#_c_1829_n 0.0101517f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_1039 N_VPWR_c_1671_n N_A_37_78#_c_1829_n 0.0121689f $X=1.01 $Y=3.33 $X2=0
+ $Y2=0
cc_1040 N_VPWR_c_1652_n N_A_37_78#_c_1829_n 0.010069f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1041 N_VPWR_M1035_d N_A_37_78#_c_1831_n 0.00231422f $X=1.04 $Y=2.54 $X2=0
+ $Y2=0
cc_1042 N_VPWR_M1010_d N_A_37_78#_c_1831_n 0.00430061f $X=2.035 $Y=1.975 $X2=0
+ $Y2=0
cc_1043 N_VPWR_c_1655_n N_A_37_78#_c_1831_n 0.0207649f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_1044 N_VPWR_c_1656_n N_A_37_78#_c_1831_n 0.0165487f $X=2.17 $Y=2.815 $X2=0
+ $Y2=0
cc_1045 N_VPWR_c_1652_n N_A_37_78#_c_1831_n 0.0526056f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1046 N_VPWR_c_1654_n N_A_37_78#_c_1834_n 0.00364316f $X=0.275 $Y=2.75 $X2=0
+ $Y2=0
cc_1047 N_VPWR_c_1671_n N_A_37_78#_c_1834_n 4.9563e-19 $X=1.01 $Y=3.33 $X2=0
+ $Y2=0
cc_1048 N_VPWR_c_1652_n N_A_37_78#_c_1834_n 0.00110836f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1049 N_VPWR_c_1673_n N_A_37_78#_c_1835_n 0.00735065f $X=4.4 $Y=3.33 $X2=0
+ $Y2=0
cc_1050 N_VPWR_c_1652_n N_A_37_78#_c_1835_n 0.00897587f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1051 N_VPWR_c_1661_n N_Q_c_1950_n 0.0366243f $X=10.7 $Y=2.19 $X2=0 $Y2=0
cc_1052 N_VPWR_c_1662_n N_Q_c_1950_n 0.0324053f $X=12.12 $Y=2.305 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1675_n N_Q_c_1950_n 0.014549f $X=11.535 $Y=3.33 $X2=0 $Y2=0
cc_1054 N_VPWR_c_1652_n N_Q_c_1950_n 0.0119743f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1055 N_VPWR_M1021_s N_Q_c_1951_n 0.00945662f $X=11.515 $Y=1.84 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1662_n N_Q_c_1951_n 0.0513372f $X=12.12 $Y=2.305 $X2=0 $Y2=0
cc_1057 N_VPWR_c_1662_n N_Q_c_1953_n 0.0324053f $X=12.12 $Y=2.305 $X2=0 $Y2=0
cc_1058 N_VPWR_c_1664_n N_Q_c_1953_n 0.0386506f $X=13.075 $Y=2.115 $X2=0 $Y2=0
cc_1059 N_VPWR_c_1676_n N_Q_c_1953_n 0.0144623f $X=12.91 $Y=3.33 $X2=0 $Y2=0
cc_1060 N_VPWR_c_1652_n N_Q_c_1953_n 0.0118344f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1061 N_VPWR_c_1664_n Q 0.0279131f $X=13.075 $Y=2.115 $X2=0 $Y2=0
cc_1062 N_A_37_78#_c_1822_n A_124_78# 0.00236678f $X=0.685 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_1063 N_A_37_78#_c_1822_n N_VGND_c_2015_n 0.00131521f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_1064 N_A_37_78#_c_1828_n N_VGND_c_2015_n 0.00434714f $X=0.33 $Y=0.6 $X2=0
+ $Y2=0
cc_1065 N_A_37_78#_c_1822_n N_VGND_c_2023_n 0.00520932f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_1066 N_A_37_78#_c_1828_n N_VGND_c_2023_n 0.0131067f $X=0.33 $Y=0.6 $X2=0
+ $Y2=0
cc_1067 N_A_37_78#_c_1822_n N_VGND_c_2038_n 0.0102476f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_1068 N_A_37_78#_c_1828_n N_VGND_c_2038_n 0.0117869f $X=0.33 $Y=0.6 $X2=0
+ $Y2=0
cc_1069 N_Q_c_1945_n N_VGND_M1023_d 0.00253871f $X=12.575 $Y=1.005 $X2=0 $Y2=0
cc_1070 N_Q_c_1943_n N_VGND_c_2019_n 0.00156718f $X=11.752 $Y=0.88 $X2=0 $Y2=0
cc_1071 N_Q_c_1944_n N_VGND_c_2019_n 3.09414e-19 $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1072 N_Q_c_1944_n N_VGND_c_2020_n 0.0130802f $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1073 N_Q_c_1945_n N_VGND_c_2020_n 0.0211572f $X=12.575 $Y=1.005 $X2=0 $Y2=0
cc_1074 N_Q_c_1946_n N_VGND_c_2020_n 0.0137341f $X=12.74 $Y=0.515 $X2=0 $Y2=0
cc_1075 N_Q_c_1946_n N_VGND_c_2022_n 0.0197239f $X=12.74 $Y=0.515 $X2=0 $Y2=0
cc_1076 Q N_VGND_c_2022_n 0.0250286f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_1077 N_Q_c_1944_n N_VGND_c_2031_n 0.0131726f $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1078 N_Q_c_1946_n N_VGND_c_2032_n 0.0109942f $X=12.74 $Y=0.515 $X2=0 $Y2=0
cc_1079 N_Q_c_1944_n N_VGND_c_2038_n 0.0114552f $X=11.76 $Y=0.53 $X2=0 $Y2=0
cc_1080 N_Q_c_1946_n N_VGND_c_2038_n 0.00904371f $X=12.74 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__clkbuf_8.spice
* Created: Wed Sep  2 12:00:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkbuf_8.pex.spice"
.subckt sky130_fd_sc_ms__clkbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_M1012_g N_A_128_74#_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.3
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_128_74#_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.08295 AS=0.0588 PD=0.815 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75004 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1015_d N_A_128_74#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.08295 AS=0.06405 PD=0.815 PS=0.725 NRD=12.852 NRS=7.14 M=1 R=2.8
+ SA=75001.3 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_128_74#_M1001_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.06405 PD=0.84 PS=0.725 NRD=19.992 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1001_d N_A_128_74#_M1006_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.0588 PD=0.84 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_128_74#_M1007_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1007_d N_A_128_74#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.1 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_128_74#_M1013_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75003.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1013_d N_A_128_74#_M1017_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75004.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_128_74#_M1019_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_128_74#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.364 AS=0.154 PD=2.89 PS=1.395 NRD=7.0329 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_128_74#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.154 PD=1.49 PS=1.395 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90004 A=0.2016 P=2.6 MULT=1
MM1002 N_X_M1002_d N_A_128_74#_M1002_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.2
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1003 N_X_M1002_d N_A_128_74#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.7
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1005_d N_A_128_74#_M1005_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1005_d N_A_128_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.6
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1009_d N_A_128_74#_M1009_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1009_d N_A_128_74#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.5
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1014 N_X_M1014_d N_A_128_74#_M1014_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.1792 PD=1.405 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1018 N_X_M1014_d N_A_128_74#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.3136 PD=1.405 PS=2.8 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90004.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ms__clkbuf_8.pxi.spice"
*
.ends
*
*

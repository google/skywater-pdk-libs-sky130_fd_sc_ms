* File: sky130_fd_sc_ms__ha_4.spice
* Created: Fri Aug 28 17:37:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__ha_4.pex.spice"
.subckt sky130_fd_sc_ms__ha_4  VNB VPB B A VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1013 N_A_27_125#_M1013_d N_A_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1022 N_A_27_125#_M1022_d N_A_M1022_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_27_125#_M1022_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1002_d N_B_M1007_g N_A_27_125#_M1007_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0992 PD=0.92 PS=0.95 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_297_392#_M1023_d N_A_435_99#_M1023_g N_A_27_125#_M1007_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1024 AS=0.0992 PD=0.96 PS=0.95 NRD=7.488 NRS=5.616 M=1
+ R=4.26667 SA=75002 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1028 N_A_297_392#_M1023_d N_A_435_99#_M1028_g N_A_27_125#_M1028_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1024 AS=0.2144 PD=0.96 PS=1.95 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75002.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_A_435_99#_M1000_d N_B_M1000_g N_A_707_119#_M1000_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1856 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_435_99#_M1000_d N_B_M1003_g N_A_707_119#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_707_119#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1004_d N_A_M1011_g N_A_707_119#_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.176 PD=0.99 PS=1.83 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A_435_99#_M1010_g N_COUT_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_435_99#_M1012_g N_COUT_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1012_d N_A_435_99#_M1032_g N_COUT_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_A_435_99#_M1033_g N_COUT_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1033_d N_A_297_392#_M1005_g N_SUM_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_297_392#_M1015_g N_SUM_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1015_d N_A_297_392#_M1026_g N_SUM_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.14985 PD=1.09 PS=1.145 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1030_d N_A_297_392#_M1030_g N_SUM_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.14985 PD=2.05 PS=1.145 NRD=0 NRS=8.916 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_27_392#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1016_d N_A_M1017_g N_A_27_392#_M1017_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1019 N_A_297_392#_M1019_d N_B_M1019_g N_A_27_392#_M1017_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1021 N_A_297_392#_M1019_d N_B_M1021_g N_A_27_392#_M1021_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_297_392#_M1001_d N_A_435_99#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2268 PD=1.11 PS=2.22 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90005.5 A=0.1512 P=2.04 MULT=1
MM1006 N_A_297_392#_M1001_d N_A_435_99#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.1134 PD=1.11 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.6 SB=90005.1 A=0.1512 P=2.04 MULT=1
MM1008 N_A_435_99#_M1008_d N_B_M1008_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=0.84
+ AD=0.209937 AS=0.1134 PD=1.55 PS=1.11 NRD=17.5724 NRS=0 M=1 R=4.66667
+ SA=90001.1 SB=90004.6 A=0.1512 P=2.04 MULT=1
MM1025 N_A_435_99#_M1008_d N_B_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=0.84
+ AD=0.209937 AS=0.1134 PD=1.55 PS=1.11 NRD=45.704 NRS=0 M=1 R=4.66667
+ SA=90001.4 SB=90004.2 A=0.1512 P=2.04 MULT=1
MM1029 N_A_435_99#_M1029_d N_A_M1029_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=0.84
+ AD=0.163275 AS=0.1134 PD=1.395 PS=1.11 NRD=32.6823 NRS=0 M=1 R=4.66667
+ SA=90001.9 SB=90003.7 A=0.1512 P=2.04 MULT=1
MM1034 N_A_435_99#_M1029_d N_A_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.18 W=0.84
+ AD=0.163275 AS=0.2214 PD=1.395 PS=1.37143 NRD=0 NRS=48.8954 M=1 R=4.66667
+ SA=90002 SB=90004.4 A=0.1512 P=2.04 MULT=1
MM1009 N_COUT_M1009_d N_A_435_99#_M1009_g N_VPWR_M1034_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2408 AS=0.2952 PD=1.55 PS=1.82857 NRD=26.3783 NRS=10.5395 M=1
+ R=6.22222 SA=90002.1 SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1014 N_COUT_M1009_d N_A_435_99#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2408 AS=0.1512 PD=1.55 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.7 SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1018 N_COUT_M1018_d N_A_435_99#_M1018_g N_VPWR_M1014_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.2 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1020 N_COUT_M1018_d N_A_435_99#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.6 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1024 N_SUM_M1024_d N_A_297_392#_M1024_g N_VPWR_M1020_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.1 SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1027 N_SUM_M1024_d N_A_297_392#_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.5 SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1031 N_SUM_M1031_d N_A_297_392#_M1031_g N_VPWR_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.1512 PD=1.65 PS=1.39 NRD=25.4918 NRS=0 M=1 R=6.22222
+ SA=90005 SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1035 N_SUM_M1031_d N_A_297_392#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.3136 PD=1.65 PS=2.8 NRD=18.4589 NRS=0 M=1 R=6.22222
+ SA=90005.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.5501 P=24.79
c_106 VNB 0 2.61855e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__ha_4.pxi.spice"
*
.ends
*
*

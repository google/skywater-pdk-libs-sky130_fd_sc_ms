* File: sky130_fd_sc_ms__o41a_4.pex.spice
* Created: Wed Sep  2 12:27:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O41A_4%A_110_48# 1 2 3 12 16 20 24 28 32 36 40 42 50
+ 51 56 60 64 75
c131 56 0 2.7959e-19 $X=3.19 $Y=0.765
c132 50 0 1.29575e-19 $X=2.945 $Y=1.6
r133 72 73 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.735 $Y=1.435
+ $X2=1.985 $Y2=1.435
r134 71 72 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.555 $Y=1.435
+ $X2=1.735 $Y2=1.435
r135 70 71 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.285 $Y=1.435
+ $X2=1.555 $Y2=1.435
r136 69 70 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.055 $Y=1.435
+ $X2=1.285 $Y2=1.435
r137 68 69 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.835 $Y=1.435
+ $X2=1.055 $Y2=1.435
r138 58 64 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=2.035
+ $X2=2.945 $Y2=2.035
r139 58 60 114.171 $w=1.68e-07 $l=1.75e-06 $layer=LI1_cond $X=3.11 $Y=2.035
+ $X2=4.86 $Y2=2.035
r140 54 62 15.2248 $w=3.31e-07 $l=4.08448e-07 $layer=LI1_cond $X=3.19 $Y=1.1
+ $X2=3.027 $Y2=1.435
r141 54 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.19 $Y=1.1
+ $X2=3.19 $Y2=0.765
r142 51 64 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=1.95
+ $X2=2.945 $Y2=2.035
r143 50 62 6.08157 $w=3.31e-07 $l=2.01879e-07 $layer=LI1_cond $X=2.945 $Y=1.6
+ $X2=3.027 $Y2=1.435
r144 50 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.945 $Y=1.6
+ $X2=2.945 $Y2=1.95
r145 49 75 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.11 $Y=1.435
+ $X2=2.185 $Y2=1.435
r146 49 73 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.11 $Y=1.435
+ $X2=1.985 $Y2=1.435
r147 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.11
+ $Y=1.435 $X2=2.11 $Y2=1.435
r148 45 68 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=0.75 $Y=1.435
+ $X2=0.835 $Y2=1.435
r149 45 65 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.75 $Y=1.435
+ $X2=0.625 $Y2=1.435
r150 44 48 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=0.75 $Y=1.435
+ $X2=2.11 $Y2=1.435
r151 44 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.75
+ $Y=1.435 $X2=0.75 $Y2=1.435
r152 42 62 0.734941 $w=3.3e-07 $l=2.47e-07 $layer=LI1_cond $X=2.78 $Y=1.435
+ $X2=3.027 $Y2=1.435
r153 42 48 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=2.78 $Y=1.435
+ $X2=2.11 $Y2=1.435
r154 38 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.185 $Y=1.6
+ $X2=2.185 $Y2=1.435
r155 38 40 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=2.185 $Y=1.6
+ $X2=2.185 $Y2=2.4
r156 34 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=1.27
+ $X2=1.985 $Y2=1.435
r157 34 36 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.985 $Y=1.27
+ $X2=1.985 $Y2=0.74
r158 30 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=1.6
+ $X2=1.735 $Y2=1.435
r159 30 32 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=1.735 $Y=1.6
+ $X2=1.735 $Y2=2.4
r160 26 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.555 $Y=1.27
+ $X2=1.555 $Y2=1.435
r161 26 28 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.555 $Y=1.27
+ $X2=1.555 $Y2=0.74
r162 22 70 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.6
+ $X2=1.285 $Y2=1.435
r163 22 24 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=1.285 $Y=1.6
+ $X2=1.285 $Y2=2.4
r164 18 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.27
+ $X2=1.055 $Y2=1.435
r165 18 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.055 $Y=1.27
+ $X2=1.055 $Y2=0.74
r166 14 68 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=1.6
+ $X2=0.835 $Y2=1.435
r167 14 16 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=0.835 $Y=1.6
+ $X2=0.835 $Y2=2.4
r168 10 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.27
+ $X2=0.625 $Y2=1.435
r169 10 12 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.625 $Y=1.27
+ $X2=0.625 $Y2=0.74
r170 3 60 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.84 $X2=4.86 $Y2=2.035
r171 2 64 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.93 $X2=2.945 $Y2=2.075
r172 1 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.05
+ $Y=0.62 $X2=3.19 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%B1 3 7 11 15 17 18 24
c55 18 0 9.69802e-20 $X=4.08 $Y=1.665
c56 15 0 2.69757e-19 $X=3.405 $Y=0.94
c57 7 0 1.93825e-19 $X=2.975 $Y=0.94
c58 3 0 1.29575e-19 $X=2.72 $Y=2.35
r59 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.605 $X2=3.445 $Y2=1.605
r60 24 26 7.80567 $w=2.47e-07 $l=4e-08 $layer=POLY_cond $X=3.405 $Y=1.605
+ $X2=3.445 $Y2=1.605
r61 23 24 45.8583 $w=2.47e-07 $l=2.35e-07 $layer=POLY_cond $X=3.17 $Y=1.605
+ $X2=3.405 $Y2=1.605
r62 17 18 16.2698 $w=3.38e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.61 $X2=4.08
+ $Y2=1.61
r63 17 27 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=1.61
+ $X2=3.445 $Y2=1.61
r64 13 24 14.4406 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.44
+ $X2=3.405 $Y2=1.605
r65 13 15 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.405 $Y=1.44
+ $X2=3.405 $Y2=0.94
r66 9 23 10.2394 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.77
+ $X2=3.17 $Y2=1.605
r67 9 11 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.17 $Y=1.77 $X2=3.17
+ $Y2=2.35
r68 5 23 38.0526 $w=2.47e-07 $l=2.64953e-07 $layer=POLY_cond $X=2.975 $Y=1.44
+ $X2=3.17 $Y2=1.605
r69 5 7 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.975 $Y=1.44 $X2=2.975
+ $Y2=0.94
r70 1 5 49.7611 $w=2.47e-07 $l=3.21364e-07 $layer=POLY_cond $X=2.72 $Y=1.59
+ $X2=2.975 $Y2=1.44
r71 1 3 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=2.72 $Y=1.59 $X2=2.72
+ $Y2=2.35
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A4 3 5 7 10 12 14 15 16 26
c49 12 0 1.44963e-19 $X=5.105 $Y=1.35
c50 3 0 9.69802e-20 $X=4.63 $Y=2.4
r51 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.09 $Y=1.515
+ $X2=5.105 $Y2=1.515
r52 23 25 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.015 $Y=1.515
+ $X2=5.09 $Y2=1.515
r53 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.015
+ $Y=1.515 $X2=5.015 $Y2=1.515
r54 21 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.675 $Y=1.515
+ $X2=5.015 $Y2=1.515
r55 19 21 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=4.63 $Y=1.515
+ $X2=4.675 $Y2=1.515
r56 16 24 0.81158 $w=3.53e-07 $l=2.5e-08 $layer=LI1_cond $X=5.04 $Y=1.602
+ $X2=5.015 $Y2=1.602
r57 15 24 14.7707 $w=3.53e-07 $l=4.55e-07 $layer=LI1_cond $X=4.56 $Y=1.602
+ $X2=5.015 $Y2=1.602
r58 12 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=1.35
+ $X2=5.105 $Y2=1.515
r59 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.105 $Y=1.35
+ $X2=5.105 $Y2=0.92
r60 8 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.68
+ $X2=5.09 $Y2=1.515
r61 8 10 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.09 $Y=1.68 $X2=5.09
+ $Y2=2.4
r62 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.35
+ $X2=4.675 $Y2=1.515
r63 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.675 $Y=1.35
+ $X2=4.675 $Y2=0.92
r64 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=1.68
+ $X2=4.63 $Y2=1.515
r65 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.63 $Y=1.68 $X2=4.63
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A3 4 5 7 9 11 13 18 24 26 30
c74 30 0 1.29962e-19 $X=4.04 $Y=0.345
c75 18 0 1.4317e-19 $X=5.535 $Y=0.92
r76 29 31 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=4.027 $Y=0.345
+ $X2=4.027 $Y2=0.51
r77 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.04
+ $Y=0.345 $X2=4.04 $Y2=0.345
r78 26 29 26.0075 $w=3.55e-07 $l=1.6e-07 $layer=POLY_cond $X=4.027 $Y=0.185
+ $X2=4.027 $Y2=0.345
r79 24 30 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.04 $Y=0.555
+ $X2=4.04 $Y2=0.345
r80 18 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.535 $Y=0.92
+ $X2=5.535 $Y2=1.315
r81 15 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.535 $Y=0.26
+ $X2=5.535 $Y2=0.92
r82 11 23 36.2738 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.54 $Y=1.405 $X2=5.54
+ $Y2=1.315
r83 11 13 386.766 $w=1.8e-07 $l=9.95e-07 $layer=POLY_cond $X=5.54 $Y=1.405
+ $X2=5.54 $Y2=2.4
r84 10 26 22.9692 $w=1.5e-07 $l=1.78e-07 $layer=POLY_cond $X=4.205 $Y=0.185
+ $X2=4.027 $Y2=0.185
r85 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.46 $Y=0.185
+ $X2=5.535 $Y2=0.26
r86 9 10 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=5.46 $Y=0.185
+ $X2=4.205 $Y2=0.185
r87 5 19 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.18 $Y=1.41
+ $X2=3.925 $Y2=1.41
r88 5 7 355.669 $w=1.8e-07 $l=9.15e-07 $layer=POLY_cond $X=4.18 $Y=1.485
+ $X2=4.18 $Y2=2.4
r89 4 31 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.925 $Y=0.94
+ $X2=3.925 $Y2=0.51
r90 2 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=1.335
+ $X2=3.925 $Y2=1.41
r91 2 4 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.925 $Y=1.335
+ $X2=3.925 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A1 1 3 6 8 10 13 15 16 24
c48 13 0 1.72297e-19 $X=6.93 $Y=2.4
c49 8 0 1.74935e-19 $X=6.835 $Y=1.35
r50 22 24 54.4452 $w=3.01e-07 $l=3.4e-07 $layer=POLY_cond $X=6.495 $Y=1.515
+ $X2=6.835 $Y2=1.515
r51 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.495
+ $Y=1.515 $X2=6.495 $Y2=1.515
r52 20 22 8.80731 $w=3.01e-07 $l=5.5e-08 $layer=POLY_cond $X=6.44 $Y=1.515
+ $X2=6.495 $Y2=1.515
r53 19 20 5.60465 $w=3.01e-07 $l=3.5e-08 $layer=POLY_cond $X=6.405 $Y=1.515
+ $X2=6.44 $Y2=1.515
r54 16 23 14.8857 $w=3.58e-07 $l=4.65e-07 $layer=LI1_cond $X=6.96 $Y=1.6
+ $X2=6.495 $Y2=1.6
r55 15 23 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=6.48 $Y=1.6
+ $X2=6.495 $Y2=1.6
r56 11 24 15.2126 $w=3.01e-07 $l=2.07123e-07 $layer=POLY_cond $X=6.93 $Y=1.68
+ $X2=6.835 $Y2=1.515
r57 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.93 $Y=1.68
+ $X2=6.93 $Y2=2.4
r58 8 24 19.0468 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.835 $Y=1.35
+ $X2=6.835 $Y2=1.515
r59 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.835 $Y=1.35
+ $X2=6.835 $Y2=0.92
r60 4 20 14.7967 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.44 $Y=1.68
+ $X2=6.44 $Y2=1.515
r61 4 6 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.44 $Y=1.68 $X2=6.44
+ $Y2=2.4
r62 1 19 19.0468 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.405 $Y=1.35
+ $X2=6.405 $Y2=1.515
r63 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.405 $Y=1.35
+ $X2=6.405 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A2 4 5 7 9 10 14 17 21 22
c63 22 0 2.99718e-20 $X=7.92 $Y=0.555
c64 4 0 3.02049e-19 $X=5.975 $Y=0.92
r65 27 29 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.447 $Y=0.34
+ $X2=7.447 $Y2=0.505
r66 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.47
+ $Y=0.34 $X2=7.47 $Y2=0.34
r67 22 28 21.2791 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=7.92 $Y=0.462
+ $X2=7.47 $Y2=0.462
r68 20 21 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.39 $Y=1.33
+ $X2=7.39 $Y2=1.48
r69 17 21 357.613 $w=1.8e-07 $l=9.2e-07 $layer=POLY_cond $X=7.43 $Y=2.4 $X2=7.43
+ $Y2=1.48
r70 14 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.335 $Y=0.935
+ $X2=7.335 $Y2=1.33
r71 14 29 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.335 $Y=0.935
+ $X2=7.335 $Y2=0.505
r72 9 27 22.9877 $w=3.75e-07 $l=1.55e-07 $layer=POLY_cond $X=7.447 $Y=0.185
+ $X2=7.447 $Y2=0.34
r73 9 10 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=7.26 $Y=0.185
+ $X2=6.05 $Y2=0.185
r74 5 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.99 $Y=1.405 $X2=5.99
+ $Y2=1.315
r75 5 7 386.766 $w=1.8e-07 $l=9.95e-07 $layer=POLY_cond $X=5.99 $Y=1.405
+ $X2=5.99 $Y2=2.4
r76 4 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.975 $Y=0.92
+ $X2=5.975 $Y2=1.315
r77 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.975 $Y=0.26
+ $X2=6.05 $Y2=0.185
r78 1 4 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.975 $Y=0.26
+ $X2=5.975 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 46 47 49 50 51 76 77
r97 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r98 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r99 73 76 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33 $X2=7.92
+ $Y2=3.33
r100 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r101 71 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 70 71 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r103 67 70 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 67 68 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 65 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r106 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r107 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 51 71 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 49 70 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.58 $Y=3.33 $X2=6.48
+ $Y2=3.33
r116 49 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.725 $Y2=3.33
r117 48 73 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.87 $Y=3.33 $X2=6.96
+ $Y2=3.33
r118 48 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.87 $Y=3.33
+ $X2=6.725 $Y2=3.33
r119 46 64 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.31 $Y=3.33
+ $X2=3.12 $Y2=3.33
r120 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.31 $Y=3.33
+ $X2=3.435 $Y2=3.33
r121 45 67 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.56 $Y=3.33 $X2=3.6
+ $Y2=3.33
r122 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=3.33
+ $X2=3.435 $Y2=3.33
r123 43 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r124 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.45 $Y2=3.33
r125 42 64 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=2.45 $Y2=3.33
r127 40 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.425 $Y=3.33
+ $X2=1.51 $Y2=3.33
r129 39 61 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.51 $Y2=3.33
r131 37 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.61 $Y2=3.33
r133 36 58 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.695 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.33
+ $X2=0.61 $Y2=3.33
r135 32 50 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.725 $Y=3.245
+ $X2=6.725 $Y2=3.33
r136 32 34 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=6.725 $Y=3.245
+ $X2=6.725 $Y2=2.815
r137 28 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.435 $Y=3.245
+ $X2=3.435 $Y2=3.33
r138 28 30 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=3.435 $Y=3.245
+ $X2=3.435 $Y2=2.54
r139 24 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=3.33
r140 24 26 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=2.075
r141 20 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=3.245
+ $X2=1.51 $Y2=3.33
r142 20 22 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.51 $Y=3.245
+ $X2=1.51 $Y2=2.275
r143 16 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=3.245
+ $X2=0.61 $Y2=3.33
r144 16 18 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.61 $Y=3.245
+ $X2=0.61 $Y2=2.275
r145 5 34 600 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=6.53
+ $Y=1.84 $X2=6.685 $Y2=2.815
r146 4 30 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.93 $X2=3.395 $Y2=2.54
r147 3 26 300 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=1.84 $X2=2.41 $Y2=2.075
r148 2 22 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=1.375
+ $Y=1.84 $X2=1.51 $Y2=2.275
r149 1 18 300 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=2 $X=0.465
+ $Y=1.84 $X2=0.61 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%X 1 2 3 4 14 15 16 17 21 25 29 31 35 39 44 45
+ 46 47 48 49
c79 14 0 1.60655e-19 $X=0.21 $Y=1.77
r80 48 49 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.775
r81 47 48 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r82 43 47 4.76009 $w=2.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.24 $Y=1.94
+ $X2=0.24 $Y2=2.035
r83 43 44 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.94 $X2=0.24
+ $Y2=1.855
r84 39 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.96 $Y=1.985
+ $X2=1.96 $Y2=2.815
r85 37 39 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.96 $Y=1.94
+ $X2=1.96 $Y2=1.985
r86 33 35 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=1.73 $Y=0.93
+ $X2=1.73 $Y2=0.515
r87 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=1.855
+ $X2=1.06 $Y2=1.855
r88 31 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=1.855
+ $X2=1.96 $Y2=1.94
r89 31 32 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.795 $Y=1.855
+ $X2=1.225 $Y2=1.855
r90 30 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.925 $Y=1.015
+ $X2=0.8 $Y2=1.015
r91 29 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.605 $Y=1.015
+ $X2=1.73 $Y2=0.93
r92 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=1.015
+ $X2=0.925 $Y2=1.015
r93 25 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.06 $Y=1.985
+ $X2=1.06 $Y2=2.815
r94 23 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=1.94 $X2=1.06
+ $Y2=1.855
r95 23 25 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.06 $Y=1.94
+ $X2=1.06 $Y2=1.985
r96 19 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.93
+ $X2=0.8 $Y2=1.015
r97 19 21 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=0.8 $Y=0.93 $X2=0.8
+ $Y2=0.515
r98 18 44 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.855
+ $X2=0.24 $Y2=1.855
r99 17 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.855
+ $X2=1.06 $Y2=1.855
r100 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.895 $Y=1.855
+ $X2=0.355 $Y2=1.855
r101 15 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.675 $Y=1.015
+ $X2=0.8 $Y2=1.015
r102 15 16 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.675 $Y=1.015
+ $X2=0.295 $Y2=1.015
r103 14 44 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.21 $Y=1.77
+ $X2=0.24 $Y2=1.855
r104 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.21 $Y=1.1
+ $X2=0.295 $Y2=1.015
r105 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.21 $Y=1.1
+ $X2=0.21 $Y2=1.77
r106 4 41 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.84 $X2=1.96 $Y2=2.815
r107 4 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.84 $X2=1.96 $Y2=1.985
r108 3 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.925
+ $Y=1.84 $X2=1.06 $Y2=2.815
r109 3 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.925
+ $Y=1.84 $X2=1.06 $Y2=1.985
r110 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.63
+ $Y=0.37 $X2=1.77 $Y2=0.515
r111 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.7
+ $Y=0.37 $X2=0.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A_762_368# 1 2 3 12 14 18 20 22 25 29
c51 14 0 1.65567e-19 $X=5.765 $Y=2.12
r52 20 31 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.705 $Y=2.12
+ $X2=7.705 $Y2=1.97
r53 20 22 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.705 $Y=2.12
+ $X2=7.705 $Y2=2.4
r54 19 27 3.40825 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=5.85 $Y=2.035
+ $X2=5.765 $Y2=1.97
r55 18 31 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=7.54 $Y=2.035
+ $X2=7.705 $Y2=1.97
r56 18 19 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=7.54 $Y=2.035
+ $X2=5.85 $Y2=2.035
r57 15 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.765 $Y=2.29
+ $X2=5.765 $Y2=2.375
r58 14 27 3.40825 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.765 $Y=2.12
+ $X2=5.765 $Y2=1.97
r59 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.765 $Y=2.12
+ $X2=5.765 $Y2=2.29
r60 13 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.04 $Y=2.375
+ $X2=3.915 $Y2=2.375
r61 12 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=2.375
+ $X2=5.765 $Y2=2.375
r62 12 13 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=5.68 $Y=2.375
+ $X2=4.04 $Y2=2.375
r63 3 31 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.52
+ $Y=1.84 $X2=7.705 $Y2=1.985
r64 3 22 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=7.52
+ $Y=1.84 $X2=7.705 $Y2=2.4
r65 2 29 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=5.63
+ $Y=1.84 $X2=5.765 $Y2=2.4
r66 2 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=1.84 $X2=5.765 $Y2=1.985
r67 1 25 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=3.81
+ $Y=1.84 $X2=3.955 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A_854_368# 1 2 11
r14 8 11 29.9635 $w=3.48e-07 $l=9.1e-07 $layer=LI1_cond $X=4.405 $Y=2.805
+ $X2=5.315 $Y2=2.805
r15 2 11 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=5.18
+ $Y=1.84 $X2=5.315 $Y2=2.805
r16 1 8 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.84 $X2=4.405 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A_1216_368# 1 2 9 14 16
c23 16 0 1.72297e-19 $X=7.205 $Y=2.455
r24 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=2.375
+ $X2=6.215 $Y2=2.375
r25 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=2.375
+ $X2=7.205 $Y2=2.375
r26 9 10 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.04 $Y=2.375
+ $X2=6.38 $Y2=2.375
r27 2 16 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=7.02
+ $Y=1.84 $X2=7.205 $Y2=2.455
r28 1 14 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.08
+ $Y=1.84 $X2=6.215 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46 50
+ 53 54 56 57 58 59 60 62 67 87 88 94 97 100
c121 1 0 1.60655e-19 $X=0.195 $Y=0.37
r122 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r123 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r124 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r126 88 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=6.96 $Y2=0
r127 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r128 85 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.135 $Y=0
+ $X2=7.01 $Y2=0
r129 85 87 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.135 $Y=0
+ $X2=7.92 $Y2=0
r130 84 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r131 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r132 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r133 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r134 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r135 74 77 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r136 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r137 72 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.2
+ $Y2=0
r138 72 74 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=0
+ $X2=2.64 $Y2=0
r139 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r140 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r141 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r142 68 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.27
+ $Y2=0
r143 68 70 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.68
+ $Y2=0
r144 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.2
+ $Y2=0
r145 67 70 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=1.68 $Y2=0
r146 66 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r147 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r148 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r149 63 91 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.252 $Y2=0
r150 63 65 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.72 $Y2=0
r151 62 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.27
+ $Y2=0
r152 62 65 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=0
+ $X2=0.72 $Y2=0
r153 60 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r154 60 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r155 60 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r156 58 83 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.025 $Y=0 $X2=6
+ $Y2=0
r157 58 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.025 $Y=0 $X2=6.15
+ $Y2=0
r158 56 80 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.04 $Y2=0
r159 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.32
+ $Y2=0
r160 55 83 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.485 $Y=0 $X2=6
+ $Y2=0
r161 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.32
+ $Y2=0
r162 53 77 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.08
+ $Y2=0
r163 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.46
+ $Y2=0
r164 52 80 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.545 $Y=0
+ $X2=5.04 $Y2=0
r165 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=0 $X2=4.46
+ $Y2=0
r166 48 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0
r167 48 50 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0.745
r168 47 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.15
+ $Y2=0
r169 46 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.885 $Y=0
+ $X2=7.01 $Y2=0
r170 46 47 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.885 $Y=0
+ $X2=6.275 $Y2=0
r171 42 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0
r172 42 44 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0.745
r173 38 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.32 $Y=0.085
+ $X2=5.32 $Y2=0
r174 38 40 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=5.32 $Y=0.085
+ $X2=5.32 $Y2=0.745
r175 34 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r176 34 36 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.75
r177 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r178 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.515
r179 26 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=0.085
+ $X2=1.27 $Y2=0
r180 26 28 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.27 $Y=0.085
+ $X2=1.27 $Y2=0.555
r181 22 91 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.252 $Y2=0
r182 22 24 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.34 $Y2=0.555
r183 7 50 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.91
+ $Y=0.6 $X2=7.05 $Y2=0.745
r184 6 44 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.05
+ $Y=0.6 $X2=6.19 $Y2=0.745
r185 5 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.6 $X2=5.32 $Y2=0.745
r186 4 36 182 $w=1.7e-07 $l=5.20961e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.62 $X2=4.46 $Y2=0.75
r187 3 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.37 $X2=2.2 $Y2=0.515
r188 2 28 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.37 $X2=1.27 $Y2=0.555
r189 1 24 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.37 $X2=0.34 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_4%A_523_124# 1 2 3 4 5 6 21 23 24 28 29 30 33
+ 35 39 41 45 47 49 52 53 54
c107 53 0 1.58878e-19 $X=5.755 $Y=1.167
c108 45 0 1.44963e-19 $X=6.62 $Y=0.745
c109 41 0 1.65567e-19 $X=6.455 $Y=1.165
c110 39 0 2.86341e-19 $X=5.755 $Y=0.745
c111 33 0 1.44963e-19 $X=4.89 $Y=0.745
c112 30 0 5.40297e-20 $X=3.705 $Y=1.17
r113 49 51 5.124 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.51 $Y=1.08 $X2=7.51
+ $Y2=0.975
r114 48 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=1.165
+ $X2=6.58 $Y2=1.165
r115 47 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.385 $Y=1.165
+ $X2=7.51 $Y2=1.08
r116 47 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.385 $Y=1.165
+ $X2=6.705 $Y2=1.165
r117 43 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=1.08
+ $X2=6.58 $Y2=1.165
r118 43 45 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.58 $Y=1.08
+ $X2=6.58 $Y2=0.745
r119 42 53 5.41628 $w=1.7e-07 $l=9.09945e-08 $layer=LI1_cond $X=5.845 $Y=1.165
+ $X2=5.755 $Y2=1.167
r120 41 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.455 $Y=1.165
+ $X2=6.58 $Y2=1.165
r121 41 42 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.455 $Y=1.165
+ $X2=5.845 $Y2=1.165
r122 37 53 1.13756 $w=1.8e-07 $l=8.7e-08 $layer=LI1_cond $X=5.755 $Y=1.08
+ $X2=5.755 $Y2=1.167
r123 37 39 20.6414 $w=1.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.755 $Y=1.08
+ $X2=5.755 $Y2=0.745
r124 36 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.975 $Y=1.17
+ $X2=4.85 $Y2=1.17
r125 35 53 5.41628 $w=1.7e-07 $l=9.14877e-08 $layer=LI1_cond $X=5.665 $Y=1.17
+ $X2=5.755 $Y2=1.167
r126 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.665 $Y=1.17
+ $X2=4.975 $Y2=1.17
r127 31 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.85 $Y=1.085
+ $X2=4.85 $Y2=1.17
r128 31 33 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.85 $Y=1.085
+ $X2=4.85 $Y2=0.745
r129 29 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.725 $Y=1.17
+ $X2=4.85 $Y2=1.17
r130 29 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.725 $Y=1.17
+ $X2=3.705 $Y2=1.17
r131 26 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.58 $Y=1.085
+ $X2=3.705 $Y2=1.17
r132 26 28 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=3.58 $Y=1.085
+ $X2=3.58 $Y2=0.765
r133 25 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.58 $Y=0.43
+ $X2=3.58 $Y2=0.765
r134 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.455 $Y=0.345
+ $X2=3.58 $Y2=0.43
r135 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.455 $Y=0.345
+ $X2=2.925 $Y2=0.345
r136 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.76 $Y=0.43
+ $X2=2.925 $Y2=0.345
r137 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.76 $Y=0.43
+ $X2=2.76 $Y2=0.765
r138 6 51 182 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.615 $X2=7.55 $Y2=0.975
r139 5 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.48
+ $Y=0.6 $X2=6.62 $Y2=0.745
r140 4 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.61
+ $Y=0.6 $X2=5.755 $Y2=0.745
r141 3 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.75
+ $Y=0.6 $X2=4.89 $Y2=0.745
r142 2 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.48
+ $Y=0.62 $X2=3.62 $Y2=0.765
r143 1 21 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.62 $X2=2.76 $Y2=0.765
.ends


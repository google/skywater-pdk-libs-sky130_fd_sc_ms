# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__einvp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.430000 1.780000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.756600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.980000 1.300000 5.650000 1.630000 ;
        RECT 5.405000 1.180000 5.650000 1.300000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.154700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.660000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 1.945000 1.180000 ;
        RECT 0.615000 1.950000 1.895000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.565000 2.120000 1.895000 2.735000 ;
        RECT 1.615000 0.660000 1.945000 1.010000 ;
        RECT 1.615000 1.180000 1.895000 1.950000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.255000 2.445000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 1.130000 ;
      RECT 0.115000  1.950000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.395000 3.075000 ;
      RECT 1.115000  0.425000 1.445000 0.800000 ;
      RECT 1.115000  2.290000 1.365000 2.905000 ;
      RECT 2.065000  1.640000 4.175000 1.810000 ;
      RECT 2.065000  1.810000 2.395000 2.905000 ;
      RECT 2.115000  0.425000 2.445000 1.300000 ;
      RECT 2.115000  1.300000 4.445000 1.470000 ;
      RECT 2.565000  1.980000 2.815000 3.245000 ;
      RECT 2.615000  0.085000 2.945000 1.130000 ;
      RECT 3.015000  1.810000 3.265000 2.980000 ;
      RECT 3.115000  0.350000 3.445000 1.300000 ;
      RECT 3.465000  1.980000 3.725000 3.245000 ;
      RECT 3.615000  0.085000 3.945000 1.130000 ;
      RECT 3.925000  1.810000 4.175000 2.980000 ;
      RECT 4.115000  0.350000 4.445000 1.300000 ;
      RECT 4.395000  1.640000 4.785000 1.820000 ;
      RECT 4.395000  1.820000 5.195000 2.980000 ;
      RECT 4.395000  2.980000 4.785000 2.990000 ;
      RECT 4.615000  0.350000 5.005000 1.130000 ;
      RECT 4.615000  1.130000 4.785000 1.640000 ;
      RECT 5.175000  0.085000 5.505000 1.010000 ;
      RECT 5.395000  1.820000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__einvp_4
END LIBRARY

* File: sky130_fd_sc_ms__o221a_4.pex.spice
* Created: Fri Aug 28 17:57:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O221A_4%C1 3 7 11 15 17 18 28
c45 11 0 1.44963e-19 $X=0.925 $Y=0.945
r46 27 28 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.61
+ $X2=0.955 $Y2=1.61
r47 25 27 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.725 $Y=1.61
+ $X2=0.925 $Y2=1.61
r48 23 25 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.505 $Y=1.61
+ $X2=0.725 $Y2=1.61
r49 21 23 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.61
+ $X2=0.505 $Y2=1.61
r50 18 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.61 $X2=0.725 $Y2=1.61
r51 17 18 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.612
+ $X2=0.72 $Y2=1.612
r52 13 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.775
+ $X2=0.955 $Y2=1.61
r53 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.775
+ $X2=0.955 $Y2=2.435
r54 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.445
+ $X2=0.925 $Y2=1.61
r55 9 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.925 $Y=1.445
+ $X2=0.925 $Y2=0.945
r56 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.445
+ $X2=0.495 $Y2=1.61
r57 5 7 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.495 $Y=1.445 $X2=0.495
+ $Y2=0.945
r58 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.775
+ $X2=0.505 $Y2=1.61
r59 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.775
+ $X2=0.505 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%B2 3 7 11 15 17 18 27
c47 27 0 8.30843e-20 $X=2.355 $Y=1.61
c48 18 0 1.5417e-19 $X=2.64 $Y=1.665
c49 3 0 1.70191e-19 $X=1.89 $Y=0.945
r50 25 27 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=1.61
+ $X2=2.355 $Y2=1.61
r51 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.61 $X2=2.28 $Y2=1.61
r52 23 25 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.905 $Y=1.61
+ $X2=2.28 $Y2=1.61
r53 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.89 $Y=1.61
+ $X2=1.905 $Y2=1.61
r54 18 26 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=2.64 $Y=1.612
+ $X2=2.28 $Y2=1.612
r55 17 26 4.12815 $w=3.33e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=1.612
+ $X2=2.28 $Y2=1.612
r56 13 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.445
+ $X2=2.355 $Y2=1.61
r57 13 15 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.355 $Y=1.445
+ $X2=2.355 $Y2=0.945
r58 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.775
+ $X2=2.355 $Y2=1.61
r59 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.355 $Y=1.775
+ $X2=2.355 $Y2=2.435
r60 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.775
+ $X2=1.905 $Y2=1.61
r61 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.905 $Y=1.775
+ $X2=1.905 $Y2=2.435
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.445
+ $X2=1.89 $Y2=1.61
r63 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.89 $Y=1.445 $X2=1.89
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%B1 1 3 8 9 10 13 17 22 24 25 26 27 34 35
c85 35 0 1.5417e-19 $X=3.3 $Y=1.61
c86 27 0 8.30843e-20 $X=4.08 $Y=1.665
r87 32 35 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.27 $Y=1.61 $X2=3.3
+ $Y2=1.61
r88 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.61
+ $X2=3.105 $Y2=1.61
r89 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.61 $X2=3.27 $Y2=1.61
r90 26 27 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.612
+ $X2=4.08 $Y2=1.612
r91 26 33 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=3.6 $Y=1.612
+ $X2=3.27 $Y2=1.612
r92 25 33 5.16019 $w=3.33e-07 $l=1.5e-07 $layer=LI1_cond $X=3.12 $Y=1.612
+ $X2=3.27 $Y2=1.612
r93 22 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.445
+ $X2=3.3 $Y2=1.61
r94 21 22 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=3.3 $Y=0.255
+ $X2=3.3 $Y2=1.445
r95 20 24 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.895 $Y=1.52
+ $X2=2.805 $Y2=1.52
r96 20 34 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.895 $Y=1.52
+ $X2=3.105 $Y2=1.52
r97 15 24 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.805 $Y=1.595
+ $X2=2.805 $Y2=1.52
r98 15 17 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=2.805 $Y=1.595
+ $X2=2.805 $Y2=2.435
r99 11 24 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.79 $Y=1.445
+ $X2=2.805 $Y2=1.52
r100 11 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.79 $Y=1.445
+ $X2=2.79 $Y2=0.945
r101 9 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.225 $Y=0.18
+ $X2=3.3 $Y2=0.255
r102 9 10 884.521 $w=1.5e-07 $l=1.725e-06 $layer=POLY_cond $X=3.225 $Y=0.18
+ $X2=1.5 $Y2=0.18
r103 8 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=0.945
+ $X2=1.425 $Y2=1.34
r104 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.425 $Y=0.255
+ $X2=1.5 $Y2=0.18
r105 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.425 $Y=0.255
+ $X2=1.425 $Y2=0.945
r106 1 23 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.41 $Y=1.43 $X2=1.41
+ $Y2=1.34
r107 1 3 390.653 $w=1.8e-07 $l=1.005e-06 $layer=POLY_cond $X=1.41 $Y=1.43
+ $X2=1.41 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A2 3 7 11 15 17 24
c48 17 0 2.66651e-19 $X=4.56 $Y=1.665
c49 11 0 3.38411e-20 $X=4.675 $Y=0.915
c50 7 0 6.92713e-20 $X=4.245 $Y=0.915
c51 3 0 6.40318e-20 $X=4.215 $Y=2.435
r52 24 25 2.23839 $w=3.23e-07 $l=1.5e-08 $layer=POLY_cond $X=4.675 $Y=1.61
+ $X2=4.69 $Y2=1.61
r53 22 24 21.6378 $w=3.23e-07 $l=1.45e-07 $layer=POLY_cond $X=4.53 $Y=1.61
+ $X2=4.675 $Y2=1.61
r54 20 22 42.5294 $w=3.23e-07 $l=2.85e-07 $layer=POLY_cond $X=4.245 $Y=1.61
+ $X2=4.53 $Y2=1.61
r55 19 20 4.47678 $w=3.23e-07 $l=3e-08 $layer=POLY_cond $X=4.215 $Y=1.61
+ $X2=4.245 $Y2=1.61
r56 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.61 $X2=4.53 $Y2=1.61
r57 13 25 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.775
+ $X2=4.69 $Y2=1.61
r58 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.69 $Y=1.775
+ $X2=4.69 $Y2=2.435
r59 9 24 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=1.61
r60 9 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=0.915
r61 5 20 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.445
+ $X2=4.245 $Y2=1.61
r62 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.245 $Y=1.445
+ $X2=4.245 $Y2=0.915
r63 1 19 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.215 $Y=1.775
+ $X2=4.215 $Y2=1.61
r64 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.215 $Y=1.775
+ $X2=4.215 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A1 3 8 9 10 14 17 20 21 24 25
c75 20 0 7.73759e-21 $X=3.767 $Y=1.46
c76 17 0 8.7589e-20 $X=5.19 $Y=2.435
c77 8 0 2.67289e-19 $X=3.81 $Y=0.915
c78 3 0 1.71325e-19 $X=3.74 $Y=2.435
r79 24 27 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.515
+ $X2=5.155 $Y2=1.68
r80 24 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.515
+ $X2=5.155 $Y2=1.35
r81 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.515 $X2=5.155 $Y2=1.515
r82 21 25 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=5.122 $Y=1.665
+ $X2=5.122 $Y2=1.515
r83 19 20 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.767 $Y=1.31
+ $X2=3.767 $Y2=1.46
r84 17 27 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=5.19 $Y=2.435
+ $X2=5.19 $Y2=1.68
r85 14 26 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.105 $Y=0.915
+ $X2=5.105 $Y2=1.35
r86 11 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.105 $Y=0.255
+ $X2=5.105 $Y2=0.915
r87 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.03 $Y=0.18
+ $X2=5.105 $Y2=0.255
r88 9 10 587.117 $w=1.5e-07 $l=1.145e-06 $layer=POLY_cond $X=5.03 $Y=0.18
+ $X2=3.885 $Y2=0.18
r89 8 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.81 $Y=0.915
+ $X2=3.81 $Y2=1.31
r90 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.81 $Y=0.255
+ $X2=3.885 $Y2=0.18
r91 5 8 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.81 $Y=0.255 $X2=3.81
+ $Y2=0.915
r92 3 20 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=3.74 $Y=2.435
+ $X2=3.74 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A_114_125# 1 2 3 4 13 15 18 20 22 25 29 31
+ 33 34 36 38 41 43 46 50 52 53 55 56 57 60 64 67 68 73 81 83 93
c176 83 0 6.40318e-20 $X=4.465 $Y=2.115
c177 68 0 1.22796e-19 $X=5.66 $Y=1.515
c178 46 0 1.44963e-19 $X=0.71 $Y=0.77
c179 20 0 1.46284e-19 $X=6.115 $Y=1.35
c180 18 0 1.23902e-19 $X=5.695 $Y=2.4
r181 92 93 14.8876 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.685 $Y=1.515
+ $X2=6.76 $Y2=1.515
r182 91 92 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.67 $Y=1.515
+ $X2=6.685 $Y2=1.515
r183 88 89 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.115 $Y=1.515
+ $X2=6.22 $Y2=1.515
r184 84 86 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.68 $Y=1.515
+ $X2=5.695 $Y2=1.515
r185 77 79 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.73 $Y=2.035
+ $X2=1.145 $Y2=2.035
r186 74 91 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=6.45 $Y=1.515
+ $X2=6.67 $Y2=1.515
r187 74 89 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=6.45 $Y=1.515
+ $X2=6.22 $Y2=1.515
r188 73 74 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.515 $X2=6.45 $Y2=1.515
r189 71 88 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=5.77 $Y=1.515
+ $X2=6.115 $Y2=1.515
r190 71 86 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.77 $Y=1.515
+ $X2=5.695 $Y2=1.515
r191 70 73 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.77 $Y=1.515
+ $X2=6.45 $Y2=1.515
r192 70 71 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.77
+ $Y=1.515 $X2=5.77 $Y2=1.515
r193 68 70 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.66 $Y=1.515
+ $X2=5.77 $Y2=1.515
r194 66 68 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.575 $Y=1.68
+ $X2=5.66 $Y2=1.515
r195 66 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.575 $Y=1.68
+ $X2=5.575 $Y2=1.95
r196 65 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=2.035
+ $X2=4.465 $Y2=2.035
r197 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.49 $Y=2.035
+ $X2=5.575 $Y2=1.95
r198 64 65 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=5.49 $Y=2.035
+ $X2=4.63 $Y2=2.035
r199 61 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=2.035
+ $X2=2.13 $Y2=2.035
r200 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=2.035
+ $X2=4.465 $Y2=2.035
r201 60 61 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=4.3 $Y=2.035
+ $X2=2.215 $Y2=2.035
r202 57 79 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.035
+ $X2=1.145 $Y2=2.035
r203 56 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.13 $Y2=2.035
r204 56 57 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.23 $Y2=2.035
r205 55 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.95
+ $X2=1.145 $Y2=2.035
r206 54 55 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.145 $Y=1.275
+ $X2=1.145 $Y2=1.95
r207 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=1.19
+ $X2=1.145 $Y2=1.275
r208 52 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.06 $Y=1.19
+ $X2=0.795 $Y2=1.19
r209 50 77 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=0.73 $Y=2.79
+ $X2=0.73 $Y2=2.12
r210 44 53 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.67 $Y=1.105
+ $X2=0.795 $Y2=1.19
r211 44 46 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.67 $Y=1.105
+ $X2=0.67 $Y2=0.77
r212 39 43 30.4925 $w=1.65e-07 $l=1.49057e-07 $layer=POLY_cond $X=7.175 $Y=1.625
+ $X2=7.152 $Y2=1.487
r213 39 41 301.25 $w=1.8e-07 $l=7.75e-07 $layer=POLY_cond $X=7.175 $Y=1.625
+ $X2=7.175 $Y2=2.4
r214 36 43 30.4925 $w=1.65e-07 $l=1.54396e-07 $layer=POLY_cond $X=7.115 $Y=1.35
+ $X2=7.152 $Y2=1.487
r215 36 38 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.115 $Y=1.35
+ $X2=7.115 $Y2=0.865
r216 34 43 1.63566 $w=2.75e-07 $l=1.12e-07 $layer=POLY_cond $X=7.04 $Y=1.487
+ $X2=7.152 $Y2=1.487
r217 34 93 61.0776 $w=2.75e-07 $l=2.8e-07 $layer=POLY_cond $X=7.04 $Y=1.487
+ $X2=6.76 $Y2=1.487
r218 31 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.685 $Y=1.35
+ $X2=6.685 $Y2=1.515
r219 31 33 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.685 $Y=1.35
+ $X2=6.685 $Y2=0.865
r220 27 91 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.67 $Y=1.68
+ $X2=6.67 $Y2=1.515
r221 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.67 $Y=1.68
+ $X2=6.67 $Y2=2.4
r222 23 89 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.22 $Y=1.68
+ $X2=6.22 $Y2=1.515
r223 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.22 $Y=1.68
+ $X2=6.22 $Y2=2.4
r224 20 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.35
+ $X2=6.115 $Y2=1.515
r225 20 22 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.115 $Y=1.35
+ $X2=6.115 $Y2=0.865
r226 16 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.68
+ $X2=5.695 $Y2=1.515
r227 16 18 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.695 $Y=1.68
+ $X2=5.695 $Y2=2.4
r228 13 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.68 $Y=1.35
+ $X2=5.68 $Y2=1.515
r229 13 15 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.68 $Y=1.35
+ $X2=5.68 $Y2=0.865
r230 4 83 300 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.935 $X2=4.465 $Y2=2.115
r231 3 81 300 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.935 $X2=2.13 $Y2=2.115
r232 2 77 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.935 $X2=0.73 $Y2=2.11
r233 2 50 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.935 $X2=0.73 $Y2=2.79
r234 1 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.625 $X2=0.71 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 41 43 47
+ 49 54 62 67 72 81 84 89 92 96
r95 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r96 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r97 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 85 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 84 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r101 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r102 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 76 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 76 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.61 $Y=3.33
+ $X2=6.485 $Y2=3.33
r107 73 75 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.61 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 72 95 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=7.497 $Y2=3.33
r109 72 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=6.96 $Y2=3.33
r110 71 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r111 71 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r112 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r113 68 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=3.33
+ $X2=5.465 $Y2=3.33
r114 68 70 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.63 $Y=3.33 $X2=6
+ $Y2=3.33
r115 67 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.36 $Y=3.33
+ $X2=6.485 $Y2=3.33
r116 67 70 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.36 $Y=3.33 $X2=6
+ $Y2=3.33
r117 66 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r118 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 63 84 13.8148 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.272 $Y2=3.33
r120 63 65 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 62 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.465 $Y2=3.33
r122 62 65 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 61 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r124 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 55 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.22 $Y2=3.33
r130 55 57 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r131 54 84 13.8148 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.272 $Y2=3.33
r132 54 60 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 53 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 53 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 50 78 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r137 50 52 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 49 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.22 $Y2=3.33
r139 49 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 47 66 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=5.04 $Y2=3.33
r141 47 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r142 43 46 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=7.44 $Y=2.115
+ $X2=7.44 $Y2=2.815
r143 41 95 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.497 $Y2=3.33
r144 41 46 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=3.245
+ $X2=7.44 $Y2=2.815
r145 37 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=3.33
r146 37 39 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=2.355
r147 33 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=3.33
r148 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.465 $Y=3.245
+ $X2=5.465 $Y2=2.415
r149 29 84 2.90666 $w=7.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=3.33
r150 29 31 13.2154 $w=7.13e-07 $l=7.9e-07 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=2.455
r151 25 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r152 25 27 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.455
r153 21 24 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=2.115
+ $X2=0.24 $Y2=2.795
r154 19 78 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r155 19 24 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.795
r156 6 46 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.84 $X2=7.4 $Y2=2.815
r157 6 43 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.84 $X2=7.4 $Y2=2.115
r158 5 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.31
+ $Y=1.84 $X2=6.445 $Y2=2.355
r159 4 35 300 $w=1.7e-07 $l=5.64978e-07 $layer=licon1_PDIFF $count=2 $X=5.28
+ $Y=1.935 $X2=5.465 $Y2=2.415
r160 3 31 150 $w=1.7e-07 $l=8.40714e-07 $layer=licon1_PDIFF $count=4 $X=2.895
+ $Y=1.935 $X2=3.515 $Y2=2.455
r161 2 27 300 $w=1.7e-07 $l=5.83609e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.935 $X2=1.18 $Y2=2.455
r162 1 24 400 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.795
r163 1 21 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A_300_387# 1 2 9 11 12 15
r24 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.58 $Y=2.905
+ $X2=2.58 $Y2=2.415
r25 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=2.99
+ $X2=2.58 $Y2=2.905
r26 11 12 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.415 $Y=2.99
+ $X2=1.845 $Y2=2.99
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.68 $Y=2.905
+ $X2=1.845 $Y2=2.99
r28 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.68 $Y=2.905 $X2=1.68
+ $Y2=2.415
r29 2 15 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=1.935 $X2=2.58 $Y2=2.415
r30 1 9 300 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.935 $X2=1.68 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A_766_387# 1 2 9 11 12 15
c24 11 0 1.23902e-19 $X=4.8 $Y=2.99
r25 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.965 $Y=2.905
+ $X2=4.965 $Y2=2.415
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.8 $Y=2.99
+ $X2=4.965 $Y2=2.905
r27 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.8 $Y=2.99 $X2=4.13
+ $Y2=2.99
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.965 $Y=2.905
+ $X2=4.13 $Y2=2.99
r29 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=3.965 $Y=2.905
+ $X2=3.965 $Y2=2.415
r30 2 15 300 $w=1.7e-07 $l=5.64978e-07 $layer=licon1_PDIFF $count=2 $X=4.78
+ $Y=1.935 $X2=4.965 $Y2=2.415
r31 1 9 300 $w=1.7e-07 $l=5.43323e-07 $layer=licon1_PDIFF $count=2 $X=3.83
+ $Y=1.935 $X2=3.965 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%X 1 2 3 4 15 17 19 21 22 23 27 33 37 38 40
+ 44
c68 15 0 1.46284e-19 $X=5.9 $Y=0.64
r69 41 43 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=6.95 $Y=1.935 $X2=6.95
+ $Y2=1.985
r70 39 44 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=1.665
+ $X2=7.44 $Y2=1.665
r71 38 41 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.95 $Y=1.665
+ $X2=6.95 $Y2=1.935
r72 38 40 4.31382 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.95 $Y=1.665
+ $X2=6.95 $Y2=1.55
r73 38 39 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=1.665
+ $X2=7.115 $Y2=1.665
r74 31 43 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.95 $Y=2.02
+ $X2=6.95 $Y2=1.985
r75 31 33 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=6.95 $Y=2.02
+ $X2=6.95 $Y2=2.815
r76 29 37 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.925 $Y=1.18
+ $X2=6.9 $Y2=1.095
r77 29 40 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.925 $Y=1.18
+ $X2=6.925 $Y2=1.55
r78 25 37 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.9 $Y=1.01 $X2=6.9
+ $Y2=1.095
r79 25 27 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.9 $Y=1.01 $X2=6.9
+ $Y2=0.64
r80 24 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.16 $Y=1.935
+ $X2=5.995 $Y2=1.935
r81 23 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=1.935
+ $X2=6.95 $Y2=1.935
r82 23 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.785 $Y=1.935
+ $X2=6.16 $Y2=1.935
r83 21 37 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.735 $Y=1.095
+ $X2=6.9 $Y2=1.095
r84 21 22 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.735 $Y=1.095
+ $X2=5.985 $Y2=1.095
r85 17 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=2.02
+ $X2=5.995 $Y2=1.935
r86 17 19 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=5.995 $Y=2.02
+ $X2=5.995 $Y2=2.815
r87 13 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.86 $Y=1.01
+ $X2=5.985 $Y2=1.095
r88 13 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=5.86 $Y=1.01
+ $X2=5.86 $Y2=0.64
r89 4 43 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=1.84 $X2=6.95 $Y2=1.985
r90 4 33 400 $w=1.7e-07 $l=1.06577e-06 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=1.84 $X2=6.95 $Y2=2.815
r91 3 36 400 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.995 $Y2=2.015
r92 3 19 400 $w=1.7e-07 $l=1.07488e-06 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.995 $Y2=2.815
r93 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.76
+ $Y=0.495 $X2=6.9 $Y2=0.64
r94 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.755
+ $Y=0.495 $X2=5.9 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A_27_125# 1 2 3 4 15 17 18 21 23 27 29 33 35
+ 36
c68 29 0 1.98018e-19 $X=2.84 $Y=0.37
r69 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.005 $Y=0.455
+ $X2=3.005 $Y2=0.77
r70 30 36 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.305 $Y=0.37
+ $X2=2.14 $Y2=0.36
r71 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.84 $Y=0.37
+ $X2=3.005 $Y2=0.455
r72 29 30 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.84 $Y=0.37
+ $X2=2.305 $Y2=0.37
r73 25 36 0.89609 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.14 $Y=0.455
+ $X2=2.14 $Y2=0.36
r74 25 27 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.14 $Y=0.455
+ $X2=2.14 $Y2=0.77
r75 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0.35
+ $X2=1.14 $Y2=0.35
r76 23 36 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=1.975 $Y=0.35
+ $X2=2.14 $Y2=0.36
r77 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=0.35
+ $X2=1.305 $Y2=0.35
r78 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.435
+ $X2=1.14 $Y2=0.35
r79 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.14 $Y=0.435
+ $X2=1.14 $Y2=0.77
r80 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0.35
+ $X2=1.14 $Y2=0.35
r81 17 18 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.975 $Y=0.35
+ $X2=0.365 $Y2=0.35
r82 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.435
+ $X2=0.365 $Y2=0.35
r83 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=0.435
+ $X2=0.24 $Y2=0.77
r84 4 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.625 $X2=3.005 $Y2=0.77
r85 3 27 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.625 $X2=2.14 $Y2=0.77
r86 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.625 $X2=1.14 $Y2=0.77
r87 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%A_300_125# 1 2 3 4 13 15 17 21 23 27 29 31
+ 33 38 39
c69 33 0 3.38411e-20 $X=4.89 $Y=0.755
c70 27 0 1.38543e-19 $X=4.025 $Y=0.75
c71 15 0 1.70191e-19 $X=1.64 $Y=0.77
r72 31 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.01 $X2=4.93
+ $Y2=1.095
r73 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.93 $Y=1.01
+ $X2=4.93 $Y2=0.755
r74 30 39 5.29182 $w=1.7e-07 $l=1.08995e-07 $layer=LI1_cond $X=4.115 $Y=1.095
+ $X2=4.027 $Y2=1.142
r75 29 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.805 $Y=1.095
+ $X2=4.93 $Y2=1.095
r76 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.805 $Y=1.095
+ $X2=4.115 $Y2=1.095
r77 25 39 1.23839 $w=1.75e-07 $l=1.32e-07 $layer=LI1_cond $X=4.027 $Y=1.01
+ $X2=4.027 $Y2=1.142
r78 25 27 16.4779 $w=1.73e-07 $l=2.6e-07 $layer=LI1_cond $X=4.027 $Y=1.01
+ $X2=4.027 $Y2=0.75
r79 24 38 4.85493 $w=2.1e-07 $l=1.51687e-07 $layer=LI1_cond $X=2.74 $Y=1.19
+ $X2=2.607 $Y2=1.15
r80 23 39 5.29182 $w=1.7e-07 $l=1.08374e-07 $layer=LI1_cond $X=3.94 $Y=1.19
+ $X2=4.027 $Y2=1.142
r81 23 24 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=3.94 $Y=1.19
+ $X2=2.74 $Y2=1.19
r82 19 38 1.61074 $w=1.95e-07 $l=1.41421e-07 $layer=LI1_cond $X=2.572 $Y=1.025
+ $X2=2.607 $Y2=1.15
r83 19 21 12.7972 $w=1.93e-07 $l=2.25e-07 $layer=LI1_cond $X=2.572 $Y=1.025
+ $X2=2.572 $Y2=0.8
r84 18 36 3.95903 $w=2.5e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.805 $Y=1.15
+ $X2=1.64 $Y2=1.155
r85 17 38 4.85493 $w=2.1e-07 $l=1.32e-07 $layer=LI1_cond $X=2.475 $Y=1.15
+ $X2=2.607 $Y2=1.15
r86 17 18 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=1.15
+ $X2=1.805 $Y2=1.15
r87 13 36 3.0275 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.64 $Y=1.025 $X2=1.64
+ $Y2=1.155
r88 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.64 $Y=1.025
+ $X2=1.64 $Y2=0.77
r89 4 41 182 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.595 $X2=4.89 $Y2=1.095
r90 4 33 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.595 $X2=4.89 $Y2=0.755
r91 3 27 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.595 $X2=4.025 $Y2=0.75
r92 2 38 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.625 $X2=2.57 $Y2=1.14
r93 2 21 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.625 $X2=2.57 $Y2=0.8
r94 1 36 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.625 $X2=1.64 $Y2=1.12
r95 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.625 $X2=1.64 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_4%VGND 1 2 3 4 5 18 22 26 32 34 36 39 40 42 43
+ 44 46 61 65 71 74 78
r91 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r92 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r93 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r94 69 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r95 69 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r96 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r97 66 74 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.565 $Y=0 $X2=6.365
+ $Y2=0
r98 66 68 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.565 $Y=0 $X2=6.96
+ $Y2=0
r99 65 77 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.235 $Y=0 $X2=7.457
+ $Y2=0
r100 65 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.235 $Y=0
+ $X2=6.96 $Y2=0
r101 64 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r102 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r103 61 74 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.165 $Y=0 $X2=6.365
+ $Y2=0
r104 61 63 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=0 $X2=6
+ $Y2=0
r105 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r106 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r107 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r108 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 54 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.595
+ $Y2=0
r110 54 56 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=4.08
+ $Y2=0
r111 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r112 52 53 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r113 49 53 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=3.12 $Y2=0
r114 48 52 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r115 48 49 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r116 46 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.595
+ $Y2=0
r117 46 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.12
+ $Y2=0
r118 44 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r119 44 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r120 42 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.235 $Y=0
+ $X2=5.04 $Y2=0
r121 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.4
+ $Y2=0
r122 41 63 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=6
+ $Y2=0
r123 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.4
+ $Y2=0
r124 39 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.08 $Y2=0
r125 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.46
+ $Y2=0
r126 38 59 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=5.04 $Y2=0
r127 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.46
+ $Y2=0
r128 34 77 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.457 $Y2=0
r129 34 36 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.4 $Y2=0.64
r130 30 74 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0
r131 30 32 15.9901 $w=3.98e-07 $l=5.55e-07 $layer=LI1_cond $X=6.365 $Y=0.085
+ $X2=6.365 $Y2=0.64
r132 26 28 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.4 $Y=0.64
+ $X2=5.4 $Y2=1.055
r133 24 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=0.085 $X2=5.4
+ $Y2=0
r134 24 26 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=5.4 $Y=0.085
+ $X2=5.4 $Y2=0.64
r135 20 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r136 20 22 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.745
r137 16 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0
r138 16 18 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0.755
r139 5 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.19
+ $Y=0.495 $X2=7.4 $Y2=0.64
r140 4 32 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.495 $X2=6.365 $Y2=0.64
r141 3 28 182 $w=1.7e-07 $l=5.59285e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.595 $X2=5.4 $Y2=1.055
r142 3 26 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.595 $X2=5.4 $Y2=0.64
r143 2 22 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.595 $X2=4.46 $Y2=0.745
r144 1 18 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.595 $X2=3.595 $Y2=0.755
.ends


* File: sky130_fd_sc_ms__dfbbn_1.spice
* Created: Fri Aug 28 17:21:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfbbn_1.pex.spice"
.subckt sky130_fd_sc_ms__dfbbn_1  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1035 N_VGND_M1035_d N_CLK_N_M1035_g N_A_27_74#_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1036 N_A_200_74#_M1036_d N_A_27_74#_M1036_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g N_A_311_119#_M1014_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.137937 AS=0.1197 PD=1.13 PS=1.41 NRD=78.12 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1010 A_523_119# N_A_474_405#_M1010_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.137937 PD=0.63 PS=1.13 NRD=14.28 NRS=78.12 M=1 R=2.8 SA=75000.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_A_595_119#_M1001_d N_A_27_74#_M1001_g A_523_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 N_A_311_119#_M1005_d N_A_200_74#_M1005_g N_A_595_119#_M1001_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.40005 AS=0.0588 PD=2.58 PS=0.7 NRD=256.428 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_474_405#_M1020_d N_A_595_119#_M1020_g N_A_867_119#_M1020_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.15675 PD=0.9 PS=1.67 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75004.8 A=0.0825 P=1.4 MULT=1
MM1032 N_A_867_119#_M1032_d N_A_978_357#_M1032_g N_A_474_405#_M1020_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.09625 PD=0.9 PS=0.9 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.7 SB=75004.3 A=0.0825 P=1.4 MULT=1
MM1027 N_VGND_M1027_d N_SET_B_M1027_g N_A_867_119#_M1032_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.09625 AS=0.09625 PD=0.9 PS=0.9 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.2 SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1024 A_1254_119# N_A_474_405#_M1024_g N_VGND_M1027_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.0915625 AS=0.09625 PD=0.9 PS=0.9 NRD=24.312 NRS=0 M=1 R=3.66667
+ SA=75001.7 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1028 N_A_1349_114#_M1028_d N_A_27_74#_M1028_g A_1254_119# VNB NLOWVT L=0.15
+ W=0.55 AD=0.356224 AS=0.0915625 PD=1.93918 PS=0.9 NRD=0 NRS=24.312 M=1
+ R=3.66667 SA=75002.1 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1022 A_1611_140# N_A_200_74#_M1022_g N_A_1349_114#_M1028_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.272026 PD=0.66 PS=1.48082 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75003.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_1534_446#_M1000_g A_1611_140# VNB NLOWVT L=0.15 W=0.42
+ AD=0.108295 AS=0.0504 PD=0.89431 PS=0.66 NRD=57.948 NRS=18.564 M=1 R=2.8
+ SA=75003.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_1818_76#_M1016_d N_SET_B_M1016_g N_VGND_M1000_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.190805 PD=1.02 PS=1.57569 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1034 N_A_1534_446#_M1034_d N_A_978_357#_M1034_g N_A_1818_76#_M1016_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=3.24 NRS=0 M=1
+ R=4.93333 SA=75003.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1033 N_A_1818_76#_M1033_d N_A_1349_114#_M1033_g N_A_1534_446#_M1034_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.296 AS=0.1184 PD=2.52 PS=1.06 NRD=55.944 NRS=0 M=1
+ R=4.93333 SA=75003.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g N_A_978_357#_M1008_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.12457 AS=0.1134 PD=1.00293 PS=1.38 NRD=69.024 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1029 N_Q_N_M1029_d N_A_1534_446#_M1029_g N_VGND_M1008_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.21948 PD=2.02 PS=1.76707 NRD=0 NRS=39.168 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_1534_446#_M1002_g N_A_2412_410#_M1002_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0837466 AS=0.1134 PD=0.78569 PS=1.38 NRD=18.564 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_Q_M1009_d N_A_2412_410#_M1009_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.147553 PD=2.02 PS=1.38431 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 N_VPWR_M1030_d N_CLK_N_M1030_g N_A_27_74#_M1030_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1031 N_A_200_74#_M1031_d N_A_27_74#_M1031_g N_VPWR_M1030_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.1512 PD=2.77 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1017_d N_D_M1017_g N_A_311_119#_M1017_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0882 AS=0.17175 PD=0.84 PS=1.72 NRD=65.6601 NRS=39.8531 M=1 R=2.33333
+ SA=90000.3 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1006 A_540_503# N_A_474_405#_M1006_g N_VPWR_M1017_d VPB PSHORT L=0.18 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=30.4759 NRS=0 M=1 R=2.33333 SA=90000.9
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1015 N_A_595_119#_M1015_d N_A_200_74#_M1015_g A_540_503# VPB PSHORT L=0.18
+ W=0.42 AD=0.0693 AS=0.0504 PD=0.75 PS=0.66 NRD=11.7215 NRS=30.4759 M=1
+ R=2.33333 SA=90001.3 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1012 N_A_311_119#_M1012_d N_A_27_74#_M1012_g N_A_595_119#_M1015_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1641 AS=0.0693 PD=1.69 PS=0.75 NRD=32.8202 NRS=11.7215 M=1
+ R=2.33333 SA=90001.8 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1021 A_936_424# N_A_595_119#_M1021_g N_A_474_405#_M1021_s VPB PSHORT L=0.18
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001 A=0.1512 P=2.04 MULT=1
MM1003 N_VPWR_M1003_d N_A_978_357#_M1003_g A_936_424# VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.0882 PD=1.11 PS=1.05 NRD=0 NRS=11.7215 M=1 R=4.66667 SA=90000.6
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1013 N_A_474_405#_M1013_d N_SET_B_M1013_g N_VPWR_M1003_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2226 AS=0.1134 PD=2.21 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667 SA=90001
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1007 A_1300_424# N_A_474_405#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1038 N_A_1349_114#_M1038_d N_A_200_74#_M1038_g A_1300_424# VPB PSHORT L=0.18
+ W=0.84 AD=0.1792 AS=0.0882 PD=1.6 PS=1.05 NRD=0 NRS=11.7215 M=1 R=4.66667
+ SA=90000.6 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1018 A_1486_508# N_A_27_74#_M1018_g N_A_1349_114#_M1038_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0896 PD=0.66 PS=0.8 NRD=30.4759 NRS=39.8531 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1023 N_VPWR_M1023_d N_A_1534_446#_M1023_g A_1486_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.244375 AS=0.0504 PD=2.11 PS=0.66 NRD=247.097 NRS=30.4759 M=1 R=2.33333
+ SA=90001.5 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1025 N_VPWR_M1025_d N_SET_B_M1025_g N_A_1534_446#_M1025_s VPB PSHORT L=0.18
+ W=1 AD=0.254075 AS=0.28 PD=1.675 PS=2.56 NRD=39.203 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1019 A_1920_392# N_A_978_357#_M1019_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.254075 PD=1.24 PS=1.675 NRD=12.7853 NRS=39.203 M=1 R=5.55556
+ SA=90000.8 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1026 N_A_1534_446#_M1026_d N_A_1349_114#_M1026_g A_1920_392# VPB PSHORT L=0.18
+ W=1 AD=0.265 AS=0.12 PD=2.53 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_RESET_B_M1011_g N_A_978_357#_M1011_s VPB PSHORT L=0.18
+ W=0.64 AD=0.127418 AS=0.1696 PD=1.06545 PS=1.81 NRD=44.3447 NRS=0 M=1
+ R=3.55556 SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1004 N_Q_N_M1004_d N_A_1534_446#_M1004_g N_VPWR_M1011_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.222982 PD=2.77 PS=1.86455 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1039 N_VPWR_M1039_d N_A_1534_446#_M1039_g N_A_2412_410#_M1039_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1566 AS=0.2268 PD=1.25571 PS=2.22 NRD=32.2292 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1037 N_Q_M1037_d N_A_2412_410#_M1037_g N_VPWR_M1039_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.2088 PD=2.78 PS=1.67429 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.7052 P=31.36
c_147 VNB 0 5.76555e-20 $X=0 $Y=0
c_278 VPB 0 4.72451e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dfbbn_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 a_195_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=7.498e+11p ps=6.7e+06u
M1001 X a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.4496e+12p ps=9.24e+06u
M1002 VPWR a_27_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_27_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 a_195_74# B1 a_117_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1005 a_317_368# A2 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.5e+11p ps=5.1e+06u
M1006 a_27_368# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C1 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_317_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_195_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_117_74# C1 a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends

* File: sky130_fd_sc_ms__o22a_2.spice
* Created: Wed Sep  2 12:23:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o22a_2.pex.spice"
.subckt sky130_fd_sc_ms__o22a_2  VNB VPB B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_A_82_48#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1004_d N_A_82_48#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19325 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_82_48#_M1003_d N_B1_M1003_g N_A_307_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1147 AS=0.195 PD=1.05 PS=2.03 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1011 N_A_307_74#_M1011_d N_B2_M1011_g N_A_82_48#_M1003_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1147 PD=1.09 PS=1.05 NRD=11.34 NRS=2.424 M=1 R=4.93333
+ SA=75000.6 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_307_74#_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_A_307_74#_M1007_d N_A1_M1007_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_82_48#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1002 N_X_M1001_d N_A_82_48#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.353011 PD=1.39 PS=1.85434 NRD=0 NRS=45.7631 M=1 R=6.22222
+ SA=90000.7 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1006 A_386_384# N_B1_M1006_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1 AD=0.135
+ AS=0.315189 PD=1.27 PS=1.65566 NRD=15.7403 NRS=51.2397 M=1 R=5.55556
+ SA=90001.5 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1008 N_A_82_48#_M1008_d N_B2_M1008_g A_386_384# VPB PSHORT L=0.18 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=0 NRS=15.7403 M=1 R=5.55556 SA=90002 SB=90001.2
+ A=0.18 P=2.36 MULT=1
MM1000 A_578_384# N_A2_M1000_g N_A_82_48#_M1008_d VPB PSHORT L=0.18 W=1 AD=0.18
+ AS=0.165 PD=1.36 PS=1.33 NRD=24.6053 NRS=10.8153 M=1 R=5.55556 SA=90002.5
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_578_384# VPB PSHORT L=0.18 W=1 AD=0.275
+ AS=0.18 PD=2.55 PS=1.36 NRD=0 NRS=24.6053 M=1 R=5.55556 SA=90003 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o22a_2.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or3_2 A B C VGND VNB VPB VPWR X
M1000 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=9.725e+11p pd=7.09e+06u as=2.072e+11p ps=2.04e+06u
M1001 VPWR A a_237_392# VPB pshort w=1e+06u l=180000u
+  ad=8.296e+11p pd=6e+06u as=3.9e+11p ps=2.78e+06u
M1002 a_237_392# B a_153_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1003 a_153_392# C a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1004 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VGND A a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.064e+11p ps=3.83e+06u
M1006 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

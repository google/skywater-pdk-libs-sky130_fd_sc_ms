* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2_4 A B VGND VNB VPB VPWR X
X0 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X1 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X7 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X12 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

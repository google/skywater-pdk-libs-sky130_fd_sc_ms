* File: sky130_fd_sc_ms__sdlclkp_4.spice
* Created: Wed Sep  2 12:32:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdlclkp_4.pex.spice"
.subckt sky130_fd_sc_ms__sdlclkp_4  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1023 N_A_119_143#_M1023_d N_SCE_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.089375 AS=0.1705 PD=0.875 PS=1.72 NRD=9.816 NRS=5.448 M=1
+ R=3.66667 SA=75000.2 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1026 N_VGND_M1026_d N_GATE_M1026_g N_A_119_143#_M1023_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.233963 AS=0.089375 PD=1.43256 PS=0.875 NRD=80.808 NRS=0 M=1
+ R=3.66667 SA=75000.7 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1021 N_A_354_105#_M1021_d N_A_324_79#_M1021_g N_VGND_M1026_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.314787 PD=2.05 PS=1.92744 NRD=0 NRS=60.06 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_634_74#_M1024_d N_A_324_79#_M1024_g N_A_119_143#_M1024_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.119214 AS=0.38225 PD=1.07732 PS=2.49 NRD=4.356 NRS=77.448
+ M=1 R=3.66667 SA=75000.6 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1017 A_744_74# N_A_354_105#_M1017_g N_A_634_74#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0910361 PD=0.66 PS=0.82268 NRD=18.564 NRS=30 M=1 R=2.8
+ SA=75001.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_792_48#_M1007_g A_744_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.136934 AS=0.0504 PD=1.05 PS=0.66 NRD=5.712 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_792_48#_M1006_d N_A_634_74#_M1006_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.241266 PD=2.05 PS=1.85 NRD=0 NRS=66.48 M=1 R=4.93333
+ SA=75001.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_CLK_M1013_g N_A_324_79#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 A_1292_74# N_CLK_M1011_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1295 PD=0.98 PS=1.09 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_1292_368#_M1012_d N_A_792_48#_M1012_g A_1292_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_1292_368#_M1000_g N_GCLK_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1221 PD=2.05 PS=1.07 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_1292_368#_M1003_g N_GCLK_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1003_d N_A_1292_368#_M1015_g N_GCLK_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_1292_368#_M1027_g N_GCLK_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 A_119_395# N_SCE_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1008 AS=0.2352 PD=1.08 PS=2.24 NRD=15.2281 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1001 N_A_119_143#_M1001_d N_GATE_M1001_g A_119_395# VPB PSHORT L=0.18 W=0.84
+ AD=0.2352 AS=0.1008 PD=2.24 PS=1.08 NRD=0 NRS=15.2281 M=1 R=4.66667 SA=90000.6
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1004 N_A_354_105#_M1004_d N_A_324_79#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18
+ W=0.84 AD=0.3907 AS=0.4746 PD=2.99 PS=2.81 NRD=96.1754 NRS=0 M=1 R=4.66667
+ SA=90000.5 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1005 N_A_634_74#_M1005_d N_A_354_105#_M1005_g N_A_119_143#_M1005_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1778 AS=0.2352 PD=1.59333 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1008 A_788_455# N_A_324_79#_M1008_g N_A_634_74#_M1005_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0889 PD=0.66 PS=0.796667 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90000.7 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1014 N_VPWR_M1014_d N_A_792_48#_M1014_g A_788_455# VPB PSHORT L=0.18 W=0.42
+ AD=0.0958364 AS=0.0504 PD=0.812727 PS=0.66 NRD=46.886 NRS=30.4759 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1022 N_A_792_48#_M1022_d N_A_634_74#_M1022_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.255564 PD=2.8 PS=2.16727 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.8 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_CLK_M1002_g N_A_324_79#_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1614 AS=0.2394 PD=1.26429 PS=2.25 NRD=32.1504 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003.4 A=0.1512 P=2.04 MULT=1
MM1020 N_A_1292_368#_M1020_d N_CLK_M1020_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2604 AS=0.2152 PD=1.585 PS=1.68571 NRD=33.4112 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1019_d N_A_792_48#_M1019_g N_A_1292_368#_M1020_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.1792 AS=0.2604 PD=1.44 PS=1.585 NRD=7.8997 NRS=0 M=1
+ R=6.22222 SA=90001.2 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1009 N_GCLK_M1009_d N_A_1292_368#_M1009_g N_VPWR_M1019_d VPB PSHORT L=0.18
+ W=1.12 AD=0.224 AS=0.1792 PD=1.52 PS=1.44 NRD=21.9852 NRS=0 M=1 R=6.22222
+ SA=90001.7 SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1010 N_GCLK_M1009_d N_A_1292_368#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.224 AS=0.1792 PD=1.52 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1016 N_GCLK_M1016_d N_A_1292_368#_M1016_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1764 AS=0.1792 PD=1.435 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.8 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1018 N_GCLK_M1016_d N_A_1292_368#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1764 AS=0.3192 PD=1.435 PS=2.81 NRD=7.0329 NRS=0 M=1 R=6.22222
+ SA=90003.3 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.6851 P=23.85
*
.include "sky130_fd_sc_ms__sdlclkp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand2_4.pxi.spice
* Created: Wed Sep  2 12:12:55 2020
* 
x_PM_SKY130_FD_SC_MS__NAND2_4%B N_B_M1004_g N_B_M1001_g N_B_M1007_g N_B_M1010_g
+ N_B_M1008_g N_B_M1011_g B B B N_B_c_72_n N_B_c_77_n N_B_c_94_p
+ PM_SKY130_FD_SC_MS__NAND2_4%B
x_PM_SKY130_FD_SC_MS__NAND2_4%A N_A_M1002_g N_A_M1000_g N_A_M1003_g N_A_c_129_n
+ N_A_c_130_n N_A_M1005_g N_A_M1009_g N_A_M1006_g N_A_c_133_n N_A_c_134_n
+ N_A_c_135_n A A A N_A_c_143_n PM_SKY130_FD_SC_MS__NAND2_4%A
x_PM_SKY130_FD_SC_MS__NAND2_4%VPWR N_VPWR_M1001_s N_VPWR_M1008_s N_VPWR_M1009_d
+ N_VPWR_c_196_n N_VPWR_c_197_n N_VPWR_c_198_n N_VPWR_c_199_n N_VPWR_c_200_n
+ N_VPWR_c_201_n N_VPWR_c_202_n VPWR N_VPWR_c_203_n N_VPWR_c_195_n
+ PM_SKY130_FD_SC_MS__NAND2_4%VPWR
x_PM_SKY130_FD_SC_MS__NAND2_4%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1001_d N_Y_M1000_s
+ N_Y_c_249_n N_Y_c_232_n N_Y_c_233_n N_Y_c_294_p N_Y_c_234_n N_Y_c_237_n
+ N_Y_c_238_n N_Y_c_246_n N_Y_c_239_n N_Y_c_235_n Y Y
+ PM_SKY130_FD_SC_MS__NAND2_4%Y
x_PM_SKY130_FD_SC_MS__NAND2_4%A_27_74# N_A_27_74#_M1004_s N_A_27_74#_M1007_s
+ N_A_27_74#_M1011_s N_A_27_74#_M1003_s N_A_27_74#_M1006_s N_A_27_74#_c_297_n
+ N_A_27_74#_c_298_n N_A_27_74#_c_299_n N_A_27_74#_c_300_n N_A_27_74#_c_301_n
+ N_A_27_74#_c_302_n N_A_27_74#_c_303_n N_A_27_74#_c_326_n N_A_27_74#_c_304_n
+ N_A_27_74#_c_305_n N_A_27_74#_c_306_n N_A_27_74#_c_307_n
+ PM_SKY130_FD_SC_MS__NAND2_4%A_27_74#
x_PM_SKY130_FD_SC_MS__NAND2_4%VGND N_VGND_M1004_d N_VGND_M1010_d N_VGND_c_365_n
+ N_VGND_c_366_n VGND N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n
+ N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n PM_SKY130_FD_SC_MS__NAND2_4%VGND
cc_1 VNB N_B_M1004_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B_M1007_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_B_M1010_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_4 VNB N_B_M1011_g 0.0235145f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.74
cc_5 VNB B 0.00341995f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_B_c_72_n 0.0764705f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.515
cc_7 VNB N_A_M1002_g 0.02421f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_A_M1003_g 0.0236518f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_9 VNB N_A_c_129_n 0.0155576f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_10 VNB N_A_c_130_n 0.0278603f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_11 VNB N_A_M1005_g 0.0249853f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.68
cc_12 VNB N_A_M1006_g 0.027911f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.515
cc_13 VNB N_A_c_133_n 0.004935f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.515
cc_14 VNB N_A_c_134_n 0.0183368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_135_n 0.0137989f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_16 VNB N_VPWR_c_195_n 0.183584f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.565
cc_17 VNB N_Y_c_232_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.4
cc_18 VNB N_Y_c_233_n 0.00579183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_234_n 0.0112196f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.515
cc_20 VNB N_Y_c_235_n 0.00281002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB Y 0.024009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_297_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.4
cc_23 VNB N_A_27_74#_c_298_n 0.00365673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_299_n 0.0116376f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_25 VNB N_A_27_74#_c_300_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_301_n 0.00628038f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.515
cc_27 VNB N_A_27_74#_c_302_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_28 VNB N_A_27_74#_c_303_n 0.00286768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_304_n 0.0133886f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_30 VNB N_A_27_74#_c_305_n 0.0148481f $X=-0.19 $Y=-0.245 $X2=1.695 $Y2=1.515
cc_31 VNB N_A_27_74#_c_306_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=1.695 $Y2=1.515
cc_32 VNB N_A_27_74#_c_307_n 0.002205f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_33 VNB N_VGND_c_365_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.35
cc_34 VNB N_VGND_c_366_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_35 VNB N_VGND_c_367_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.68
cc_36 VNB N_VGND_c_368_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.74
cc_37 VNB N_VGND_c_369_n 0.0621234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_370_n 0.253463f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_39 VNB N_VGND_c_371_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_372_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_41 VPB N_B_M1001_g 0.0341735f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_42 VPB N_B_M1008_g 0.0274958f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=2.4
cc_43 VPB B 0.00451804f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_44 VPB N_B_c_72_n 0.0296283f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.515
cc_45 VPB N_B_c_77_n 0.00549802f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.565
cc_46 VPB N_A_M1000_g 0.0278208f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_47 VPB N_A_c_129_n 0.0106787f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.35
cc_48 VPB N_A_c_130_n 0.0113002f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_49 VPB N_A_M1009_g 0.0295127f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.35
cc_50 VPB N_A_c_133_n 0.00459923f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.515
cc_51 VPB N_A_c_134_n 0.00921362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_c_135_n 8.9025e-19 $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_53 VPB N_A_c_143_n 0.0120703f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.515
cc_54 VPB N_VPWR_c_196_n 0.0120013f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_55 VPB N_VPWR_c_197_n 0.0524677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_198_n 0.00635448f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=2.4
cc_57 VPB N_VPWR_c_199_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_200_n 0.0391645f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.74
cc_59 VPB N_VPWR_c_201_n 0.0355463f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.515
cc_60 VPB N_VPWR_c_202_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.515
cc_61 VPB N_VPWR_c_203_n 0.0437907f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_62 VPB N_VPWR_c_195_n 0.0681937f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.565
cc_63 VPB N_Y_c_237_n 0.00707089f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.515
cc_64 VPB N_Y_c_238_n 0.0099111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_Y_c_239_n 0.0119707f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.515
cc_66 VPB Y 0.012933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 N_B_M1011_g N_A_M1002_g 0.018445f $X=1.785 $Y=0.74 $X2=0 $Y2=0
cc_68 N_B_M1008_g N_A_M1000_g 0.018445f $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_69 B N_A_M1000_g 0.00422776f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_70 B N_A_c_130_n 0.0167617f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_71 N_B_c_72_n N_A_c_130_n 0.018445f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_72 B N_A_c_143_n 0.0366331f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_73 N_B_M1001_g N_VPWR_c_197_n 0.0250669f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_74 N_B_M1008_g N_VPWR_c_198_n 0.0153892f $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_75 N_B_M1001_g N_VPWR_c_201_n 0.00475445f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_76 N_B_M1008_g N_VPWR_c_201_n 0.00460063f $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_77 N_B_M1001_g N_VPWR_c_195_n 0.00943794f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_78 N_B_M1008_g N_VPWR_c_195_n 0.00913687f $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_79 N_B_M1001_g N_Y_c_238_n 4.72675e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_80 N_B_M1008_g N_Y_c_238_n 4.69668e-19 $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_81 N_B_c_72_n N_Y_c_238_n 0.0129542f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B_c_77_n N_Y_c_238_n 0.0456966f $X=1.515 $Y=1.565 $X2=0 $Y2=0
cc_83 N_B_c_94_p N_Y_c_238_n 0.0257641f $X=1.085 $Y=1.565 $X2=0 $Y2=0
cc_84 N_B_M1008_g N_Y_c_246_n 0.0132456f $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_85 B N_Y_c_246_n 0.0456966f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_86 N_B_M1008_g N_Y_c_239_n 5.44639e-19 $X=1.77 $Y=2.4 $X2=0 $Y2=0
cc_87 N_B_M1004_g N_A_27_74#_c_297_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_88 N_B_M1004_g N_A_27_74#_c_298_n 0.0160671f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B_M1007_g N_A_27_74#_c_298_n 0.0131257f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_90 N_B_c_72_n N_A_27_74#_c_298_n 0.00236025f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_91 N_B_c_94_p N_A_27_74#_c_298_n 0.0401403f $X=1.085 $Y=1.565 $X2=0 $Y2=0
cc_92 N_B_M1007_g N_A_27_74#_c_300_n 3.92313e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_93 N_B_M1010_g N_A_27_74#_c_300_n 3.92313e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B_M1010_g N_A_27_74#_c_301_n 0.0131257f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_95 N_B_M1011_g N_A_27_74#_c_301_n 0.0130879f $X=1.785 $Y=0.74 $X2=0 $Y2=0
cc_96 B N_A_27_74#_c_301_n 0.0225421f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_97 N_B_c_72_n N_A_27_74#_c_301_n 0.00236025f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_98 N_B_c_77_n N_A_27_74#_c_301_n 0.0519295f $X=1.515 $Y=1.565 $X2=0 $Y2=0
cc_99 N_B_M1011_g N_A_27_74#_c_303_n 0.00100872f $X=1.785 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B_c_72_n N_A_27_74#_c_306_n 0.00232957f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B_c_94_p N_A_27_74#_c_306_n 0.0145185f $X=1.085 $Y=1.565 $X2=0 $Y2=0
cc_102 N_B_M1004_g N_VGND_c_365_n 0.0127698f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B_M1007_g N_VGND_c_365_n 0.0097465f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_104 N_B_M1010_g N_VGND_c_365_n 4.61192e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_105 N_B_M1007_g N_VGND_c_366_n 4.61192e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B_M1010_g N_VGND_c_366_n 0.0097465f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_107 N_B_M1011_g N_VGND_c_366_n 0.0091452f $X=1.785 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VGND_c_367_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B_M1007_g N_VGND_c_368_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_110 N_B_M1010_g N_VGND_c_368_n 0.00383152f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_111 N_B_M1011_g N_VGND_c_369_n 0.00383152f $X=1.785 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B_M1004_g N_VGND_c_370_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B_M1007_g N_VGND_c_370_n 0.0075754f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B_M1010_g N_VGND_c_370_n 0.0075754f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B_M1011_g N_VGND_c_370_n 0.00757998f $X=1.785 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_M1000_g N_VPWR_c_198_n 0.00339365f $X=2.27 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_M1009_g N_VPWR_c_200_n 0.00546942f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_M1000_g N_VPWR_c_203_n 0.00519794f $X=2.27 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_M1009_g N_VPWR_c_203_n 0.00519794f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_M1000_g N_VPWR_c_195_n 0.00983645f $X=2.27 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_M1009_g N_VPWR_c_195_n 0.00986983f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_M1003_g N_Y_c_249_n 0.00673416f $X=2.715 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_M1005_g N_Y_c_249_n 6.07762e-19 $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_M1003_g N_Y_c_232_n 0.0093986f $X=2.715 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_c_129_n N_Y_c_232_n 0.00381149f $X=3.14 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_M1005_g N_Y_c_232_n 0.0132585f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_c_143_n N_Y_c_232_n 0.0501792f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_M1002_g N_Y_c_233_n 0.00116487f $X=2.255 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_M1003_g N_Y_c_233_n 0.00264402f $X=2.715 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_c_130_n N_Y_c_233_n 0.00362741f $X=2.79 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_c_143_n N_Y_c_233_n 0.0185202f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_M1006_g N_Y_c_234_n 0.0137226f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_c_143_n N_Y_c_234_n 0.0065328f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_M1009_g N_Y_c_237_n 0.0162996f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_M1000_g N_Y_c_246_n 0.0130369f $X=2.27 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_M1000_g N_Y_c_239_n 0.0140606f $X=2.27 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_c_130_n N_Y_c_239_n 0.00693896f $X=2.79 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_M1009_g N_Y_c_239_n 0.0178797f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_c_143_n N_Y_c_239_n 0.114637f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A_M1006_g N_Y_c_235_n 0.0027366f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_c_134_n N_Y_c_235_n 0.00555564f $X=3.675 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_c_143_n N_Y_c_235_n 0.0312938f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_M1006_g Y 0.024494f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_c_143_n Y 0.0349192f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A_M1002_g N_A_27_74#_c_301_n 6.49072e-19 $X=2.255 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_A_27_74#_c_302_n 0.0131021f $X=2.255 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_M1003_g N_A_27_74#_c_302_n 0.011414f $X=2.715 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_A_27_74#_c_326_n 0.00610666f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_A_27_74#_c_326_n 8.34587e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_M1005_g N_A_27_74#_c_304_n 0.00862423f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_A_27_74#_c_304_n 0.013369f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_M1005_g N_A_27_74#_c_307_n 0.00294698f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_VGND_c_369_n 0.00278271f $X=2.255 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_M1003_g N_VGND_c_369_n 0.00278271f $X=2.715 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_M1005_g N_VGND_c_369_n 0.00278247f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_M1006_g N_VGND_c_369_n 0.00278271f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_VGND_c_370_n 0.00354179f $X=2.255 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_VGND_c_370_n 0.0035438f $X=2.715 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_M1005_g N_VGND_c_370_n 0.0035528f $X=3.215 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_M1006_g N_VGND_c_370_n 0.00358426f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_161 N_VPWR_M1009_d N_Y_c_237_n 0.0063718f $X=3.855 $Y=1.84 $X2=0 $Y2=0
cc_162 N_VPWR_c_200_n N_Y_c_237_n 0.0249562f $X=4.04 $Y=2.42 $X2=0 $Y2=0
cc_163 N_VPWR_c_197_n N_Y_c_238_n 0.0395953f $X=0.28 $Y=2.015 $X2=0 $Y2=0
cc_164 N_VPWR_c_198_n N_Y_c_238_n 0.0268148f $X=1.995 $Y=2.42 $X2=0 $Y2=0
cc_165 N_VPWR_c_201_n N_Y_c_238_n 0.0464425f $X=1.83 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VPWR_c_195_n N_Y_c_238_n 0.0385721f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_167 N_VPWR_M1008_s N_Y_c_246_n 0.00438498f $X=1.86 $Y=1.84 $X2=0 $Y2=0
cc_168 N_VPWR_c_198_n N_Y_c_246_n 0.0189268f $X=1.995 $Y=2.42 $X2=0 $Y2=0
cc_169 N_VPWR_c_198_n N_Y_c_239_n 0.0297756f $X=1.995 $Y=2.42 $X2=0 $Y2=0
cc_170 N_VPWR_c_200_n N_Y_c_239_n 0.0297756f $X=4.04 $Y=2.42 $X2=0 $Y2=0
cc_171 N_VPWR_c_203_n N_Y_c_239_n 0.0609295f $X=3.875 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_195_n N_Y_c_239_n 0.0504633f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_M1009_d Y 0.00217208f $X=3.855 $Y=1.84 $X2=0 $Y2=0
cc_174 N_VPWR_c_197_n N_A_27_74#_c_298_n 0.00134655f $X=0.28 $Y=2.015 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_197_n N_A_27_74#_c_299_n 0.00842269f $X=0.28 $Y=2.015 $X2=0
+ $Y2=0
cc_176 N_Y_c_232_n N_A_27_74#_M1003_s 0.00271958f $X=3.335 $Y=1.095 $X2=0 $Y2=0
cc_177 N_Y_c_234_n N_A_27_74#_M1006_s 0.00407071f $X=3.965 $Y=1.095 $X2=0 $Y2=0
cc_178 N_Y_c_233_n N_A_27_74#_c_301_n 0.00646046f $X=2.665 $Y=1.095 $X2=0 $Y2=0
cc_179 N_Y_M1002_d N_A_27_74#_c_302_n 0.00215923f $X=2.33 $Y=0.37 $X2=0 $Y2=0
cc_180 N_Y_c_249_n N_A_27_74#_c_302_n 0.0152139f $X=2.5 $Y=0.785 $X2=0 $Y2=0
cc_181 N_Y_c_232_n N_A_27_74#_c_302_n 0.00304353f $X=3.335 $Y=1.095 $X2=0 $Y2=0
cc_182 N_Y_c_232_n N_A_27_74#_c_326_n 0.0179263f $X=3.335 $Y=1.095 $X2=0 $Y2=0
cc_183 N_Y_M1005_d N_A_27_74#_c_304_n 0.00348036f $X=3.29 $Y=0.37 $X2=0 $Y2=0
cc_184 N_Y_c_232_n N_A_27_74#_c_304_n 0.00304353f $X=3.335 $Y=1.095 $X2=0 $Y2=0
cc_185 N_Y_c_294_p N_A_27_74#_c_304_n 0.0210188f $X=3.52 $Y=0.785 $X2=0 $Y2=0
cc_186 N_Y_c_234_n N_A_27_74#_c_304_n 0.00365468f $X=3.965 $Y=1.095 $X2=0 $Y2=0
cc_187 N_Y_c_234_n N_A_27_74#_c_305_n 0.0214359f $X=3.965 $Y=1.095 $X2=0 $Y2=0
cc_188 N_A_27_74#_c_298_n N_VGND_M1004_d 0.00191292f $X=1.055 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_27_74#_c_301_n N_VGND_M1010_d 0.00191292f $X=1.915 $Y=1.095 $X2=0
+ $Y2=0
cc_190 N_A_27_74#_c_297_n N_VGND_c_365_n 0.0170358f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_191 N_A_27_74#_c_298_n N_VGND_c_365_n 0.0148206f $X=1.055 $Y=1.095 $X2=0
+ $Y2=0
cc_192 N_A_27_74#_c_300_n N_VGND_c_365_n 0.0169944f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_193 N_A_27_74#_c_300_n N_VGND_c_366_n 0.0169944f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_194 N_A_27_74#_c_301_n N_VGND_c_366_n 0.0148206f $X=1.915 $Y=1.095 $X2=0
+ $Y2=0
cc_195 N_A_27_74#_c_303_n N_VGND_c_366_n 0.0112234f $X=2.165 $Y=0.34 $X2=0 $Y2=0
cc_196 N_A_27_74#_c_297_n N_VGND_c_367_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_197 N_A_27_74#_c_300_n N_VGND_c_368_n 0.00749631f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_198 N_A_27_74#_c_302_n N_VGND_c_369_n 0.0422287f $X=2.835 $Y=0.34 $X2=0 $Y2=0
cc_199 N_A_27_74#_c_303_n N_VGND_c_369_n 0.0179217f $X=2.165 $Y=0.34 $X2=0 $Y2=0
cc_200 N_A_27_74#_c_304_n N_VGND_c_369_n 0.0681649f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_201 N_A_27_74#_c_307_n N_VGND_c_369_n 0.0231983f $X=3 $Y=0.34 $X2=0 $Y2=0
cc_202 N_A_27_74#_c_297_n N_VGND_c_370_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_203 N_A_27_74#_c_300_n N_VGND_c_370_n 0.0062048f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_204 N_A_27_74#_c_302_n N_VGND_c_370_n 0.0238173f $X=2.835 $Y=0.34 $X2=0 $Y2=0
cc_205 N_A_27_74#_c_303_n N_VGND_c_370_n 0.00971942f $X=2.165 $Y=0.34 $X2=0
+ $Y2=0
cc_206 N_A_27_74#_c_304_n N_VGND_c_370_n 0.0381951f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_207 N_A_27_74#_c_307_n N_VGND_c_370_n 0.0126453f $X=3 $Y=0.34 $X2=0 $Y2=0

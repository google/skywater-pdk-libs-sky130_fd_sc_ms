* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_368_74# B1 a_260_74# VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=2.886e+11p ps=2.26e+06u
M1001 VPWR A1 a_493_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1872e+12p pd=8.84e+06u as=3.08e+11p ps=2.79e+06u
M1002 VGND A2 a_368_74# VNB nlowvt w=740000u l=150000u
+  ad=3.256e+11p pd=2.36e+06u as=0p ps=0u
M1003 a_493_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.328e+11p ps=5.61e+06u
M1004 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_368_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_182_74# D1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=4.625e+11p ps=2.73e+06u
M1007 a_260_74# C1 a_182_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y D1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__a221oi_2.pxi.spice
* Created: Wed Sep  2 11:52:24 2020
* 
x_PM_SKY130_FD_SC_MS__A221OI_2%C1 N_C1_M1016_g N_C1_M1015_g N_C1_M1017_g
+ N_C1_M1019_g C1 N_C1_c_103_n N_C1_c_104_n PM_SKY130_FD_SC_MS__A221OI_2%C1
x_PM_SKY130_FD_SC_MS__A221OI_2%B1 N_B1_M1012_g N_B1_M1003_g N_B1_M1018_g
+ N_B1_M1014_g N_B1_c_153_n N_B1_c_170_p N_B1_c_215_p N_B1_c_147_n N_B1_c_148_n
+ B1 N_B1_c_150_n PM_SKY130_FD_SC_MS__A221OI_2%B1
x_PM_SKY130_FD_SC_MS__A221OI_2%B2 N_B2_M1001_g N_B2_M1010_g N_B2_M1011_g
+ N_B2_M1008_g B2 N_B2_c_245_n N_B2_c_242_n PM_SKY130_FD_SC_MS__A221OI_2%B2
x_PM_SKY130_FD_SC_MS__A221OI_2%A1 N_A1_M1006_g N_A1_M1000_g N_A1_M1013_g
+ N_A1_M1009_g N_A1_c_298_n N_A1_c_316_p N_A1_c_309_n N_A1_c_292_n N_A1_c_300_n
+ A1 A1 N_A1_c_294_n N_A1_c_295_n PM_SKY130_FD_SC_MS__A221OI_2%A1
x_PM_SKY130_FD_SC_MS__A221OI_2%A2 N_A2_M1004_g N_A2_M1002_g N_A2_M1007_g
+ N_A2_M1005_g A2 A2 N_A2_c_373_n PM_SKY130_FD_SC_MS__A221OI_2%A2
x_PM_SKY130_FD_SC_MS__A221OI_2%A_29_368# N_A_29_368#_M1016_s N_A_29_368#_M1017_s
+ N_A_29_368#_M1010_d N_A_29_368#_M1018_d N_A_29_368#_c_422_n
+ N_A_29_368#_c_423_n N_A_29_368#_c_424_n N_A_29_368#_c_433_n
+ N_A_29_368#_c_425_n N_A_29_368#_c_426_n N_A_29_368#_c_427_n
+ N_A_29_368#_c_428_n PM_SKY130_FD_SC_MS__A221OI_2%A_29_368#
x_PM_SKY130_FD_SC_MS__A221OI_2%Y N_Y_M1015_d N_Y_M1019_d N_Y_M1014_s N_Y_M1013_d
+ N_Y_M1016_d N_Y_c_464_n N_Y_c_465_n N_Y_c_482_n N_Y_c_475_n N_Y_c_466_n
+ N_Y_c_467_n N_Y_c_468_n N_Y_c_469_n N_Y_c_470_n N_Y_c_471_n N_Y_c_484_n
+ N_Y_c_472_n N_Y_c_473_n Y Y PM_SKY130_FD_SC_MS__A221OI_2%Y
x_PM_SKY130_FD_SC_MS__A221OI_2%A_297_368# N_A_297_368#_M1012_s
+ N_A_297_368#_M1011_s N_A_297_368#_M1000_d N_A_297_368#_M1005_s
+ N_A_297_368#_c_554_n N_A_297_368#_c_581_n N_A_297_368#_c_566_n
+ N_A_297_368#_c_555_n N_A_297_368#_c_556_n
+ PM_SKY130_FD_SC_MS__A221OI_2%A_297_368#
x_PM_SKY130_FD_SC_MS__A221OI_2%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_M1009_s
+ N_VPWR_c_612_n N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n
+ N_VPWR_c_617_n N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_620_n N_VPWR_c_621_n
+ VPWR N_VPWR_c_611_n PM_SKY130_FD_SC_MS__A221OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A221OI_2%VGND N_VGND_M1015_s N_VGND_M1001_d N_VGND_M1004_s
+ N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n N_VGND_c_679_n N_VGND_c_680_n
+ VGND N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n
+ N_VGND_c_685_n N_VGND_c_686_n PM_SKY130_FD_SC_MS__A221OI_2%VGND
x_PM_SKY130_FD_SC_MS__A221OI_2%A_293_74# N_A_293_74#_M1003_d N_A_293_74#_M1008_s
+ N_A_293_74#_c_752_n N_A_293_74#_c_750_n N_A_293_74#_c_754_n
+ N_A_293_74#_c_751_n PM_SKY130_FD_SC_MS__A221OI_2%A_293_74#
x_PM_SKY130_FD_SC_MS__A221OI_2%A_675_74# N_A_675_74#_M1006_s N_A_675_74#_M1007_d
+ N_A_675_74#_c_783_n N_A_675_74#_c_780_n N_A_675_74#_c_778_n
+ N_A_675_74#_c_779_n PM_SKY130_FD_SC_MS__A221OI_2%A_675_74#
cc_1 VNB N_C1_M1015_g 0.0277392f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_2 VNB N_C1_M1019_g 0.0232324f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_3 VNB N_C1_c_103_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_4 VNB N_C1_c_104_n 0.0377928f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.515
cc_5 VNB N_B1_M1003_g 0.0237005f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_6 VNB N_B1_M1014_g 0.0235923f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_7 VNB N_B1_c_147_n 0.0224717f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_8 VNB N_B1_c_148_n 0.00376742f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.515
cc_9 VNB B1 0.00702307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_150_n 0.0229795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_M1001_g 0.0249084f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_12 VNB N_B2_M1008_g 0.0241114f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_13 VNB N_B2_c_242_n 0.0396205f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_14 VNB N_A1_M1006_g 0.0275773f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_15 VNB N_A1_M1013_g 0.03089f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_16 VNB N_A1_c_292_n 0.00226868f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_17 VNB A1 0.0194528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_294_n 0.0408708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_295_n 0.0299403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_M1004_g 0.0278279f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_21 VNB N_A2_M1007_g 0.0238434f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_22 VNB A2 0.00226937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_373_n 0.0371993f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_24 VNB N_Y_c_464_n 0.0273059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_465_n 0.00532838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_466_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_27 VNB N_Y_c_467_n 0.0164284f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.665
cc_28 VNB N_Y_c_468_n 0.0023323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_469_n 0.0295057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_470_n 0.0300805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_471_n 0.00742669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_472_n 0.00346528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_473_n 0.00228751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB Y 0.0244824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_611_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_676_n 0.00396654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_677_n 0.00978606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_678_n 0.00965695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_679_n 0.0498315f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_40 VNB N_VGND_c_680_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.515
cc_41 VNB N_VGND_c_681_n 0.0178292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_682_n 0.0280335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_683_n 0.0363163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_684_n 0.330714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_685_n 0.00640853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_686_n 0.00651315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_293_74#_c_750_n 0.00280031f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.68
cc_48 VNB N_A_293_74#_c_751_n 0.0023154f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_49 VNB N_A_675_74#_c_778_n 0.00262401f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_50 VNB N_A_675_74#_c_779_n 0.0063328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_C1_M1016_g 0.0233737f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_52 VPB N_C1_M1017_g 0.020351f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_53 VPB N_C1_c_103_n 0.00311867f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_54 VPB N_C1_c_104_n 0.00472173f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.515
cc_55 VPB N_B1_M1012_g 0.0204786f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_56 VPB N_B1_M1018_g 0.0241615f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_57 VPB N_B1_c_153_n 0.00141536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_147_n 0.00648034f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_59 VPB N_B1_c_148_n 3.51482e-19 $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.515
cc_60 VPB B1 0.00665779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_B1_c_150_n 0.00544857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B2_M1010_g 0.0206583f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_63 VPB N_B2_M1011_g 0.0208836f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_64 VPB N_B2_c_245_n 0.0025068f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_65 VPB N_B2_c_242_n 0.00461649f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_66 VPB N_A1_M1000_g 0.0242972f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_67 VPB N_A1_M1009_g 0.0245513f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_68 VPB N_A1_c_298_n 0.00117995f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_69 VPB N_A1_c_292_n 7.88439e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_70 VPB N_A1_c_300_n 5.62538e-19 $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.515
cc_71 VPB A1 0.0153918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A1_c_294_n 0.0152512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A1_c_295_n 0.00579103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A2_M1002_g 0.0207886f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_75 VPB N_A2_M1005_g 0.0213541f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_76 VPB A2 0.00460632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A2_c_373_n 0.00631576f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_78 VPB N_A_29_368#_c_422_n 0.0239548f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_79 VPB N_A_29_368#_c_423_n 0.0026202f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_80 VPB N_A_29_368#_c_424_n 0.00933537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_29_368#_c_425_n 0.00840775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_29_368#_c_426_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_29_368#_c_427_n 0.0028338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_29_368#_c_428_n 0.00159264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_Y_c_475_n 0.00722749f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_86 VPB Y 0.0131016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_297_368#_c_554_n 0.0122146f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.35
cc_88 VPB N_A_297_368#_c_555_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_297_368#_c_556_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_612_n 0.0126417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_613_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_614_n 0.0505116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_615_n 0.0809436f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.515
cc_94 VPB N_VPWR_c_616_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.515
cc_95 VPB N_VPWR_c_617_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.515
cc_96 VPB N_VPWR_c_618_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_619_n 0.0108943f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.665
cc_98 VPB N_VPWR_c_620_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_621_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_611_n 0.0861515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 N_C1_M1017_g N_B1_M1012_g 0.014198f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_102 N_C1_c_103_n N_B1_M1012_g 2.99605e-19 $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_103 N_C1_M1019_g N_B1_M1003_g 0.0187145f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_104 N_C1_M1017_g N_B1_c_153_n 6.63946e-19 $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_105 N_C1_c_103_n N_B1_c_153_n 0.00288203f $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_106 N_C1_c_103_n N_B1_c_147_n 7.03909e-19 $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_107 N_C1_c_104_n N_B1_c_147_n 0.022351f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_108 N_C1_c_103_n N_B1_c_148_n 0.011021f $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_109 N_C1_c_104_n N_B1_c_148_n 0.00105611f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_110 N_C1_M1016_g N_A_29_368#_c_423_n 0.0149887f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_111 N_C1_M1017_g N_A_29_368#_c_423_n 0.0139961f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_112 N_C1_M1015_g N_Y_c_464_n 0.00159347f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_113 N_C1_M1015_g N_Y_c_465_n 0.0183358f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_114 N_C1_M1019_g N_Y_c_465_n 0.0168873f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_115 N_C1_c_103_n N_Y_c_465_n 0.025176f $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_116 N_C1_c_104_n N_Y_c_465_n 0.0020883f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_117 N_C1_M1016_g N_Y_c_482_n 0.0188125f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_118 N_C1_M1019_g N_Y_c_466_n 3.92313e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_119 N_C1_M1016_g N_Y_c_484_n 0.0173251f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_120 N_C1_M1017_g N_Y_c_484_n 0.0120614f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_121 N_C1_c_103_n N_Y_c_484_n 0.0212074f $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_122 N_C1_c_104_n N_Y_c_484_n 5.53536e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_123 N_C1_M1019_g N_Y_c_472_n 0.00253148f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_124 N_C1_M1015_g Y 0.0068844f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_125 N_C1_c_103_n Y 0.0293891f $X=0.75 $Y=1.515 $X2=0 $Y2=0
cc_126 N_C1_c_104_n Y 0.0175901f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_127 N_C1_M1016_g N_VPWR_c_615_n 0.00333926f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_128 N_C1_M1017_g N_VPWR_c_615_n 0.00333926f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_129 N_C1_M1016_g N_VPWR_c_611_n 0.00426394f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_130 N_C1_M1017_g N_VPWR_c_611_n 0.00422798f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_131 N_C1_M1015_g N_VGND_c_676_n 0.0139204f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_132 N_C1_M1019_g N_VGND_c_676_n 0.0109872f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_133 N_C1_M1015_g N_VGND_c_681_n 0.00383152f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_134 N_C1_M1019_g N_VGND_c_682_n 0.00383152f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_135 N_C1_M1015_g N_VGND_c_684_n 0.00761248f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_136 N_C1_M1019_g N_VGND_c_684_n 0.00757637f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B1_M1003_g N_B2_M1001_g 0.0179748f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B1_M1012_g N_B2_M1010_g 0.041604f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_139 N_B1_c_153_n N_B2_M1010_g 0.00422939f $X=1.51 $Y=1.95 $X2=0 $Y2=0
cc_140 N_B1_c_170_p N_B2_M1010_g 0.0167024f $X=2.525 $Y=2.035 $X2=0 $Y2=0
cc_141 N_B1_M1018_g N_B2_M1011_g 0.028262f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_142 N_B1_c_170_p N_B2_M1011_g 0.0159295f $X=2.525 $Y=2.035 $X2=0 $Y2=0
cc_143 N_B1_M1014_g N_B2_M1008_g 0.0209473f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_144 N_B1_c_153_n N_B2_c_245_n 0.00436071f $X=1.51 $Y=1.95 $X2=0 $Y2=0
cc_145 N_B1_c_170_p N_B2_c_245_n 0.0212727f $X=2.525 $Y=2.035 $X2=0 $Y2=0
cc_146 N_B1_c_147_n N_B2_c_245_n 2.42155e-19 $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_147 N_B1_c_148_n N_B2_c_245_n 0.0115507f $X=1.51 $Y=1.555 $X2=0 $Y2=0
cc_148 B1 N_B2_c_245_n 0.0190033f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B1_c_150_n N_B2_c_245_n 3.08121e-19 $X=2.85 $Y=1.515 $X2=0 $Y2=0
cc_150 N_B1_c_170_p N_B2_c_242_n 0.00160815f $X=2.525 $Y=2.035 $X2=0 $Y2=0
cc_151 N_B1_c_147_n N_B2_c_242_n 0.0228036f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_152 N_B1_c_148_n N_B2_c_242_n 0.00203997f $X=1.51 $Y=1.555 $X2=0 $Y2=0
cc_153 B1 N_B2_c_242_n 0.00772723f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_154 N_B1_c_150_n N_B2_c_242_n 0.039212f $X=2.85 $Y=1.515 $X2=0 $Y2=0
cc_155 N_B1_M1014_g N_A1_M1006_g 0.0167344f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_156 B1 N_A1_M1000_g 0.00202324f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B1_M1018_g N_A1_c_298_n 9.28333e-19 $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_158 B1 N_A1_c_298_n 0.0387978f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B1_c_150_n N_A1_c_298_n 2.02035e-19 $X=2.85 $Y=1.515 $X2=0 $Y2=0
cc_160 N_B1_M1018_g N_A1_c_309_n 6.29387e-19 $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_161 B1 N_A1_c_309_n 0.0156277f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_162 B1 N_A1_c_294_n 0.00413846f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_163 N_B1_c_150_n N_A1_c_294_n 0.0226f $X=2.85 $Y=1.515 $X2=0 $Y2=0
cc_164 N_B1_c_170_p N_A_29_368#_M1010_d 0.00314436f $X=2.525 $Y=2.035 $X2=0
+ $Y2=0
cc_165 B1 N_A_29_368#_M1018_d 0.00339717f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_166 N_B1_c_148_n N_A_29_368#_c_433_n 4.59812e-19 $X=1.51 $Y=1.555 $X2=0 $Y2=0
cc_167 N_B1_M1018_g N_A_29_368#_c_425_n 0.0144876f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_168 N_B1_M1012_g N_A_29_368#_c_427_n 0.0141334f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_169 N_B1_M1018_g N_A_29_368#_c_428_n 4.43424e-19 $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B1_M1003_g N_Y_c_466_n 3.92313e-19 $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B1_M1003_g N_Y_c_467_n 0.013957f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B1_M1014_g N_Y_c_467_n 0.0141288f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B1_c_147_n N_Y_c_467_n 0.00419315f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_174 N_B1_c_148_n N_Y_c_467_n 0.0241329f $X=1.51 $Y=1.555 $X2=0 $Y2=0
cc_175 B1 N_Y_c_467_n 0.0297803f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_176 N_B1_c_150_n N_Y_c_467_n 0.00313112f $X=2.85 $Y=1.515 $X2=0 $Y2=0
cc_177 N_B1_M1014_g N_Y_c_468_n 4.44013e-19 $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_178 B1 N_Y_c_469_n 0.00304394f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B1_c_147_n N_Y_c_472_n 3.85139e-19 $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_180 N_B1_c_148_n N_Y_c_472_n 0.0012413f $X=1.51 $Y=1.555 $X2=0 $Y2=0
cc_181 B1 N_Y_c_473_n 0.0162955f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_182 N_B1_c_150_n N_Y_c_473_n 0.00166767f $X=2.85 $Y=1.515 $X2=0 $Y2=0
cc_183 N_B1_c_153_n N_A_297_368#_M1012_s 0.00128176f $X=1.51 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_184 N_B1_c_170_p N_A_297_368#_M1012_s 0.00643972f $X=2.525 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_185 N_B1_c_215_p N_A_297_368#_M1012_s 5.67855e-19 $X=1.595 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_186 N_B1_c_170_p N_A_297_368#_M1011_s 0.00242374f $X=2.525 $Y=2.035 $X2=0
+ $Y2=0
cc_187 B1 N_A_297_368#_M1011_s 0.00260088f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B1_M1018_g N_A_297_368#_c_554_n 0.0117919f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_189 N_B1_c_170_p N_A_297_368#_c_554_n 0.0374777f $X=2.525 $Y=2.035 $X2=0
+ $Y2=0
cc_190 B1 N_A_297_368#_c_554_n 0.0475085f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_191 N_B1_c_150_n N_A_297_368#_c_554_n 3.74849e-19 $X=2.85 $Y=1.515 $X2=0
+ $Y2=0
cc_192 N_B1_M1012_g N_A_297_368#_c_566_n 0.0067764f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_193 N_B1_c_170_p N_A_297_368#_c_566_n 0.0125531f $X=2.525 $Y=2.035 $X2=0
+ $Y2=0
cc_194 N_B1_c_215_p N_A_297_368#_c_566_n 0.00674079f $X=1.595 $Y=2.035 $X2=0
+ $Y2=0
cc_195 N_B1_c_147_n N_A_297_368#_c_566_n 2.11515e-19 $X=1.41 $Y=1.515 $X2=0
+ $Y2=0
cc_196 N_B1_M1018_g N_VPWR_c_612_n 0.00340447f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_197 N_B1_M1012_g N_VPWR_c_615_n 0.00333926f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_198 N_B1_M1018_g N_VPWR_c_615_n 0.00349978f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_199 N_B1_M1012_g N_VPWR_c_611_n 0.00423187f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_200 N_B1_M1018_g N_VPWR_c_611_n 0.00434762f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_201 N_B1_M1003_g N_VGND_c_676_n 6.96322e-19 $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B1_M1014_g N_VGND_c_679_n 0.00433834f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B1_M1003_g N_VGND_c_682_n 0.00434272f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B1_M1003_g N_VGND_c_684_n 0.00821825f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B1_M1014_g N_VGND_c_684_n 0.00821519f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B1_M1003_g N_A_293_74#_c_752_n 0.00209548f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B1_M1003_g N_A_293_74#_c_750_n 0.00457794f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B1_M1014_g N_A_293_74#_c_754_n 0.0020603f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B1_M1014_g N_A_293_74#_c_751_n 0.00507972f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B2_M1011_g N_A_29_368#_c_425_n 0.0124097f $X=2.325 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B2_M1010_g N_A_29_368#_c_427_n 0.0109859f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_212 N_B2_M1011_g N_A_29_368#_c_428_n 0.00477264f $X=2.325 $Y=2.4 $X2=0 $Y2=0
cc_213 N_B2_M1001_g N_Y_c_467_n 0.0158392f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B2_M1008_g N_Y_c_467_n 0.0153251f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B2_c_245_n N_Y_c_467_n 0.0248845f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_216 N_B2_c_242_n N_Y_c_467_n 0.00568876f $X=2.325 $Y=1.515 $X2=0 $Y2=0
cc_217 N_B2_M1010_g N_A_297_368#_c_554_n 0.0103548f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_218 N_B2_M1011_g N_A_297_368#_c_554_n 0.00967619f $X=2.325 $Y=2.4 $X2=0 $Y2=0
cc_219 N_B2_M1010_g N_A_297_368#_c_566_n 0.00700376f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_220 N_B2_M1011_g N_A_297_368#_c_566_n 8.44031e-19 $X=2.325 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B2_M1010_g N_VPWR_c_615_n 0.00333926f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B2_M1011_g N_VPWR_c_615_n 0.00347303f $X=2.325 $Y=2.4 $X2=0 $Y2=0
cc_223 N_B2_M1010_g N_VPWR_c_611_n 0.00423076f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_224 N_B2_M1011_g N_VPWR_c_611_n 0.00428491f $X=2.325 $Y=2.4 $X2=0 $Y2=0
cc_225 N_B2_M1001_g N_VGND_c_677_n 0.00352921f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B2_M1008_g N_VGND_c_677_n 0.0041419f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B2_M1008_g N_VGND_c_679_n 0.00331f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B2_M1001_g N_VGND_c_682_n 0.00338063f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B2_M1001_g N_VGND_c_684_n 0.00441436f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B2_M1008_g N_VGND_c_684_n 0.00426874f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B2_M1001_g N_A_293_74#_c_754_n 0.0107174f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B2_M1008_g N_A_293_74#_c_754_n 0.0100699f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B2_M1001_g N_A_293_74#_c_751_n 5.73516e-19 $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B2_M1008_g N_A_293_74#_c_751_n 0.00660389f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1006_g N_A2_M1004_g 0.00761807f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1000_g N_A2_M1002_g 0.0321961f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A1_c_298_n N_A2_M1002_g 9.79029e-19 $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A1_c_316_p N_A2_M1002_g 0.0116236f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_239 N_A1_M1013_g N_A2_M1007_g 0.0207249f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A1_M1009_g N_A2_M1005_g 0.0309771f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A1_c_316_p N_A2_M1005_g 0.0133855f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_242 N_A1_c_300_n N_A2_M1005_g 0.00352898f $X=4.98 $Y=1.95 $X2=0 $Y2=0
cc_243 N_A1_c_298_n A2 0.0234621f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A1_c_316_p A2 0.0474282f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_245 N_A1_c_292_n A2 0.0255769f $X=4.98 $Y=1.78 $X2=0 $Y2=0
cc_246 N_A1_c_294_n A2 0.00282684f $X=3.745 $Y=1.515 $X2=0 $Y2=0
cc_247 N_A1_c_295_n A2 2.49009e-19 $X=5.14 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A1_c_298_n N_A2_c_373_n 2.31553e-19 $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A1_c_316_p N_A2_c_373_n 7.10058e-19 $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_250 N_A1_c_292_n N_A2_c_373_n 0.00280724f $X=4.98 $Y=1.78 $X2=0 $Y2=0
cc_251 N_A1_c_294_n N_A2_c_373_n 0.022927f $X=3.745 $Y=1.515 $X2=0 $Y2=0
cc_252 N_A1_c_295_n N_A2_c_373_n 0.0194633f $X=5.14 $Y=1.515 $X2=0 $Y2=0
cc_253 N_A1_M1006_g N_Y_c_468_n 4.43702e-19 $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A1_M1006_g N_Y_c_469_n 0.0194738f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A1_M1013_g N_Y_c_469_n 0.0151964f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A1_c_298_n N_Y_c_469_n 0.0262406f $X=3.57 $Y=1.515 $X2=0 $Y2=0
cc_257 N_A1_c_292_n N_Y_c_469_n 0.0136292f $X=4.98 $Y=1.78 $X2=0 $Y2=0
cc_258 A1 N_Y_c_469_n 0.030069f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_259 N_A1_c_294_n N_Y_c_469_n 0.0142629f $X=3.745 $Y=1.515 $X2=0 $Y2=0
cc_260 N_A1_c_295_n N_Y_c_469_n 0.00482041f $X=5.14 $Y=1.515 $X2=0 $Y2=0
cc_261 N_A1_M1013_g N_Y_c_470_n 0.00159319f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A1_c_316_p N_A_297_368#_M1000_d 0.00529615f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_263 N_A1_c_316_p N_A_297_368#_M1005_s 0.00555185f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_264 N_A1_c_300_n N_A_297_368#_M1005_s 0.00125604f $X=4.98 $Y=1.95 $X2=0 $Y2=0
cc_265 N_A1_M1000_g N_A_297_368#_c_554_n 0.0148021f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_266 N_A1_c_316_p N_A_297_368#_c_554_n 0.00467684f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_267 N_A1_c_309_n N_A_297_368#_c_554_n 0.0217353f $X=3.735 $Y=2.035 $X2=0
+ $Y2=0
cc_268 N_A1_c_294_n N_A_297_368#_c_554_n 0.00510021f $X=3.745 $Y=1.515 $X2=0
+ $Y2=0
cc_269 N_A1_c_316_p N_A_297_368#_c_581_n 0.0315971f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_270 N_A1_M1000_g N_A_297_368#_c_555_n 0.013595f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A1_c_316_p N_A_297_368#_c_555_n 0.0171986f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_272 N_A1_M1009_g N_A_297_368#_c_556_n 0.00994386f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A1_c_316_p N_A_297_368#_c_556_n 0.0178456f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_274 N_A1_c_298_n N_VPWR_M1000_s 0.0014039f $X=3.57 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_275 N_A1_c_309_n N_VPWR_M1000_s 0.00448191f $X=3.735 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A1_c_316_p N_VPWR_M1002_d 0.0031478f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_277 N_A1_M1000_g N_VPWR_c_612_n 0.00501904f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A1_M1009_g N_VPWR_c_614_n 0.00501904f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_279 A1 N_VPWR_c_614_n 0.0213917f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_280 N_A1_c_295_n N_VPWR_c_614_n 4.10279e-19 $X=5.14 $Y=1.515 $X2=0 $Y2=0
cc_281 N_A1_M1000_g N_VPWR_c_617_n 0.005209f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_282 N_A1_M1009_g N_VPWR_c_620_n 0.005209f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A1_M1000_g N_VPWR_c_611_n 0.00987509f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A1_M1009_g N_VPWR_c_611_n 0.0098656f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_285 N_A1_M1006_g N_VGND_c_679_n 0.00432706f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A1_M1013_g N_VGND_c_683_n 0.00433834f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A1_M1006_g N_VGND_c_684_n 0.00820461f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A1_M1013_g N_VGND_c_684_n 0.00825261f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A1_M1013_g N_A_675_74#_c_780_n 0.00219352f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A1_M1013_g N_A_675_74#_c_778_n 0.00581668f $X=5.05 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A1_M1006_g N_A_675_74#_c_779_n 0.00750072f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A2_M1004_g N_Y_c_469_n 0.0122883f $X=4.12 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A2_M1007_g N_Y_c_469_n 0.0114501f $X=4.62 $Y=0.74 $X2=0 $Y2=0
cc_294 A2 N_Y_c_469_n 0.0528884f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_295 N_A2_c_373_n N_Y_c_469_n 0.00638803f $X=4.645 $Y=1.515 $X2=0 $Y2=0
cc_296 N_A2_M1002_g N_A_297_368#_c_581_n 0.012696f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A2_M1005_g N_A_297_368#_c_581_n 0.012696f $X=4.645 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A2_M1002_g N_A_297_368#_c_555_n 0.00916709f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A2_M1005_g N_A_297_368#_c_555_n 5.64228e-19 $X=4.645 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A2_M1002_g N_A_297_368#_c_556_n 5.64228e-19 $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_301 N_A2_M1005_g N_A_297_368#_c_556_n 0.00916709f $X=4.645 $Y=2.4 $X2=0 $Y2=0
cc_302 N_A2_M1002_g N_VPWR_c_613_n 0.0027763f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A2_M1005_g N_VPWR_c_613_n 0.0027763f $X=4.645 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A2_M1002_g N_VPWR_c_617_n 0.005209f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A2_M1005_g N_VPWR_c_620_n 0.005209f $X=4.645 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A2_M1002_g N_VPWR_c_611_n 0.00982376f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_307 N_A2_M1005_g N_VPWR_c_611_n 0.00982376f $X=4.645 $Y=2.4 $X2=0 $Y2=0
cc_308 N_A2_M1004_g N_VGND_c_678_n 0.00304942f $X=4.12 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A2_M1007_g N_VGND_c_678_n 0.00298683f $X=4.62 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A2_M1004_g N_VGND_c_679_n 0.00338063f $X=4.12 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A2_M1007_g N_VGND_c_683_n 0.00338063f $X=4.62 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A2_M1004_g N_VGND_c_684_n 0.00443346f $X=4.12 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A2_M1007_g N_VGND_c_684_n 0.00440962f $X=4.62 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A2_M1004_g N_A_675_74#_c_783_n 0.0105237f $X=4.12 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A2_M1007_g N_A_675_74#_c_783_n 0.0105237f $X=4.62 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A2_M1007_g N_A_675_74#_c_778_n 3.24493e-19 $X=4.62 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A2_M1004_g N_A_675_74#_c_779_n 5.19636e-19 $X=4.12 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_29_368#_c_423_n N_Y_M1016_d 0.00165831f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_319 N_A_29_368#_M1016_s N_Y_c_475_n 0.00299921f $X=0.145 $Y=1.84 $X2=0 $Y2=0
cc_320 N_A_29_368#_c_422_n N_Y_c_475_n 0.0201299f $X=0.27 $Y=2.455 $X2=0 $Y2=0
cc_321 N_A_29_368#_c_423_n N_Y_c_484_n 0.0159318f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_322 N_A_29_368#_c_433_n N_Y_c_472_n 0.00574789f $X=1.17 $Y=2.015 $X2=0 $Y2=0
cc_323 N_A_29_368#_M1016_s Y 4.82655e-19 $X=0.145 $Y=1.84 $X2=0 $Y2=0
cc_324 N_A_29_368#_c_427_n N_A_297_368#_M1012_s 0.00197722f $X=2.015 $Y=2.852
+ $X2=-0.19 $Y2=1.66
cc_325 N_A_29_368#_c_425_n N_A_297_368#_M1011_s 0.00169972f $X=3 $Y=2.805 $X2=0
+ $Y2=0
cc_326 N_A_29_368#_M1010_d N_A_297_368#_c_554_n 0.00324479f $X=1.965 $Y=1.84
+ $X2=0 $Y2=0
cc_327 N_A_29_368#_M1018_d N_A_297_368#_c_554_n 0.00498276f $X=2.865 $Y=1.84
+ $X2=0 $Y2=0
cc_328 N_A_29_368#_c_427_n N_A_297_368#_c_554_n 0.00464895f $X=2.015 $Y=2.852
+ $X2=0 $Y2=0
cc_329 N_A_29_368#_c_428_n N_A_297_368#_c_554_n 0.0686462f $X=2.265 $Y=2.852
+ $X2=0 $Y2=0
cc_330 N_A_29_368#_c_427_n N_A_297_368#_c_566_n 0.0177055f $X=2.015 $Y=2.852
+ $X2=0 $Y2=0
cc_331 N_A_29_368#_c_425_n N_VPWR_c_612_n 0.0279004f $X=3 $Y=2.805 $X2=0 $Y2=0
cc_332 N_A_29_368#_c_423_n N_VPWR_c_615_n 0.0459191f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_333 N_A_29_368#_c_424_n N_VPWR_c_615_n 0.0179217f $X=0.355 $Y=2.99 $X2=0
+ $Y2=0
cc_334 N_A_29_368#_c_425_n N_VPWR_c_615_n 0.0372208f $X=3 $Y=2.805 $X2=0 $Y2=0
cc_335 N_A_29_368#_c_426_n N_VPWR_c_615_n 0.0121867f $X=1.17 $Y=2.99 $X2=0 $Y2=0
cc_336 N_A_29_368#_c_427_n N_VPWR_c_615_n 0.0650004f $X=2.015 $Y=2.852 $X2=0
+ $Y2=0
cc_337 N_A_29_368#_c_423_n N_VPWR_c_611_n 0.0258001f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_338 N_A_29_368#_c_424_n N_VPWR_c_611_n 0.00971942f $X=0.355 $Y=2.99 $X2=0
+ $Y2=0
cc_339 N_A_29_368#_c_425_n N_VPWR_c_611_n 0.0309148f $X=3 $Y=2.805 $X2=0 $Y2=0
cc_340 N_A_29_368#_c_426_n N_VPWR_c_611_n 0.00660921f $X=1.17 $Y=2.99 $X2=0
+ $Y2=0
cc_341 N_A_29_368#_c_427_n N_VPWR_c_611_n 0.0363998f $X=2.015 $Y=2.852 $X2=0
+ $Y2=0
cc_342 N_Y_c_465_n N_VGND_M1015_s 0.00197722f $X=1.09 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_343 N_Y_c_467_n N_VGND_M1001_d 0.00297264f $X=2.95 $Y=1.175 $X2=0 $Y2=0
cc_344 N_Y_c_469_n N_VGND_M1004_s 0.00251484f $X=5.18 $Y=1.175 $X2=0 $Y2=0
cc_345 N_Y_c_464_n N_VGND_c_676_n 0.0184513f $X=0.295 $Y=0.515 $X2=0 $Y2=0
cc_346 N_Y_c_465_n N_VGND_c_676_n 0.0187049f $X=1.09 $Y=1.095 $X2=0 $Y2=0
cc_347 N_Y_c_466_n N_VGND_c_676_n 0.0184077f $X=1.175 $Y=0.515 $X2=0 $Y2=0
cc_348 N_Y_c_468_n N_VGND_c_679_n 0.0101736f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_349 N_Y_c_464_n N_VGND_c_681_n 0.0112891f $X=0.295 $Y=0.515 $X2=0 $Y2=0
cc_350 N_Y_c_466_n N_VGND_c_682_n 0.00749631f $X=1.175 $Y=0.515 $X2=0 $Y2=0
cc_351 N_Y_c_470_n N_VGND_c_683_n 0.011066f $X=5.265 $Y=0.515 $X2=0 $Y2=0
cc_352 N_Y_c_464_n N_VGND_c_684_n 0.00934413f $X=0.295 $Y=0.515 $X2=0 $Y2=0
cc_353 N_Y_c_466_n N_VGND_c_684_n 0.0062048f $X=1.175 $Y=0.515 $X2=0 $Y2=0
cc_354 N_Y_c_468_n N_VGND_c_684_n 0.0084208f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_355 N_Y_c_470_n N_VGND_c_684_n 0.00915947f $X=5.265 $Y=0.515 $X2=0 $Y2=0
cc_356 N_Y_c_467_n N_A_293_74#_M1003_d 0.00218982f $X=2.95 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_357 N_Y_c_467_n N_A_293_74#_M1008_s 0.00176461f $X=2.95 $Y=1.175 $X2=0 $Y2=0
cc_358 N_Y_c_467_n N_A_293_74#_c_752_n 0.0183576f $X=2.95 $Y=1.175 $X2=0 $Y2=0
cc_359 N_Y_c_466_n N_A_293_74#_c_750_n 0.0149873f $X=1.175 $Y=0.515 $X2=0 $Y2=0
cc_360 N_Y_c_467_n N_A_293_74#_c_754_n 0.055652f $X=2.95 $Y=1.175 $X2=0 $Y2=0
cc_361 N_Y_c_468_n N_A_293_74#_c_751_n 0.0157199f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_362 N_Y_c_469_n N_A_675_74#_M1006_s 0.00625081f $X=5.18 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_363 N_Y_c_469_n N_A_675_74#_M1007_d 0.00176461f $X=5.18 $Y=1.175 $X2=0 $Y2=0
cc_364 N_Y_c_469_n N_A_675_74#_c_780_n 0.0151918f $X=5.18 $Y=1.175 $X2=0 $Y2=0
cc_365 N_Y_c_470_n N_A_675_74#_c_778_n 0.0148214f $X=5.265 $Y=0.515 $X2=0 $Y2=0
cc_366 N_Y_c_468_n N_A_675_74#_c_779_n 0.0247202f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_367 N_Y_c_469_n N_A_675_74#_c_779_n 0.0837462f $X=5.18 $Y=1.175 $X2=0 $Y2=0
cc_368 N_A_297_368#_c_554_n N_VPWR_M1000_s 0.00494201f $X=3.805 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_369 N_A_297_368#_c_581_n N_VPWR_M1002_d 0.00324075f $X=4.705 $Y=2.375 $X2=0
+ $Y2=0
cc_370 N_A_297_368#_c_554_n N_VPWR_c_612_n 0.0198097f $X=3.805 $Y=2.375 $X2=0
+ $Y2=0
cc_371 N_A_297_368#_c_555_n N_VPWR_c_612_n 0.0122069f $X=3.97 $Y=2.39 $X2=0
+ $Y2=0
cc_372 N_A_297_368#_c_581_n N_VPWR_c_613_n 0.0126919f $X=4.705 $Y=2.375 $X2=0
+ $Y2=0
cc_373 N_A_297_368#_c_555_n N_VPWR_c_613_n 0.0121684f $X=3.97 $Y=2.39 $X2=0
+ $Y2=0
cc_374 N_A_297_368#_c_556_n N_VPWR_c_613_n 0.0121684f $X=4.87 $Y=2.39 $X2=0
+ $Y2=0
cc_375 N_A_297_368#_c_556_n N_VPWR_c_614_n 0.0177747f $X=4.87 $Y=2.39 $X2=0
+ $Y2=0
cc_376 N_A_297_368#_c_555_n N_VPWR_c_617_n 0.0144776f $X=3.97 $Y=2.39 $X2=0
+ $Y2=0
cc_377 N_A_297_368#_c_556_n N_VPWR_c_620_n 0.0144776f $X=4.87 $Y=2.39 $X2=0
+ $Y2=0
cc_378 N_A_297_368#_c_555_n N_VPWR_c_611_n 0.0118404f $X=3.97 $Y=2.39 $X2=0
+ $Y2=0
cc_379 N_A_297_368#_c_556_n N_VPWR_c_611_n 0.0118404f $X=4.87 $Y=2.39 $X2=0
+ $Y2=0
cc_380 N_VGND_c_677_n N_A_293_74#_c_750_n 0.00158453f $X=2.11 $Y=0.495 $X2=0
+ $Y2=0
cc_381 N_VGND_c_682_n N_A_293_74#_c_750_n 0.0143793f $X=1.94 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_684_n N_A_293_74#_c_750_n 0.0119266f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_M1001_d N_A_293_74#_c_754_n 0.0057943f $X=1.935 $Y=0.37 $X2=0
+ $Y2=0
cc_384 N_VGND_c_677_n N_A_293_74#_c_754_n 0.0217251f $X=2.11 $Y=0.495 $X2=0
+ $Y2=0
cc_385 N_VGND_c_679_n N_A_293_74#_c_754_n 0.00189877f $X=4.2 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_682_n N_A_293_74#_c_754_n 0.00203359f $X=1.94 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_c_684_n N_A_293_74#_c_754_n 0.0088132f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_677_n N_A_293_74#_c_751_n 0.0110105f $X=2.11 $Y=0.495 $X2=0
+ $Y2=0
cc_389 N_VGND_c_679_n N_A_293_74#_c_751_n 0.0155998f $X=4.2 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_684_n N_A_293_74#_c_751_n 0.0119723f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_M1004_s N_A_675_74#_c_783_n 0.00472947f $X=4.195 $Y=0.37 $X2=0
+ $Y2=0
cc_392 N_VGND_c_678_n N_A_675_74#_c_783_n 0.0185765f $X=4.365 $Y=0.495 $X2=0
+ $Y2=0
cc_393 N_VGND_c_679_n N_A_675_74#_c_783_n 0.00203359f $X=4.2 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_683_n N_A_675_74#_c_783_n 0.00203359f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_684_n N_A_675_74#_c_783_n 0.00864073f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_678_n N_A_675_74#_c_778_n 0.00322188f $X=4.365 $Y=0.495 $X2=0
+ $Y2=0
cc_397 N_VGND_c_683_n N_A_675_74#_c_778_n 0.0142325f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_398 N_VGND_c_684_n N_A_675_74#_c_778_n 0.0109709f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_678_n N_A_675_74#_c_779_n 0.00335908f $X=4.365 $Y=0.495 $X2=0
+ $Y2=0
cc_400 N_VGND_c_679_n N_A_675_74#_c_779_n 0.032418f $X=4.2 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_684_n N_A_675_74#_c_779_n 0.0251588f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_402 N_A_293_74#_c_751_n N_A_675_74#_c_779_n 5.5809e-19 $X=2.615 $Y=0.495
+ $X2=0 $Y2=0

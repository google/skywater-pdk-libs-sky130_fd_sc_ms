* File: sky130_fd_sc_ms__and3_2.pex.spice
* Created: Wed Sep  2 11:57:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND3_2%A 1 3 5 8 10 11 12 16
c34 3 0 1.80268e-19 $X=0.575 $Y=2.34
r35 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=0.405 $X2=0.63 $Y2=0.405
r36 19 23 9.4417 $w=4.13e-07 $l=3.4e-07 $layer=LI1_cond $X=0.29 $Y=0.462
+ $X2=0.63 $Y2=0.462
r37 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=0.405 $X2=0.29 $Y2=0.405
r38 16 22 12.1753 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=0.515 $Y=0.405
+ $X2=0.655 $Y2=0.405
r39 16 18 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.515 $Y=0.405
+ $X2=0.29 $Y2=0.405
r40 11 12 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=0.462
+ $X2=1.2 $Y2=0.462
r41 11 23 2.49927 $w=4.13e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=0.462 $X2=0.63
+ $Y2=0.462
r42 10 19 1.38849 $w=4.13e-07 $l=5e-08 $layer=LI1_cond $X=0.24 $Y=0.462 $X2=0.29
+ $Y2=0.462
r43 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.59 $Y=1 $X2=0.59
+ $Y2=1.395
r44 5 22 20.0022 $w=1.5e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.59 $Y=0.57
+ $X2=0.655 $Y2=0.405
r45 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.59 $Y=0.57 $X2=0.59
+ $Y2=1
r46 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.575 $Y=1.485 $X2=0.575
+ $Y2=1.395
r47 1 3 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=0.575 $Y=1.485
+ $X2=0.575 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_2%B 3 7 8 9 13 15
c37 15 0 2.89246e-20 $X=1.07 $Y=1.43
c38 8 0 2.4843e-19 $X=1.2 $Y=1.295
c39 3 0 5.69497e-20 $X=1.145 $Y=2.34
r40 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.595
+ $X2=1.07 $Y2=1.76
r41 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.595
+ $X2=1.07 $Y2=1.43
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.595 $X2=1.07 $Y2=1.595
r43 9 14 1.96759 $w=4.08e-07 $l=7e-08 $layer=LI1_cond $X=1.11 $Y=1.665 $X2=1.11
+ $Y2=1.595
r44 8 14 8.43251 $w=4.08e-07 $l=3e-07 $layer=LI1_cond $X=1.11 $Y=1.295 $X2=1.11
+ $Y2=1.595
r45 7 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.16 $Y=1 $X2=1.16
+ $Y2=1.43
r46 3 16 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.145 $Y=2.34
+ $X2=1.145 $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_2%C 3 6 8 11 13
c38 8 0 5.69497e-20 $X=1.68 $Y=1.665
c39 6 0 1.80646e-19 $X=1.595 $Y=2.34
r40 11 14 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.645 $Y=1.595
+ $X2=1.645 $Y2=1.76
r41 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.645 $Y=1.595
+ $X2=1.645 $Y2=1.43
r42 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.595 $X2=1.65 $Y2=1.595
r43 6 14 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.595 $Y=2.34
+ $X2=1.595 $Y2=1.76
r44 3 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.55 $Y=1 $X2=1.55
+ $Y2=1.43
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_2%A_41_384# 1 2 3 12 16 20 24 27 30 34 37 39 43
+ 45 49 57
c95 49 0 1.15e-19 $X=2.22 $Y=1.505
c96 27 0 2.89246e-20 $X=0.35 $Y=1.95
r97 56 57 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.505
+ $X2=2.765 $Y2=1.505
r98 55 56 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.315 $Y=1.505
+ $X2=2.6 $Y2=1.505
r99 50 55 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.22 $Y=1.505
+ $X2=2.315 $Y2=1.505
r100 50 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.22 $Y=1.505
+ $X2=2.13 $Y2=1.505
r101 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.505 $X2=2.22 $Y2=1.505
r102 46 49 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.12 $Y=1.505
+ $X2=2.22 $Y2=1.505
r103 39 41 8.19036 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=0.362 $Y=1.09
+ $X2=0.362 $Y2=1.34
r104 36 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=1.67
+ $X2=2.12 $Y2=1.505
r105 36 37 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.12 $Y=1.67
+ $X2=2.12 $Y2=1.95
r106 35 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.37 $Y2=2.035
r107 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=2.12 $Y2=1.95
r108 34 35 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=1.535 $Y2=2.035
r109 31 43 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.035
+ $X2=0.35 $Y2=2.035
r110 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=1.37 $Y2=2.035
r111 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.205 $Y=2.035
+ $X2=0.515 $Y2=2.035
r112 27 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.95
+ $X2=0.35 $Y2=2.035
r113 27 41 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.35 $Y=1.95
+ $X2=0.35 $Y2=1.34
r114 22 57 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.67
+ $X2=2.765 $Y2=1.505
r115 22 24 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=2.765 $Y=1.67
+ $X2=2.765 $Y2=2.4
r116 18 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.34
+ $X2=2.6 $Y2=1.505
r117 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.6 $Y=1.34 $X2=2.6
+ $Y2=0.78
r118 14 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.67
+ $X2=2.315 $Y2=1.505
r119 14 16 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=2.315 $Y=1.67
+ $X2=2.315 $Y2=2.4
r120 10 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.34
+ $X2=2.13 $Y2=1.505
r121 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.13 $Y=1.34
+ $X2=2.13 $Y2=0.78
r122 3 45 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=1.235
+ $Y=1.92 $X2=1.37 $Y2=2.115
r123 2 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.205
+ $Y=1.92 $X2=0.35 $Y2=2.065
r124 1 39 182 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_NDIFF $count=1 $X=0.23
+ $Y=0.68 $X2=0.375 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_2%VPWR 1 2 3 14 18 20 22 27 28 29 35 40 44
r43 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 35 43 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.127 $Y2=3.33
r48 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.85 $Y2=3.33
r50 31 33 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 29 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 29 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 29 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 27 33 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.04 $Y2=3.33
r56 26 37 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.205 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=3.33
+ $X2=2.04 $Y2=3.33
r58 22 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.06 $Y=1.985
+ $X2=3.06 $Y2=2.815
r59 20 43 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.127 $Y2=3.33
r60 20 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.815
r61 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=3.245
+ $X2=2.04 $Y2=3.33
r62 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.04 $Y=3.245
+ $X2=2.04 $Y2=2.455
r63 12 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=3.33
r64 12 14 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=2.455
r65 3 25 400 $w=1.7e-07 $l=1.07261e-06 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.84 $X2=3.06 $Y2=2.815
r66 3 22 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.84 $X2=3.06 $Y2=1.985
r67 2 18 300 $w=1.7e-07 $l=6.90036e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=1.92 $X2=2.04 $Y2=2.455
r68 1 14 600 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.92 $X2=0.85 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_2%X 1 2 9 13 18 19 20
c39 18 0 1.12484e-19 $X=2.54 $Y=2.005
r40 20 24 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.64 $Y=0.99
+ $X2=2.345 $Y2=0.99
r41 18 19 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=2.005
+ $X2=2.55 $Y2=1.84
r42 15 20 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.17 $X2=2.64
+ $Y2=0.99
r43 15 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.64 $Y=1.17
+ $X2=2.64 $Y2=1.84
r44 11 18 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=2.55 $Y=2.015
+ $X2=2.55 $Y2=2.005
r45 11 13 26.3416 $w=3.48e-07 $l=8e-07 $layer=LI1_cond $X=2.55 $Y=2.015 $X2=2.55
+ $Y2=2.815
r46 7 24 1.2416 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=2.345 $Y=0.81 $X2=2.345
+ $Y2=0.99
r47 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.345 $Y=0.81
+ $X2=2.345 $Y2=0.555
r48 2 18 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.84 $X2=2.54 $Y2=2.005
r49 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=1.84 $X2=2.54 $Y2=2.815
r50 1 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.205
+ $Y=0.41 $X2=2.345 $Y2=1.005
r51 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.205
+ $Y=0.41 $X2=2.345 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__AND3_2%VGND 1 2 9 11 13 15 17 22 28 32
r37 31 34 11.4569 $w=5.91e-07 $l=5.55e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.02
+ $Y2=0.555
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r40 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.845
+ $Y2=0
r42 23 25 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.64
+ $Y2=0
r43 22 31 8.21944 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=3.02
+ $Y2=0
r44 22 25 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.64
+ $Y2=0
r45 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.845
+ $Y2=0
r47 17 19 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r48 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r49 15 20 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r50 15 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 11 34 4.30265 $w=5.91e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.085 $Y=0.64
+ $X2=3.02 $Y2=0.555
r52 11 13 13.1451 $w=3.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0.64
+ $X2=3.085 $Y2=1.005
r53 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0
r54 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0.555
r55 2 34 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.41 $X2=2.96 $Y2=0.555
r56 2 13 182 $w=1.7e-07 $l=7.43875e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.41 $X2=3.01 $Y2=1.005
r57 1 9 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=1.625 $Y=0.68
+ $X2=1.845 $Y2=0.555
.ends


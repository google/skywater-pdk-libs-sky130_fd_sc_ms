* File: sky130_fd_sc_ms__and4b_1.spice
* Created: Wed Sep  2 11:58:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4b_1.pex.spice"
.subckt sky130_fd_sc_ms__and4b_1  VNB VPB A_N B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_N_M1007_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.15675 PD=1.63 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 A_353_124# N_A_27_74#_M1003_g N_A_229_424#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.110562 AS=0.1824 PD=1.04 PS=1.85 NRD=22.068 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002 A=0.096 P=1.58 MULT=1
MM1001 A_448_139# N_B_M1001_g A_353_124# VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.110562 PD=0.88 PS=1.04 NRD=12.18 NRS=22.068 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 A_526_139# N_C_M1011_g A_448_139# VNB NLOWVT L=0.15 W=0.64 AD=0.1709
+ AS=0.0768 PD=1.275 PS=0.88 NRD=39.744 NRS=12.18 M=1 R=4.26667 SA=75001
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_526_139# VNB NLOWVT L=0.15 W=0.64
+ AD=0.144093 AS=0.1709 PD=1.08522 PS=1.275 NRD=14.988 NRS=39.744 M=1 R=4.26667
+ SA=75001.5 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_229_424#_M1005_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.166607 PD=2.05 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_27_74#_M1004_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90003.5 A=0.1512 P=2.04 MULT=1
MM1002 N_A_229_424#_M1002_d N_A_27_74#_M1002_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=0.84 AD=0.147 AS=0.1554 PD=1.19 PS=1.21 NRD=2.3443 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_229_424#_M1002_d VPB PSHORT L=0.18 W=0.84
+ AD=0.3738 AS=0.147 PD=1.73 PS=1.19 NRD=0 NRS=14.0658 M=1 R=4.66667 SA=90001.3
+ SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1009 N_A_229_424#_M1009_d N_C_M1009_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.3738 PD=1.16 PS=1.73 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90002.3
+ SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_229_424#_M1009_d VPB PSHORT L=0.18 W=0.84
+ AD=0.2028 AS=0.1344 PD=1.37143 PS=1.16 NRD=26.9693 NRS=0 M=1 R=4.66667
+ SA=90002.8 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1010 N_X_M1010_d N_A_229_424#_M1010_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2704 PD=2.8 PS=1.82857 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90002.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.224 P=13.68
*
.include "sky130_fd_sc_ms__and4b_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a221o_1.pxi.spice
* Created: Wed Sep  2 11:51:58 2020
* 
x_PM_SKY130_FD_SC_MS__A221O_1%A_148_260# N_A_148_260#_M1005_d
+ N_A_148_260#_M1003_d N_A_148_260#_M1006_d N_A_148_260#_M1000_g
+ N_A_148_260#_M1007_g N_A_148_260#_c_74_n N_A_148_260#_c_75_n
+ N_A_148_260#_c_76_n N_A_148_260#_c_77_n N_A_148_260#_c_78_n
+ N_A_148_260#_c_79_n N_A_148_260#_c_80_n N_A_148_260#_c_81_n
+ PM_SKY130_FD_SC_MS__A221O_1%A_148_260#
x_PM_SKY130_FD_SC_MS__A221O_1%A2 N_A2_c_159_n N_A2_M1001_g N_A2_c_160_n
+ N_A2_c_161_n N_A2_M1004_g A2 PM_SKY130_FD_SC_MS__A221O_1%A2
x_PM_SKY130_FD_SC_MS__A221O_1%A1 N_A1_M1002_g N_A1_M1005_g A1 N_A1_c_203_n
+ PM_SKY130_FD_SC_MS__A221O_1%A1
x_PM_SKY130_FD_SC_MS__A221O_1%B1 N_B1_M1010_g N_B1_M1008_g B1 N_B1_c_239_n
+ N_B1_c_240_n PM_SKY130_FD_SC_MS__A221O_1%B1
x_PM_SKY130_FD_SC_MS__A221O_1%B2 N_B2_M1009_g N_B2_M1011_g B2 N_B2_c_276_n
+ PM_SKY130_FD_SC_MS__A221O_1%B2
x_PM_SKY130_FD_SC_MS__A221O_1%C1 N_C1_M1003_g N_C1_c_312_n N_C1_M1006_g C1
+ N_C1_c_314_n N_C1_c_315_n PM_SKY130_FD_SC_MS__A221O_1%C1
x_PM_SKY130_FD_SC_MS__A221O_1%X N_X_M1007_s N_X_M1000_s N_X_c_338_n X X X
+ N_X_c_340_n N_X_c_339_n PM_SKY130_FD_SC_MS__A221O_1%X
x_PM_SKY130_FD_SC_MS__A221O_1%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_c_360_n
+ N_VPWR_c_361_n VPWR N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n
+ N_VPWR_c_359_n N_VPWR_c_366_n N_VPWR_c_367_n PM_SKY130_FD_SC_MS__A221O_1%VPWR
x_PM_SKY130_FD_SC_MS__A221O_1%A_313_392# N_A_313_392#_M1001_d
+ N_A_313_392#_M1010_d N_A_313_392#_c_405_n N_A_313_392#_c_406_n
+ N_A_313_392#_c_407_n N_A_313_392#_c_408_n
+ PM_SKY130_FD_SC_MS__A221O_1%A_313_392#
x_PM_SKY130_FD_SC_MS__A221O_1%A_509_392# N_A_509_392#_M1010_s
+ N_A_509_392#_M1011_d N_A_509_392#_c_438_n N_A_509_392#_c_439_n
+ N_A_509_392#_c_440_n N_A_509_392#_c_441_n
+ PM_SKY130_FD_SC_MS__A221O_1%A_509_392#
x_PM_SKY130_FD_SC_MS__A221O_1%VGND N_VGND_M1007_d N_VGND_M1009_d N_VGND_c_461_n
+ VGND N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n
+ N_VGND_c_466_n N_VGND_c_467_n PM_SKY130_FD_SC_MS__A221O_1%VGND
cc_1 VNB N_A_148_260#_M1000_g 0.00182816f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_2 VNB N_A_148_260#_M1007_g 0.0272723f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_148_260#_c_74_n 0.00606973f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_4 VNB N_A_148_260#_c_75_n 0.0146376f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.095
cc_5 VNB N_A_148_260#_c_76_n 0.00351237f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.52
cc_6 VNB N_A_148_260#_c_77_n 0.0155437f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=1.2
cc_7 VNB N_A_148_260#_c_78_n 0.016015f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.105
cc_8 VNB N_A_148_260#_c_79_n 0.0340198f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.465
cc_9 VNB N_A_148_260#_c_80_n 0.00697255f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.01
cc_10 VNB N_A_148_260#_c_81_n 0.018536f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=1.005
cc_11 VNB N_A2_c_159_n 0.0427169f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=0.395
cc_12 VNB N_A2_c_160_n 0.0278546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_161_n 0.0158993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2 0.00382554f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.63
cc_15 VNB N_A1_M1005_g 0.0360321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A1 0.00325885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_203_n 0.0280862f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_18 VNB N_B1_M1008_g 0.0314209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_239_n 0.0161022f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_20 VNB N_B1_c_240_n 0.00393964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B2_M1009_g 0.0312467f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=1.96
cc_22 VNB B2 0.00431791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_c_276_n 0.0162243f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_24 VNB N_C1_M1003_g 0.0117153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_312_n 0.00721267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_M1006_g 0.015492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_c_314_n 0.0650756f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_28 VNB N_C1_c_315_n 0.00655821f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_29 VNB N_X_c_338_n 0.0653482f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_30 VNB N_X_c_339_n 0.0329591f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.105
cc_31 VNB N_VPWR_c_359_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.465
cc_32 VNB N_VGND_c_461_n 0.00920632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_462_n 0.0397973f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_34 VNB N_VGND_c_463_n 0.0188832f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.105
cc_35 VNB N_VGND_c_464_n 0.269269f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.815
cc_36 VNB N_VGND_c_465_n 0.0294689f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.465
cc_37 VNB N_VGND_c_466_n 0.0280769f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.465
cc_38 VNB N_VGND_c_467_n 0.00711538f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.63
cc_39 VPB N_A_148_260#_M1000_g 0.0289433f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_40 VPB N_A_148_260#_c_78_n 0.0546103f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.105
cc_41 VPB N_A2_c_159_n 0.00605454f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=0.395
cc_42 VPB N_A2_M1001_g 0.0288679f $X=-0.19 $Y=1.66 $X2=3.915 $Y2=1.96
cc_43 VPB A2 0.00443472f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.63
cc_44 VPB N_A1_M1002_g 0.0281837f $X=-0.19 $Y=1.66 $X2=3.915 $Y2=1.96
cc_45 VPB A1 0.00258775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A1_c_203_n 0.0260758f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_47 VPB N_B1_M1010_g 0.0288619f $X=-0.19 $Y=1.66 $X2=3.915 $Y2=1.96
cc_48 VPB N_B1_c_239_n 0.0102925f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_49 VPB N_B1_c_240_n 0.00281847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B2_M1011_g 0.0225099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB B2 0.00411652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_B2_c_276_n 0.0117386f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_53 VPB N_C1_M1006_g 0.0367049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_X_c_340_n 0.0851171f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.105
cc_55 VPB N_X_c_339_n 0.0102058f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.105
cc_56 VPB N_VPWR_c_360_n 0.00872052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_361_n 0.0117473f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_58 VPB N_VPWR_c_362_n 0.0311089f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.095
cc_59 VPB N_VPWR_c_363_n 0.018048f $X=-0.19 $Y=1.66 $X2=3.86 $Y2=1.2
cc_60 VPB N_VPWR_c_364_n 0.052003f $X=-0.19 $Y=1.66 $X2=0.905 $Y2=1.465
cc_61 VPB N_VPWR_c_359_n 0.0771127f $X=-0.19 $Y=1.66 $X2=0.905 $Y2=1.465
cc_62 VPB N_VPWR_c_366_n 0.0047828f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.005
cc_63 VPB N_VPWR_c_367_n 0.0061274f $X=-0.19 $Y=1.66 $X2=4.037 $Y2=1.285
cc_64 VPB N_A_313_392#_c_405_n 0.00174321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_313_392#_c_406_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_313_392#_c_407_n 0.0134249f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_67 VPB N_A_313_392#_c_408_n 0.00399729f $X=-0.19 $Y=1.66 $X2=2.42 $Y2=1.095
cc_68 VPB N_A_509_392#_c_438_n 0.00564696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_509_392#_c_439_n 0.00529952f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_70 VPB N_A_509_392#_c_440_n 0.00391319f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_71 VPB N_A_509_392#_c_441_n 0.00184217f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_72 N_A_148_260#_M1000_g N_A2_c_159_n 0.00278253f $X=0.96 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_73 N_A_148_260#_M1007_g N_A2_c_159_n 0.0250238f $X=0.995 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_148_260#_c_74_n N_A2_c_159_n 0.0128633f $X=2.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A_148_260#_c_75_n N_A2_c_159_n 0.00598031f $X=1.205 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_148_260#_M1000_g N_A2_M1001_g 0.0271163f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_148_260#_c_74_n N_A2_c_160_n 0.0141544f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_78 N_A_148_260#_c_74_n N_A2_c_161_n 0.0103411f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_79 N_A_148_260#_c_76_n N_A2_c_161_n 0.00210649f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_80 N_A_148_260#_M1000_g A2 0.00237085f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A_148_260#_c_74_n A2 0.031704f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_82 N_A_148_260#_c_75_n A2 0.0233111f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_148_260#_c_79_n A2 2.39791e-19 $X=0.905 $Y=1.465 $X2=0 $Y2=0
cc_84 N_A_148_260#_c_74_n N_A1_M1005_g 0.0142322f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_85 N_A_148_260#_c_76_n N_A1_M1005_g 0.0109036f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_86 N_A_148_260#_c_80_n N_A1_M1005_g 0.00743095f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_87 N_A_148_260#_c_74_n A1 0.0161399f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_88 N_A_148_260#_c_74_n N_A1_c_203_n 0.00229257f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_89 N_A_148_260#_c_76_n N_B1_M1008_g 0.0107522f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_90 N_A_148_260#_c_77_n N_B1_M1008_g 0.0106483f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_91 N_A_148_260#_c_80_n N_B1_M1008_g 0.00634212f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_92 N_A_148_260#_c_80_n N_B1_c_239_n 0.00433744f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_93 N_A_148_260#_c_77_n N_B1_c_240_n 0.00888173f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_94 N_A_148_260#_c_80_n N_B1_c_240_n 0.0286449f $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_95 N_A_148_260#_c_76_n N_B2_M1009_g 0.00186941f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_96 N_A_148_260#_c_77_n N_B2_M1009_g 0.0143581f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_97 N_A_148_260#_c_78_n N_B2_M1009_g 5.28813e-19 $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_98 N_A_148_260#_c_80_n N_B2_M1009_g 5.21288e-19 $X=2.42 $Y=1.01 $X2=0 $Y2=0
cc_99 N_A_148_260#_c_81_n N_B2_M1009_g 6.52731e-19 $X=4.025 $Y=1.005 $X2=0 $Y2=0
cc_100 N_A_148_260#_c_78_n N_B2_M1011_g 0.00110831f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_101 N_A_148_260#_c_77_n B2 0.0392571f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_102 N_A_148_260#_c_78_n B2 0.0266398f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_103 N_A_148_260#_c_77_n N_B2_c_276_n 0.0044159f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_104 N_A_148_260#_c_78_n N_B2_c_276_n 2.58616e-19 $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_105 N_A_148_260#_c_77_n N_C1_M1003_g 0.0160911f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_106 N_A_148_260#_c_78_n N_C1_M1003_g 0.00196628f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_107 N_A_148_260#_c_81_n N_C1_M1003_g 0.00871597f $X=4.025 $Y=1.005 $X2=0
+ $Y2=0
cc_108 N_A_148_260#_c_78_n N_C1_c_312_n 0.00434931f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_109 N_A_148_260#_c_78_n N_C1_M1006_g 0.031427f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_110 N_A_148_260#_c_81_n N_C1_c_314_n 0.00152775f $X=4.025 $Y=1.005 $X2=0
+ $Y2=0
cc_111 N_A_148_260#_M1003_d N_C1_c_315_n 0.00226737f $X=3.885 $Y=0.615 $X2=0
+ $Y2=0
cc_112 N_A_148_260#_c_81_n N_C1_c_315_n 0.0229409f $X=4.025 $Y=1.005 $X2=0 $Y2=0
cc_113 N_A_148_260#_M1007_g N_X_c_338_n 0.00202121f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_148_260#_c_75_n N_X_c_338_n 0.0164255f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_115 N_A_148_260#_c_79_n N_X_c_338_n 9.8857e-19 $X=0.905 $Y=1.465 $X2=0 $Y2=0
cc_116 N_A_148_260#_M1000_g N_X_c_340_n 0.0180358f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_148_260#_c_75_n N_X_c_340_n 0.0122545f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_118 N_A_148_260#_c_79_n N_X_c_340_n 0.00101434f $X=0.905 $Y=1.465 $X2=0 $Y2=0
cc_119 N_A_148_260#_M1000_g N_X_c_339_n 0.00587143f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_148_260#_M1007_g N_X_c_339_n 0.00297287f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_148_260#_c_75_n N_X_c_339_n 0.0266447f $X=1.205 $Y=1.095 $X2=0 $Y2=0
cc_122 N_A_148_260#_c_79_n N_X_c_339_n 0.00233547f $X=0.905 $Y=1.465 $X2=0 $Y2=0
cc_123 N_A_148_260#_M1000_g N_VPWR_c_360_n 0.00309378f $X=0.96 $Y=2.4 $X2=0
+ $Y2=0
cc_124 N_A_148_260#_c_75_n N_VPWR_c_360_n 0.005852f $X=1.205 $Y=1.095 $X2=0
+ $Y2=0
cc_125 N_A_148_260#_M1000_g N_VPWR_c_362_n 0.005209f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_148_260#_c_78_n N_VPWR_c_364_n 0.014549f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_127 N_A_148_260#_M1000_g N_VPWR_c_359_n 0.00988094f $X=0.96 $Y=2.4 $X2=0
+ $Y2=0
cc_128 N_A_148_260#_c_78_n N_VPWR_c_359_n 0.0119743f $X=4.05 $Y=2.105 $X2=0
+ $Y2=0
cc_129 N_A_148_260#_c_77_n N_A_313_392#_c_408_n 0.00682195f $X=3.86 $Y=1.2 $X2=0
+ $Y2=0
cc_130 N_A_148_260#_c_78_n N_A_509_392#_c_439_n 0.00327031f $X=4.05 $Y=2.105
+ $X2=0 $Y2=0
cc_131 N_A_148_260#_c_78_n N_A_509_392#_c_441_n 0.0317724f $X=4.05 $Y=2.105
+ $X2=0 $Y2=0
cc_132 N_A_148_260#_c_74_n N_VGND_M1007_d 0.00740749f $X=2.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_148_260#_c_75_n N_VGND_M1007_d 8.62855e-19 $X=1.205 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_134 N_A_148_260#_c_77_n N_VGND_M1009_d 0.00228244f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_135 N_A_148_260#_c_76_n N_VGND_c_461_n 0.0196681f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_136 N_A_148_260#_c_77_n N_VGND_c_461_n 0.0265066f $X=3.86 $Y=1.2 $X2=0 $Y2=0
cc_137 N_A_148_260#_c_76_n N_VGND_c_462_n 0.0176208f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_138 N_A_148_260#_M1007_g N_VGND_c_464_n 0.00757924f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_148_260#_c_76_n N_VGND_c_464_n 0.0158894f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_140 N_A_148_260#_c_81_n N_VGND_c_464_n 0.0015257f $X=4.025 $Y=1.005 $X2=0
+ $Y2=0
cc_141 N_A_148_260#_M1007_g N_VGND_c_465_n 0.00383152f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_148_260#_M1007_g N_VGND_c_466_n 0.0170948f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_148_260#_c_74_n N_VGND_c_466_n 0.0567101f $X=2.42 $Y=1.095 $X2=0
+ $Y2=0
cc_144 N_A_148_260#_c_75_n N_VGND_c_466_n 0.00900333f $X=1.205 $Y=1.095 $X2=0
+ $Y2=0
cc_145 N_A_148_260#_c_76_n N_VGND_c_466_n 0.0169741f $X=2.64 $Y=0.52 $X2=0 $Y2=0
cc_146 N_A_148_260#_c_74_n A_417_79# 0.00366293f $X=2.42 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A2_c_159_n N_A1_M1005_g 0.00353069f $X=1.475 $Y=1.68 $X2=0 $Y2=0
cc_148 N_A2_c_161_n N_A1_M1005_g 0.0598892f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_149 A2 N_A1_M1005_g 0.00226541f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A2_c_160_n A1 5.06846e-19 $X=1.935 $Y=1.185 $X2=0 $Y2=0
cc_151 A2 A1 0.0250482f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_152 N_A2_c_159_n N_A1_c_203_n 0.0135515f $X=1.475 $Y=1.68 $X2=0 $Y2=0
cc_153 N_A2_M1001_g N_A1_c_203_n 0.0199788f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_154 N_A2_c_160_n N_A1_c_203_n 0.0171365f $X=1.935 $Y=1.185 $X2=0 $Y2=0
cc_155 A2 N_A1_c_203_n 0.00263634f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A2_M1001_g N_X_c_340_n 8.68815e-19 $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_157 N_A2_c_159_n N_VPWR_c_360_n 0.00221155f $X=1.475 $Y=1.68 $X2=0 $Y2=0
cc_158 N_A2_M1001_g N_VPWR_c_360_n 0.00723475f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_159 N_A2_M1001_g N_VPWR_c_361_n 5.51905e-19 $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_160 N_A2_M1001_g N_VPWR_c_363_n 0.005209f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_161 N_A2_M1001_g N_VPWR_c_359_n 0.00982736f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_162 N_A2_c_159_n N_A_313_392#_c_405_n 3.6687e-19 $X=1.475 $Y=1.68 $X2=0 $Y2=0
cc_163 N_A2_M1001_g N_A_313_392#_c_405_n 0.00273589f $X=1.475 $Y=2.46 $X2=0
+ $Y2=0
cc_164 A2 N_A_313_392#_c_405_n 0.0222779f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_A_313_392#_c_406_n 0.010224f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_166 N_A2_c_161_n N_VGND_c_462_n 0.00446421f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_167 N_A2_c_161_n N_VGND_c_464_n 0.00430282f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_168 N_A2_c_159_n N_VGND_c_466_n 0.00269777f $X=1.475 $Y=1.68 $X2=0 $Y2=0
cc_169 N_A2_c_161_n N_VGND_c_466_n 0.0158598f $X=2.01 $Y=1.11 $X2=0 $Y2=0
cc_170 N_A1_c_203_n N_B1_M1010_g 7.9776e-19 $X=2.37 $Y=1.635 $X2=0 $Y2=0
cc_171 N_A1_M1005_g N_B1_M1008_g 0.0176935f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_172 N_A1_M1005_g N_B1_c_239_n 0.0212847f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_173 A1 N_B1_c_239_n 2.50009e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A1_M1005_g N_B1_c_240_n 0.00303956f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_175 A1 N_B1_c_240_n 0.0201161f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A1_M1002_g N_VPWR_c_361_n 0.0137532f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_177 N_A1_M1002_g N_VPWR_c_363_n 0.00460063f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_178 N_A1_M1002_g N_VPWR_c_359_n 0.00908665f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_179 N_A1_M1002_g N_A_313_392#_c_405_n 2.38006e-19 $X=1.925 $Y=2.46 $X2=0
+ $Y2=0
cc_180 N_A1_M1002_g N_A_313_392#_c_407_n 0.0200282f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_181 A1 N_A_313_392#_c_407_n 0.0221682f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_182 N_A1_c_203_n N_A_313_392#_c_407_n 0.00810593f $X=2.37 $Y=1.635 $X2=0
+ $Y2=0
cc_183 N_A1_M1002_g N_A_509_392#_c_440_n 5.89323e-19 $X=1.925 $Y=2.46 $X2=0
+ $Y2=0
cc_184 N_A1_M1005_g N_VGND_c_462_n 0.00534051f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_185 N_A1_M1005_g N_VGND_c_464_n 0.00537853f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_186 N_A1_M1005_g N_VGND_c_466_n 0.00181914f $X=2.37 $Y=0.715 $X2=0 $Y2=0
cc_187 N_B1_M1008_g N_B2_M1009_g 0.0463342f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_188 N_B1_M1010_g N_B2_M1011_g 0.0279266f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_189 N_B1_c_239_n B2 4.06298e-19 $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_190 N_B1_c_240_n B2 0.0219204f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_191 N_B1_c_239_n N_B2_c_276_n 0.0463342f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_192 N_B1_c_240_n N_B2_c_276_n 4.06919e-19 $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_193 N_B1_M1010_g N_VPWR_c_361_n 8.96399e-19 $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_194 N_B1_M1010_g N_VPWR_c_364_n 0.00333926f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_195 N_B1_M1010_g N_VPWR_c_359_n 0.00427931f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_196 N_B1_M1010_g N_A_313_392#_c_407_n 0.0151751f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_197 N_B1_c_239_n N_A_313_392#_c_407_n 0.0031865f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_198 N_B1_c_240_n N_A_313_392#_c_407_n 0.0273703f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_199 N_B1_M1010_g N_A_313_392#_c_408_n 0.0160507f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_200 N_B1_c_240_n N_A_313_392#_c_408_n 0.0023921f $X=2.82 $Y=1.615 $X2=0 $Y2=0
cc_201 N_B1_M1010_g N_A_509_392#_c_439_n 0.01495f $X=2.895 $Y=2.46 $X2=0 $Y2=0
cc_202 N_B1_M1008_g N_VGND_c_461_n 0.00210079f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_203 N_B1_M1008_g N_VGND_c_462_n 0.00534051f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_204 N_B1_M1008_g N_VGND_c_464_n 0.00537853f $X=2.91 $Y=0.715 $X2=0 $Y2=0
cc_205 N_B2_M1011_g N_C1_M1006_g 0.0127441f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_206 B2 N_C1_M1006_g 0.0024298f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_207 N_B2_c_276_n N_C1_M1006_g 0.0195527f $X=3.36 $Y=1.615 $X2=0 $Y2=0
cc_208 N_B2_M1009_g N_C1_c_314_n 0.0241579f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_209 N_B2_M1011_g N_VPWR_c_364_n 0.00333926f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_210 N_B2_M1011_g N_VPWR_c_359_n 0.00423187f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_211 N_B2_M1011_g N_A_313_392#_c_408_n 0.0116181f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_212 B2 N_A_313_392#_c_408_n 0.00744682f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B2_c_276_n N_A_313_392#_c_408_n 0.00163439f $X=3.36 $Y=1.615 $X2=0
+ $Y2=0
cc_214 N_B2_M1011_g N_A_509_392#_c_439_n 0.013807f $X=3.345 $Y=2.46 $X2=0 $Y2=0
cc_215 B2 N_A_509_392#_c_441_n 0.0173356f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_216 N_B2_c_276_n N_A_509_392#_c_441_n 9.08531e-19 $X=3.36 $Y=1.615 $X2=0
+ $Y2=0
cc_217 N_B2_M1009_g N_VGND_c_461_n 0.0135704f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_218 N_B2_M1009_g N_VGND_c_462_n 0.00465077f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_219 N_B2_M1009_g N_VGND_c_464_n 0.00451796f $X=3.27 $Y=0.715 $X2=0 $Y2=0
cc_220 N_C1_M1006_g N_VPWR_c_364_n 0.005209f $X=3.825 $Y=2.46 $X2=0 $Y2=0
cc_221 N_C1_M1006_g N_VPWR_c_359_n 0.00987459f $X=3.825 $Y=2.46 $X2=0 $Y2=0
cc_222 N_C1_M1006_g N_A_509_392#_c_439_n 0.00324857f $X=3.825 $Y=2.46 $X2=0
+ $Y2=0
cc_223 N_C1_c_314_n N_VGND_c_461_n 0.0089245f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_224 N_C1_c_315_n N_VGND_c_461_n 0.0300657f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_225 N_C1_c_314_n N_VGND_c_463_n 0.0108828f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_226 N_C1_c_315_n N_VGND_c_463_n 0.0215843f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_227 N_C1_c_314_n N_VGND_c_464_n 0.0176737f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_228 N_C1_c_315_n N_VGND_c_464_n 0.0110944f $X=4.03 $Y=0.34 $X2=0 $Y2=0
cc_229 N_X_c_340_n N_VPWR_c_360_n 0.0385914f $X=0.735 $Y=1.985 $X2=0 $Y2=0
cc_230 N_X_c_340_n N_VPWR_c_362_n 0.0344053f $X=0.735 $Y=1.985 $X2=0 $Y2=0
cc_231 N_X_c_340_n N_VPWR_c_359_n 0.0284096f $X=0.735 $Y=1.985 $X2=0 $Y2=0
cc_232 N_X_c_338_n N_VGND_c_464_n 0.0273142f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_233 N_X_c_338_n N_VGND_c_465_n 0.0328875f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_234 N_X_c_338_n N_VGND_c_466_n 0.0205275f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_235 N_VPWR_c_360_n N_A_313_392#_c_405_n 0.00770452f $X=1.185 $Y=2.115 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_360_n N_A_313_392#_c_406_n 0.0289071f $X=1.185 $Y=2.115 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_361_n N_A_313_392#_c_406_n 0.0227494f $X=2.15 $Y=2.475 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_363_n N_A_313_392#_c_406_n 0.0109793f $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_359_n N_A_313_392#_c_406_n 0.00901959f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_VPWR_M1002_d N_A_313_392#_c_407_n 0.00455718f $X=2.015 $Y=1.96 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_361_n N_A_313_392#_c_407_n 0.0219767f $X=2.15 $Y=2.475 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_361_n N_A_509_392#_c_438_n 0.0452161f $X=2.15 $Y=2.475 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_364_n N_A_509_392#_c_439_n 0.0583239f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_359_n N_A_509_392#_c_439_n 0.0324477f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_361_n N_A_509_392#_c_440_n 0.0139f $X=2.15 $Y=2.475 $X2=0 $Y2=0
cc_246 N_VPWR_c_364_n N_A_509_392#_c_440_n 0.0200723f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_359_n N_A_509_392#_c_440_n 0.0108858f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_248 N_A_313_392#_c_407_n N_A_509_392#_M1010_s 0.00494823f $X=2.955 $Y=2.055
+ $X2=-0.19 $Y2=1.66
cc_249 N_A_313_392#_c_407_n N_A_509_392#_c_438_n 0.0198097f $X=2.955 $Y=2.055
+ $X2=0 $Y2=0
cc_250 N_A_313_392#_M1010_d N_A_509_392#_c_439_n 0.00165831f $X=2.985 $Y=1.96
+ $X2=0 $Y2=0
cc_251 N_A_313_392#_c_408_n N_A_509_392#_c_439_n 0.0159318f $X=3.12 $Y=2.115
+ $X2=0 $Y2=0
cc_252 N_A_313_392#_c_408_n N_A_509_392#_c_441_n 0.00725578f $X=3.12 $Y=2.115
+ $X2=0 $Y2=0

* File: sky130_fd_sc_ms__or4b_4.pex.spice
* Created: Fri Aug 28 18:09:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR4B_4%B 3 7 10 12 14 18 20 21 25 27 32 39
c71 18 0 1.33875e-19 $X=1.87 $Y=1.385
c72 10 0 1.72297e-19 $X=1.905 $Y=2.46
c73 3 0 1.47716e-19 $X=0.505 $Y=2.46
r74 26 32 4.8455 $w=4.38e-07 $l=1.85e-07 $layer=LI1_cond $X=0.43 $Y=1.33
+ $X2=0.615 $Y2=1.33
r75 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.385
+ $X2=0.43 $Y2=1.55
r76 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.385
+ $X2=0.43 $Y2=1.22
r77 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.385 $X2=0.43 $Y2=1.385
r78 21 39 7.52572 $w=4.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.33
+ $X2=0.835 $Y2=1.33
r79 21 32 2.75015 $w=4.38e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=1.33
+ $X2=0.615 $Y2=1.33
r80 20 26 4.97646 $w=4.38e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.33
+ $X2=0.43 $Y2=1.33
r81 18 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.385
+ $X2=1.87 $Y2=1.55
r82 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.87
+ $Y=1.385 $X2=1.87 $Y2=1.385
r83 14 17 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=1.195
+ $X2=1.87 $Y2=1.385
r84 12 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=1.195
+ $X2=1.87 $Y2=1.195
r85 12 39 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.705 $Y=1.195
+ $X2=0.835 $Y2=1.195
r86 10 31 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=1.905 $Y=2.46
+ $X2=1.905 $Y2=1.55
r87 7 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.22
r88 3 28 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.505 $Y=2.46
+ $X2=0.505 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%A 3 7 11 13 21
c45 11 0 1.72297e-19 $X=1.405 $Y=2.46
c46 3 0 1.95399e-19 $X=0.955 $Y=2.46
r47 19 21 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.405 $Y2=1.615
r48 17 19 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.065 $Y=1.615
+ $X2=1.17 $Y2=1.615
r49 15 17 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.955 $Y=1.615
+ $X2=1.065 $Y2=1.615
r50 13 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r51 9 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.78
+ $X2=1.405 $Y2=1.615
r52 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.405 $Y=1.78
+ $X2=1.405 $Y2=2.46
r53 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.45
+ $X2=1.065 $Y2=1.615
r54 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.065 $Y=1.45
+ $X2=1.065 $Y2=0.74
r55 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.78
+ $X2=0.955 $Y2=1.615
r56 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.955 $Y=1.78
+ $X2=0.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%C 3 6 10 12 13 15 16 18 21 23 28 34
c87 23 0 2.8262e-20 $X=2.41 $Y=1.22
c88 16 0 9.18809e-20 $X=4.08 $Y=1.295
c89 10 0 6.86532e-20 $X=3.805 $Y=2.46
c90 6 0 3.08277e-19 $X=2.405 $Y=2.46
r91 25 28 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.805 $Y=1.345
+ $X2=4.03 $Y2=1.345
r92 22 34 4.58497 $w=5.98e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=1.48
+ $X2=2.64 $Y2=1.48
r93 21 24 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.385
+ $X2=2.41 $Y2=1.55
r94 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.385
+ $X2=2.41 $Y2=1.22
r95 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.385 $X2=2.41 $Y2=1.385
r96 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.295
r97 16 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.345 $X2=4.03 $Y2=1.345
r98 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r99 13 18 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.295
+ $X2=2.64 $Y2=1.295
r100 12 15 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=4.08 $Y2=1.295
r101 12 13 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=2.785 $Y2=1.295
r102 8 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.51
+ $X2=3.805 $Y2=1.345
r103 8 10 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=3.805 $Y=1.51
+ $X2=3.805 $Y2=2.46
r104 6 24 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=2.405 $Y=2.46
+ $X2=2.405 $Y2=1.55
r105 3 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.32 $Y=0.74 $X2=2.32
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%A_563_48# 1 2 9 13 17 20 23 26 28 29 32 44
c91 44 0 2.89917e-19 $X=3.4 $Y=1.635
r92 43 44 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.355 $Y=1.635
+ $X2=3.4 $Y2=1.635
r93 39 41 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.89 $Y=1.635
+ $X2=2.905 $Y2=1.635
r94 38 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.34 $Y=1.635
+ $X2=3.355 $Y2=1.635
r95 38 41 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=1.635
+ $X2=2.905 $Y2=1.635
r96 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.34
+ $Y=1.635 $X2=3.34 $Y2=1.635
r97 32 34 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.59 $Y=1.985
+ $X2=4.59 $Y2=2.695
r98 30 32 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.59 $Y=1.89
+ $X2=4.59 $Y2=1.985
r99 29 37 13.3429 $w=3.68e-07 $l=3.51994e-07 $layer=LI1_cond $X=3.635 $Y=1.805
+ $X2=3.34 $Y2=1.68
r100 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.425 $Y=1.805
+ $X2=4.59 $Y2=1.89
r101 28 29 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.425 $Y=1.805
+ $X2=3.635 $Y2=1.805
r102 23 46 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.605 $Y=0.505
+ $X2=3.4 $Y2=0.505
r103 22 26 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=3.605 $Y=0.505
+ $X2=4.4 $Y2=0.505
r104 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.605
+ $Y=0.505 $X2=3.605 $Y2=0.505
r105 20 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.47
+ $X2=3.4 $Y2=1.635
r106 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=0.67
+ $X2=3.4 $Y2=0.505
r107 19 20 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.4 $Y=0.67 $X2=3.4
+ $Y2=1.47
r108 15 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.8
+ $X2=3.355 $Y2=1.635
r109 15 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.355 $Y=1.8
+ $X2=3.355 $Y2=2.46
r110 11 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.8
+ $X2=2.905 $Y2=1.635
r111 11 13 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.905 $Y=1.8
+ $X2=2.905 $Y2=2.46
r112 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.89 $Y=1.47
+ $X2=2.89 $Y2=1.635
r113 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.89 $Y=1.47 $X2=2.89
+ $Y2=0.74
r114 2 34 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.84 $X2=4.59 $Y2=2.695
r115 2 32 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.84 $X2=4.59 $Y2=1.985
r116 1 26 91 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.36 $X2=4.4 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%D_N 1 3 6 8 15
c38 1 0 5.98002e-20 $X=4.695 $Y=1.22
r39 14 15 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=4.695 $Y=1.385
+ $X2=4.815 $Y2=1.385
r40 11 14 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=4.65 $Y=1.385
+ $X2=4.695 $Y2=1.385
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.65
+ $Y=1.385 $X2=4.65 $Y2=1.385
r42 8 12 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=4.63 $Y=1.295 $X2=4.63
+ $Y2=1.385
r43 4 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.55
+ $X2=4.815 $Y2=1.385
r44 4 6 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=4.815 $Y=1.55
+ $X2=4.815 $Y2=2.34
r45 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.695 $Y=1.22
+ $X2=4.695 $Y2=1.385
r46 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.695 $Y=1.22
+ $X2=4.695 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%A_27_74# 1 2 3 4 15 19 23 27 31 35 37 39 43
+ 47 50 51 52 55 59 62 63 66 67 72 75 78 85
c192 63 0 1.67773e-19 $X=4.985 $Y=0.925
c193 62 0 9.69152e-20 $X=2.98 $Y=2.02
r194 93 94 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=6.25 $Y=1.485
+ $X2=6.275 $Y2=1.485
r195 90 91 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=5.775 $Y=1.485
+ $X2=5.8 $Y2=1.485
r196 89 90 63.2253 $w=3.24e-07 $l=4.25e-07 $layer=POLY_cond $X=5.35 $Y=1.485
+ $X2=5.775 $Y2=1.485
r197 82 85 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.98 $Y=2.105
+ $X2=3.13 $Y2=2.105
r198 80 81 9.78374 $w=3.73e-07 $l=2.05e-07 $layer=LI1_cond $X=3.082 $Y=0.925
+ $X2=3.082 $Y2=1.13
r199 77 78 10.0909 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0.645
+ $X2=2.2 $Y2=0.645
r200 73 93 38.679 $w=3.24e-07 $l=2.6e-07 $layer=POLY_cond $X=5.99 $Y=1.485
+ $X2=6.25 $Y2=1.485
r201 73 91 28.2654 $w=3.24e-07 $l=1.9e-07 $layer=POLY_cond $X=5.99 $Y=1.485
+ $X2=5.8 $Y2=1.485
r202 72 73 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.99
+ $Y=1.485 $X2=5.99 $Y2=1.485
r203 70 89 5.95062 $w=3.24e-07 $l=4e-08 $layer=POLY_cond $X=5.31 $Y=1.485
+ $X2=5.35 $Y2=1.485
r204 70 87 13.3889 $w=3.24e-07 $l=9e-08 $layer=POLY_cond $X=5.31 $Y=1.485
+ $X2=5.22 $Y2=1.485
r205 69 72 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.31 $Y=1.485
+ $X2=5.99 $Y2=1.485
r206 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.31
+ $Y=1.485 $X2=5.31 $Y2=1.485
r207 67 69 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.155 $Y=1.485
+ $X2=5.31 $Y2=1.485
r208 66 67 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.07 $Y=1.32
+ $X2=5.155 $Y2=1.485
r209 65 66 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.07 $Y=1.01
+ $X2=5.07 $Y2=1.32
r210 64 80 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.27 $Y=0.925
+ $X2=3.082 $Y2=0.925
r211 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.985 $Y=0.925
+ $X2=5.07 $Y2=1.01
r212 63 64 111.888 $w=1.68e-07 $l=1.715e-06 $layer=LI1_cond $X=4.985 $Y=0.925
+ $X2=3.27 $Y2=0.925
r213 62 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.02
+ $X2=2.98 $Y2=2.105
r214 62 81 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.98 $Y=2.02
+ $X2=2.98 $Y2=1.13
r215 57 59 7.83661 $w=3.73e-07 $l=2.55e-07 $layer=LI1_cond $X=3.082 $Y=0.77
+ $X2=3.082 $Y2=0.515
r216 55 80 2.15123 $w=3.73e-07 $l=7e-08 $layer=LI1_cond $X=3.082 $Y=0.855
+ $X2=3.082 $Y2=0.925
r217 55 57 2.6122 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=3.082 $Y=0.855
+ $X2=3.082 $Y2=0.77
r218 55 78 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.895 $Y=0.855
+ $X2=2.2 $Y2=0.855
r219 52 75 12.7264 $w=5.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.41 $Y=0.645
+ $X2=1.115 $Y2=0.645
r220 52 54 4.96677 $w=5.88e-07 $l=2.45e-07 $layer=LI1_cond $X=1.41 $Y=0.645
+ $X2=1.655 $Y2=0.645
r221 51 77 2.63543 $w=5.88e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=0.645
+ $X2=2.035 $Y2=0.645
r222 51 54 5.06813 $w=5.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.905 $Y=0.645
+ $X2=1.655 $Y2=0.645
r223 50 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.445 $Y=0.855
+ $X2=1.115 $Y2=0.855
r224 45 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.77
+ $X2=0.445 $Y2=0.855
r225 45 47 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.28 $Y=0.77
+ $X2=0.28 $Y2=0.515
r226 41 96 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.705 $Y=1.32
+ $X2=6.705 $Y2=1.485
r227 41 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.705 $Y=1.32
+ $X2=6.705 $Y2=0.74
r228 37 96 0.743827 $w=3.24e-07 $l=5e-09 $layer=POLY_cond $X=6.7 $Y=1.485
+ $X2=6.705 $Y2=1.485
r229 37 94 63.2253 $w=3.24e-07 $l=4.25e-07 $layer=POLY_cond $X=6.7 $Y=1.485
+ $X2=6.275 $Y2=1.485
r230 37 39 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=6.7 $Y=1.635
+ $X2=6.7 $Y2=2.4
r231 33 94 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.275 $Y=1.32
+ $X2=6.275 $Y2=1.485
r232 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.275 $Y=1.32
+ $X2=6.275 $Y2=0.74
r233 29 93 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.65
+ $X2=6.25 $Y2=1.485
r234 29 31 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.25 $Y=1.65
+ $X2=6.25 $Y2=2.4
r235 25 91 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=1.65
+ $X2=5.8 $Y2=1.485
r236 25 27 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.8 $Y=1.65 $X2=5.8
+ $Y2=2.4
r237 21 90 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=1.32
+ $X2=5.775 $Y2=1.485
r238 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.775 $Y=1.32
+ $X2=5.775 $Y2=0.74
r239 17 89 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.35 $Y=1.65
+ $X2=5.35 $Y2=1.485
r240 17 19 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.35 $Y=1.65
+ $X2=5.35 $Y2=2.4
r241 13 87 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.22 $Y=1.32
+ $X2=5.22 $Y2=1.485
r242 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.22 $Y=1.32
+ $X2=5.22 $Y2=0.74
r243 4 85 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.995
+ $Y=1.96 $X2=3.13 $Y2=2.105
r244 3 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.965
+ $Y=0.37 $X2=3.105 $Y2=0.515
r245 2 77 91 $w=1.7e-07 $l=9.6478e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=2.035 $Y2=0.515
r246 2 54 45.5 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_NDIFF $count=4 $X=1.14
+ $Y=0.37 $X2=1.655 $Y2=0.515
r247 1 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%A_27_392# 1 2 3 10 12 14 16 17 20 22 26 30 36
+ 37
c71 22 0 9.00629e-20 $X=3.945 $Y=2.445
c72 20 0 1.72297e-19 $X=2.18 $Y=2.815
c73 16 0 1.33875e-19 $X=2.18 $Y=2.12
c74 10 0 4.76839e-20 $X=0.28 $Y=2.12
r75 28 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.53 $X2=4.07
+ $Y2=2.445
r76 28 30 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.07 $Y=2.53
+ $X2=4.07 $Y2=2.815
r77 24 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.36 $X2=4.07
+ $Y2=2.445
r78 24 26 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=4.07 $Y=2.36
+ $X2=4.07 $Y2=2.225
r79 23 36 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.445
+ $X2=2.18 $Y2=2.445
r80 22 37 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=2.445
+ $X2=4.07 $Y2=2.445
r81 22 23 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=3.945 $Y=2.445
+ $X2=2.345 $Y2=2.445
r82 18 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.53 $X2=2.18
+ $Y2=2.445
r83 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.18 $Y=2.53
+ $X2=2.18 $Y2=2.815
r84 17 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.36 $X2=2.18
+ $Y2=2.445
r85 16 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.12 $X2=2.18
+ $Y2=2.035
r86 16 17 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.18 $Y=2.12 $X2=2.18
+ $Y2=2.36
r87 15 33 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.03
r88 14 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.18 $Y2=2.035
r89 14 15 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=0.445 $Y2=2.035
r90 10 33 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.03
r91 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r92 3 30 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.96 $X2=4.03 $Y2=2.815
r93 3 26 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.96 $X2=4.03 $Y2=2.225
r94 2 35 400 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.96 $X2=2.18 $Y2=2.115
r95 2 20 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.96 $X2=2.18 $Y2=2.815
r96 1 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
r97 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%A_119_392# 1 2 9 14 16
c20 16 0 3.0476e-19 $X=1.68 $Y=2.455
c21 14 0 2.95431e-19 $X=0.73 $Y=2.455
r22 10 14 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.375
+ $X2=0.73 $Y2=2.375
r23 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=1.68 $Y2=2.375
r24 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.515 $Y=2.375
+ $X2=0.815 $Y2=2.375
r25 2 16 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.96 $X2=1.68 $Y2=2.455
r26 1 14 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%VPWR 1 2 3 4 15 19 25 27 29 31 33 38 43 48 54
+ 57 60 64
r90 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r92 57 58 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r94 52 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r95 52 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r96 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r97 49 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.025 $Y2=3.33
r98 49 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.48 $Y2=3.33
r99 48 63 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=6.76 $Y=3.33 $X2=6.98
+ $Y2=3.33
r100 48 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r102 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r104 44 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.085 $Y2=3.33
r105 44 46 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 43 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=6.025 $Y2=3.33
r107 43 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 41 42 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r111 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 38 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=5.085 $Y2=3.33
r113 38 41 213.989 $w=1.68e-07 $l=3.28e-06 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 33 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r117 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 31 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 31 42 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 27 63 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=6.925 $Y=3.245
+ $X2=6.98 $Y2=3.33
r121 27 29 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.925 $Y=3.245
+ $X2=6.925 $Y2=2.405
r122 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=3.245
+ $X2=6.025 $Y2=3.33
r123 23 25 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=6.025 $Y=3.245
+ $X2=6.025 $Y2=2.405
r124 19 22 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.085 $Y=1.985
+ $X2=5.085 $Y2=2.815
r125 17 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=3.245
+ $X2=5.085 $Y2=3.33
r126 17 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.085 $Y=3.245
+ $X2=5.085 $Y2=2.815
r127 13 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r128 13 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.805
r129 4 29 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=6.79
+ $Y=1.84 $X2=6.925 $Y2=2.405
r130 3 25 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=5.89
+ $Y=1.84 $X2=6.025 $Y2=2.405
r131 2 22 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.84 $X2=5.125 $Y2=2.815
r132 2 19 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=4.905
+ $Y=1.84 $X2=5.125 $Y2=1.985
r133 1 15 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.96 $X2=1.18 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%A_499_392# 1 2 11
c12 11 0 1.75814e-19 $X=3.58 $Y=2.8
r13 8 11 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=2.68 $Y=2.84 $X2=3.58
+ $Y2=2.84
r14 2 11 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.96 $X2=3.58 $Y2=2.8
r15 1 8 600 $w=1.7e-07 $l=9.27901e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.96 $X2=2.68 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%X 1 2 3 4 15 17 19 21 22 23 27 33 36 39 40 41
+ 42 43
c75 42 0 4.99714e-20 $X=6.48 $Y=2.035
c76 36 0 1.8329e-19 $X=6.51 $Y=1.82
r77 43 46 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.96 $Y=1.985
+ $X2=6.655 $Y2=1.985
r78 42 46 2.3561 $w=3.3e-07 $l=1.48e-07 $layer=LI1_cond $X=6.507 $Y=1.985
+ $X2=6.655 $Y2=1.985
r79 40 41 7.00677 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.49 $Y=1.3 $X2=6.49
+ $Y2=1.47
r80 36 42 3.80668 $w=2.9e-07 $l=1.66493e-07 $layer=LI1_cond $X=6.51 $Y=1.82
+ $X2=6.507 $Y2=1.985
r81 36 41 13.9088 $w=2.88e-07 $l=3.5e-07 $layer=LI1_cond $X=6.51 $Y=1.82
+ $X2=6.51 $Y2=1.47
r82 31 42 3.80668 $w=2.3e-07 $l=1.80291e-07 $layer=LI1_cond $X=6.475 $Y=2.15
+ $X2=6.507 $Y2=1.985
r83 31 33 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.475 $Y=2.15
+ $X2=6.475 $Y2=2.4
r84 29 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=1.15 $X2=6.45
+ $Y2=1.065
r85 29 40 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=6.45 $Y=1.15
+ $X2=6.45 $Y2=1.3
r86 25 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=0.98 $X2=6.45
+ $Y2=1.065
r87 25 27 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=6.45 $Y=0.98
+ $X2=6.45 $Y2=0.515
r88 24 38 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=5.69 $Y=1.985 $X2=5.55
+ $Y2=1.985
r89 23 42 2.3561 $w=3.3e-07 $l=1.47e-07 $layer=LI1_cond $X=6.36 $Y=1.985
+ $X2=6.507 $Y2=1.985
r90 23 24 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=6.36 $Y=1.985
+ $X2=5.69 $Y2=1.985
r91 21 39 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.325 $Y=1.065
+ $X2=6.45 $Y2=1.065
r92 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.325 $Y=1.065
+ $X2=5.655 $Y2=1.065
r93 17 38 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.55 $Y=2.15
+ $X2=5.55 $Y2=1.985
r94 17 19 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=5.55 $Y=2.15
+ $X2=5.55 $Y2=2.4
r95 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.49 $Y=0.98
+ $X2=5.655 $Y2=1.065
r96 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.49 $Y=0.98
+ $X2=5.49 $Y2=0.515
r97 4 42 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.34
+ $Y=1.84 $X2=6.475 $Y2=1.985
r98 4 33 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=6.34
+ $Y=1.84 $X2=6.475 $Y2=2.4
r99 3 38 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=1.84 $X2=5.575 $Y2=1.985
r100 3 19 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.84 $X2=5.575 $Y2=2.4
r101 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.35
+ $Y=0.37 $X2=6.49 $Y2=0.515
r102 1 15 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.37 $X2=5.49 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 51
+ 59 64 70 73 76 79 83
r83 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r84 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r85 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r86 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r87 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r88 68 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r89 68 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r91 65 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=5.99
+ $Y2=0
r92 65 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.48
+ $Y2=0
r93 64 82 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r94 64 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r95 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r96 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r97 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r98 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=4.99
+ $Y2=0
r99 60 62 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.52
+ $Y2=0
r100 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0 $X2=5.99
+ $Y2=0
r101 59 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.52 $Y2=0
r102 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r103 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r104 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r105 54 57 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r106 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r107 52 73 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=2.547 $Y2=0
r108 52 54 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=3.12 $Y2=0
r109 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.99
+ $Y2=0
r110 51 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.56 $Y2=0
r111 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r112 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r113 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r115 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r116 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r118 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r119 43 73 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.547
+ $Y2=0
r120 43 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.16
+ $Y2=0
r121 41 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r124 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r125 36 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r126 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r127 32 82 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r128 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r129 28 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0
r130 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.99 $Y=0.085
+ $X2=5.99 $Y2=0.58
r131 24 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0
r132 24 26 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0.55
r133 20 73 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.547 $Y=0.085
+ $X2=2.547 $Y2=0
r134 20 22 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=2.547 $Y=0.085
+ $X2=2.547 $Y2=0.515
r135 16 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r136 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.515
r137 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.78
+ $Y=0.37 $X2=6.92 $Y2=0.515
r138 4 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.85
+ $Y=0.37 $X2=5.99 $Y2=0.58
r139 3 26 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.47 $X2=4.99 $Y2=0.55
r140 2 22 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.37 $X2=2.545 $Y2=0.515
r141 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__clkinv_4.spice
* Created: Wed Sep  2 12:01:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkinv_4.pex.spice"
.subckt sky130_fd_sc_ms__clkinv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.14805 AS=0.3066 PD=1.125 PS=2.3 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.7
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.14805 AS=0.0882 PD=1.125 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.5
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.06405 AS=0.0882 PD=0.725 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1008_d N_A_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.06405 AS=0.1386 PD=0.725 PS=1.5 NRD=7.14 NRS=12.852 M=1 R=2.8 SA=75002.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90002.5
+ A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6 SB=90002.1
+ A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90001.6
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5 SB=90001.2
+ A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.5 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__clkinv_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__and3_4.spice
* Created: Fri Aug 28 17:12:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and3_4.pex.spice"
.subckt sky130_fd_sc_ms__and3_4  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_83_260#_M1011_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_83_260#_M1015_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1015_d N_A_83_260#_M1017_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_83_260#_M1018_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.133522 AS=0.1036 PD=1.16899 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1009 N_A_489_74#_M1009_d N_C_M1009_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.115478 PD=0.92 PS=1.01101 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_489_74#_M1009_d N_C_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_686_74#_M1000_d N_B_M1000_g N_A_489_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1024 PD=1.85 PS=0.96 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_686_74#_M1002_d N_B_M1002_g N_A_489_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75000.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1010 N_A_83_260#_M1010_d N_A_M1010_g N_A_686_74#_M1002_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1184 AS=0.0896 PD=1.01 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_83_260#_M1010_d N_A_M1019_g N_A_686_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1184 AS=0.2144 PD=1.01 PS=1.95 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_83_260#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004.1 A=0.2016 P=2.6 MULT=1
MM1004 N_X_M1003_d N_A_83_260#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1005_d N_A_83_260#_M1005_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.2
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1005_d N_A_83_260#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2176 PD=1.39 PS=1.70286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.6 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1007 N_A_83_260#_M1007_d N_C_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1632 PD=1.11 PS=1.27714 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90002.2 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1008 N_A_83_260#_M1007_d N_C_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2604 PD=1.11 PS=1.46 NRD=0 NRS=0 M=1 R=4.66667 SA=90002.6
+ SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1008_s N_B_M1001_g N_A_83_260#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2604 AS=0.1302 PD=1.46 PS=1.15 NRD=0 NRS=0 M=1 R=4.66667 SA=90003.4
+ SB=90001.7 A=0.1512 P=2.04 MULT=1
MM1013 N_VPWR_M1013_d N_B_M1013_g N_A_83_260#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1386 AS=0.1302 PD=1.17 PS=1.15 NRD=1.1623 NRS=8.1952 M=1 R=4.66667
+ SA=90003.9 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1012 N_A_83_260#_M1012_d N_A_M1012_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1386 PD=1.11 PS=1.17 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90004.4
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1016 N_A_83_260#_M1012_d N_A_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2772 PD=1.11 PS=2.34 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90004.9
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
c_57 VNB 0 1.52826e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__and3_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__and3_4.pxi.spice
* Created: Wed Sep  2 11:57:51 2020
* 
x_PM_SKY130_FD_SC_MS__AND3_4%A_83_260# N_A_83_260#_M1010_d N_A_83_260#_M1007_d
+ N_A_83_260#_M1001_s N_A_83_260#_M1012_d N_A_83_260#_M1003_g
+ N_A_83_260#_M1011_g N_A_83_260#_M1015_g N_A_83_260#_M1004_g
+ N_A_83_260#_M1017_g N_A_83_260#_M1005_g N_A_83_260#_M1018_g
+ N_A_83_260#_M1006_g N_A_83_260#_c_115_n N_A_83_260#_c_116_n
+ N_A_83_260#_c_127_n N_A_83_260#_c_193_p N_A_83_260#_c_128_n
+ N_A_83_260#_c_129_n N_A_83_260#_c_130_n N_A_83_260#_c_131_n
+ N_A_83_260#_c_117_n N_A_83_260#_c_132_n N_A_83_260#_c_118_n
+ N_A_83_260#_c_119_n N_A_83_260#_c_133_n N_A_83_260#_c_120_n
+ N_A_83_260#_c_135_n N_A_83_260#_c_136_n N_A_83_260#_c_172_p
+ N_A_83_260#_c_121_n PM_SKY130_FD_SC_MS__AND3_4%A_83_260#
x_PM_SKY130_FD_SC_MS__AND3_4%C N_C_M1009_g N_C_M1007_g N_C_M1014_g N_C_M1008_g C
+ C N_C_c_281_n PM_SKY130_FD_SC_MS__AND3_4%C
x_PM_SKY130_FD_SC_MS__AND3_4%B N_B_M1001_g N_B_M1000_g N_B_M1013_g N_B_M1002_g B
+ B N_B_c_338_n N_B_c_339_n PM_SKY130_FD_SC_MS__AND3_4%B
x_PM_SKY130_FD_SC_MS__AND3_4%A N_A_M1010_g N_A_c_396_n N_A_M1012_g N_A_c_397_n
+ N_A_M1016_g N_A_M1019_g A N_A_c_395_n PM_SKY130_FD_SC_MS__AND3_4%A
x_PM_SKY130_FD_SC_MS__AND3_4%VPWR N_VPWR_M1003_s N_VPWR_M1004_s N_VPWR_M1006_s
+ N_VPWR_M1008_s N_VPWR_M1013_d N_VPWR_M1016_s N_VPWR_c_447_n N_VPWR_c_448_n
+ N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n VPWR N_VPWR_c_456_n N_VPWR_c_457_n
+ N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n
+ N_VPWR_c_463_n N_VPWR_c_446_n PM_SKY130_FD_SC_MS__AND3_4%VPWR
x_PM_SKY130_FD_SC_MS__AND3_4%X N_X_M1011_s N_X_M1017_s N_X_M1003_d N_X_M1005_d
+ N_X_c_528_n N_X_c_533_n N_X_c_529_n N_X_c_534_n X X X X X X X X X
+ PM_SKY130_FD_SC_MS__AND3_4%X
x_PM_SKY130_FD_SC_MS__AND3_4%VGND N_VGND_M1011_d N_VGND_M1015_d N_VGND_M1018_d
+ N_VGND_M1014_s N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n
+ N_VGND_c_600_n VGND N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n
+ N_VGND_c_604_n N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n
+ PM_SKY130_FD_SC_MS__AND3_4%VGND
x_PM_SKY130_FD_SC_MS__AND3_4%A_489_74# N_A_489_74#_M1009_d N_A_489_74#_M1000_s
+ N_A_489_74#_c_668_n N_A_489_74#_c_669_n N_A_489_74#_c_670_n
+ N_A_489_74#_c_683_n PM_SKY130_FD_SC_MS__AND3_4%A_489_74#
x_PM_SKY130_FD_SC_MS__AND3_4%A_686_74# N_A_686_74#_M1000_d N_A_686_74#_M1002_d
+ N_A_686_74#_M1019_s N_A_686_74#_c_699_n N_A_686_74#_c_700_n
+ N_A_686_74#_c_701_n N_A_686_74#_c_702_n N_A_686_74#_c_703_n
+ N_A_686_74#_c_704_n N_A_686_74#_c_705_n PM_SKY130_FD_SC_MS__AND3_4%A_686_74#
cc_1 VNB N_A_83_260#_M1003_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_260#_M1011_g 0.0260209f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_3 VNB N_A_83_260#_M1015_g 0.0217361f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_4 VNB N_A_83_260#_M1004_g 0.00164813f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_5 VNB N_A_83_260#_M1017_g 0.0217567f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_6 VNB N_A_83_260#_M1005_g 0.00165414f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_7 VNB N_A_83_260#_M1018_g 0.0217125f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_8 VNB N_A_83_260#_M1006_g 0.00168415f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_9 VNB N_A_83_260#_c_115_n 0.00583139f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.465
cc_10 VNB N_A_83_260#_c_116_n 4.80171e-19 $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.95
cc_11 VNB N_A_83_260#_c_117_n 0.00138548f $X=-0.19 $Y=-0.245 $X2=4.975 $Y2=0.76
cc_12 VNB N_A_83_260#_c_118_n 0.0142609f $X=-0.19 $Y=-0.245 $X2=5.455 $Y2=1.195
cc_13 VNB N_A_83_260#_c_119_n 0.00504352f $X=-0.19 $Y=-0.245 $X2=5.14 $Y2=1.195
cc_14 VNB N_A_83_260#_c_120_n 0.0181243f $X=-0.19 $Y=-0.245 $X2=5.54 $Y2=1.95
cc_15 VNB N_A_83_260#_c_121_n 0.10247f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.465
cc_16 VNB N_C_M1009_g 0.0350062f $X=-0.19 $Y=-0.245 $X2=3.845 $Y2=2.12
cc_17 VNB N_C_M1014_g 0.0428859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB C 0.00209752f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_19 VNB N_C_c_281_n 0.0427034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1000_g 0.0352995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_M1002_g 0.0277135f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_22 VNB N_B_c_338_n 0.00843288f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_23 VNB N_B_c_339_n 0.0439585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_M1010_g 0.0354336f $X=-0.19 $Y=-0.245 $X2=3.845 $Y2=2.12
cc_25 VNB N_A_M1019_g 0.041601f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_26 VNB A 0.00356694f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_27 VNB N_A_c_395_n 0.028603f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_28 VNB N_VPWR_c_446_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_29 VNB N_X_c_528_n 0.00478873f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_30 VNB N_X_c_529_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_31 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_32 VNB X 4.55249e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB X 0.0019078f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.3
cc_34 VNB N_VGND_c_596_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_35 VNB N_VGND_c_597_n 0.0505972f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_36 VNB N_VGND_c_598_n 0.00805556f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_37 VNB N_VGND_c_599_n 0.00610839f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_38 VNB N_VGND_c_600_n 0.00986029f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_39 VNB N_VGND_c_601_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_40 VNB N_VGND_c_602_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_603_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.63
cc_42 VNB N_VGND_c_604_n 0.0626662f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_43 VNB N_VGND_c_605_n 0.329024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_606_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=2.035
cc_45 VNB N_VGND_c_607_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=2.265
cc_46 VNB N_VGND_c_608_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.815 $Y2=2.035
cc_47 VNB N_A_489_74#_c_668_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_489_74#_c_669_n 0.0286475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_489_74#_c_670_n 0.00457226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_686_74#_c_699_n 0.00361938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_686_74#_c_700_n 0.00227843f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_52 VNB N_A_686_74#_c_701_n 0.00417796f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_53 VNB N_A_686_74#_c_702_n 0.0114037f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_54 VNB N_A_686_74#_c_703_n 0.0129442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_686_74#_c_704_n 0.0201348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_686_74#_c_705_n 0.00203831f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_57 VPB N_A_83_260#_M1003_g 0.0274066f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_58 VPB N_A_83_260#_M1004_g 0.0231904f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_59 VPB N_A_83_260#_M1005_g 0.0231975f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_60 VPB N_A_83_260#_M1006_g 0.0237939f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_61 VPB N_A_83_260#_c_116_n 0.00315544f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=1.95
cc_62 VPB N_A_83_260#_c_127_n 0.00296888f $X=-0.19 $Y=1.66 $X2=2.565 $Y2=2.035
cc_63 VPB N_A_83_260#_c_128_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=2.265
cc_64 VPB N_A_83_260#_c_129_n 0.0199499f $X=-0.19 $Y=1.66 $X2=3.815 $Y2=2.035
cc_65 VPB N_A_83_260#_c_130_n 0.00275632f $X=-0.19 $Y=1.66 $X2=3.98 $Y2=2.265
cc_66 VPB N_A_83_260#_c_131_n 0.0138658f $X=-0.19 $Y=1.66 $X2=4.815 $Y2=2.035
cc_67 VPB N_A_83_260#_c_132_n 0.00231613f $X=-0.19 $Y=1.66 $X2=4.98 $Y2=2.265
cc_68 VPB N_A_83_260#_c_133_n 0.0122709f $X=-0.19 $Y=1.66 $X2=5.455 $Y2=2.035
cc_69 VPB N_A_83_260#_c_120_n 0.0139038f $X=-0.19 $Y=1.66 $X2=5.54 $Y2=1.95
cc_70 VPB N_A_83_260#_c_135_n 0.00224287f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=2.035
cc_71 VPB N_A_83_260#_c_136_n 0.00244814f $X=-0.19 $Y=1.66 $X2=3.98 $Y2=2.035
cc_72 VPB N_C_M1007_g 0.0315807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_C_M1008_g 0.0347207f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_74 VPB C 0.00129072f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_75 VPB N_C_c_281_n 0.0209856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_B_M1001_g 0.0419075f $X=-0.19 $Y=1.66 $X2=3.845 $Y2=2.12
cc_77 VPB N_B_M1013_g 0.0367643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_B_c_338_n 0.00637526f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_79 VPB N_A_c_396_n 0.016822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_c_397_n 0.018002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB A 0.00203094f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_82 VPB N_A_c_395_n 0.0475825f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.74
cc_83 VPB N_VPWR_c_447_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_84 VPB N_VPWR_c_448_n 0.0645562f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.3
cc_85 VPB N_VPWR_c_449_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_86 VPB N_VPWR_c_450_n 0.0083004f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=0.74
cc_87 VPB N_VPWR_c_451_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.63
cc_88 VPB N_VPWR_c_452_n 0.0109286f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.3
cc_89 VPB N_VPWR_c_453_n 0.00521399f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.63
cc_90 VPB N_VPWR_c_454_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_91 VPB N_VPWR_c_455_n 0.0387928f $X=-0.19 $Y=1.66 $X2=2.065 $Y2=1.465
cc_92 VPB N_VPWR_c_456_n 0.0196104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_457_n 0.0186948f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=1.95
cc_94 VPB N_VPWR_c_458_n 0.0185368f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=2.265
cc_95 VPB N_VPWR_c_459_n 0.0186948f $X=-0.19 $Y=1.66 $X2=3.98 $Y2=2.265
cc_96 VPB N_VPWR_c_460_n 0.00632158f $X=-0.19 $Y=1.66 $X2=4.98 $Y2=2.12
cc_97 VPB N_VPWR_c_461_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_462_n 0.0111303f $X=-0.19 $Y=1.66 $X2=5.455 $Y2=2.035
cc_99 VPB N_VPWR_c_463_n 0.00613664f $X=-0.19 $Y=1.66 $X2=5.54 $Y2=1.95
cc_100 VPB N_VPWR_c_446_n 0.0647f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_101 VPB N_X_c_533_n 0.00504941f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_102 VPB N_X_c_534_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.74
cc_103 VPB X 0.00133258f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.3
cc_104 VPB X 4.55249e-19 $X=-0.19 $Y=1.66 $X2=1.44 $Y2=0.74
cc_105 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 N_A_83_260#_M1018_g N_C_M1009_g 0.0217513f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_83_260#_c_115_n N_C_M1009_g 0.00640814f $X=2.065 $Y=1.465 $X2=0 $Y2=0
cc_108 N_A_83_260#_c_121_n N_C_M1009_g 0.0148765f $X=1.955 $Y=1.465 $X2=0 $Y2=0
cc_109 N_A_83_260#_M1006_g N_C_M1007_g 0.0105747f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_83_260#_c_127_n N_C_M1007_g 0.0165444f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A_83_260#_c_128_n N_C_M1007_g 0.0137865f $X=2.73 $Y=2.265 $X2=0 $Y2=0
cc_112 N_A_83_260#_c_135_n N_C_M1007_g 0.00287083f $X=2.73 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_83_260#_c_128_n N_C_M1008_g 0.017935f $X=2.73 $Y=2.265 $X2=0 $Y2=0
cc_114 N_A_83_260#_c_129_n N_C_M1008_g 0.0142918f $X=3.815 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_83_260#_c_135_n N_C_M1008_g 0.00287083f $X=2.73 $Y=2.035 $X2=0 $Y2=0
cc_116 N_A_83_260#_c_115_n C 0.0107061f $X=2.065 $Y=1.465 $X2=0 $Y2=0
cc_117 N_A_83_260#_c_116_n C 0.00795969f $X=2.15 $Y=1.95 $X2=0 $Y2=0
cc_118 N_A_83_260#_c_127_n C 0.00282261f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_119 N_A_83_260#_c_129_n C 0.0247265f $X=3.815 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A_83_260#_c_135_n C 0.0275631f $X=2.73 $Y=2.035 $X2=0 $Y2=0
cc_121 N_A_83_260#_c_115_n N_C_c_281_n 3.25203e-19 $X=2.065 $Y=1.465 $X2=0 $Y2=0
cc_122 N_A_83_260#_c_116_n N_C_c_281_n 0.00506611f $X=2.15 $Y=1.95 $X2=0 $Y2=0
cc_123 N_A_83_260#_c_127_n N_C_c_281_n 0.00411291f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_124 N_A_83_260#_c_129_n N_C_c_281_n 0.00336308f $X=3.815 $Y=2.035 $X2=0 $Y2=0
cc_125 N_A_83_260#_c_135_n N_C_c_281_n 0.00245159f $X=2.73 $Y=2.035 $X2=0 $Y2=0
cc_126 N_A_83_260#_c_121_n N_C_c_281_n 0.0105747f $X=1.955 $Y=1.465 $X2=0 $Y2=0
cc_127 N_A_83_260#_c_129_n N_B_M1001_g 0.0142918f $X=3.815 $Y=2.035 $X2=0 $Y2=0
cc_128 N_A_83_260#_c_130_n N_B_M1001_g 0.0178457f $X=3.98 $Y=2.265 $X2=0 $Y2=0
cc_129 N_A_83_260#_c_136_n N_B_M1001_g 0.00311233f $X=3.98 $Y=2.035 $X2=0 $Y2=0
cc_130 N_A_83_260#_c_130_n N_B_M1013_g 0.00101582f $X=3.98 $Y=2.265 $X2=0 $Y2=0
cc_131 N_A_83_260#_c_131_n N_B_M1013_g 0.0171201f $X=4.815 $Y=2.035 $X2=0 $Y2=0
cc_132 N_A_83_260#_c_132_n N_B_M1013_g 6.23974e-19 $X=4.98 $Y=2.265 $X2=0 $Y2=0
cc_133 N_A_83_260#_c_129_n N_B_c_338_n 0.0256056f $X=3.815 $Y=2.035 $X2=0 $Y2=0
cc_134 N_A_83_260#_c_131_n N_B_c_338_n 0.0139703f $X=4.815 $Y=2.035 $X2=0 $Y2=0
cc_135 N_A_83_260#_c_136_n N_B_c_338_n 0.0296131f $X=3.98 $Y=2.035 $X2=0 $Y2=0
cc_136 N_A_83_260#_c_136_n N_B_c_339_n 7.57032e-19 $X=3.98 $Y=2.035 $X2=0 $Y2=0
cc_137 N_A_83_260#_c_117_n N_A_M1010_g 0.00470593f $X=4.975 $Y=0.76 $X2=0 $Y2=0
cc_138 N_A_83_260#_c_119_n N_A_M1010_g 0.00564493f $X=5.14 $Y=1.195 $X2=0 $Y2=0
cc_139 N_A_83_260#_c_131_n N_A_c_396_n 0.00858962f $X=4.815 $Y=2.035 $X2=0 $Y2=0
cc_140 N_A_83_260#_c_132_n N_A_c_396_n 0.0137058f $X=4.98 $Y=2.265 $X2=0 $Y2=0
cc_141 N_A_83_260#_c_172_p N_A_c_396_n 0.00105382f $X=4.98 $Y=2.035 $X2=0 $Y2=0
cc_142 N_A_83_260#_c_132_n N_A_c_397_n 0.017935f $X=4.98 $Y=2.265 $X2=0 $Y2=0
cc_143 N_A_83_260#_c_133_n N_A_c_397_n 0.00911633f $X=5.455 $Y=2.035 $X2=0 $Y2=0
cc_144 N_A_83_260#_c_172_p N_A_c_397_n 0.00105382f $X=4.98 $Y=2.035 $X2=0 $Y2=0
cc_145 N_A_83_260#_c_117_n N_A_M1019_g 0.0122187f $X=4.975 $Y=0.76 $X2=0 $Y2=0
cc_146 N_A_83_260#_c_118_n N_A_M1019_g 0.0140437f $X=5.455 $Y=1.195 $X2=0 $Y2=0
cc_147 N_A_83_260#_c_119_n N_A_M1019_g 0.00224308f $X=5.14 $Y=1.195 $X2=0 $Y2=0
cc_148 N_A_83_260#_c_120_n N_A_M1019_g 0.00582711f $X=5.54 $Y=1.95 $X2=0 $Y2=0
cc_149 N_A_83_260#_c_131_n A 0.0144358f $X=4.815 $Y=2.035 $X2=0 $Y2=0
cc_150 N_A_83_260#_c_118_n A 0.0103209f $X=5.455 $Y=1.195 $X2=0 $Y2=0
cc_151 N_A_83_260#_c_119_n A 0.027827f $X=5.14 $Y=1.195 $X2=0 $Y2=0
cc_152 N_A_83_260#_c_133_n A 0.00996387f $X=5.455 $Y=2.035 $X2=0 $Y2=0
cc_153 N_A_83_260#_c_120_n A 0.0261813f $X=5.54 $Y=1.95 $X2=0 $Y2=0
cc_154 N_A_83_260#_c_172_p A 0.0263422f $X=4.98 $Y=2.035 $X2=0 $Y2=0
cc_155 N_A_83_260#_c_131_n N_A_c_395_n 0.00590257f $X=4.815 $Y=2.035 $X2=0 $Y2=0
cc_156 N_A_83_260#_c_119_n N_A_c_395_n 0.00507634f $X=5.14 $Y=1.195 $X2=0 $Y2=0
cc_157 N_A_83_260#_c_133_n N_A_c_395_n 0.00533945f $X=5.455 $Y=2.035 $X2=0 $Y2=0
cc_158 N_A_83_260#_c_120_n N_A_c_395_n 0.00925512f $X=5.54 $Y=1.95 $X2=0 $Y2=0
cc_159 N_A_83_260#_c_172_p N_A_c_395_n 0.00998644f $X=4.98 $Y=2.035 $X2=0 $Y2=0
cc_160 N_A_83_260#_c_116_n N_VPWR_M1006_s 0.00206918f $X=2.15 $Y=1.95 $X2=0
+ $Y2=0
cc_161 N_A_83_260#_c_127_n N_VPWR_M1006_s 0.00287836f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_162 N_A_83_260#_c_193_p N_VPWR_M1006_s 0.00271221f $X=2.235 $Y=2.035 $X2=0
+ $Y2=0
cc_163 N_A_83_260#_c_133_n N_VPWR_M1016_s 0.00188126f $X=5.455 $Y=2.035 $X2=0
+ $Y2=0
cc_164 N_A_83_260#_M1003_g N_VPWR_c_448_n 0.00648878f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_165 N_A_83_260#_M1004_g N_VPWR_c_449_n 0.00415677f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_166 N_A_83_260#_M1005_g N_VPWR_c_449_n 0.00275958f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_167 N_A_83_260#_M1006_g N_VPWR_c_450_n 0.00203999f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_168 N_A_83_260#_c_127_n N_VPWR_c_450_n 0.0114156f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_169 N_A_83_260#_c_193_p N_VPWR_c_450_n 0.0119464f $X=2.235 $Y=2.035 $X2=0
+ $Y2=0
cc_170 N_A_83_260#_c_128_n N_VPWR_c_450_n 0.0266809f $X=2.73 $Y=2.265 $X2=0
+ $Y2=0
cc_171 N_A_83_260#_c_128_n N_VPWR_c_451_n 0.0144623f $X=2.73 $Y=2.265 $X2=0
+ $Y2=0
cc_172 N_A_83_260#_c_128_n N_VPWR_c_452_n 0.0267512f $X=2.73 $Y=2.265 $X2=0
+ $Y2=0
cc_173 N_A_83_260#_c_129_n N_VPWR_c_452_n 0.0445631f $X=3.815 $Y=2.035 $X2=0
+ $Y2=0
cc_174 N_A_83_260#_c_130_n N_VPWR_c_452_n 0.0267512f $X=3.98 $Y=2.265 $X2=0
+ $Y2=0
cc_175 N_A_83_260#_c_130_n N_VPWR_c_453_n 0.0266809f $X=3.98 $Y=2.265 $X2=0
+ $Y2=0
cc_176 N_A_83_260#_c_131_n N_VPWR_c_453_n 0.0227823f $X=4.815 $Y=2.035 $X2=0
+ $Y2=0
cc_177 N_A_83_260#_c_132_n N_VPWR_c_453_n 0.0266809f $X=4.98 $Y=2.265 $X2=0
+ $Y2=0
cc_178 N_A_83_260#_c_132_n N_VPWR_c_455_n 0.0266809f $X=4.98 $Y=2.265 $X2=0
+ $Y2=0
cc_179 N_A_83_260#_c_133_n N_VPWR_c_455_n 0.0251678f $X=5.455 $Y=2.035 $X2=0
+ $Y2=0
cc_180 N_A_83_260#_M1003_g N_VPWR_c_456_n 0.00515235f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_181 N_A_83_260#_M1004_g N_VPWR_c_456_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_83_260#_M1005_g N_VPWR_c_457_n 0.005209f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_83_260#_M1006_g N_VPWR_c_457_n 0.005209f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_83_260#_c_130_n N_VPWR_c_458_n 0.014549f $X=3.98 $Y=2.265 $X2=0 $Y2=0
cc_185 N_A_83_260#_c_132_n N_VPWR_c_459_n 0.0144623f $X=4.98 $Y=2.265 $X2=0
+ $Y2=0
cc_186 N_A_83_260#_M1003_g N_VPWR_c_446_n 0.00967664f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_187 N_A_83_260#_M1004_g N_VPWR_c_446_n 0.00982526f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_188 N_A_83_260#_M1005_g N_VPWR_c_446_n 0.00982526f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_189 N_A_83_260#_M1006_g N_VPWR_c_446_n 0.00982576f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_190 N_A_83_260#_c_128_n N_VPWR_c_446_n 0.0118344f $X=2.73 $Y=2.265 $X2=0
+ $Y2=0
cc_191 N_A_83_260#_c_130_n N_VPWR_c_446_n 0.0119743f $X=3.98 $Y=2.265 $X2=0
+ $Y2=0
cc_192 N_A_83_260#_c_132_n N_VPWR_c_446_n 0.0118344f $X=4.98 $Y=2.265 $X2=0
+ $Y2=0
cc_193 N_A_83_260#_M1015_g N_X_c_528_n 0.0132575f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_83_260#_M1017_g N_X_c_528_n 0.0124641f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_83_260#_M1018_g N_X_c_528_n 3.20368e-19 $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_83_260#_c_115_n N_X_c_528_n 0.0546701f $X=2.065 $Y=1.465 $X2=0 $Y2=0
cc_197 N_A_83_260#_c_121_n N_X_c_528_n 0.00657479f $X=1.955 $Y=1.465 $X2=0 $Y2=0
cc_198 N_A_83_260#_M1004_g N_X_c_533_n 0.0155352f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_83_260#_M1005_g N_X_c_533_n 0.0148403f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_83_260#_M1006_g N_X_c_533_n 0.00281733f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_83_260#_c_115_n N_X_c_533_n 0.0667661f $X=2.065 $Y=1.465 $X2=0 $Y2=0
cc_202 N_A_83_260#_c_116_n N_X_c_533_n 0.00779205f $X=2.15 $Y=1.95 $X2=0 $Y2=0
cc_203 N_A_83_260#_c_121_n N_X_c_533_n 0.0068296f $X=1.955 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_83_260#_M1015_g N_X_c_529_n 5.56443e-19 $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_83_260#_M1017_g N_X_c_529_n 0.00865504f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_83_260#_M1018_g N_X_c_529_n 3.97481e-19 $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_83_260#_M1004_g N_X_c_534_n 6.31736e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_83_260#_M1005_g N_X_c_534_n 0.0142049f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_83_260#_M1006_g N_X_c_534_n 0.0142026f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_83_260#_c_128_n N_X_c_534_n 0.00403964f $X=2.73 $Y=2.265 $X2=0 $Y2=0
cc_211 N_A_83_260#_M1011_g X 0.00783249f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_83_260#_M1015_g X 0.0089867f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_83_260#_M1017_g X 6.30851e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_83_260#_M1011_g X 0.00209097f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_83_260#_M1015_g X 0.00132257f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_83_260#_M1003_g X 0.0088815f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A_83_260#_M1011_g X 0.00875215f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_83_260#_M1015_g X 0.00456408f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_83_260#_M1004_g X 0.0045713f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_83_260#_c_115_n X 0.022673f $X=2.065 $Y=1.465 $X2=0 $Y2=0
cc_221 N_A_83_260#_c_121_n X 0.0315269f $X=1.955 $Y=1.465 $X2=0 $Y2=0
cc_222 N_A_83_260#_M1003_g X 0.00333871f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_83_260#_M1004_g X 0.00177091f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A_83_260#_M1003_g X 0.0139967f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_83_260#_M1004_g X 0.0142049f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A_83_260#_M1005_g X 6.31623e-19 $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_83_260#_M1011_g N_VGND_c_597_n 0.00647381f $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_A_83_260#_M1015_g N_VGND_c_598_n 0.00337101f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_229 N_A_83_260#_M1017_g N_VGND_c_598_n 0.00391054f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_230 N_A_83_260#_M1017_g N_VGND_c_599_n 5.74413e-19 $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_83_260#_M1018_g N_VGND_c_599_n 0.0115166f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_83_260#_c_115_n N_VGND_c_599_n 0.0177405f $X=2.065 $Y=1.465 $X2=0
+ $Y2=0
cc_233 N_A_83_260#_c_121_n N_VGND_c_599_n 0.00233853f $X=1.955 $Y=1.465 $X2=0
+ $Y2=0
cc_234 N_A_83_260#_M1011_g N_VGND_c_601_n 0.00434272f $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_83_260#_M1015_g N_VGND_c_601_n 0.00434272f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_236 N_A_83_260#_M1017_g N_VGND_c_602_n 0.00434272f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_237 N_A_83_260#_M1018_g N_VGND_c_602_n 0.00383152f $X=1.87 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_83_260#_M1011_g N_VGND_c_605_n 0.00823992f $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_239 N_A_83_260#_M1015_g N_VGND_c_605_n 0.00820942f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_83_260#_M1017_g N_VGND_c_605_n 0.00820718f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_83_260#_M1018_g N_VGND_c_605_n 0.0075754f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_83_260#_M1018_g N_A_489_74#_c_670_n 3.6056e-19 $X=1.87 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_83_260#_c_117_n N_A_686_74#_c_702_n 0.0171127f $X=4.975 $Y=0.76 $X2=0
+ $Y2=0
cc_244 N_A_83_260#_M1010_d N_A_686_74#_c_703_n 0.00275122f $X=4.765 $Y=0.37
+ $X2=0 $Y2=0
cc_245 N_A_83_260#_c_117_n N_A_686_74#_c_703_n 0.0197439f $X=4.975 $Y=0.76 $X2=0
+ $Y2=0
cc_246 N_A_83_260#_c_118_n N_A_686_74#_c_704_n 0.0261289f $X=5.455 $Y=1.195
+ $X2=0 $Y2=0
cc_247 N_C_M1008_g N_B_M1001_g 0.0113206f $X=2.955 $Y=2.54 $X2=0 $Y2=0
cc_248 N_C_M1014_g N_B_c_338_n 0.00321894f $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_249 C N_B_c_338_n 0.0231613f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_250 N_C_c_281_n N_B_c_338_n 0.00146345f $X=2.955 $Y=1.615 $X2=0 $Y2=0
cc_251 C N_B_c_339_n 0.00109256f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_252 N_C_c_281_n N_B_c_339_n 0.00716622f $X=2.955 $Y=1.615 $X2=0 $Y2=0
cc_253 N_C_M1007_g N_VPWR_c_450_n 0.00203999f $X=2.505 $Y=2.54 $X2=0 $Y2=0
cc_254 N_C_M1007_g N_VPWR_c_451_n 0.005209f $X=2.505 $Y=2.54 $X2=0 $Y2=0
cc_255 N_C_M1008_g N_VPWR_c_451_n 0.005209f $X=2.955 $Y=2.54 $X2=0 $Y2=0
cc_256 N_C_M1008_g N_VPWR_c_452_n 0.00260425f $X=2.955 $Y=2.54 $X2=0 $Y2=0
cc_257 N_C_M1007_g N_VPWR_c_446_n 0.00982576f $X=2.505 $Y=2.54 $X2=0 $Y2=0
cc_258 N_C_M1008_g N_VPWR_c_446_n 0.00984174f $X=2.955 $Y=2.54 $X2=0 $Y2=0
cc_259 N_C_M1007_g N_X_c_534_n 6.99364e-19 $X=2.505 $Y=2.54 $X2=0 $Y2=0
cc_260 N_C_M1009_g N_VGND_c_599_n 0.00529194f $X=2.37 $Y=0.69 $X2=0 $Y2=0
cc_261 N_C_M1009_g N_VGND_c_600_n 4.83116e-19 $X=2.37 $Y=0.69 $X2=0 $Y2=0
cc_262 N_C_M1014_g N_VGND_c_600_n 0.0120095f $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_263 N_C_M1009_g N_VGND_c_603_n 0.00434272f $X=2.37 $Y=0.69 $X2=0 $Y2=0
cc_264 N_C_M1014_g N_VGND_c_603_n 0.00383152f $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_265 N_C_M1009_g N_VGND_c_605_n 0.00820772f $X=2.37 $Y=0.69 $X2=0 $Y2=0
cc_266 N_C_M1014_g N_VGND_c_605_n 0.0075754f $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_267 N_C_M1009_g N_A_489_74#_c_668_n 0.00688879f $X=2.37 $Y=0.69 $X2=0 $Y2=0
cc_268 N_C_M1014_g N_A_489_74#_c_669_n 0.0167483f $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_269 C N_A_489_74#_c_669_n 0.0274448f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_270 N_C_c_281_n N_A_489_74#_c_669_n 0.00716132f $X=2.955 $Y=1.615 $X2=0 $Y2=0
cc_271 N_C_M1009_g N_A_489_74#_c_670_n 0.00603115f $X=2.37 $Y=0.69 $X2=0 $Y2=0
cc_272 C N_A_489_74#_c_670_n 0.00811578f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_273 N_C_c_281_n N_A_489_74#_c_670_n 0.00251351f $X=2.955 $Y=1.615 $X2=0 $Y2=0
cc_274 N_C_M1014_g N_A_686_74#_c_699_n 7.40886e-19 $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_275 N_C_M1014_g N_A_686_74#_c_701_n 7.24903e-19 $X=2.8 $Y=0.69 $X2=0 $Y2=0
cc_276 N_B_M1002_g N_A_M1010_g 0.0202091f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_277 N_B_c_338_n N_A_M1010_g 7.74814e-19 $X=4.17 $Y=1.49 $X2=0 $Y2=0
cc_278 N_B_c_338_n A 0.0185151f $X=4.17 $Y=1.49 $X2=0 $Y2=0
cc_279 N_B_c_339_n A 4.16811e-19 $X=4.26 $Y=1.49 $X2=0 $Y2=0
cc_280 N_B_M1013_g N_A_c_395_n 0.0237937f $X=4.245 $Y=2.54 $X2=0 $Y2=0
cc_281 N_B_c_338_n N_A_c_395_n 4.13836e-19 $X=4.17 $Y=1.49 $X2=0 $Y2=0
cc_282 N_B_c_339_n N_A_c_395_n 0.0202091f $X=4.26 $Y=1.49 $X2=0 $Y2=0
cc_283 N_B_M1001_g N_VPWR_c_452_n 0.00260425f $X=3.755 $Y=2.54 $X2=0 $Y2=0
cc_284 N_B_M1001_g N_VPWR_c_453_n 5.73041e-19 $X=3.755 $Y=2.54 $X2=0 $Y2=0
cc_285 N_B_M1013_g N_VPWR_c_453_n 0.0116424f $X=4.245 $Y=2.54 $X2=0 $Y2=0
cc_286 N_B_M1001_g N_VPWR_c_458_n 0.005209f $X=3.755 $Y=2.54 $X2=0 $Y2=0
cc_287 N_B_M1013_g N_VPWR_c_458_n 0.00490827f $X=4.245 $Y=2.54 $X2=0 $Y2=0
cc_288 N_B_M1001_g N_VPWR_c_446_n 0.00984568f $X=3.755 $Y=2.54 $X2=0 $Y2=0
cc_289 N_B_M1013_g N_VPWR_c_446_n 0.00969162f $X=4.245 $Y=2.54 $X2=0 $Y2=0
cc_290 N_B_M1000_g N_VGND_c_600_n 0.00174555f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_291 N_B_M1000_g N_VGND_c_604_n 0.00278247f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_292 N_B_M1002_g N_VGND_c_604_n 0.00278247f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_293 N_B_M1000_g N_VGND_c_605_n 0.00358812f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_294 N_B_M1002_g N_VGND_c_605_n 0.00353911f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_295 N_B_M1000_g N_A_489_74#_c_669_n 0.0135492f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_296 N_B_M1002_g N_A_489_74#_c_669_n 0.00413855f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_297 N_B_c_338_n N_A_489_74#_c_669_n 0.0481273f $X=4.17 $Y=1.49 $X2=0 $Y2=0
cc_298 N_B_c_339_n N_A_489_74#_c_669_n 0.00453879f $X=4.26 $Y=1.49 $X2=0 $Y2=0
cc_299 N_B_M1002_g N_A_489_74#_c_683_n 0.00134389f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_300 N_B_M1000_g N_A_686_74#_c_699_n 0.00630099f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_301 N_B_M1002_g N_A_686_74#_c_699_n 5.72812e-19 $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_302 N_B_M1000_g N_A_686_74#_c_700_n 0.00808403f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_303 N_B_M1002_g N_A_686_74#_c_700_n 0.0103048f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_304 N_B_M1000_g N_A_686_74#_c_701_n 0.00395315f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_305 N_B_M1000_g N_A_686_74#_c_702_n 6.65971e-19 $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_306 N_B_M1002_g N_A_686_74#_c_702_n 0.008708f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_307 N_B_c_338_n N_A_686_74#_c_702_n 0.0012598f $X=4.17 $Y=1.49 $X2=0 $Y2=0
cc_308 N_B_M1002_g N_A_686_74#_c_705_n 0.00184834f $X=4.26 $Y=0.69 $X2=0 $Y2=0
cc_309 N_A_c_396_n N_VPWR_c_453_n 0.00196833f $X=4.755 $Y=2.045 $X2=0 $Y2=0
cc_310 N_A_c_397_n N_VPWR_c_455_n 0.00394849f $X=5.205 $Y=2.045 $X2=0 $Y2=0
cc_311 N_A_c_396_n N_VPWR_c_459_n 0.005209f $X=4.755 $Y=2.045 $X2=0 $Y2=0
cc_312 N_A_c_397_n N_VPWR_c_459_n 0.005209f $X=5.205 $Y=2.045 $X2=0 $Y2=0
cc_313 N_A_c_396_n N_VPWR_c_446_n 0.00982246f $X=4.755 $Y=2.045 $X2=0 $Y2=0
cc_314 N_A_c_397_n N_VPWR_c_446_n 0.00985497f $X=5.205 $Y=2.045 $X2=0 $Y2=0
cc_315 N_A_M1010_g N_VGND_c_604_n 0.00278247f $X=4.69 $Y=0.69 $X2=0 $Y2=0
cc_316 N_A_M1019_g N_VGND_c_604_n 0.00278271f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_317 N_A_M1010_g N_VGND_c_605_n 0.00354355f $X=4.69 $Y=0.69 $X2=0 $Y2=0
cc_318 N_A_M1019_g N_VGND_c_605_n 0.00354455f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_319 N_A_M1010_g N_A_686_74#_c_702_n 0.00865041f $X=4.69 $Y=0.69 $X2=0 $Y2=0
cc_320 N_A_M1019_g N_A_686_74#_c_702_n 5.9419e-19 $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_321 A N_A_686_74#_c_702_n 9.20473e-19 $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_322 N_A_M1010_g N_A_686_74#_c_703_n 0.0105638f $X=4.69 $Y=0.69 $X2=0 $Y2=0
cc_323 N_A_M1019_g N_A_686_74#_c_703_n 0.0143926f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_324 N_A_M1010_g N_A_686_74#_c_705_n 0.00184834f $X=4.69 $Y=0.69 $X2=0 $Y2=0
cc_325 N_VPWR_M1004_s N_X_c_533_n 0.00279273f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_326 N_VPWR_c_449_n N_X_c_533_n 0.0208278f $X=1.23 $Y=2.305 $X2=0 $Y2=0
cc_327 N_VPWR_c_449_n N_X_c_534_n 0.0323093f $X=1.23 $Y=2.305 $X2=0 $Y2=0
cc_328 N_VPWR_c_450_n N_X_c_534_n 0.0266809f $X=2.23 $Y=2.455 $X2=0 $Y2=0
cc_329 N_VPWR_c_457_n N_X_c_534_n 0.0144623f $X=2.065 $Y=3.33 $X2=0 $Y2=0
cc_330 N_VPWR_c_446_n N_X_c_534_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_331 N_VPWR_c_448_n X 0.00634826f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_332 N_VPWR_c_448_n X 0.0346872f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_333 N_VPWR_c_449_n X 0.0323819f $X=1.23 $Y=2.305 $X2=0 $Y2=0
cc_334 N_VPWR_c_456_n X 0.0146704f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_446_n X 0.0119949f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_336 N_X_c_528_n N_VGND_M1015_d 0.00250873f $X=1.49 $Y=1.045 $X2=0 $Y2=0
cc_337 X N_VGND_c_597_n 0.0225553f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_338 X N_VGND_c_597_n 0.00756924f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_339 N_X_c_528_n N_VGND_c_598_n 0.0192006f $X=1.49 $Y=1.045 $X2=0 $Y2=0
cc_340 N_X_c_529_n N_VGND_c_598_n 0.0165801f $X=1.655 $Y=0.515 $X2=0 $Y2=0
cc_341 X N_VGND_c_598_n 0.0164981f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_342 N_X_c_529_n N_VGND_c_599_n 0.0225912f $X=1.655 $Y=0.515 $X2=0 $Y2=0
cc_343 X N_VGND_c_601_n 0.0144922f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_344 N_X_c_529_n N_VGND_c_602_n 0.0109942f $X=1.655 $Y=0.515 $X2=0 $Y2=0
cc_345 N_X_c_529_n N_VGND_c_605_n 0.00904371f $X=1.655 $Y=0.515 $X2=0 $Y2=0
cc_346 X N_VGND_c_605_n 0.0118826f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_347 N_X_c_528_n N_A_489_74#_c_670_n 0.00164421f $X=1.49 $Y=1.045 $X2=0 $Y2=0
cc_348 N_VGND_c_599_n N_A_489_74#_c_668_n 0.0235888f $X=2.085 $Y=0.515 $X2=0
+ $Y2=0
cc_349 N_VGND_c_600_n N_A_489_74#_c_668_n 0.0173942f $X=3.015 $Y=0.65 $X2=0
+ $Y2=0
cc_350 N_VGND_c_603_n N_A_489_74#_c_668_n 0.0109942f $X=2.85 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_605_n N_A_489_74#_c_668_n 0.00904371f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_M1014_s N_A_489_74#_c_669_n 0.00256317f $X=2.875 $Y=0.37 $X2=0
+ $Y2=0
cc_353 N_VGND_c_600_n N_A_489_74#_c_669_n 0.0219406f $X=3.015 $Y=0.65 $X2=0
+ $Y2=0
cc_354 N_VGND_c_599_n N_A_489_74#_c_670_n 0.0026894f $X=2.085 $Y=0.515 $X2=0
+ $Y2=0
cc_355 N_VGND_c_600_n N_A_686_74#_c_699_n 0.0262595f $X=3.015 $Y=0.65 $X2=0
+ $Y2=0
cc_356 N_VGND_c_604_n N_A_686_74#_c_700_n 0.0359382f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_605_n N_A_686_74#_c_700_n 0.0202862f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_600_n N_A_686_74#_c_701_n 0.0121616f $X=3.015 $Y=0.65 $X2=0
+ $Y2=0
cc_359 N_VGND_c_604_n N_A_686_74#_c_701_n 0.0232293f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_605_n N_A_686_74#_c_701_n 0.0126511f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_604_n N_A_686_74#_c_703_n 0.0659741f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_605_n N_A_686_74#_c_703_n 0.0367637f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_604_n N_A_686_74#_c_705_n 0.0234809f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_605_n N_A_686_74#_c_705_n 0.0126009f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_365 N_A_489_74#_c_669_n N_A_686_74#_M1000_d 0.00256317f $X=3.92 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_366 N_A_489_74#_c_669_n N_A_686_74#_c_699_n 0.0215964f $X=3.92 $Y=1.07 $X2=0
+ $Y2=0
cc_367 N_A_489_74#_M1000_s N_A_686_74#_c_700_n 0.00322515f $X=3.865 $Y=0.37
+ $X2=0 $Y2=0
cc_368 N_A_489_74#_c_669_n N_A_686_74#_c_700_n 0.00315383f $X=3.92 $Y=1.07 $X2=0
+ $Y2=0
cc_369 N_A_489_74#_c_683_n N_A_686_74#_c_700_n 0.012523f $X=4.005 $Y=0.81 $X2=0
+ $Y2=0
cc_370 N_A_489_74#_c_669_n N_A_686_74#_c_702_n 0.0030826f $X=3.92 $Y=1.07 $X2=0
+ $Y2=0
cc_371 N_A_489_74#_c_683_n N_A_686_74#_c_702_n 0.0235816f $X=4.005 $Y=0.81 $X2=0
+ $Y2=0

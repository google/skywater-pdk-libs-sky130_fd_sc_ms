* File: sky130_fd_sc_ms__sdfrtn_1.spice
* Created: Fri Aug 28 18:12:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfrtn_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfrtn_1  VNB VPB SCE D SCD CLK_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK_N	CLK_N
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1037 N_VGND_M1037_d N_SCE_M1037_g N_A_27_88#_M1037_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1491 AS=0.1197 PD=1.55 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1018 noxref_25 N_A_27_88#_M1018_g N_noxref_24_M1018_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=1.39 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1020 N_A_287_464#_M1020_d N_D_M1020_g noxref_25 VNB NLOWVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=0.98 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1006 noxref_26 N_SCE_M1006_g N_A_287_464#_M1020_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1176 PD=0.66 PS=0.98 NRD=18.564 NRS=39.996 M=1 R=2.8 SA=75001.3
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1032 N_noxref_24_M1032_d N_SCD_M1032_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0609 AS=0.0504 PD=0.71 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_RESET_B_M1023_g N_noxref_24_M1032_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.2226 AS=0.0609 PD=1.9 PS=0.71 NRD=45.708 NRS=1.428 M=1 R=2.8
+ SA=75002.1 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_CLK_N_M1007_g N_A_859_347#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.14615 AS=0.2442 PD=1.135 PS=2.14 NRD=9.72 NRS=3.24 M=1 R=4.93333
+ SA=75000.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1008 N_A_1069_74#_M1008_d N_A_859_347#_M1008_g N_VGND_M1007_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2257 AS=0.14615 PD=2.09 PS=1.135 NRD=6.48 NRS=8.916 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_A_1273_131#_M1021_d N_A_1069_74#_M1021_g N_A_287_464#_M1021_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1028 A_1409_131# N_A_859_347#_M1028_g N_A_1273_131#_M1021_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0462 AS=0.1113 PD=0.64 PS=0.95 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1016 A_1483_131# N_A_1417_294#_M1016_g A_1409_131# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0462 PD=0.63 PS=0.64 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75001.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_1483_131# VNB NLOWVT L=0.15 W=0.42
+ AD=0.139957 AS=0.0441 PD=1.16491 PS=0.63 NRD=79.488 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1035 N_A_1417_294#_M1035_d N_A_1273_131#_M1035_g N_VGND_M1003_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1792 AS=0.213268 PD=1.2 PS=1.77509 NRD=46.872 NRS=52.164
+ M=1 R=4.26667 SA=75001.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1039 N_A_1827_144#_M1039_d N_A_859_347#_M1039_g N_A_1417_294#_M1035_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.397902 AS=0.1792 PD=2.57208 PS=1.2 NRD=106.26
+ NRS=0.312 M=1 R=4.26667 SA=75002 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1026 A_2073_74# N_A_1069_74#_M1026_g N_A_1827_144#_M1039_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0525 AS=0.261123 PD=0.67 PS=1.68792 NRD=19.992 NRS=161.916 M=1
+ R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_2087_410#_M1004_g A_2073_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0861 AS=0.0525 PD=0.83 PS=0.67 NRD=17.136 NRS=19.992 M=1 R=2.8 SA=75001.9
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 A_2265_74# N_RESET_B_M1009_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0861 PD=0.66 PS=0.83 NRD=18.564 NRS=19.992 M=1 R=2.8 SA=75002.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_2087_410#_M1010_d N_A_1827_144#_M1010_g A_2265_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.21 AS=0.0504 PD=1.84 PS=0.66 NRD=30 NRS=18.564 M=1 R=2.8
+ SA=75002.8 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_A_1827_144#_M1027_g N_A_2492_424#_M1027_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=25.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1017 N_Q_M1017_d N_A_2492_424#_M1017_g N_VGND_M1027_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_SCE_M1011_g N_A_27_88#_M1011_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.1792 PD=0.91 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90003 A=0.1152 P=1.64 MULT=1
MM1012 A_209_464# N_SCE_M1012_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.6
+ SB=90002.5 A=0.1152 P=1.64 MULT=1
MM1034 N_A_287_464#_M1034_d N_D_M1034_g A_209_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.2416 AS=0.0672 PD=1.395 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556 SA=90001
+ SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1015 A_474_464# N_A_27_88#_M1015_g N_A_287_464#_M1034_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0672 AS=0.2416 PD=0.85 PS=1.395 NRD=15.3857 NRS=0 M=1 R=3.55556
+ SA=90002 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1036 N_VPWR_M1036_d N_SCD_M1036_g A_474_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.174875 AS=0.0672 PD=1.315 PS=0.85 NRD=67.177 NRS=15.3857 M=1 R=3.55556
+ SA=90002.4 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1002 N_A_287_464#_M1002_d N_RESET_B_M1002_g N_VPWR_M1036_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.174875 PD=1.84 PS=1.315 NRD=0 NRS=67.177 M=1 R=3.55556
+ SA=90003 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1000 N_VPWR_M1000_d N_CLK_N_M1000_g N_A_859_347#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.210787 AS=0.325 PD=1.47 PS=2.65 NRD=12.7853 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1029 N_A_1069_74#_M1029_d N_A_859_347#_M1029_g N_VPWR_M1000_d VPB PSHORT
+ L=0.18 W=1 AD=0.265 AS=0.210787 PD=2.53 PS=1.47 NRD=0 NRS=11.8003 M=1
+ R=5.55556 SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_1273_131#_M1001_d N_A_859_347#_M1001_g N_A_287_464#_M1001_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1024 A_1381_457# N_A_1069_74#_M1024_g N_A_1273_131#_M1001_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1033 N_VPWR_M1033_d N_A_1417_294#_M1033_g A_1381_457# VPB PSHORT L=0.18 W=0.42
+ AD=0.063 AS=0.0504 PD=0.72 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90001.1
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1030 N_A_1273_131#_M1030_d N_RESET_B_M1030_g N_VPWR_M1033_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1092 AS=0.063 PD=1.36 PS=0.72 NRD=0 NRS=11.7215 M=1 R=2.33333
+ SA=90001.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1038 N_A_1417_294#_M1038_d N_A_1273_131#_M1038_g N_VPWR_M1038_s VPB PSHORT
+ L=0.18 W=1 AD=0.3775 AS=0.26 PD=1.755 PS=2.52 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002 A=0.18 P=2.36 MULT=1
MM1031 N_A_1827_144#_M1031_d N_A_1069_74#_M1031_g N_A_1417_294#_M1038_d VPB
+ PSHORT L=0.18 W=1 AD=0.205282 AS=0.3775 PD=1.88028 PS=1.755 NRD=2.6201 NRS=0
+ M=1 R=5.55556 SA=90001.1 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 A_2045_508# N_A_859_347#_M1005_g N_A_1827_144#_M1031_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0483 AS=0.0862183 PD=0.65 PS=0.789718 NRD=28.1316 NRS=16.4101 M=1
+ R=2.33333 SA=90001.6 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1013 N_VPWR_M1013_d N_A_2087_410#_M1013_g A_2045_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.12495 AS=0.0483 PD=1.015 PS=0.65 NRD=60.9715 NRS=28.1316 M=1 R=2.33333
+ SA=90002 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1019 N_A_2087_410#_M1019_d N_RESET_B_M1019_g N_VPWR_M1013_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.12495 PD=0.69 PS=1.015 NRD=0 NRS=86.7588 M=1 R=2.33333
+ SA=90002.8 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1022 N_VPWR_M1022_d N_A_1827_144#_M1022_g N_A_2087_410#_M1019_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1386 AS=0.0567 PD=1.5 PS=0.69 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90003.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1025 N_VPWR_M1025_d N_A_1827_144#_M1025_g N_A_2492_424#_M1025_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.183 AS=0.2352 PD=1.30286 PS=2.24 NRD=18.7544 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1014 N_Q_M1014_d N_A_2492_424#_M1014_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3192 AS=0.244 PD=2.81 PS=1.73714 NRD=0 NRS=7.0329 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=26.3107 P=32.77
c_137 VNB 0 1.94919e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sdfrtn_1.pxi.spice"
*
.ends
*
*

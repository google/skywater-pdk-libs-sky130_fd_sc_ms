* File: sky130_fd_sc_ms__dfxtp_4.pex.spice
* Created: Fri Aug 28 17:25:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFXTP_4%CLK 3 7 9 13 16
c36 3 0 1.52766e-19 $X=0.505 $Y=2.4
r37 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r38 12 15 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.34 $Y=1.465
+ $X2=0.495 $Y2=1.465
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.465 $X2=0.34 $Y2=1.465
r40 9 13 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.465
r41 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r42 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r43 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r44 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_27_74# 1 2 9 13 16 21 25 27 28 32 33 34 37
+ 39 41 43 44 45 48 51 52 54 55 56 58 59 60 61 64 67 69 70 73 75 78 79 82 86 87
+ 88 91 94
c274 86 0 6.73668e-20 $X=5.83 $Y=0.345
c275 70 0 1.76602e-19 $X=4.51 $Y=0.775
c276 28 0 5.53797e-20 $X=5.185 $Y=1.765
c277 27 0 1.11025e-19 $X=5.74 $Y=1.765
c278 25 0 1.80422e-19 $X=5.095 $Y=2.54
c279 9 0 6.77311e-20 $X=0.955 $Y=2.4
r280 87 98 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=0.345
+ $X2=5.83 $Y2=0.51
r281 86 88 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.83 $Y=0.382
+ $X2=5.665 $Y2=0.382
r282 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.83
+ $Y=0.345 $X2=5.83 $Y2=0.345
r283 82 92 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.385 $X2=1
+ $Y2=1.55
r284 82 91 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.385 $X2=1
+ $Y2=1.22
r285 81 83 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.385
+ $X2=0.905 $Y2=1.55
r286 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.385 $X2=0.97 $Y2=1.385
r287 78 81 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=1.385
r288 78 79 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=0.96
r289 75 88 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=4.68 $Y=0.34
+ $X2=5.665 $Y2=0.34
r290 72 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.595 $Y=0.425
+ $X2=4.68 $Y2=0.34
r291 72 73 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.595 $Y=0.425
+ $X2=4.595 $Y2=0.69
r292 71 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=0.775
+ $X2=3.79 $Y2=0.775
r293 70 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.51 $Y=0.775
+ $X2=4.595 $Y2=0.69
r294 70 71 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.51 $Y=0.775
+ $X2=3.875 $Y2=0.775
r295 68 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.86
+ $X2=3.79 $Y2=0.775
r296 68 69 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.79 $Y=0.86
+ $X2=3.79 $Y2=1.75
r297 67 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.69
+ $X2=3.79 $Y2=0.775
r298 66 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.79 $Y=0.425
+ $X2=3.79 $Y2=0.69
r299 64 95 39.8861 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=3.287 $Y=1.915
+ $X2=3.287 $Y2=2.08
r300 64 94 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=3.287 $Y=1.915
+ $X2=3.287 $Y2=1.75
r301 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.915 $X2=3.32 $Y2=1.915
r302 61 69 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.705 $Y=1.915
+ $X2=3.79 $Y2=1.75
r303 61 63 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.705 $Y=1.915
+ $X2=3.32 $Y2=1.915
r304 59 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=0.34
+ $X2=3.79 $Y2=0.425
r305 59 60 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.705 $Y=0.34
+ $X2=2.655 $Y2=0.34
r306 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.57 $Y=0.425
+ $X2=2.655 $Y2=0.34
r307 57 58 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.57 $Y=0.425
+ $X2=2.57 $Y2=0.73
r308 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.485 $Y=0.815
+ $X2=2.57 $Y2=0.73
r309 55 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.485 $Y=0.815
+ $X2=1.815 $Y2=0.815
r310 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=0.73
+ $X2=1.815 $Y2=0.815
r311 53 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.73 $Y=0.425
+ $X2=1.73 $Y2=0.73
r312 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.73 $Y2=0.425
r313 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.135 $Y2=0.34
r314 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.135 $Y2=0.34
r315 49 79 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.05 $Y2=0.96
r316 48 83 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.76 $Y=1.95 $X2=0.76
+ $Y2=1.55
r317 46 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r318 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.76 $Y2=1.95
r319 45 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.445 $Y2=2.035
r320 43 78 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.905 $Y2=1.045
r321 43 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.445 $Y2=1.045
r322 39 77 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r323 39 41 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r324 35 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.445 $Y2=1.045
r325 35 37 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.515
r326 34 94 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.165 $Y=1.24
+ $X2=3.165 $Y2=1.75
r327 33 34 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=3.145 $Y=1.09
+ $X2=3.145 $Y2=1.24
r328 32 98 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.815 $Y=0.83
+ $X2=5.815 $Y2=0.51
r329 30 32 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.815 $Y=1.69
+ $X2=5.815 $Y2=0.83
r330 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.74 $Y=1.765
+ $X2=5.815 $Y2=1.69
r331 27 28 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.74 $Y=1.765
+ $X2=5.185 $Y2=1.765
r332 23 28 33.7919 $w=1.32e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.095 $Y=1.84
+ $X2=5.185 $Y2=1.765
r333 23 25 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=5.095 $Y=1.84
+ $X2=5.095 $Y2=2.54
r334 21 95 250.718 $w=1.8e-07 $l=6.45e-07 $layer=POLY_cond $X=3.18 $Y=2.725
+ $X2=3.18 $Y2=2.08
r335 16 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.125 $Y=0.805
+ $X2=3.125 $Y2=1.09
r336 13 91 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.12 $Y=0.74
+ $X2=1.12 $Y2=1.22
r337 9 92 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.955 $Y=2.4
+ $X2=0.955 $Y2=1.55
r338 2 77 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r339 2 41 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r340 1 37 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%D 3 5 7 9 13 15 17 18 24 26 38
c62 38 0 1.17955e-19 $X=2.16 $Y=1.665
c63 13 0 1.60912e-19 $X=1.95 $Y=2.19
c64 7 0 1.63132e-19 $X=2.695 $Y=1.125
c65 5 0 1.82072e-19 $X=2.62 $Y=1.2
r66 32 38 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=2.125 $Y=1.6
+ $X2=2.125 $Y2=1.665
r67 26 29 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.14 $Y=1.2 $X2=2.14
+ $Y2=1.29
r68 18 40 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.125 $Y=1.675
+ $X2=2.125 $Y2=1.78
r69 18 38 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=2.125 $Y=1.675
+ $X2=2.125 $Y2=1.665
r70 18 32 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=2.125 $Y=1.59
+ $X2=2.125 $Y2=1.6
r71 17 18 9.60369 $w=3.58e-07 $l=3e-07 $layer=LI1_cond $X=2.125 $Y=1.29
+ $X2=2.125 $Y2=1.59
r72 17 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.29 $X2=2.14 $Y2=1.29
r73 15 40 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.03 $Y=2.025
+ $X2=2.03 $Y2=1.78
r74 14 24 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.95 $Y=2.19
+ $X2=2.11 $Y2=2.19
r75 13 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=2.19
+ $X2=1.95 $Y2=2.025
r76 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=2.19 $X2=1.95 $Y2=2.19
r77 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.695 $Y=1.125
+ $X2=2.695 $Y2=0.805
r78 6 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.2
+ $X2=2.14 $Y2=1.2
r79 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.62 $Y=1.2
+ $X2=2.695 $Y2=1.125
r80 5 6 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.62 $Y=1.2 $X2=2.305
+ $Y2=1.2
r81 1 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=2.355
+ $X2=2.11 $Y2=2.19
r82 1 3 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.11 $Y=2.355 $X2=2.11
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_209_368# 1 2 8 9 10 11 15 19 21 23 26 30
+ 33 37 40 41 42 44 45 46 48 49 50 51 52 53 57 58 61 62 63 70 71 76 77
c238 76 0 3.86493e-19 $X=5.355 $Y=1.315
c239 61 0 1.52766e-19 $X=1.18 $Y=1.985
c240 48 0 1.34159e-19 $X=4.3 $Y=2.905
c241 45 0 4.62629e-20 $X=4.215 $Y=2.675
c242 37 0 6.77311e-20 $X=1.995 $Y=2.61
c243 21 0 9.7909e-20 $X=5.23 $Y=1.15
c244 15 0 1.60912e-19 $X=2.645 $Y=2.635
r245 76 80 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.355 $Y=1.315
+ $X2=5.23 $Y2=1.315
r246 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.355
+ $Y=1.315 $X2=5.355 $Y2=1.315
r247 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.385 $X2=1.6 $Y2=1.385
r248 67 70 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.39 $Y=1.385
+ $X2=1.6 $Y2=1.385
r249 63 65 5.33035 $w=4.58e-07 $l=2.05e-07 $layer=LI1_cond $X=1.245 $Y=2.61
+ $X2=1.245 $Y2=2.815
r250 61 62 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=1.985
+ $X2=1.245 $Y2=1.82
r251 58 84 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.79 $Y=2.215
+ $X2=5.63 $Y2=2.215
r252 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.79
+ $Y=2.215 $X2=5.79 $Y2=2.215
r253 55 57 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.79 $Y=2.905
+ $X2=5.79 $Y2=2.215
r254 54 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.99
+ $X2=4.98 $Y2=2.99
r255 53 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.625 $Y=2.99
+ $X2=5.79 $Y2=2.905
r256 53 54 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.625 $Y=2.99
+ $X2=5.065 $Y2=2.99
r257 52 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.905
+ $X2=4.98 $Y2=2.99
r258 51 75 15.9965 $w=2.86e-07 $l=4.62331e-07 $layer=LI1_cond $X=4.98 $Y=1.54
+ $X2=5.355 $Y2=1.345
r259 51 52 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.98 $Y=1.54
+ $X2=4.98 $Y2=2.905
r260 49 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=2.99
+ $X2=4.98 $Y2=2.99
r261 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.895 $Y=2.99
+ $X2=4.385 $Y2=2.99
r262 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.3 $Y=2.905
+ $X2=4.385 $Y2=2.99
r263 47 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.3 $Y=2.76
+ $X2=4.3 $Y2=2.905
r264 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.215 $Y=2.675
+ $X2=4.3 $Y2=2.76
r265 45 46 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.215 $Y=2.675
+ $X2=3.375 $Y2=2.675
r266 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.29 $Y=2.76
+ $X2=3.375 $Y2=2.675
r267 43 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.29 $Y=2.76
+ $X2=3.29 $Y2=2.905
r268 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.205 $Y=2.99
+ $X2=3.29 $Y2=2.905
r269 41 42 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.205 $Y=2.99
+ $X2=2.165 $Y2=2.99
r270 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.165 $Y2=2.99
r271 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.08 $Y=2.695
+ $X2=2.08 $Y2=2.905
r272 38 63 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.475 $Y=2.61
+ $X2=1.245 $Y2=2.61
r273 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.995 $Y=2.61
+ $X2=2.08 $Y2=2.695
r274 37 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.995 $Y=2.61
+ $X2=1.475 $Y2=2.61
r275 35 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.55
+ $X2=1.39 $Y2=1.385
r276 35 62 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.39 $Y=1.55
+ $X2=1.39 $Y2=1.82
r277 31 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.22
+ $X2=1.39 $Y2=1.385
r278 31 33 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.39 $Y=1.22
+ $X2=1.39 $Y2=0.86
r279 30 63 2.21014 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=2.525
+ $X2=1.245 $Y2=2.61
r280 29 61 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.245 $Y=2.05
+ $X2=1.245 $Y2=1.985
r281 29 30 12.3508 $w=4.58e-07 $l=4.75e-07 $layer=LI1_cond $X=1.245 $Y=2.05
+ $X2=1.245 $Y2=2.525
r282 24 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=2.38
+ $X2=5.63 $Y2=2.215
r283 24 26 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.63 $Y=2.38
+ $X2=5.63 $Y2=2.75
r284 21 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.23 $Y=1.15
+ $X2=5.23 $Y2=1.315
r285 21 23 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.23 $Y=1.15
+ $X2=5.23 $Y2=0.765
r286 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.6 $Y=0.255
+ $X2=3.6 $Y2=0.72
r287 13 28 0.70609 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.645 $Y=1.845
+ $X2=2.645 $Y2=1.755
r288 13 15 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.645 $Y=1.845
+ $X2=2.645 $Y2=2.635
r289 12 71 68.7189 $w=2.49e-07 $l=4.29651e-07 $layer=POLY_cond $X=1.765 $Y=1.74
+ $X2=1.6 $Y2=1.385
r290 11 28 60.3792 $w=1.65e-07 $l=2.12368e-07 $layer=POLY_cond $X=2.44 $Y=1.74
+ $X2=2.645 $Y2=1.755
r291 11 12 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.44 $Y=1.74
+ $X2=1.765 $Y2=1.74
r292 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.525 $Y=0.18
+ $X2=3.6 $Y2=0.255
r293 9 10 902.468 $w=1.5e-07 $l=1.76e-06 $layer=POLY_cond $X=3.525 $Y=0.18
+ $X2=1.765 $Y2=0.18
r294 8 71 39.5011 $w=2.49e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.69 $Y=1.22
+ $X2=1.6 $Y2=1.385
r295 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.765 $Y2=0.18
r296 7 8 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.69 $Y2=1.22
r297 2 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r298 2 61 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r299 1 33 182 $w=1.7e-07 $l=5.79353e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.37 $X2=1.39 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_696_458# 1 2 7 9 10 11 12 14 17 21 24 26
+ 28
c82 28 0 8.37878e-20 $X=4.64 $Y=2.46
c83 26 0 5.53797e-20 $X=4.64 $Y=1.37
c84 12 0 1.7945e-19 $X=3.96 $Y=1.04
r85 31 32 17.0325 $w=3.08e-07 $l=4.3e-07 $layer=LI1_cond $X=4.867 $Y=0.77
+ $X2=4.867 $Y2=1.2
r86 26 32 9.16445 $w=3.08e-07 $l=3.00198e-07 $layer=LI1_cond $X=4.64 $Y=1.37
+ $X2=4.867 $Y2=1.2
r87 26 28 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.64 $Y=1.37
+ $X2=4.64 $Y2=2.46
r88 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.205 $X2=4.21 $Y2=1.205
r89 21 32 0.104369 $w=3.4e-07 $l=3.12e-07 $layer=LI1_cond $X=4.555 $Y=1.2
+ $X2=4.867 $Y2=1.2
r90 21 23 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=4.555 $Y=1.2
+ $X2=4.21 $Y2=1.2
r91 20 24 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.035 $Y=1.205
+ $X2=4.21 $Y2=1.205
r92 12 20 40.7148 $w=2.25e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.96 $Y=1.04
+ $X2=3.885 $Y2=1.205
r93 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.96 $Y=1.04
+ $X2=3.96 $Y2=0.72
r94 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=2.29
+ $X2=3.77 $Y2=2.365
r95 10 20 51.4259 $w=2.25e-07 $l=2.66364e-07 $layer=POLY_cond $X=3.77 $Y=1.42
+ $X2=3.885 $Y2=1.205
r96 10 11 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.77 $Y=1.42
+ $X2=3.77 $Y2=2.29
r97 7 17 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.57 $Y=2.365 $X2=3.77
+ $Y2=2.365
r98 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.57 $Y=2.44 $X2=3.57
+ $Y2=2.725
r99 2 28 600 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.12 $X2=4.64 $Y2=2.46
r100 1 31 182 $w=1.7e-07 $l=4.7355e-07 $layer=licon1_NDIFF $count=1 $X=4.83
+ $Y=0.38 $X2=5.015 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_547_485# 1 2 9 12 15 18 20 21 22 23 26 29
+ 32 38 43
c107 38 0 1.7945e-19 $X=3.355 $Y=0.785
c108 26 0 3.15687e-19 $X=3.26 $Y=1.41
c109 18 0 1.76602e-19 $X=4.722 $Y=1.45
r110 42 43 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=4.415 $Y=1.795
+ $X2=4.69 $Y2=1.795
r111 35 38 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.26 $Y=0.785
+ $X2=3.355 $Y2=0.785
r112 32 34 13.9239 $w=2.76e-07 $l=3.15e-07 $layer=LI1_cond $X=2.87 $Y=2.335
+ $X2=2.87 $Y2=2.65
r113 30 42 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.22 $Y=1.795
+ $X2=4.415 $Y2=1.795
r114 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=1.795 $X2=4.22 $Y2=1.795
r115 27 29 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.22 $Y=2.25
+ $X2=4.22 $Y2=1.795
r116 25 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=0.95
+ $X2=3.26 $Y2=0.785
r117 25 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.26 $Y=0.95
+ $X2=3.26 $Y2=1.41
r118 24 32 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=2.335
+ $X2=2.87 $Y2=2.335
r119 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.055 $Y=2.335
+ $X2=4.22 $Y2=2.25
r120 23 24 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.055 $Y=2.335
+ $X2=3.035 $Y2=2.335
r121 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.175 $Y=1.495
+ $X2=3.26 $Y2=1.41
r122 21 22 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.175 $Y=1.495
+ $X2=2.985 $Y2=1.495
r123 20 32 5.54508 $w=2.76e-07 $l=9.88686e-08 $layer=LI1_cond $X=2.9 $Y=2.25
+ $X2=2.87 $Y2=2.335
r124 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.9 $Y=1.58
+ $X2=2.985 $Y2=1.495
r125 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.9 $Y=1.58 $X2=2.9
+ $Y2=2.25
r126 17 18 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=4.722 $Y=1.3
+ $X2=4.722 $Y2=1.45
r127 15 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.755 $Y=0.655
+ $X2=4.755 $Y2=1.3
r128 12 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.63
+ $X2=4.69 $Y2=1.795
r129 12 18 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.69 $Y=1.63
+ $X2=4.69 $Y2=1.45
r130 7 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.96
+ $X2=4.415 $Y2=1.795
r131 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.415 $Y=1.96
+ $X2=4.415 $Y2=2.54
r132 2 34 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=2.425 $X2=2.87 $Y2=2.65
r133 1 38 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.595 $X2=3.355 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_1226_296# 1 2 9 13 17 21 25 29 33 37 41 45
+ 47 51 53 55 58 59 64 68 69 86
c165 86 0 1.97011e-19 $X=9.08 $Y=1.465
c166 69 0 1.21137e-19 $X=6.295 $Y=1.645
c167 68 0 2.00281e-19 $X=6.295 $Y=1.645
c168 51 0 3.64416e-20 $X=6.985 $Y=2.265
c169 13 0 6.73668e-20 $X=6.28 $Y=0.83
r170 85 86 65.1761 $w=3.18e-07 $l=4.3e-07 $layer=POLY_cond $X=8.65 $Y=1.465
+ $X2=9.08 $Y2=1.465
r171 84 85 0.757862 $w=3.18e-07 $l=5e-09 $layer=POLY_cond $X=8.645 $Y=1.465
+ $X2=8.65 $Y2=1.465
r172 81 82 0.757862 $w=3.18e-07 $l=5e-09 $layer=POLY_cond $X=8.195 $Y=1.465
+ $X2=8.2 $Y2=1.465
r173 78 79 2.27358 $w=3.18e-07 $l=1.5e-08 $layer=POLY_cond $X=7.73 $Y=1.465
+ $X2=7.745 $Y2=1.465
r174 69 77 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.645
+ $X2=6.295 $Y2=1.81
r175 69 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.645
+ $X2=6.295 $Y2=1.48
r176 68 70 6.55034 $w=2.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.295 $Y=1.645
+ $X2=6.295 $Y2=1.805
r177 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.295
+ $Y=1.645 $X2=6.295 $Y2=1.645
r178 65 84 21.978 $w=3.18e-07 $l=1.45e-07 $layer=POLY_cond $X=8.5 $Y=1.465
+ $X2=8.645 $Y2=1.465
r179 65 82 45.4717 $w=3.18e-07 $l=3e-07 $layer=POLY_cond $X=8.5 $Y=1.465 $X2=8.2
+ $Y2=1.465
r180 64 65 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.5
+ $Y=1.465 $X2=8.5 $Y2=1.465
r181 62 81 56.8396 $w=3.18e-07 $l=3.75e-07 $layer=POLY_cond $X=7.82 $Y=1.465
+ $X2=8.195 $Y2=1.465
r182 62 79 11.3679 $w=3.18e-07 $l=7.5e-08 $layer=POLY_cond $X=7.82 $Y=1.465
+ $X2=7.745 $Y2=1.465
r183 61 64 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.82 $Y=1.465
+ $X2=8.5 $Y2=1.465
r184 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.82
+ $Y=1.465 $X2=7.82 $Y2=1.465
r185 59 72 3.46916 $w=3.3e-07 $l=2.94449e-07 $layer=LI1_cond $X=7.47 $Y=1.465
+ $X2=7.385 $Y2=1.72
r186 59 61 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=7.47 $Y=1.465
+ $X2=7.82 $Y2=1.465
r187 58 72 3.63555 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=7.385 $Y=1.3
+ $X2=7.385 $Y2=1.72
r188 57 74 0.265075 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=1.05
+ $X2=7.385 $Y2=0.965
r189 57 58 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.385 $Y=1.05
+ $X2=7.385 $Y2=1.3
r190 53 74 28.5696 $w=1.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.015 $Y=0.965
+ $X2=7.385 $Y2=0.965
r191 53 55 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=7.015 $Y=0.88
+ $X2=7.015 $Y2=0.515
r192 49 72 17.491 $w=2.79e-07 $l=4e-07 $layer=LI1_cond $X=6.985 $Y=1.72
+ $X2=7.385 $Y2=1.72
r193 49 51 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.985 $Y=1.89
+ $X2=6.985 $Y2=2.265
r194 48 70 4.02169 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=1.805
+ $X2=6.295 $Y2=1.805
r195 47 49 9.06394 $w=2.79e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.82 $Y=1.805
+ $X2=6.985 $Y2=1.72
r196 47 48 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.82 $Y=1.805
+ $X2=6.46 $Y2=1.805
r197 43 86 2.27358 $w=3.18e-07 $l=1.5e-08 $layer=POLY_cond $X=9.095 $Y=1.465
+ $X2=9.08 $Y2=1.465
r198 43 45 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=9.095 $Y=1.6
+ $X2=9.095 $Y2=2.4
r199 39 86 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.08 $Y=1.3
+ $X2=9.08 $Y2=1.465
r200 39 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.08 $Y=1.3
+ $X2=9.08 $Y2=0.74
r201 35 85 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.65 $Y=1.3
+ $X2=8.65 $Y2=1.465
r202 35 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.65 $Y=1.3
+ $X2=8.65 $Y2=0.74
r203 31 84 16.0701 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.63
+ $X2=8.645 $Y2=1.465
r204 31 33 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.645 $Y=1.63
+ $X2=8.645 $Y2=2.4
r205 27 82 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=1.3 $X2=8.2
+ $Y2=1.465
r206 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.2 $Y=1.3 $X2=8.2
+ $Y2=0.74
r207 23 81 16.0701 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=1.63
+ $X2=8.195 $Y2=1.465
r208 23 25 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.195 $Y=1.63
+ $X2=8.195 $Y2=2.4
r209 19 79 16.0701 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.745 $Y=1.63
+ $X2=7.745 $Y2=1.465
r210 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.745 $Y=1.63
+ $X2=7.745 $Y2=2.4
r211 15 78 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.73 $Y=1.3
+ $X2=7.73 $Y2=1.465
r212 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.73 $Y=1.3
+ $X2=7.73 $Y2=0.74
r213 13 76 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=6.28 $Y=0.83
+ $X2=6.28 $Y2=1.48
r214 9 77 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=6.255 $Y=2.75
+ $X2=6.255 $Y2=1.81
r215 2 51 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.85
+ $Y=2.12 $X2=6.985 $Y2=2.265
r216 1 55 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.91
+ $Y=0.37 $X2=7.055 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_1037_424# 1 2 7 9 11 12 14 16 17 19 20 23
+ 25 29 30 32 34 35 37 40
c101 40 0 8.92564e-20 $X=6.965 $Y=1.385
c102 37 0 9.7909e-20 $X=5.775 $Y=1.225
c103 35 0 1.97011e-19 $X=6.63 $Y=1.225
c104 30 0 1.79413e-19 $X=5.405 $Y=1.795
c105 29 0 2.44429e-19 $X=5.69 $Y=1.795
c106 11 0 3.64416e-20 $X=6.875 $Y=1.895
r107 40 41 16.814 $w=2.58e-07 $l=9e-08 $layer=POLY_cond $X=6.965 $Y=1.385
+ $X2=6.875 $Y2=1.385
r108 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.965
+ $Y=1.385 $X2=6.965 $Y2=1.385
r109 36 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.86 $Y=1.225
+ $X2=5.775 $Y2=1.225
r110 35 39 15.8449 $w=3.02e-07 $l=3.90416e-07 $layer=LI1_cond $X=6.63 $Y=1.225
+ $X2=6.965 $Y2=1.345
r111 35 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.63 $Y=1.225
+ $X2=5.86 $Y2=1.225
r112 33 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=1.31
+ $X2=5.775 $Y2=1.225
r113 33 34 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.775 $Y=1.31
+ $X2=5.775 $Y2=1.71
r114 32 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=1.14
+ $X2=5.775 $Y2=1.225
r115 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.775 $Y=0.97
+ $X2=5.775 $Y2=1.14
r116 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.69 $Y=1.795
+ $X2=5.775 $Y2=1.71
r117 29 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.69 $Y=1.795
+ $X2=5.405 $Y2=1.795
r118 25 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.69 $Y=0.845
+ $X2=5.775 $Y2=0.97
r119 25 27 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.69 $Y=0.845
+ $X2=5.555 $Y2=0.845
r120 21 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.32 $Y=1.88
+ $X2=5.405 $Y2=1.795
r121 21 23 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=5.32 $Y=1.88
+ $X2=5.32 $Y2=2.46
r122 17 40 56.9806 $w=2.58e-07 $l=3.78616e-07 $layer=POLY_cond $X=7.27 $Y=1.22
+ $X2=6.965 $Y2=1.385
r123 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.27 $Y=1.22
+ $X2=7.27 $Y2=0.74
r124 14 16 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.21 $Y=2.045
+ $X2=7.21 $Y2=2.54
r125 13 20 6.66866 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=6.95 $Y=1.97
+ $X2=6.81 $Y2=1.97
r126 12 14 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.12 $Y=1.97
+ $X2=7.21 $Y2=2.045
r127 12 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.12 $Y=1.97
+ $X2=6.95 $Y2=1.97
r128 11 20 18.8402 $w=1.65e-07 $l=1.0247e-07 $layer=POLY_cond $X=6.875 $Y=1.895
+ $X2=6.81 $Y2=1.97
r129 10 41 15.449 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.875 $Y=1.55
+ $X2=6.875 $Y2=1.385
r130 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.875 $Y=1.55
+ $X2=6.875 $Y2=1.895
r131 7 20 18.8402 $w=1.65e-07 $l=9.68246e-08 $layer=POLY_cond $X=6.76 $Y=2.045
+ $X2=6.81 $Y2=1.97
r132 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=6.76 $Y=2.045
+ $X2=6.76 $Y2=2.54
r133 2 23 600 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=2.12 $X2=5.32 $Y2=2.46
r134 1 27 182 $w=1.7e-07 $l=4.21871e-07 $layer=licon1_NDIFF $count=1 $X=5.305
+ $Y=0.49 $X2=5.555 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%VPWR 1 2 3 4 5 6 7 26 28 32 36 40 42 46 48
+ 50 55 58 61 70 77 82 88 91 94 97 100 104
r126 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r127 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r129 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r130 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r131 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r132 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 86 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r135 86 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r136 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r137 83 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.42 $Y2=3.33
r138 83 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.505 $Y=3.33
+ $X2=8.88 $Y2=3.33
r139 82 103 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.235 $Y=3.33
+ $X2=9.417 $Y2=3.33
r140 82 85 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.235 $Y=3.33
+ $X2=8.88 $Y2=3.33
r141 81 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r142 81 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r143 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r144 78 94 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.482 $Y2=3.33
r145 78 80 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.96 $Y2=3.33
r146 77 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.355 $Y=3.33
+ $X2=7.48 $Y2=3.33
r147 77 80 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.355 $Y=3.33
+ $X2=6.96 $Y2=3.33
r148 76 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r149 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r150 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r151 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r152 70 94 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=6.315 $Y=3.33
+ $X2=6.482 $Y2=3.33
r153 70 75 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.315 $Y=3.33
+ $X2=6 $Y2=3.33
r154 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r155 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 66 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r157 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r158 65 68 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r160 63 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.74 $Y2=3.33
r161 63 65 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=2.16 $Y2=3.33
r162 61 76 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=3.33 $X2=6
+ $Y2=3.33
r163 61 73 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.08 $Y2=3.33
r164 59 72 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.08 $Y2=3.33
r165 58 68 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.6 $Y2=3.33
r166 57 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=4.045 $Y2=3.33
r167 57 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=3.715 $Y2=3.33
r168 55 57 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.88 $Y=3.015
+ $X2=3.88 $Y2=3.33
r169 50 53 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.36 $Y=1.985
+ $X2=9.36 $Y2=2.815
r170 48 103 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.36 $Y=3.245
+ $X2=9.417 $Y2=3.33
r171 48 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.36 $Y=3.245
+ $X2=9.36 $Y2=2.815
r172 44 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=3.33
r173 44 46 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=2.305
r174 43 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.48 $Y2=3.33
r175 42 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=3.33
+ $X2=8.42 $Y2=3.33
r176 42 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.335 $Y=3.33
+ $X2=7.605 $Y2=3.33
r177 38 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.48 $Y=3.245
+ $X2=7.48 $Y2=3.33
r178 38 40 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=7.48 $Y=3.245
+ $X2=7.48 $Y2=2.225
r179 34 94 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.482 $Y=3.245
+ $X2=6.482 $Y2=3.33
r180 34 36 19.9527 $w=3.33e-07 $l=5.8e-07 $layer=LI1_cond $X=6.482 $Y=3.245
+ $X2=6.482 $Y2=2.665
r181 30 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r182 30 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.03
r183 29 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r184 28 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=3.33
+ $X2=1.74 $Y2=3.33
r185 28 29 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.655 $Y=3.33
+ $X2=0.815 $Y2=3.33
r186 24 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r187 24 26 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r188 7 53 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.185
+ $Y=1.84 $X2=9.32 $Y2=2.815
r189 7 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.185
+ $Y=1.84 $X2=9.32 $Y2=1.985
r190 6 46 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=8.285
+ $Y=1.84 $X2=8.42 $Y2=2.305
r191 5 40 300 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_PDIFF $count=2 $X=7.3
+ $Y=2.12 $X2=7.52 $Y2=2.225
r192 4 36 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=2.54 $X2=6.485 $Y2=2.665
r193 3 55 600 $w=1.7e-07 $l=6e-07 $layer=licon1_PDIFF $count=1 $X=3.66 $Y=2.515
+ $X2=3.88 $Y2=3.015
r194 2 32 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.515 $X2=1.74 $Y2=3.03
r195 1 26 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%A_440_503# 1 2 9 12 13 14 17 21
c48 21 0 2.95165e-20 $X=2.56 $Y=2.035
r49 19 21 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.42 $Y=2.035
+ $X2=2.56 $Y2=2.035
r50 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.91 $Y=1.07
+ $X2=2.91 $Y2=0.815
r51 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.825 $Y=1.155
+ $X2=2.91 $Y2=1.07
r52 13 14 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.825 $Y=1.155
+ $X2=2.645 $Y2=1.155
r53 12 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=1.95
+ $X2=2.56 $Y2=2.035
r54 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=1.24
+ $X2=2.645 $Y2=1.155
r55 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.56 $Y=1.24
+ $X2=2.56 $Y2=1.95
r56 7 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=2.12 $X2=2.42
+ $Y2=2.035
r57 7 9 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.42 $Y=2.12 $X2=2.42
+ $Y2=2.57
r58 2 9 600 $w=1.7e-07 $l=2.45967e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=2.515 $X2=2.42 $Y2=2.57
r59 1 17 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.595 $X2=2.91 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%Q 1 2 3 4 15 21 23 24 25 26 29 32 33 34 35
+ 36 44
r79 41 44 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.87 $Y=1.97
+ $X2=8.87 $Y2=1.985
r80 35 36 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.87 $Y=2.405
+ $X2=8.87 $Y2=2.775
r81 34 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=1.885
+ $X2=8.87 $Y2=1.97
r82 34 35 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.87 $Y=2.045
+ $X2=8.87 $Y2=2.405
r83 34 44 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=8.87 $Y=2.045 $X2=8.87
+ $Y2=1.985
r84 32 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.95 $Y=1.8
+ $X2=8.87 $Y2=1.885
r85 31 33 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=8.95 $Y=1.13
+ $X2=8.867 $Y2=1.045
r86 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.95 $Y=1.13
+ $X2=8.95 $Y2=1.8
r87 27 33 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=8.867 $Y=0.96
+ $X2=8.867 $Y2=1.045
r88 27 29 15.3086 $w=3.33e-07 $l=4.45e-07 $layer=LI1_cond $X=8.867 $Y=0.96
+ $X2=8.867 $Y2=0.515
r89 25 33 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=8.7 $Y=1.045
+ $X2=8.867 $Y2=1.045
r90 25 26 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.7 $Y=1.045
+ $X2=8.15 $Y2=1.045
r91 23 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.885
+ $X2=8.87 $Y2=1.885
r92 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.705 $Y=1.885
+ $X2=8.135 $Y2=1.885
r93 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.985 $Y=0.96
+ $X2=8.15 $Y2=1.045
r94 19 21 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.985 $Y=0.96
+ $X2=7.985 $Y2=0.515
r95 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.97 $Y=1.985
+ $X2=7.97 $Y2=2.815
r96 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.97 $Y=1.97
+ $X2=8.135 $Y2=1.885
r97 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.97 $Y=1.97
+ $X2=7.97 $Y2=1.985
r98 4 36 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.735
+ $Y=1.84 $X2=8.87 $Y2=2.815
r99 4 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.735
+ $Y=1.84 $X2=8.87 $Y2=1.985
r100 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.835
+ $Y=1.84 $X2=7.97 $Y2=2.815
r101 3 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.835
+ $Y=1.84 $X2=7.97 $Y2=1.985
r102 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.725
+ $Y=0.37 $X2=8.865 $Y2=0.515
r103 1 21 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=7.805
+ $Y=0.37 $X2=7.985 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 46 48
+ 50 53 54 55 57 62 74 78 83 89 92 95 98 101 105
r132 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r133 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r134 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r135 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r136 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r137 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r138 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r139 87 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r140 87 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r141 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r142 84 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.5 $Y=0 $X2=8.415
+ $Y2=0
r143 84 86 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.5 $Y=0 $X2=8.88
+ $Y2=0
r144 83 104 3.97976 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=9.21 $Y=0
+ $X2=9.405 $Y2=0
r145 83 86 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.21 $Y=0 $X2=8.88
+ $Y2=0
r146 82 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r147 82 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r148 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r149 79 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=0 $X2=6.535
+ $Y2=0
r150 79 81 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.66 $Y=0 $X2=6.96
+ $Y2=0
r151 78 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=0 $X2=7.485
+ $Y2=0
r152 78 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.32 $Y=0 $X2=6.96
+ $Y2=0
r153 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r154 74 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.535
+ $Y2=0
r155 74 76 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=6.41 $Y=0 $X2=4.56
+ $Y2=0
r156 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r157 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r158 70 73 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.08 $Y2=0
r159 70 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r160 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r161 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r162 67 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r163 67 69 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.64 $Y2=0
r164 66 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r165 66 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r166 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r167 63 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.71
+ $Y2=0
r168 63 65 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r169 62 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r170 62 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.68 $Y2=0
r171 60 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r173 57 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.71
+ $Y2=0
r174 57 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r175 55 96 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6.48
+ $Y2=0
r176 55 77 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r177 53 72 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.08
+ $Y2=0
r178 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.215
+ $Y2=0
r179 52 76 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.34 $Y=0 $X2=4.56
+ $Y2=0
r180 52 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.34 $Y=0 $X2=4.215
+ $Y2=0
r181 48 104 3.1634 $w=2.5e-07 $l=1.14782e-07 $layer=LI1_cond $X=9.335 $Y=0.085
+ $X2=9.405 $Y2=0
r182 48 50 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.335 $Y=0.085
+ $X2=9.335 $Y2=0.515
r183 44 101 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.415 $Y=0.085
+ $X2=8.415 $Y2=0
r184 44 46 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.415 $Y=0.085
+ $X2=8.415 $Y2=0.57
r185 43 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=0 $X2=7.485
+ $Y2=0
r186 42 101 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=0 $X2=8.415
+ $Y2=0
r187 42 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.33 $Y=0 $X2=7.65
+ $Y2=0
r188 38 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0
r189 38 40 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0.53
r190 34 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=0.085
+ $X2=6.535 $Y2=0
r191 34 36 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=6.535 $Y=0.085
+ $X2=6.535 $Y2=0.785
r192 30 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r193 30 32 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.355
r194 26 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r195 26 28 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.475
r196 22 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r197 22 24 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.57
r198 7 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.155
+ $Y=0.37 $X2=9.295 $Y2=0.515
r199 6 46 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=8.275
+ $Y=0.37 $X2=8.415 $Y2=0.57
r200 5 40 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.37 $X2=7.485 $Y2=0.53
r201 4 36 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.62 $X2=6.495 $Y2=0.785
r202 3 32 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.51 $X2=4.255 $Y2=0.355
r203 2 28 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.33 $X2=2.15 $Y2=0.475
r204 1 24 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.57
.ends


* File: sky130_fd_sc_ms__and2_2.pxi.spice
* Created: Wed Sep  2 11:57:05 2020
* 
x_PM_SKY130_FD_SC_MS__AND2_2%A N_A_M1002_g N_A_M1006_g A N_A_c_53_n N_A_c_54_n
+ PM_SKY130_FD_SC_MS__AND2_2%A
x_PM_SKY130_FD_SC_MS__AND2_2%B N_B_M1003_g N_B_M1000_g B N_B_c_78_n N_B_c_79_n
+ PM_SKY130_FD_SC_MS__AND2_2%B
x_PM_SKY130_FD_SC_MS__AND2_2%A_31_74# N_A_31_74#_M1006_s N_A_31_74#_M1002_d
+ N_A_31_74#_c_118_n N_A_31_74#_M1005_g N_A_31_74#_M1001_g N_A_31_74#_c_120_n
+ N_A_31_74#_M1007_g N_A_31_74#_M1004_g N_A_31_74#_c_122_n N_A_31_74#_c_123_n
+ N_A_31_74#_c_124_n N_A_31_74#_c_130_n N_A_31_74#_c_131_n N_A_31_74#_c_132_n
+ N_A_31_74#_c_125_n N_A_31_74#_c_126_n N_A_31_74#_c_127_n
+ PM_SKY130_FD_SC_MS__AND2_2%A_31_74#
x_PM_SKY130_FD_SC_MS__AND2_2%VPWR N_VPWR_M1002_s N_VPWR_M1000_d N_VPWR_M1004_s
+ N_VPWR_c_210_n N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_214_n
+ VPWR N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_209_n
+ PM_SKY130_FD_SC_MS__AND2_2%VPWR
x_PM_SKY130_FD_SC_MS__AND2_2%X N_X_M1005_d N_X_M1001_d N_X_c_247_n N_X_c_248_n
+ N_X_c_250_n X X X PM_SKY130_FD_SC_MS__AND2_2%X
x_PM_SKY130_FD_SC_MS__AND2_2%VGND N_VGND_M1003_d N_VGND_M1007_s N_VGND_c_281_n
+ N_VGND_c_282_n N_VGND_c_283_n VGND N_VGND_c_284_n N_VGND_c_285_n
+ N_VGND_c_286_n N_VGND_c_287_n PM_SKY130_FD_SC_MS__AND2_2%VGND
cc_1 VNB N_A_M1002_g 0.00192204f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_2 VNB N_A_M1006_g 0.0297549f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A_c_53_n 0.0050357f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A_c_54_n 0.0582209f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_5 VNB N_B_M1003_g 0.0215375f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_6 VNB N_B_M1000_g 0.00136699f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_7 VNB N_B_c_78_n 0.0291241f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_8 VNB N_B_c_79_n 0.00419749f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_9 VNB N_A_31_74#_c_118_n 0.0174733f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_10 VNB N_A_31_74#_M1001_g 0.00527962f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_11 VNB N_A_31_74#_c_120_n 0.0188592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_31_74#_M1004_g 0.0070533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_31_74#_c_122_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_31_74#_c_123_n 0.00780948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_31_74#_c_124_n 0.00898165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_31_74#_c_125_n 0.00473431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_31_74#_c_126_n 6.4908e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_31_74#_c_127_n 0.0442792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_209_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_247_n 0.00239236f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_21 VNB N_X_c_248_n 0.0188945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_281_n 0.006479f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_VGND_c_282_n 0.0118321f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_24 VNB N_VGND_c_283_n 0.0255459f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_25 VNB N_VGND_c_284_n 0.029813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_285_n 0.0193156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_286_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_287_n 0.166974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VPB N_A_M1002_g 0.0377146f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.46
cc_30 VPB N_A_c_53_n 0.00745299f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_31 VPB N_B_M1000_g 0.0295524f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_32 VPB N_B_c_79_n 0.00533013f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_33 VPB N_A_31_74#_M1001_g 0.021717f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_34 VPB N_A_31_74#_M1004_g 0.0246413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_31_74#_c_130_n 0.00197168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_31_74#_c_131_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_31_74#_c_132_n 6.18427e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_31_74#_c_126_n 0.00133441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_210_n 0.0117348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_211_n 0.0498848f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_41 VPB N_VPWR_c_212_n 0.00505006f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_42 VPB N_VPWR_c_213_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_43 VPB N_VPWR_c_214_n 0.0461845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_215_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_216_n 0.0186844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_217_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_209_n 0.0545021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_X_c_248_n 0.00210119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_X_c_250_n 0.00957709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB X 0.00202446f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_51 N_A_M1006_g N_B_M1003_g 0.0550561f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_52 N_A_M1002_g N_B_M1000_g 0.0212009f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_53 N_A_c_53_n N_B_c_78_n 2.28826e-19 $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_54 N_A_c_54_n N_B_c_78_n 0.0209293f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_55 N_A_c_53_n N_B_c_79_n 0.0391299f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_56 N_A_c_54_n N_B_c_79_n 0.00404395f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_57 N_A_M1006_g N_A_31_74#_c_122_n 0.012125f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_58 N_A_M1006_g N_A_31_74#_c_123_n 0.0146407f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_59 N_A_M1006_g N_A_31_74#_c_124_n 0.00206782f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_60 N_A_c_53_n N_A_31_74#_c_124_n 0.0260039f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_61 N_A_c_54_n N_A_31_74#_c_124_n 0.00265455f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_VPWR_c_211_n 0.0183728f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_63 N_A_c_53_n N_VPWR_c_211_n 0.0292783f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_64 N_A_c_54_n N_VPWR_c_211_n 0.00165041f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_65 N_A_M1002_g N_VPWR_c_215_n 0.00460063f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_66 N_A_M1002_g N_VPWR_c_209_n 0.00908665f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_67 N_A_M1006_g N_VGND_c_281_n 0.00180653f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A_M1006_g N_VGND_c_284_n 0.00434272f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_69 N_A_M1006_g N_VGND_c_287_n 0.00824704f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_70 N_B_M1003_g N_A_31_74#_c_118_n 0.0259185f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_71 N_B_M1000_g N_A_31_74#_M1001_g 0.0270014f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_72 N_B_c_78_n N_A_31_74#_M1001_g 0.00425961f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_73 N_B_c_79_n N_A_31_74#_M1001_g 5.21976e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_74 N_B_M1003_g N_A_31_74#_c_122_n 0.00208517f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_75 N_B_M1003_g N_A_31_74#_c_123_n 0.0144246f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_76 N_B_c_78_n N_A_31_74#_c_123_n 0.00495365f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_77 N_B_c_79_n N_A_31_74#_c_123_n 0.0374224f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_78 N_B_M1000_g N_A_31_74#_c_130_n 9.78681e-19 $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_79 N_B_c_78_n N_A_31_74#_c_130_n 3.30055e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_80 N_B_c_79_n N_A_31_74#_c_130_n 0.0224585f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_81 N_B_M1000_g N_A_31_74#_c_131_n 0.0115053f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_82 N_B_M1000_g N_A_31_74#_c_132_n 0.0132049f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_83 N_B_c_78_n N_A_31_74#_c_132_n 0.00166044f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_84 N_B_c_79_n N_A_31_74#_c_132_n 0.0146867f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_85 N_B_M1003_g N_A_31_74#_c_125_n 0.00350413f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_86 N_B_c_78_n N_A_31_74#_c_125_n 0.00159524f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_87 N_B_c_79_n N_A_31_74#_c_125_n 0.0208197f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_88 N_B_M1000_g N_A_31_74#_c_126_n 0.00386696f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_89 N_B_c_78_n N_A_31_74#_c_126_n 4.8742e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_90 N_B_c_79_n N_A_31_74#_c_126_n 0.0184081f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_91 N_B_c_78_n N_A_31_74#_c_127_n 0.0155883f $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_92 N_B_c_79_n N_A_31_74#_c_127_n 2.4048e-19 $X=0.965 $Y=1.465 $X2=0 $Y2=0
cc_93 N_B_M1000_g N_VPWR_c_211_n 6.67731e-19 $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_94 N_B_M1000_g N_VPWR_c_212_n 0.0018933f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_95 N_B_M1000_g N_VPWR_c_215_n 0.005209f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_96 N_B_M1000_g N_VPWR_c_209_n 0.00982314f $X=0.95 $Y=2.46 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_VGND_c_281_n 0.0120683f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B_M1003_g N_VGND_c_284_n 0.00383152f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B_M1003_g N_VGND_c_287_n 0.0075725f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_31_74#_c_132_n N_VPWR_M1000_d 0.00717204f $X=1.255 $Y=2.035 $X2=0
+ $Y2=0
cc_101 N_A_31_74#_c_126_n N_VPWR_M1000_d 0.00130575f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_102 N_A_31_74#_c_130_n N_VPWR_c_211_n 0.00599715f $X=0.765 $Y=2.12 $X2=0
+ $Y2=0
cc_103 N_A_31_74#_c_131_n N_VPWR_c_211_n 0.029009f $X=0.725 $Y=2.815 $X2=0 $Y2=0
cc_104 N_A_31_74#_M1001_g N_VPWR_c_212_n 0.012533f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_31_74#_M1004_g N_VPWR_c_212_n 5.69853e-19 $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_31_74#_c_131_n N_VPWR_c_212_n 0.0256025f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_107 N_A_31_74#_c_132_n N_VPWR_c_212_n 0.019541f $X=1.255 $Y=2.035 $X2=0 $Y2=0
cc_108 N_A_31_74#_M1004_g N_VPWR_c_214_n 0.00772239f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_31_74#_c_131_n N_VPWR_c_215_n 0.0109793f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_110 N_A_31_74#_M1001_g N_VPWR_c_216_n 0.00475445f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_31_74#_M1004_g N_VPWR_c_216_n 0.005209f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_31_74#_M1001_g N_VPWR_c_209_n 0.00938661f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_31_74#_M1004_g N_VPWR_c_209_n 0.00985972f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_31_74#_c_131_n N_VPWR_c_209_n 0.00901959f $X=0.725 $Y=2.815 $X2=0
+ $Y2=0
cc_115 N_A_31_74#_c_118_n N_X_c_247_n 0.0105697f $X=1.415 $Y=1.22 $X2=0 $Y2=0
cc_116 N_A_31_74#_c_120_n N_X_c_247_n 0.0249871f $X=1.845 $Y=1.22 $X2=0 $Y2=0
cc_117 N_A_31_74#_c_125_n N_X_c_247_n 0.0126837f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_118 N_A_31_74#_c_127_n N_X_c_247_n 0.0010614f $X=1.905 $Y=1.385 $X2=0 $Y2=0
cc_119 N_A_31_74#_c_118_n N_X_c_248_n 6.22718e-19 $X=1.415 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A_31_74#_M1001_g N_X_c_248_n 5.98575e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_31_74#_c_120_n N_X_c_248_n 0.00695403f $X=1.845 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A_31_74#_M1004_g N_X_c_248_n 0.00706636f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_31_74#_c_125_n N_X_c_248_n 0.0311249f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_124 N_A_31_74#_c_126_n N_X_c_248_n 0.00557352f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_125 N_A_31_74#_c_127_n N_X_c_248_n 0.0155244f $X=1.905 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_31_74#_M1001_g N_X_c_250_n 9.17904e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_31_74#_M1004_g N_X_c_250_n 0.0146393f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_31_74#_c_125_n N_X_c_250_n 0.00566518f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_129 N_A_31_74#_c_126_n N_X_c_250_n 0.0108281f $X=1.34 $Y=1.95 $X2=0 $Y2=0
cc_130 N_A_31_74#_c_127_n N_X_c_250_n 0.00249017f $X=1.905 $Y=1.385 $X2=0 $Y2=0
cc_131 N_A_31_74#_M1001_g X 3.6964e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_31_74#_M1004_g X 0.0197415f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_31_74#_c_123_n A_118_74# 0.0048076f $X=1.255 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_31_74#_c_123_n N_VGND_M1003_d 0.00230675f $X=1.255 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_31_74#_c_125_n N_VGND_M1003_d 3.09855e-19 $X=1.34 $Y=1.55 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_31_74#_c_118_n N_VGND_c_281_n 0.00543307f $X=1.415 $Y=1.22 $X2=0
+ $Y2=0
cc_137 N_A_31_74#_c_122_n N_VGND_c_281_n 0.0139395f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_138 N_A_31_74#_c_123_n N_VGND_c_281_n 0.0195279f $X=1.255 $Y=1.045 $X2=0
+ $Y2=0
cc_139 N_A_31_74#_c_125_n N_VGND_c_281_n 0.00252453f $X=1.34 $Y=1.55 $X2=0 $Y2=0
cc_140 N_A_31_74#_c_120_n N_VGND_c_283_n 0.00500034f $X=1.845 $Y=1.22 $X2=0
+ $Y2=0
cc_141 N_A_31_74#_c_122_n N_VGND_c_284_n 0.0145639f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_142 N_A_31_74#_c_118_n N_VGND_c_285_n 0.00433139f $X=1.415 $Y=1.22 $X2=0
+ $Y2=0
cc_143 N_A_31_74#_c_120_n N_VGND_c_285_n 0.00433139f $X=1.845 $Y=1.22 $X2=0
+ $Y2=0
cc_144 N_A_31_74#_c_118_n N_VGND_c_287_n 0.00817409f $X=1.415 $Y=1.22 $X2=0
+ $Y2=0
cc_145 N_A_31_74#_c_120_n N_VGND_c_287_n 0.00451721f $X=1.845 $Y=1.22 $X2=0
+ $Y2=0
cc_146 N_A_31_74#_c_122_n N_VGND_c_287_n 0.0119984f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_147 N_VPWR_c_212_n X 0.022953f $X=1.225 $Y=2.455 $X2=0 $Y2=0
cc_148 N_VPWR_c_214_n X 0.0297232f $X=2.13 $Y=2.225 $X2=0 $Y2=0
cc_149 N_VPWR_c_216_n X 0.0109793f $X=2.045 $Y=3.33 $X2=0 $Y2=0
cc_150 N_VPWR_c_209_n X 0.00901959f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_151 N_X_c_247_n N_VGND_M1007_s 0.00752423f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_152 N_X_c_248_n N_VGND_M1007_s 0.00339584f $X=1.925 $Y=1.72 $X2=0 $Y2=0
cc_153 N_X_c_247_n N_VGND_c_281_n 0.0166176f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_154 N_X_c_247_n N_VGND_c_283_n 0.0155529f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_155 N_X_c_247_n N_VGND_c_285_n 0.0143518f $X=1.925 $Y=1.02 $X2=0 $Y2=0
cc_156 N_X_c_247_n N_VGND_c_287_n 0.0179048f $X=1.925 $Y=1.02 $X2=0 $Y2=0

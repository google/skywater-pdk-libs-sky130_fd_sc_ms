* File: sky130_fd_sc_ms__or4bb_1.spice
* Created: Wed Sep  2 12:29:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4bb_1.pex.spice"
.subckt sky130_fd_sc_ms__or4bb_1  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_C_N_M1004_g N_A_27_424#_M1004_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.1155 AS=0.15675 PD=0.97 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1008 N_A_219_424#_M1008_d N_D_N_M1008_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.15675 AS=0.1155 PD=1.67 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.8 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_357_378#_M1000_d N_A_219_424#_M1000_g N_VGND_M1000_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.092125 AS=0.165 PD=0.885 PS=1.7 NRD=11.988 NRS=3.264 M=1
+ R=3.66667 SA=75000.2 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1013 N_VGND_M1013_d N_A_27_424#_M1013_g N_A_357_378#_M1000_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.114125 AS=0.092125 PD=0.965 PS=0.885 NRD=21.816 NRS=0 M=1
+ R=3.66667 SA=75000.7 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1010 N_A_357_378#_M1010_d N_B_M1010_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.114125 PD=0.9 PS=0.965 NRD=15.264 NRS=7.632 M=1 R=3.66667
+ SA=75001.3 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_357_378#_M1010_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.126948 AS=0.09625 PD=1.01899 PS=0.9 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.8 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1011 N_X_M1011_d N_A_357_378#_M1011_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.170802 PD=2.05 PS=1.37101 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_C_N_M1005_g N_A_27_424#_M1005_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2352 PD=1.16 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1003 N_A_219_424#_M1003_d N_D_N_M1003_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=0.84 AD=0.42525 AS=0.1344 PD=2.94 PS=1.16 NRD=105.828 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1012 A_449_378# N_A_219_424#_M1012_g N_A_357_378#_M1012_s VPB PSHORT L=0.18
+ W=1 AD=0.12 AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1002 A_533_378# N_A_27_424#_M1002_g A_449_378# VPB PSHORT L=0.18 W=1 AD=0.15
+ AS=0.12 PD=1.3 PS=1.24 NRD=18.6953 NRS=12.7853 M=1 R=5.55556 SA=90000.6
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1001 A_629_378# N_B_M1001_g A_533_378# VPB PSHORT L=0.18 W=1 AD=0.18 AS=0.15
+ PD=1.36 PS=1.3 NRD=24.6053 NRS=18.6953 M=1 R=5.55556 SA=90001.1 SB=90001.3
+ A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_629_378# VPB PSHORT L=0.18 W=1 AD=0.20783
+ AS=0.18 PD=1.43868 PS=1.36 NRD=16.0752 NRS=24.6053 M=1 R=5.55556 SA=90001.6
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1007_d N_A_357_378#_M1007_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.23277 PD=2.8 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__or4bb_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor2_4.pxi.spice
* Created: Fri Aug 28 17:46:40 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2_4%A N_A_M1000_g N_A_c_57_n N_A_M1002_g N_A_M1001_g
+ N_A_M1003_g N_A_c_60_n N_A_M1004_g N_A_M1006_g A A A A N_A_c_63_n
+ PM_SKY130_FD_SC_MS__NOR2_4%A
x_PM_SKY130_FD_SC_MS__NOR2_4%B N_B_c_127_n N_B_M1005_g N_B_M1007_g N_B_c_129_n
+ N_B_M1011_g N_B_M1008_g N_B_M1009_g N_B_M1010_g B B B N_B_c_134_n
+ PM_SKY130_FD_SC_MS__NOR2_4%B
x_PM_SKY130_FD_SC_MS__NOR2_4%A_27_368# N_A_27_368#_M1000_s N_A_27_368#_M1001_s
+ N_A_27_368#_M1006_s N_A_27_368#_M1008_s N_A_27_368#_M1010_s
+ N_A_27_368#_c_193_n N_A_27_368#_c_194_n N_A_27_368#_c_195_n
+ N_A_27_368#_c_196_n N_A_27_368#_c_197_n N_A_27_368#_c_220_n
+ N_A_27_368#_c_198_n N_A_27_368#_c_199_n N_A_27_368#_c_230_n
+ N_A_27_368#_c_200_n N_A_27_368#_c_201_n N_A_27_368#_c_202_n
+ N_A_27_368#_c_203_n PM_SKY130_FD_SC_MS__NOR2_4%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR2_4%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_c_267_n
+ N_VPWR_c_268_n VPWR N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_266_n
+ N_VPWR_c_272_n N_VPWR_c_273_n PM_SKY130_FD_SC_MS__NOR2_4%VPWR
x_PM_SKY130_FD_SC_MS__NOR2_4%Y N_Y_M1002_s N_Y_M1005_d N_Y_M1007_d N_Y_M1009_d
+ N_Y_c_314_n N_Y_c_321_n N_Y_c_315_n N_Y_c_324_n N_Y_c_327_n N_Y_c_329_n
+ N_Y_c_317_n N_Y_c_351_n N_Y_c_316_n N_Y_c_352_n Y PM_SKY130_FD_SC_MS__NOR2_4%Y
x_PM_SKY130_FD_SC_MS__NOR2_4%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_M1011_s
+ N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n
+ VGND N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n
+ PM_SKY130_FD_SC_MS__NOR2_4%VGND
cc_1 VNB N_A_M1000_g 0.00916985f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_c_57_n 0.0266014f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_3 VNB N_A_M1001_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_4 VNB N_A_M1003_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_5 VNB N_A_c_60_n 0.0227304f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.22
cc_6 VNB N_A_M1006_g 0.00599174f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_7 VNB A 0.0340492f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_8 VNB N_A_c_63_n 0.105395f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.385
cc_9 VNB N_B_c_127_n 0.0176155f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_10 VNB N_B_M1007_g 0.00554239f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_11 VNB N_B_c_129_n 0.0197009f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.55
cc_12 VNB N_B_M1008_g 0.00556397f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_13 VNB N_B_M1009_g 0.00623425f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_14 VNB N_B_M1010_g 0.0093909f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_15 VNB B 0.0270754f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_16 VNB N_B_c_134_n 0.147128f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.385
cc_17 VNB N_VPWR_c_266_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_314_n 0.00695126f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_19 VNB N_Y_c_315_n 0.00257348f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_20 VNB N_Y_c_316_n 0.00334407f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.385
cc_21 VNB N_VGND_c_373_n 0.0125081f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_22 VNB N_VGND_c_374_n 0.0352733f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.55
cc_23 VNB N_VGND_c_375_n 0.00571115f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.22
cc_24 VNB N_VGND_c_376_n 0.0355045f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.55
cc_25 VNB N_VGND_c_377_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_26 VNB N_VGND_c_378_n 0.0186748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_379_n 0.082553f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_28 VNB N_VGND_c_380_n 0.244311f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_29 VPB N_A_M1000_g 0.0287755f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_30 VPB N_A_M1001_g 0.0213904f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_31 VPB N_A_M1003_g 0.0213904f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_32 VPB N_A_M1006_g 0.0211395f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_33 VPB N_B_M1007_g 0.0211133f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_34 VPB N_B_M1008_g 0.0208881f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_35 VPB N_B_M1009_g 0.0217507f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_36 VPB N_B_M1010_g 0.0289426f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_37 VPB N_A_27_368#_c_193_n 0.0439896f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_38 VPB N_A_27_368#_c_194_n 0.00219429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_368#_c_195_n 0.0106238f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_40 VPB N_A_27_368#_c_196_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_41 VPB N_A_27_368#_c_197_n 0.0133415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_368#_c_198_n 0.00219299f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.385
cc_43 VPB N_A_27_368#_c_199_n 0.00181992f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.385
cc_44 VPB N_A_27_368#_c_200_n 0.0096461f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_45 VPB N_A_27_368#_c_201_n 0.00313635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_368#_c_202_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_368#_c_203_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_267_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_268_n 0.00768031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_269_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.55
cc_51 VPB N_VPWR_c_270_n 0.0633787f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_52 VPB N_VPWR_c_266_n 0.0711036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_272_n 0.0233502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_273_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_55 VPB N_Y_c_317_n 0.0075476f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_56 N_A_c_60_n N_B_c_127_n 0.0145322f $X=1.81 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_57 A N_B_c_127_n 0.0014455f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_58 N_A_M1006_g N_B_M1007_g 0.0148975f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_59 N_A_c_63_n N_B_c_134_n 0.0294297f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_A_27_368#_c_193_n 0.0158419f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_A_27_368#_c_193_n 7.23242e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_A_27_368#_c_194_n 0.012931f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A_M1001_g N_A_27_368#_c_194_n 0.012931f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_64 A N_A_27_368#_c_194_n 0.042029f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_c_63_n N_A_27_368#_c_194_n 0.00201785f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_66 N_A_M1000_g N_A_27_368#_c_195_n 0.00330546f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_67 A N_A_27_368#_c_195_n 0.0282802f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_M1000_g N_A_27_368#_c_196_n 7.23242e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A_M1001_g N_A_27_368#_c_196_n 0.0152527f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_A_27_368#_c_196_n 0.0152527f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_71 N_A_M1006_g N_A_27_368#_c_196_n 7.23242e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_A_27_368#_c_197_n 0.0128923f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_M1006_g N_A_27_368#_c_197_n 0.019448f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_74 A N_A_27_368#_c_197_n 0.0334139f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_63_n N_A_27_368#_c_197_n 0.00213605f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_A_27_368#_c_220_n 7.0088e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_A_27_368#_c_220_n 0.0137286f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_78 N_A_M1006_g N_A_27_368#_c_199_n 0.00347836f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_A_27_368#_c_202_n 0.00228751f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_M1003_g N_A_27_368#_c_202_n 0.00228751f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_81 A N_A_27_368#_c_202_n 0.0277828f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_63_n N_A_27_368#_c_202_n 0.00209661f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_VPWR_c_267_n 0.00363491f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_M1001_g N_VPWR_c_267_n 0.00363491f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_VPWR_c_268_n 0.00363491f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_VPWR_c_268_n 0.00206481f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_VPWR_c_269_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VPWR_c_269_n 0.005209f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_VPWR_c_270_n 0.00517089f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_M1000_g N_VPWR_c_266_n 0.00986008f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_M1001_g N_VPWR_c_266_n 0.00982266f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_M1003_g N_VPWR_c_266_n 0.00982266f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_VPWR_c_266_n 0.00977588f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_VPWR_c_272_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A_c_57_n N_Y_c_314_n 6.72669e-19 $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_96 A N_Y_c_314_n 0.0963567f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A_c_63_n N_Y_c_314_n 0.00672026f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A_c_60_n N_Y_c_321_n 0.0125972f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_99 N_A_c_63_n N_Y_c_321_n 0.00118967f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_100 N_A_c_60_n N_Y_c_315_n 4.29877e-19 $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A_c_60_n N_Y_c_324_n 8.96662e-19 $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_102 A N_Y_c_324_n 0.00679233f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A_c_63_n N_Y_c_324_n 7.28848e-19 $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_104 A N_Y_c_327_n 0.00406857f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A_c_63_n N_Y_c_327_n 0.00132231f $X=1.81 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A_M1006_g N_Y_c_329_n 2.50368e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_c_60_n N_Y_c_316_n 6.72669e-19 $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A_c_57_n N_VGND_c_374_n 0.0148927f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_109 A N_VGND_c_374_n 0.0273236f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A_c_60_n N_VGND_c_375_n 0.0100967f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_111 N_A_c_57_n N_VGND_c_376_n 0.00383152f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_112 N_A_c_60_n N_VGND_c_376_n 0.00383152f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A_c_57_n N_VGND_c_380_n 0.00762539f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A_c_60_n N_VGND_c_380_n 0.00388966f $X=1.81 $Y=1.22 $X2=0 $Y2=0
cc_115 N_B_M1007_g N_A_27_368#_c_197_n 0.00104222f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_A_27_368#_c_198_n 0.0139468f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_117 N_B_M1008_g N_A_27_368#_c_198_n 0.0142213f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_118 N_B_M1009_g N_A_27_368#_c_230_n 0.0115473f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_119 N_B_M1010_g N_A_27_368#_c_230_n 2.72638e-19 $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_120 N_B_M1009_g N_A_27_368#_c_200_n 0.0119307f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_121 N_B_M1010_g N_A_27_368#_c_200_n 0.0152849f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B_M1010_g N_A_27_368#_c_201_n 0.00151632f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_123 B N_A_27_368#_c_201_n 0.0167379f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B_c_134_n N_A_27_368#_c_201_n 0.00612431f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_125 N_B_M1009_g N_A_27_368#_c_203_n 0.00214324f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_126 N_B_M1007_g N_VPWR_c_270_n 0.00333926f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B_M1008_g N_VPWR_c_270_n 0.00333926f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_128 N_B_M1009_g N_VPWR_c_270_n 0.00333896f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B_M1010_g N_VPWR_c_270_n 0.00333926f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_130 N_B_M1007_g N_VPWR_c_266_n 0.00422798f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_131 N_B_M1008_g N_VPWR_c_266_n 0.00423176f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_132 N_B_M1009_g N_VPWR_c_266_n 0.00423662f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_133 N_B_M1010_g N_VPWR_c_266_n 0.00427109f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_134 N_B_c_127_n N_Y_c_321_n 0.0142112f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_135 N_B_c_127_n N_Y_c_315_n 0.00694939f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_136 N_B_c_129_n N_Y_c_315_n 0.00644058f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_137 N_B_c_127_n N_Y_c_324_n 0.00476825f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_138 N_B_c_129_n N_Y_c_324_n 0.0142151f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_139 B N_Y_c_324_n 0.0137784f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B_c_134_n N_Y_c_324_n 0.0174866f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_141 N_B_M1007_g N_Y_c_327_n 0.00516617f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_142 N_B_M1008_g N_Y_c_327_n 0.00529131f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_143 N_B_M1009_g N_Y_c_327_n 7.87895e-19 $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_144 B N_Y_c_327_n 0.00682348f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_145 N_B_c_134_n N_Y_c_327_n 0.0114759f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_146 N_B_M1007_g N_Y_c_329_n 0.009838f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_147 N_B_M1008_g N_Y_c_329_n 0.0115411f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_148 N_B_M1009_g N_Y_c_329_n 2.72638e-19 $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_149 N_B_M1008_g N_Y_c_317_n 0.0161316f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_150 N_B_M1009_g N_Y_c_317_n 0.0161508f $X=3.255 $Y=2.4 $X2=0 $Y2=0
cc_151 N_B_M1010_g N_Y_c_317_n 0.00764667f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_152 B N_Y_c_317_n 0.0545029f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B_c_134_n N_Y_c_317_n 0.00746047f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_154 N_B_M1010_g N_Y_c_351_n 0.0103108f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_155 N_B_M1007_g N_Y_c_352_n 0.00329352f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_156 N_B_M1008_g N_Y_c_352_n 0.00185263f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_157 N_B_c_127_n N_VGND_c_375_n 0.00191937f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_158 N_B_c_127_n N_VGND_c_378_n 0.00456932f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_159 N_B_c_129_n N_VGND_c_378_n 0.00434272f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_160 N_B_c_129_n N_VGND_c_379_n 0.00394517f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_161 B N_VGND_c_379_n 0.104047f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B_c_134_n N_VGND_c_379_n 0.0144509f $X=4.01 $Y=1.385 $X2=0 $Y2=0
cc_163 N_B_c_127_n N_VGND_c_380_n 0.00455422f $X=2.29 $Y=1.22 $X2=0 $Y2=0
cc_164 N_B_c_129_n N_VGND_c_380_n 0.00825234f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_27_368#_c_194_n N_VPWR_M1000_d 0.00165831f $X=1.015 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_166 N_A_27_368#_c_197_n N_VPWR_M1003_d 0.00165831f $X=1.915 $Y=1.805 $X2=0
+ $Y2=0
cc_167 N_A_27_368#_c_193_n N_VPWR_c_267_n 0.0309473f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_27_368#_c_194_n N_VPWR_c_267_n 0.0126919f $X=1.015 $Y=1.805 $X2=0
+ $Y2=0
cc_169 N_A_27_368#_c_196_n N_VPWR_c_267_n 0.0309473f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_27_368#_c_196_n N_VPWR_c_268_n 0.0309473f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_27_368#_c_197_n N_VPWR_c_268_n 0.0126919f $X=1.915 $Y=1.805 $X2=0
+ $Y2=0
cc_172 N_A_27_368#_c_199_n N_VPWR_c_268_n 0.0101219f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_173 N_A_27_368#_c_196_n N_VPWR_c_269_n 0.0144623f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_368#_c_198_n N_VPWR_c_270_n 0.0420278f $X=2.865 $Y=2.99 $X2=0
+ $Y2=0
cc_175 N_A_27_368#_c_199_n N_VPWR_c_270_n 0.0199669f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_176 N_A_27_368#_c_200_n N_VPWR_c_270_n 0.0622165f $X=3.865 $Y=2.99 $X2=0
+ $Y2=0
cc_177 N_A_27_368#_c_203_n N_VPWR_c_270_n 0.0235512f $X=3.03 $Y=2.99 $X2=0 $Y2=0
cc_178 N_A_27_368#_c_193_n N_VPWR_c_266_n 0.0119743f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_27_368#_c_196_n N_VPWR_c_266_n 0.0118344f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_27_368#_c_198_n N_VPWR_c_266_n 0.0235408f $X=2.865 $Y=2.99 $X2=0
+ $Y2=0
cc_181 N_A_27_368#_c_199_n N_VPWR_c_266_n 0.0107485f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_182 N_A_27_368#_c_200_n N_VPWR_c_266_n 0.0345671f $X=3.865 $Y=2.99 $X2=0
+ $Y2=0
cc_183 N_A_27_368#_c_203_n N_VPWR_c_266_n 0.0126924f $X=3.03 $Y=2.99 $X2=0 $Y2=0
cc_184 N_A_27_368#_c_193_n N_VPWR_c_272_n 0.014549f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_27_368#_c_198_n N_Y_M1007_d 0.00165831f $X=2.865 $Y=2.99 $X2=0 $Y2=0
cc_186 N_A_27_368#_c_200_n N_Y_M1009_d 0.00218982f $X=3.865 $Y=2.99 $X2=0 $Y2=0
cc_187 N_A_27_368#_c_198_n N_Y_c_329_n 0.0159318f $X=2.865 $Y=2.99 $X2=0 $Y2=0
cc_188 N_A_27_368#_M1008_s N_Y_c_317_n 0.00218982f $X=2.845 $Y=1.84 $X2=0 $Y2=0
cc_189 N_A_27_368#_c_230_n N_Y_c_317_n 0.0189268f $X=3.03 $Y=2.145 $X2=0 $Y2=0
cc_190 N_A_27_368#_c_201_n N_Y_c_317_n 0.00372299f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_27_368#_c_200_n N_Y_c_351_n 0.0177084f $X=3.865 $Y=2.99 $X2=0 $Y2=0
cc_192 N_A_27_368#_c_197_n N_Y_c_352_n 0.0127663f $X=1.915 $Y=1.805 $X2=0 $Y2=0
cc_193 N_Y_c_321_n N_VGND_M1004_d 0.0103921f $X=2.36 $Y=0.925 $X2=0 $Y2=0
cc_194 N_Y_c_314_n N_VGND_c_374_n 0.0267724f $X=1.355 $Y=0.675 $X2=0 $Y2=0
cc_195 N_Y_c_321_n N_VGND_c_375_n 0.0189346f $X=2.36 $Y=0.925 $X2=0 $Y2=0
cc_196 N_Y_c_315_n N_VGND_c_375_n 0.0127976f $X=2.525 $Y=0.515 $X2=0 $Y2=0
cc_197 N_Y_c_316_n N_VGND_c_375_n 0.0137088f $X=1.69 $Y=0.675 $X2=0 $Y2=0
cc_198 N_Y_c_314_n N_VGND_c_376_n 0.0485195f $X=1.355 $Y=0.675 $X2=0 $Y2=0
cc_199 N_Y_c_315_n N_VGND_c_378_n 0.014552f $X=2.525 $Y=0.515 $X2=0 $Y2=0
cc_200 N_Y_c_315_n N_VGND_c_379_n 0.0193213f $X=2.525 $Y=0.515 $X2=0 $Y2=0
cc_201 N_Y_c_314_n N_VGND_c_380_n 0.0389588f $X=1.355 $Y=0.675 $X2=0 $Y2=0
cc_202 N_Y_c_321_n N_VGND_c_380_n 0.0108653f $X=2.36 $Y=0.925 $X2=0 $Y2=0
cc_203 N_Y_c_315_n N_VGND_c_380_n 0.0119791f $X=2.525 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dlrtp_1.pex.spice
* Created: Fri Aug 28 17:28:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRTP_1%D 3 7 9 13 14
r27 12 14 33.413 $w=3.39e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.54
+ $X2=0.505 $Y2=1.54
r28 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r29 9 13 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=0.24 $Y=1.665 $X2=0.24
+ $Y2=1.465
r30 5 14 13.5074 $w=3.39e-07 $l=2.83549e-07 $layer=POLY_cond $X=0.6 $Y=1.3
+ $X2=0.505 $Y2=1.54
r31 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.6 $Y=1.3 $X2=0.6
+ $Y2=0.835
r32 1 14 17.5597 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=1.54
r33 1 3 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%GATE 3 7 9 16
c37 7 0 7.12951e-20 $X=1.185 $Y=0.74
r38 14 16 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.095 $Y=1.615
+ $X2=1.185 $Y2=1.615
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.615 $X2=1.095 $Y2=1.615
r40 11 14 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.005 $Y=1.615
+ $X2=1.095 $Y2=1.615
r41 9 15 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.095 $Y2=1.615
r42 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.45
+ $X2=1.185 $Y2=1.615
r43 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.185 $Y=1.45
+ $X2=1.185 $Y2=0.74
r44 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.78
+ $X2=1.005 $Y2=1.615
r45 1 3 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=1.005 $Y=1.78
+ $X2=1.005 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%A_219_424# 1 2 7 11 15 17 19 20 21 24 26 27
+ 33 38 39 43 44 47 50 52 55 56 57 59
c147 56 0 1.3812e-19 $X=3.93 $Y=1.39
c148 55 0 6.93786e-20 $X=3.93 $Y=1.39
c149 42 0 5.47968e-20 $X=2.935 $Y=0.77
c150 21 0 2.77549e-19 $X=3.275 $Y=1.765
r151 55 57 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=1.39
+ $X2=3.965 $Y2=1.225
r152 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.39 $X2=3.93 $Y2=1.39
r153 51 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.665 $Y=1.615
+ $X2=1.665 $Y2=1.525
r154 50 53 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.642 $Y=1.615
+ $X2=1.642 $Y2=1.78
r155 50 52 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.642 $Y=1.615
+ $X2=1.642 $Y2=1.45
r156 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.615 $X2=1.665 $Y2=1.615
r157 48 52 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.54 $Y=1.13
+ $X2=1.54 $Y2=1.45
r158 47 48 11.8581 $w=3.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.43 $Y=0.855
+ $X2=1.43 $Y2=1.13
r159 45 57 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.92 $Y=0.425
+ $X2=3.92 $Y2=1.225
r160 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.835 $Y=0.34
+ $X2=3.92 $Y2=0.425
r161 43 44 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.835 $Y=0.34
+ $X2=3.02 $Y2=0.34
r162 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.935 $Y=0.425
+ $X2=3.02 $Y2=0.34
r163 41 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.935 $Y=0.425
+ $X2=2.935 $Y2=0.77
r164 40 47 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.625 $Y=0.855
+ $X2=1.43 $Y2=0.855
r165 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.85 $Y=0.855
+ $X2=2.935 $Y2=0.77
r166 39 40 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=2.85 $Y=0.855
+ $X2=1.625 $Y2=0.855
r167 38 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=1.97
+ $X2=1.54 $Y2=1.78
r168 31 47 2.51173 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.43 $Y=0.77
+ $X2=1.43 $Y2=0.855
r169 31 33 7.5352 $w=3.88e-07 $l=2.55e-07 $layer=LI1_cond $X=1.43 $Y=0.77
+ $X2=1.43 $Y2=0.515
r170 27 38 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.455 $Y=2.095
+ $X2=1.54 $Y2=1.97
r171 27 29 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=1.455 $Y=2.095
+ $X2=1.355 $Y2=2.095
r172 22 56 38.6777 $w=2.84e-07 $l=2.18746e-07 $layer=POLY_cond $X=3.77 $Y=1.225
+ $X2=3.895 $Y2=1.39
r173 22 24 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.77 $Y=1.225
+ $X2=3.77 $Y2=0.58
r174 20 56 63.6444 $w=2.84e-07 $l=4.64354e-07 $layer=POLY_cond $X=3.695 $Y=1.765
+ $X2=3.895 $Y2=1.39
r175 20 21 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.695 $Y=1.765
+ $X2=3.275 $Y2=1.765
r176 17 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.185 $Y=1.84
+ $X2=3.275 $Y2=1.765
r177 17 19 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.185 $Y=1.84
+ $X2=3.185 $Y2=2.46
r178 13 26 18.8402 $w=1.65e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.24 $Y=1.45
+ $X2=2.205 $Y2=1.525
r179 13 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.24 $Y=1.45
+ $X2=2.24 $Y2=0.74
r180 9 26 18.8402 $w=1.65e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.185 $Y=1.6
+ $X2=2.205 $Y2=1.525
r181 9 11 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=2.185 $Y=1.6
+ $X2=2.185 $Y2=2.38
r182 8 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.525
+ $X2=1.665 $Y2=1.525
r183 7 26 6.66866 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.095 $Y=1.525
+ $X2=2.205 $Y2=1.525
r184 7 8 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.095 $Y=1.525
+ $X2=1.83 $Y2=1.525
r185 2 29 600 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=2.12 $X2=1.355 $Y2=2.135
r186 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.26
+ $Y=0.37 $X2=1.4 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%A_27_424# 1 2 9 13 18 19 22 24 27 31 34 35
c86 34 0 1.20405e-19 $X=2.69 $Y=1.635
c87 22 0 2.0421e-19 $X=2.61 $Y=2.39
c88 13 0 1.81055e-19 $X=2.765 $Y=2.46
c89 9 0 1.71716e-19 $X=2.75 $Y=0.69
r90 35 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.635
+ $X2=2.69 $Y2=1.8
r91 35 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.635
+ $X2=2.69 $Y2=1.47
r92 34 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.635
+ $X2=2.69 $Y2=1.8
r93 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.635 $X2=2.69 $Y2=1.635
r94 29 31 4.96677 $w=5.88e-07 $l=2.45e-07 $layer=LI1_cond $X=0.385 $Y=0.835
+ $X2=0.63 $Y2=0.835
r95 26 27 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=2.33
+ $X2=0.715 $Y2=2.33
r96 24 26 9.1006 $w=4.58e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=2.33 $X2=0.63
+ $Y2=2.33
r97 22 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.61 $Y=2.39 $X2=2.61
+ $Y2=1.8
r98 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.525 $Y=2.475
+ $X2=2.61 $Y2=2.39
r99 19 27 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.525 $Y=2.475
+ $X2=0.715 $Y2=2.475
r100 18 26 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.63 $Y=2.1 $X2=0.63
+ $Y2=2.33
r101 17 31 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.63 $Y=1.13
+ $X2=0.63 $Y2=0.835
r102 17 18 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.63 $Y=1.13
+ $X2=0.63 $Y2=2.1
r103 13 40 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.765 $Y=2.46
+ $X2=2.765 $Y2=1.8
r104 9 39 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.75 $Y=0.69
+ $X2=2.75 $Y2=1.47
r105 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r106 1 29 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.24
+ $Y=0.56 $X2=0.385 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%A_363_74# 1 2 9 12 15 16 17 19 21 22 23 26
+ 27 36 40 42 46 49
c109 46 0 1.95222e-19 $X=3.23 $Y=1.285
c110 36 0 1.81055e-19 $X=2.085 $Y=2.12
c111 26 0 1.3812e-19 $X=3.88 $Y=2.215
c112 21 0 1.45332e-19 $X=3.11 $Y=1.97
c113 17 0 7.12951e-20 $X=2.17 $Y=1.195
r114 46 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.285
+ $X2=3.23 $Y2=1.12
r115 45 47 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=1.285
+ $X2=3.175 $Y2=1.45
r116 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.285 $X2=3.23 $Y2=1.285
r117 42 45 3.45733 $w=2.98e-07 $l=9e-08 $layer=LI1_cond $X=3.175 $Y=1.195
+ $X2=3.175 $Y2=1.285
r118 38 40 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.99 $Y=2.055
+ $X2=3.11 $Y2=2.055
r119 34 36 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=1.96 $Y=2.12
+ $X2=2.085 $Y2=2.12
r120 30 32 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.96 $Y=1.195
+ $X2=2.085 $Y2=1.195
r121 27 51 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.88 $Y=2.215
+ $X2=3.72 $Y2=2.215
r122 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.88
+ $Y=2.215 $X2=3.88 $Y2=2.215
r123 24 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.88 $Y=2.905
+ $X2=3.88 $Y2=2.215
r124 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.715 $Y=2.99
+ $X2=3.88 $Y2=2.905
r125 22 23 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.715 $Y=2.99
+ $X2=3.075 $Y2=2.99
r126 21 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=1.97
+ $X2=3.11 $Y2=2.055
r127 21 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.11 $Y=1.97
+ $X2=3.11 $Y2=1.45
r128 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=2.905
+ $X2=3.075 $Y2=2.99
r129 18 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.14
+ $X2=2.99 $Y2=2.055
r130 18 19 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.99 $Y=2.14
+ $X2=2.99 $Y2=2.905
r131 17 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=1.195
+ $X2=2.085 $Y2=1.195
r132 16 42 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.025 $Y=1.195
+ $X2=3.175 $Y2=1.195
r133 16 17 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.025 $Y=1.195
+ $X2=2.17 $Y2=1.195
r134 15 36 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.085 $Y=2.02
+ $X2=2.085 $Y2=2.12
r135 14 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.28
+ $X2=2.085 $Y2=1.195
r136 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.085 $Y=1.28
+ $X2=2.085 $Y2=2.02
r137 10 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=2.38
+ $X2=3.72 $Y2=2.215
r138 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.72 $Y=2.38
+ $X2=3.72 $Y2=2.75
r139 9 49 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.14 $Y=0.69
+ $X2=3.14 $Y2=1.12
r140 2 34 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=1.96 $X2=1.96 $Y2=2.12
r141 1 30 182 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.37 $X2=1.96 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%A_817_48# 1 2 7 9 10 12 15 18 21 25 27 34 40
+ 42 46 47 49 51 52 57
c116 40 0 1.72297e-19 $X=5.41 $Y=2.465
c117 25 0 6.93786e-20 $X=4.38 $Y=0.94
c118 15 0 1.44303e-19 $X=4.38 $Y=2.05
r119 53 54 5.11481 $w=4.78e-07 $l=1.58e-07 $layer=LI1_cond $X=5.335 $Y=2.222
+ $X2=5.335 $Y2=2.38
r120 51 53 2.66626 $w=4.78e-07 $l=1.07e-07 $layer=LI1_cond $X=5.335 $Y=2.115
+ $X2=5.335 $Y2=2.222
r121 51 52 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.115
+ $X2=5.335 $Y2=1.95
r122 47 58 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.385
+ $X2=6.14 $Y2=1.55
r123 47 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.385
+ $X2=6.14 $Y2=1.22
r124 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.14
+ $Y=1.385 $X2=6.14 $Y2=1.385
r125 44 46 7.38284 $w=3.18e-07 $l=2.05e-07 $layer=LI1_cond $X=6.135 $Y=1.18
+ $X2=6.135 $Y2=1.385
r126 43 49 2.76166 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=5.265 $Y=1.095
+ $X2=5.017 $Y2=1.095
r127 42 44 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=5.975 $Y=1.095
+ $X2=6.135 $Y2=1.18
r128 42 43 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.975 $Y=1.095
+ $X2=5.265 $Y2=1.095
r129 40 54 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=2.465
+ $X2=5.41 $Y2=2.38
r130 36 49 3.70735 $w=2.5e-07 $l=2.01057e-07 $layer=LI1_cond $X=5.18 $Y=1.18
+ $X2=5.017 $Y2=1.095
r131 36 52 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.18 $Y=1.18
+ $X2=5.18 $Y2=1.95
r132 32 49 3.70735 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=4.935 $Y=1.01
+ $X2=5.017 $Y2=1.095
r133 32 34 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.935 $Y=1.01
+ $X2=4.935 $Y2=0.515
r134 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.47
+ $Y=2.215 $X2=4.47 $Y2=2.215
r135 27 53 3.21507 $w=3.15e-07 $l=2.4e-07 $layer=LI1_cond $X=5.095 $Y=2.222
+ $X2=5.335 $Y2=2.222
r136 27 29 22.8659 $w=3.13e-07 $l=6.25e-07 $layer=LI1_cond $X=5.095 $Y=2.222
+ $X2=4.47 $Y2=2.222
r137 23 25 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.16 $Y=0.94
+ $X2=4.38 $Y2=0.94
r138 21 58 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.215 $Y=2.4
+ $X2=6.215 $Y2=1.55
r139 18 57 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.05 $Y=0.74
+ $X2=6.05 $Y2=1.22
r140 15 30 38.6704 $w=3.39e-07 $l=2.0106e-07 $layer=POLY_cond $X=4.38 $Y=2.05
+ $X2=4.46 $Y2=2.215
r141 14 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.38 $Y=1.015
+ $X2=4.38 $Y2=0.94
r142 14 15 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=4.38 $Y=1.015
+ $X2=4.38 $Y2=2.05
r143 10 30 34.0041 $w=3.39e-07 $l=2.03101e-07 $layer=POLY_cond $X=4.375 $Y=2.38
+ $X2=4.46 $Y2=2.215
r144 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.375 $Y=2.38
+ $X2=4.375 $Y2=2.75
r145 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.16 $Y=0.865
+ $X2=4.16 $Y2=0.94
r146 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.16 $Y=0.865 $X2=4.16
+ $Y2=0.58
r147 2 51 600 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=5.225
+ $Y=1.96 $X2=5.41 $Y2=2.115
r148 2 40 300 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=2 $X=5.225
+ $Y=1.96 $X2=5.41 $Y2=2.465
r149 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.79
+ $Y=0.37 $X2=4.935 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%A_643_74# 1 2 9 13 15 16 20 21 22 26 29 30
+ 36
c81 30 0 4.70657e-20 $X=3.39 $Y=2.405
c82 26 0 1.71716e-19 $X=3.58 $Y=0.76
c83 22 0 1.95222e-19 $X=3.665 $Y=1.81
c84 20 0 1.44303e-19 $X=3.58 $Y=1.725
c85 9 0 1.72297e-19 $X=5.135 $Y=2.46
r86 36 39 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=4.795 $Y=1.635
+ $X2=4.795 $Y2=1.81
r87 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.83
+ $Y=1.635 $X2=4.83 $Y2=1.635
r88 32 34 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.45 $Y=1.81
+ $X2=3.58 $Y2=1.81
r89 29 30 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=2.57
+ $X2=3.39 $Y2=2.405
r90 24 26 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0.76
+ $X2=3.58 $Y2=0.76
r91 22 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=1.81
+ $X2=3.58 $Y2=1.81
r92 21 39 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.665 $Y=1.81
+ $X2=4.795 $Y2=1.81
r93 21 22 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.665 $Y=1.81
+ $X2=3.665 $Y2=1.81
r94 20 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=1.725
+ $X2=3.58 $Y2=1.81
r95 19 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=0.925
+ $X2=3.58 $Y2=0.76
r96 19 20 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.58 $Y=0.925 $X2=3.58
+ $Y2=1.725
r97 17 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=1.895
+ $X2=3.45 $Y2=1.81
r98 17 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.45 $Y=1.895
+ $X2=3.45 $Y2=2.405
r99 15 37 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.045 $Y=1.635
+ $X2=4.83 $Y2=1.635
r100 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.045 $Y=1.635
+ $X2=5.135 $Y2=1.635
r101 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.15 $Y=1.47
+ $X2=5.135 $Y2=1.635
r102 11 13 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.15 $Y=1.47
+ $X2=5.15 $Y2=0.74
r103 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.135 $Y=1.8
+ $X2=5.135 $Y2=1.635
r104 7 9 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.135 $Y=1.8
+ $X2=5.135 $Y2=2.46
r105 2 29 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.96 $X2=3.41 $Y2=2.57
r106 1 24 182 $w=1.7e-07 $l=4.79687e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.37 $X2=3.415 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%RESET_B 3 7 9 12 13
c41 12 0 1.10707e-19 $X=5.6 $Y=1.515
c42 3 0 1.77844e-19 $X=5.54 $Y=0.74
r43 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.6 $Y=1.515
+ $X2=5.6 $Y2=1.68
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.6 $Y=1.515
+ $X2=5.6 $Y2=1.35
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=1.515 $X2=5.6 $Y2=1.515
r46 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.6 $Y=1.665 $X2=5.6
+ $Y2=1.515
r47 7 15 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=5.635 $Y=2.46
+ $X2=5.635 $Y2=1.68
r48 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.54 $Y=0.74 $X2=5.54
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%VPWR 1 2 3 4 15 19 23 28 29 30 32 37 45 55
+ 56 59 62 65
c76 23 0 1.10707e-19 $X=5.91 $Y=2.115
r77 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 65 68 9.62469 $w=6.38e-07 $l=5.15e-07 $layer=LI1_cond $X=4.755 $Y=2.815
+ $X2=4.755 $Y2=3.33
r79 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r82 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r83 53 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 50 68 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=5.075 $Y=3.33
+ $X2=4.755 $Y2=3.33
r86 50 52 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.075 $Y=3.33
+ $X2=5.52 $Y2=3.33
r87 49 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 46 62 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.517 $Y2=3.33
r90 46 48 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 45 68 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.755 $Y2=3.33
r92 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 44 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 41 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r98 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r99 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r100 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r101 37 62 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.517 $Y2=3.33
r102 37 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 35 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 32 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r106 32 34 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r107 30 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 30 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 28 52 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.745 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=3.33
+ $X2=5.91 $Y2=3.33
r111 27 55 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.075 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=3.33
+ $X2=5.91 $Y2=3.33
r113 23 26 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.91 $Y=2.115
+ $X2=5.91 $Y2=2.815
r114 21 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=3.245
+ $X2=5.91 $Y2=3.33
r115 21 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.91 $Y=3.245
+ $X2=5.91 $Y2=2.815
r116 17 62 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.517 $Y=3.245
+ $X2=2.517 $Y2=3.33
r117 17 19 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=2.517 $Y=3.245
+ $X2=2.517 $Y2=2.815
r118 13 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r119 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.815
r120 4 26 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=5.725
+ $Y=1.96 $X2=5.91 $Y2=2.815
r121 4 23 400 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=5.725
+ $Y=1.96 $X2=5.91 $Y2=2.115
r122 3 65 600 $w=1.7e-07 $l=4.04784e-07 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=2.54 $X2=4.755 $Y2=2.815
r123 2 19 600 $w=1.7e-07 $l=9.67587e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.96 $X2=2.515 $Y2=2.815
r124 1 15 600 $w=1.7e-07 $l=7.82049e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.12 $X2=0.78 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%Q 1 2 9 14 15 16
c23 16 0 1.77844e-19 $X=6.48 $Y=0.555
r24 22 23 9.7361 $w=5.33e-07 $l=1.65e-07 $layer=LI1_cond $X=6.367 $Y=0.675
+ $X2=6.367 $Y2=0.84
r25 16 22 2.68279 $w=5.33e-07 $l=1.2e-07 $layer=LI1_cond $X=6.367 $Y=0.555
+ $X2=6.367 $Y2=0.675
r26 15 23 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.55 $Y=1.82
+ $X2=6.55 $Y2=0.84
r27 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=1.985
+ $X2=6.455 $Y2=1.82
r28 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=6.455 $Y=2 $X2=6.455
+ $Y2=1.985
r29 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=6.455 $Y=2 $X2=6.455
+ $Y2=2.815
r30 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.84 $X2=6.44 $Y2=1.985
r31 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.84 $X2=6.44 $Y2=2.815
r32 1 22 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.125
+ $Y=0.37 $X2=6.265 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTP_1%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 44 62 63 66
r74 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r75 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r76 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r77 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r78 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r79 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r80 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r81 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r82 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r83 51 66 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.487
+ $Y2=0
r84 51 53 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.68 $Y=0 $X2=4.08
+ $Y2=0
r85 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r87 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r88 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r89 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r90 44 66 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.487
+ $Y2=0
r91 44 49 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.16
+ $Y2=0
r92 42 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r93 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 38 54 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r95 38 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.64
+ $Y2=0
r96 36 59 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.52
+ $Y2=0
r97 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.755
+ $Y2=0
r98 35 62 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=6.48
+ $Y2=0
r99 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=5.755
+ $Y2=0
r100 33 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.08
+ $Y2=0
r101 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.375
+ $Y2=0
r102 32 56 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.56
+ $Y2=0
r103 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.375
+ $Y2=0
r104 30 41 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0
+ $X2=0.72 $Y2=0
r105 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.97
+ $Y2=0
r106 29 46 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.2
+ $Y2=0
r107 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.97
+ $Y2=0
r108 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0
r109 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0.675
r110 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=0.085
+ $X2=4.375 $Y2=0
r111 21 23 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.375 $Y=0.085
+ $X2=4.375 $Y2=0.58
r112 17 66 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.487 $Y=0.085
+ $X2=2.487 $Y2=0
r113 17 19 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=2.487 $Y=0.085
+ $X2=2.487 $Y2=0.515
r114 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0
r115 13 15 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0.515
r116 4 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=5.615
+ $Y=0.37 $X2=5.755 $Y2=0.675
r117 3 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.235
+ $Y=0.37 $X2=4.375 $Y2=0.58
r118 2 19 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.37 $X2=2.485 $Y2=0.515
r119 1 15 91 $w=1.7e-07 $l=3.16702e-07 $layer=licon1_NDIFF $count=2 $X=0.675
+ $Y=0.56 $X2=0.97 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__nor3b_1.pxi.spice
* Created: Fri Aug 28 17:48:36 2020
* 
x_PM_SKY130_FD_SC_MS__NOR3B_1%C_N N_C_N_M1006_g N_C_N_M1004_g C_N N_C_N_c_53_n
+ N_C_N_c_54_n PM_SKY130_FD_SC_MS__NOR3B_1%C_N
x_PM_SKY130_FD_SC_MS__NOR3B_1%A N_A_M1003_g N_A_M1007_g A N_A_c_85_n N_A_c_86_n
+ PM_SKY130_FD_SC_MS__NOR3B_1%A
x_PM_SKY130_FD_SC_MS__NOR3B_1%B N_B_M1002_g N_B_M1005_g B N_B_c_120_n
+ N_B_c_121_n PM_SKY130_FD_SC_MS__NOR3B_1%B
x_PM_SKY130_FD_SC_MS__NOR3B_1%A_27_112# N_A_27_112#_M1004_s N_A_27_112#_M1006_s
+ N_A_27_112#_M1001_g N_A_27_112#_M1000_g N_A_27_112#_c_168_n
+ N_A_27_112#_c_191_n N_A_27_112#_c_158_n N_A_27_112#_c_163_n
+ N_A_27_112#_c_159_n N_A_27_112#_c_165_n N_A_27_112#_c_160_n
+ N_A_27_112#_c_161_n PM_SKY130_FD_SC_MS__NOR3B_1%A_27_112#
x_PM_SKY130_FD_SC_MS__NOR3B_1%VPWR N_VPWR_M1006_d N_VPWR_c_229_n N_VPWR_c_230_n
+ N_VPWR_c_231_n VPWR N_VPWR_c_232_n N_VPWR_c_228_n
+ PM_SKY130_FD_SC_MS__NOR3B_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR3B_1%Y N_Y_M1007_d N_Y_M1000_d N_Y_M1001_d N_Y_c_254_n
+ N_Y_c_255_n N_Y_c_256_n N_Y_c_260_n N_Y_c_257_n Y Y N_Y_c_258_n N_Y_c_259_n
+ PM_SKY130_FD_SC_MS__NOR3B_1%Y
x_PM_SKY130_FD_SC_MS__NOR3B_1%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_c_302_n
+ N_VGND_c_303_n N_VGND_c_304_n N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n
+ VGND N_VGND_c_308_n N_VGND_c_309_n PM_SKY130_FD_SC_MS__NOR3B_1%VGND
cc_1 VNB N_C_N_M1006_g 0.00667774f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.26
cc_2 VNB C_N 0.0104207f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_C_N_c_53_n 0.0343932f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_4 VNB N_C_N_c_54_n 0.0224251f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_5 VNB N_A_M1007_g 0.0268153f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_6 VNB N_A_c_85_n 0.0267839f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_7 VNB N_A_c_86_n 0.0023516f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_8 VNB N_B_M1005_g 0.026332f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_9 VNB N_B_c_120_n 0.0270072f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_10 VNB N_B_c_121_n 0.00165701f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_11 VNB N_A_27_112#_M1000_g 0.0321102f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_12 VNB N_A_27_112#_c_158_n 0.0138636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_112#_c_159_n 0.0299402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_112#_c_160_n 0.00165828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_112#_c_161_n 0.0289662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_228_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_254_n 0.00280874f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_18 VNB N_Y_c_255_n 0.00951425f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.55
cc_19 VNB N_Y_c_256_n 0.0107024f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_20 VNB N_Y_c_257_n 0.0227107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_258_n 0.0332097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_259_n 0.0157047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_302_n 0.0162763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_303_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_25 VNB N_VGND_c_304_n 0.0263417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_305_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_27 VNB N_VGND_c_306_n 0.0186436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_307_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_308_n 0.0214382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_309_n 0.188982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_C_N_M1006_g 0.0288699f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_32 VPB N_A_M1003_g 0.0233129f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_33 VPB N_A_c_85_n 0.00567706f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_34 VPB N_A_c_86_n 0.00248627f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.22
cc_35 VPB N_B_M1002_g 0.022787f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_36 VPB N_B_c_120_n 0.00567158f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_37 VPB N_B_c_121_n 0.00209172f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.22
cc_38 VPB N_A_27_112#_M1001_g 0.027993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_112#_c_163_n 0.0216239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_112#_c_159_n 0.00810758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_112#_c_165_n 0.032593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_112#_c_160_n 0.00241918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_27_112#_c_161_n 0.00579797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_229_n 0.0169528f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.835
cc_45 VPB N_VPWR_c_230_n 0.0265205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_231_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_47 VPB N_VPWR_c_232_n 0.0525134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_228_n 0.0850314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_Y_c_260_n 0.038413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_Y_c_257_n 0.0307877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 N_C_N_M1006_g N_A_M1003_g 0.0244596f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_52 C_N N_A_M1007_g 0.00343954f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_53 N_C_N_c_54_n N_A_M1007_g 0.014565f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_54 N_C_N_M1006_g N_A_c_85_n 0.00732394f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_55 C_N N_A_c_85_n 0.00113494f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_C_N_c_53_n N_A_c_85_n 0.0125126f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_57 N_C_N_M1006_g N_A_c_86_n 0.00313503f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_58 C_N N_A_c_86_n 0.0159708f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_59 N_C_N_c_53_n N_A_c_86_n 2.28995e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_60 N_C_N_M1006_g N_A_27_112#_c_168_n 0.0153541f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_61 C_N N_A_27_112#_c_168_n 0.00719058f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 C_N N_A_27_112#_c_158_n 0.014413f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_C_N_c_53_n N_A_27_112#_c_158_n 0.00105729f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_64 N_C_N_c_54_n N_A_27_112#_c_158_n 0.00429074f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_65 N_C_N_M1006_g N_A_27_112#_c_163_n 0.00477439f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_66 C_N N_A_27_112#_c_163_n 0.00883508f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_C_N_c_53_n N_A_27_112#_c_163_n 0.00264359f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_68 N_C_N_M1006_g N_A_27_112#_c_159_n 0.0082703f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_69 C_N N_A_27_112#_c_159_n 0.0282012f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_C_N_c_53_n N_A_27_112#_c_159_n 0.00231928f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_71 N_C_N_c_54_n N_A_27_112#_c_159_n 0.00459385f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_72 N_C_N_M1006_g N_A_27_112#_c_165_n 0.0134806f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_73 N_C_N_M1006_g N_VPWR_c_229_n 0.00693742f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_74 N_C_N_M1006_g N_VPWR_c_230_n 0.00465228f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_75 N_C_N_M1006_g N_VPWR_c_228_n 0.00555093f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_76 N_C_N_c_54_n N_VGND_c_302_n 0.00619988f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_77 N_C_N_c_54_n N_VGND_c_304_n 0.00434489f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_78 N_C_N_c_54_n N_VGND_c_309_n 0.00487769f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_B_M1002_g 0.0478249f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_M1007_g N_B_M1005_g 0.0165331f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_c_85_n N_B_c_120_n 0.0478249f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A_c_86_n N_B_c_120_n 0.00154051f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A_c_85_n N_B_c_121_n 0.00154051f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A_c_86_n N_B_c_121_n 0.0244404f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_A_27_112#_c_168_n 0.0165696f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_c_85_n N_A_27_112#_c_168_n 7.08634e-19 $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A_c_86_n N_A_27_112#_c_168_n 0.0229716f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_A_27_112#_c_163_n 0.00136424f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VPWR_c_229_n 0.0185439f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_M1003_g N_VPWR_c_232_n 0.00460063f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VPWR_c_228_n 0.00908371f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_Y_c_254_n 4.78065e-19 $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_M1007_g N_Y_c_256_n 0.00233828f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_M1007_g N_VGND_c_302_n 0.00395387f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_c_85_n N_VGND_c_302_n 0.00104145f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_c_86_n N_VGND_c_302_n 0.00718896f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A_M1007_g N_VGND_c_306_n 0.00461464f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A_M1007_g N_VGND_c_309_n 0.00912669f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B_M1002_g N_A_27_112#_M1001_g 0.0469965f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_100 N_B_c_121_n N_A_27_112#_M1001_g 7.09387e-19 $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B_M1005_g N_A_27_112#_M1000_g 0.0260254f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B_M1002_g N_A_27_112#_c_168_n 0.0174565f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_103 N_B_c_120_n N_A_27_112#_c_168_n 7.05107e-19 $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B_c_121_n N_A_27_112#_c_168_n 0.0229716f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B_M1002_g N_A_27_112#_c_191_n 0.00111344f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_106 N_B_c_120_n N_A_27_112#_c_160_n 0.00121489f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B_c_121_n N_A_27_112#_c_160_n 0.0246187f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B_c_120_n N_A_27_112#_c_161_n 0.017083f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_109 N_B_c_121_n N_A_27_112#_c_161_n 0.00121489f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_110 N_B_M1002_g N_VPWR_c_229_n 0.00385865f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_111 N_B_M1002_g N_VPWR_c_232_n 0.00553757f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_112 N_B_M1002_g N_VPWR_c_228_n 0.0109071f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_113 N_B_M1005_g N_Y_c_254_n 0.00963749f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B_M1005_g N_Y_c_255_n 0.0117933f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B_c_120_n N_Y_c_255_n 6.97898e-19 $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_116 N_B_c_121_n N_Y_c_255_n 0.0167639f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_117 N_B_M1005_g N_Y_c_256_n 0.00153788f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B_c_120_n N_Y_c_256_n 6.17801e-19 $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B_c_121_n N_Y_c_256_n 0.00886294f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_120 N_B_M1002_g N_Y_c_260_n 0.00311738f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_121 N_B_M1005_g N_Y_c_258_n 6.27049e-19 $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_122 N_B_M1005_g N_VGND_c_303_n 0.00484409f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B_M1005_g N_VGND_c_306_n 0.00434272f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_124 N_B_M1005_g N_VGND_c_309_n 0.0082177f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_27_112#_c_168_n N_VPWR_M1006_d 0.0116797f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_27_112#_c_168_n N_VPWR_c_229_n 0.0218557f $X=2.125 $Y=2.035 $X2=0
+ $Y2=0
cc_127 N_A_27_112#_c_165_n N_VPWR_c_229_n 0.0251858f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_128 N_A_27_112#_c_165_n N_VPWR_c_230_n 0.00991858f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_129 N_A_27_112#_M1001_g N_VPWR_c_232_n 0.005209f $X=2.215 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A_27_112#_M1001_g N_VPWR_c_228_n 0.00988686f $X=2.215 $Y=2.4 $X2=0
+ $Y2=0
cc_131 N_A_27_112#_c_165_n N_VPWR_c_228_n 0.0148286f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_27_112#_c_168_n A_263_368# 0.0096152f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_27_112#_c_168_n A_347_368# 0.0186283f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_27_112#_M1000_g N_Y_c_254_n 6.28869e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_27_112#_M1000_g N_Y_c_255_n 0.0117933f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_27_112#_c_160_n N_Y_c_255_n 0.0156476f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A_27_112#_c_161_n N_Y_c_255_n 5.49471e-19 $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_27_112#_M1001_g N_Y_c_260_n 0.0163551f $X=2.215 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_27_112#_c_168_n N_Y_c_260_n 0.00161016f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_140 N_A_27_112#_c_160_n N_Y_c_260_n 0.00379786f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_27_112#_c_161_n N_Y_c_260_n 6.79589e-19 $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_27_112#_M1001_g N_Y_c_257_n 0.0114868f $X=2.215 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_27_112#_M1000_g N_Y_c_257_n 0.00367585f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_27_112#_c_168_n N_Y_c_257_n 0.00824932f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_145 N_A_27_112#_c_191_n N_Y_c_257_n 0.0117569f $X=2.21 $Y=1.95 $X2=0 $Y2=0
cc_146 N_A_27_112#_c_160_n N_Y_c_257_n 0.0248017f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A_27_112#_c_161_n N_Y_c_257_n 0.00739878f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_27_112#_M1000_g N_Y_c_258_n 0.0104715f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_27_112#_M1000_g N_Y_c_259_n 0.002266f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_27_112#_c_160_n N_Y_c_259_n 0.0103958f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A_27_112#_c_161_n N_Y_c_259_n 7.83559e-19 $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A_27_112#_M1000_g N_VGND_c_303_n 0.00622602f $X=2.28 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_27_112#_c_158_n N_VGND_c_304_n 0.00858362f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_154 N_A_27_112#_M1000_g N_VGND_c_308_n 0.00434272f $X=2.28 $Y=0.74 $X2=0
+ $Y2=0
cc_155 N_A_27_112#_M1000_g N_VGND_c_309_n 0.00825279f $X=2.28 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_27_112#_c_158_n N_VGND_c_309_n 0.0154187f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_157 N_VPWR_c_232_n N_Y_c_260_n 0.0230434f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_158 N_VPWR_c_228_n N_Y_c_260_n 0.018998f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_159 N_Y_c_255_n N_VGND_M1005_d 0.00358162f $X=2.33 $Y=1.095 $X2=0 $Y2=0
cc_160 N_Y_c_254_n N_VGND_c_302_n 0.00158095f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_161 N_Y_c_254_n N_VGND_c_303_n 0.0191765f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_162 N_Y_c_255_n N_VGND_c_303_n 0.0248957f $X=2.33 $Y=1.095 $X2=0 $Y2=0
cc_163 N_Y_c_258_n N_VGND_c_303_n 0.0201667f $X=2.495 $Y=0.515 $X2=0 $Y2=0
cc_164 N_Y_c_254_n N_VGND_c_306_n 0.0145639f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_165 N_Y_c_258_n N_VGND_c_308_n 0.0205877f $X=2.495 $Y=0.515 $X2=0 $Y2=0
cc_166 N_Y_c_254_n N_VGND_c_309_n 0.0119984f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_167 N_Y_c_258_n N_VGND_c_309_n 0.0169844f $X=2.495 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o31ai_2.pex.spice
* Created: Wed Sep  2 12:25:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O31AI_2%A1 3 7 11 13 15 16 17 18 27
r49 25 27 53.0059 $w=3.41e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.432
+ $X2=0.96 $Y2=1.432
r50 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r51 23 25 10.6012 $w=3.41e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.432
+ $X2=0.585 $Y2=1.432
r52 17 18 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r53 17 26 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r54 16 26 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r55 13 27 14.8416 $w=3.41e-07 $l=2.94863e-07 $layer=POLY_cond $X=1.065 $Y=1.185
+ $X2=0.96 $Y2=1.432
r56 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.065 $Y=1.185
+ $X2=1.065 $Y2=0.74
r57 9 27 17.6972 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=1.432
r58 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.96 $Y=1.68 $X2=0.96
+ $Y2=2.4
r59 5 23 17.6972 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=0.51 $Y=1.68
+ $X2=0.51 $Y2=1.432
r60 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.51 $Y=1.68 $X2=0.51
+ $Y2=2.4
r61 1 23 2.12023 $w=3.41e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.432
+ $X2=0.51 $Y2=1.432
r62 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%A2 1 3 6 8 10 13 15 16 24
c55 24 0 1.15611e-19 $X=1.86 $Y=1.537
c56 13 0 3.67831e-20 $X=2.065 $Y=0.74
r57 22 24 21.2407 $w=2.95e-07 $l=1.3e-07 $layer=POLY_cond $X=1.73 $Y=1.537
+ $X2=1.86 $Y2=1.537
r58 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.515 $X2=1.73 $Y2=1.515
r59 20 22 38.3966 $w=2.95e-07 $l=2.35e-07 $layer=POLY_cond $X=1.495 $Y=1.537
+ $X2=1.73 $Y2=1.537
r60 16 23 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.73 $Y2=1.565
r61 15 23 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.73
+ $Y2=1.565
r62 11 24 33.4949 $w=2.95e-07 $l=2.83478e-07 $layer=POLY_cond $X=2.065 $Y=1.35
+ $X2=1.86 $Y2=1.537
r63 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.065 $Y=1.35
+ $X2=2.065 $Y2=0.74
r64 8 24 14.3312 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=1.86 $Y=1.725
+ $X2=1.86 $Y2=1.537
r65 8 10 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.86 $Y=1.725
+ $X2=1.86 $Y2=2.4
r66 4 20 18.5736 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.537
r67 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r68 1 20 13.8881 $w=2.95e-07 $l=2.26548e-07 $layer=POLY_cond $X=1.41 $Y=1.725
+ $X2=1.495 $Y2=1.537
r69 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.41 $Y=1.725 $X2=1.41
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%A3 3 6 9 13 17 19 22 25 27
c63 13 0 2.42806e-19 $X=3.345 $Y=2.4
r64 26 27 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.345 $Y=1.515
+ $X2=3.37 $Y2=1.515
r65 24 26 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.28 $Y=1.515
+ $X2=3.345 $Y2=1.515
r66 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.28
+ $Y=1.515 $X2=3.28 $Y2=1.515
r67 21 24 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=2.895 $Y=1.515
+ $X2=3.28 $Y2=1.515
r68 21 22 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.895 $Y=1.515
+ $X2=2.805 $Y2=1.515
r69 19 25 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.28 $Y2=1.565
r70 15 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=1.35
+ $X2=3.37 $Y2=1.515
r71 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.37 $Y=1.35
+ $X2=3.37 $Y2=0.74
r72 11 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.68
+ $X2=3.345 $Y2=1.515
r73 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.345 $Y=1.68
+ $X2=3.345 $Y2=2.4
r74 7 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=1.68
+ $X2=2.895 $Y2=1.515
r75 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.895 $Y=1.68
+ $X2=2.895 $Y2=2.4
r76 6 22 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.57 $Y=1.425
+ $X2=2.805 $Y2=1.425
r77 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.495 $Y=1.35
+ $X2=2.57 $Y2=1.425
r78 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.495 $Y=1.35
+ $X2=2.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%B1 3 7 11 15 17 22 28
c55 17 0 1.34959e-19 $X=4.365 $Y=1.515
r56 31 36 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=4.53 $Y=1.465 $X2=4.53
+ $Y2=1.515
r57 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.465 $X2=4.53 $Y2=1.465
r58 28 30 31.1181 $w=3.64e-07 $l=2.35e-07 $layer=POLY_cond $X=4.295 $Y=1.49
+ $X2=4.53 $Y2=1.49
r59 27 28 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=4.28 $Y=1.49
+ $X2=4.295 $Y2=1.49
r60 24 25 5.95879 $w=3.64e-07 $l=4.5e-08 $layer=POLY_cond $X=3.8 $Y=1.49
+ $X2=3.845 $Y2=1.49
r61 22 31 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.53 $Y=1.295
+ $X2=4.53 $Y2=1.465
r62 20 27 11.9176 $w=3.64e-07 $l=9e-08 $layer=POLY_cond $X=4.19 $Y=1.49 $X2=4.28
+ $Y2=1.49
r63 20 25 45.6841 $w=3.64e-07 $l=3.45e-07 $layer=POLY_cond $X=4.19 $Y=1.49
+ $X2=3.845 $Y2=1.49
r64 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.19
+ $Y=1.515 $X2=4.19 $Y2=1.515
r65 17 36 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=1.515
+ $X2=4.53 $Y2=1.515
r66 17 19 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.365 $Y=1.515
+ $X2=4.19 $Y2=1.515
r67 13 28 19.2285 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=4.295 $Y=1.68
+ $X2=4.295 $Y2=1.49
r68 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.295 $Y=1.68
+ $X2=4.295 $Y2=2.4
r69 9 27 23.572 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.28 $Y=1.3 $X2=4.28
+ $Y2=1.49
r70 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.28 $Y=1.3 $X2=4.28
+ $Y2=0.74
r71 5 25 19.2285 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=3.845 $Y=1.68
+ $X2=3.845 $Y2=1.49
r72 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.845 $Y=1.68
+ $X2=3.845 $Y2=2.4
r73 1 24 23.572 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=1.49
r74 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%A_28_368# 1 2 3 10 12 14 18 20 27 29
r40 21 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=2.035
+ $X2=1.185 $Y2=2.035
r41 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=2.085 $Y2=2.035
r42 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.35 $Y2=2.035
r43 16 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r44 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r45 15 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.37 $Y=2.035
+ $X2=0.245 $Y2=2.035
r46 14 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.185 $Y2=2.035
r47 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.37 $Y2=2.035
r48 10 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.035
r49 10 12 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.815
r50 3 29 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=1.95
+ $Y=1.84 $X2=2.085 $Y2=2.115
r51 2 27 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.115
r52 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.815
r53 1 25 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r54 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r52 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 27 30 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 25 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.695 $Y2=3.33
r57 25 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.695 $Y2=3.33
r61 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r63 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 16 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r65 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.07 $Y2=3.33
r66 15 33 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.56 $Y2=3.33
r67 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.07 $Y2=3.33
r68 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=3.33
r69 11 13 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=2.355
r70 7 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r71 7 9 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.455
r72 2 13 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.935
+ $Y=1.84 $X2=4.07 $Y2=2.355
r73 1 9 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%A_300_368# 1 2 9 11 12 15
r23 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.12 $Y=2.905
+ $X2=3.12 $Y2=2.455
r24 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=3.12 $Y2=2.905
r25 11 12 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=1.72 $Y2=2.99
r26 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.635 $Y=2.905
+ $X2=1.72 $Y2=2.99
r27 7 9 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.635 $Y=2.905
+ $X2=1.635 $Y2=2.455
r28 2 15 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.84 $X2=3.12 $Y2=2.455
r29 1 9 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%Y 1 2 3 4 15 19 20 21 23 27 29 31 34 35 40
+ 43 44
c75 43 0 1.71942e-19 $X=3.6 $Y=2.405
c76 35 0 1.15611e-19 $X=2.67 $Y=1.82
c77 34 0 7.08642e-20 $X=2.67 $Y=1.985
r78 43 44 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.62 $Y=2.405
+ $X2=3.62 $Y2=2.775
r79 38 43 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.62 $Y=2.12
+ $X2=3.62 $Y2=2.405
r80 38 40 0.89609 $w=3.3e-07 $l=2.38642e-07 $layer=LI1_cond $X=3.62 $Y=2.12
+ $X2=3.455 $Y2=1.95
r81 36 37 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.035
+ $X2=2.67 $Y2=2.12
r82 34 36 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.67 $Y=1.985 $X2=2.67
+ $Y2=2.035
r83 34 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=1.985
+ $X2=2.67 $Y2=1.82
r84 29 42 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.52 $Y=2.02 $X2=4.52
+ $Y2=1.935
r85 29 31 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=4.52 $Y=2.02
+ $X2=4.52 $Y2=2.815
r86 25 27 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.015 $Y=1.01
+ $X2=4.015 $Y2=0.775
r87 24 40 8.61065 $w=1.7e-07 $l=3.37417e-07 $layer=LI1_cond $X=3.785 $Y=1.935
+ $X2=3.455 $Y2=1.95
r88 23 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.935
+ $X2=4.52 $Y2=1.935
r89 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.355 $Y=1.935
+ $X2=3.785 $Y2=1.935
r90 22 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=2.035
+ $X2=2.67 $Y2=2.035
r91 21 40 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=2.035
+ $X2=3.455 $Y2=1.95
r92 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.455 $Y=2.035
+ $X2=2.835 $Y2=2.035
r93 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.85 $Y=1.095
+ $X2=4.015 $Y2=1.01
r94 19 20 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=3.85 $Y=1.095
+ $X2=2.835 $Y2=1.095
r95 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.75 $Y=1.18
+ $X2=2.835 $Y2=1.095
r96 17 35 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.75 $Y=1.18 $X2=2.75
+ $Y2=1.82
r97 15 37 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.63 $Y=2.57 $X2=2.63
+ $Y2=2.12
r98 4 42 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.015
r99 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.815
r100 3 44 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.84 $X2=3.62 $Y2=2.815
r101 3 40 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.84 $X2=3.62 $Y2=2.115
r102 2 34 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.84 $X2=2.67 $Y2=1.985
r103 2 15 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.84 $X2=2.67 $Y2=2.57
r104 1 27 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.37 $X2=4.015 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%A_27_74# 1 2 3 4 5 18 20 21 24 26 29 30 35
+ 36 37 40 42 44
c81 30 0 3.67831e-20 $X=3.42 $Y=0.755
r82 44 46 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.28 $Y=0.515
+ $X2=2.28 $Y2=0.755
r83 38 40 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.515 $Y=0.425
+ $X2=4.515 $Y2=0.515
r84 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=4.515 $Y2=0.425
r85 36 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=3.67 $Y2=0.34
r86 33 35 3.45733 $w=2.48e-07 $l=7.5e-08 $layer=LI1_cond $X=3.545 $Y=0.67
+ $X2=3.545 $Y2=0.595
r87 32 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.545 $Y=0.425
+ $X2=3.67 $Y2=0.34
r88 32 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.545 $Y=0.425
+ $X2=3.545 $Y2=0.595
r89 31 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0.755
+ $X2=2.28 $Y2=0.755
r90 30 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.42 $Y=0.755
+ $X2=3.545 $Y2=0.67
r91 30 31 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=3.42 $Y=0.755
+ $X2=2.445 $Y2=0.755
r92 28 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.84
+ $X2=2.28 $Y2=0.755
r93 28 29 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.28 $Y=0.84
+ $X2=2.28 $Y2=1.01
r94 27 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.095
+ $X2=1.28 $Y2=1.095
r95 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=1.095
+ $X2=2.28 $Y2=1.01
r96 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=1.095
+ $X2=1.445 $Y2=1.095
r97 22 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.01 $X2=1.28
+ $Y2=1.095
r98 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.515
r99 20 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.28 $Y2=1.095
r100 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.445 $Y2=1.095
r101 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r102 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r103 5 40 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.37 $X2=4.515 $Y2=0.515
r104 4 35 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.37 $X2=3.585 $Y2=0.595
r105 3 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.14
+ $Y=0.37 $X2=2.28 $Y2=0.515
r106 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r107 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_2%VGND 1 2 3 12 14 18 22 24 34 35 38 41 46 52
r59 50 52 9.13833 $w=5.83e-07 $l=1.2e-07 $layer=LI1_cond $X=3.12 $Y=0.207
+ $X2=3.24 $Y2=0.207
r60 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 48 50 3.8847 $w=5.83e-07 $l=1.9e-07 $layer=LI1_cond $X=2.93 $Y=0.207
+ $X2=3.12 $Y2=0.207
r62 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r63 44 48 5.92928 $w=5.83e-07 $l=2.9e-07 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=2.93 $Y2=0.207
r64 44 46 6.99152 $w=5.83e-07 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=2.625 $Y2=0.207
r65 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r68 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r70 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r71 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r72 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r73 31 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.24
+ $Y2=0
r74 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r75 27 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r76 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r78 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r79 22 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r80 22 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r81 21 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r82 21 46 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.625
+ $Y2=0
r83 16 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r84 16 18 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.66
r85 15 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r86 14 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r87 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=0.945
+ $Y2=0
r88 10 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r89 10 12 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.66
r90 3 48 182 $w=1.7e-07 $l=3.77094e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.37 $X2=2.93 $Y2=0.335
r91 2 18 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.66
r92 1 12 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.66
.ends


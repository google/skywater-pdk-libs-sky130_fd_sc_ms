* File: sky130_fd_sc_ms__o32ai_2.pex.spice
* Created: Fri Aug 28 18:04:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O32AI_2%B2 3 7 11 15 17 18 19 30
c45 30 0 1.94533e-19 $X=0.955 $Y=1.515
c46 19 0 6.22621e-20 $X=1.2 $Y=1.665
c47 15 0 1.87992e-19 $X=0.955 $Y=2.4
r48 29 30 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.515
+ $X2=0.955 $Y2=1.515
r49 27 29 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.835 $Y=1.515
+ $X2=0.925 $Y2=1.515
r50 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.835
+ $Y=1.515 $X2=0.835 $Y2=1.515
r51 25 27 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.835 $Y2=1.515
r52 23 25 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.505 $Y2=1.515
r53 19 28 9.78236 $w=4.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.835 $Y2=1.565
r54 18 28 3.08211 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.835 $Y2=1.565
r55 17 18 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r56 13 30 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.515
r57 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r58 9 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.515
r59 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
r60 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r61 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
r62 1 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.515
r63 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%B1 3 7 11 15 17 23 24
c54 11 0 6.22621e-20 $X=1.855 $Y=2.4
r55 24 25 10.7111 $w=3.15e-07 $l=7e-08 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.925 $Y2=1.515
r56 22 24 31.3683 $w=3.15e-07 $l=2.05e-07 $layer=POLY_cond $X=1.65 $Y=1.515
+ $X2=1.855 $Y2=1.515
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r58 20 22 34.4286 $w=3.15e-07 $l=2.25e-07 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.65 $Y2=1.515
r59 19 20 3.06032 $w=3.15e-07 $l=2e-08 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.425 $Y2=1.515
r60 17 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r61 13 25 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.515
r62 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.74
r63 9 24 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=1.515
r64 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=2.4
r65 5 20 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.515
r66 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r67 1 19 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=1.515
r68 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A3 3 7 11 15 17 18 26
c59 7 0 1.72955e-19 $X=2.865 $Y=2.4
r60 26 27 9.12303 $w=3.17e-07 $l=6e-08 $layer=POLY_cond $X=3.255 $Y=1.515
+ $X2=3.315 $Y2=1.515
r61 25 26 59.2997 $w=3.17e-07 $l=3.9e-07 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=3.255 $Y2=1.515
r62 23 25 53.2177 $w=3.17e-07 $l=3.5e-07 $layer=POLY_cond $X=2.515 $Y=1.515
+ $X2=2.865 $Y2=1.515
r63 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.515 $X2=2.515 $Y2=1.515
r64 21 23 13.6845 $w=3.17e-07 $l=9e-08 $layer=POLY_cond $X=2.425 $Y=1.515
+ $X2=2.515 $Y2=1.515
r65 18 24 3.35013 $w=4.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.515 $Y2=1.565
r66 17 24 9.51435 $w=4.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.515 $Y2=1.565
r67 13 27 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.68
+ $X2=3.315 $Y2=1.515
r68 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.315 $Y=1.68
+ $X2=3.315 $Y2=2.4
r69 9 26 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=1.515
r70 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=0.74
r71 5 25 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.68
+ $X2=2.865 $Y2=1.515
r72 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.865 $Y=1.68
+ $X2=2.865 $Y2=2.4
r73 1 21 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=1.515
r74 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A2 3 7 11 15 17 18 28
r49 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.215 $Y=1.515
+ $X2=4.23 $Y2=1.515
r50 25 27 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.84 $Y=1.515
+ $X2=4.215 $Y2=1.515
r51 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.515 $X2=3.84 $Y2=1.515
r52 23 25 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.515
+ $X2=3.84 $Y2=1.515
r53 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.75 $Y=1.515
+ $X2=3.765 $Y2=1.515
r54 18 26 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.84 $Y2=1.565
r55 17 26 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.84 $Y2=1.565
r56 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.35
+ $X2=4.23 $Y2=1.515
r57 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.23 $Y=1.35
+ $X2=4.23 $Y2=0.74
r58 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.215 $Y=1.68
+ $X2=4.215 $Y2=1.515
r59 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.215 $Y=1.68
+ $X2=4.215 $Y2=2.4
r60 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.68
+ $X2=3.765 $Y2=1.515
r61 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.765 $Y=1.68
+ $X2=3.765 $Y2=2.4
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.75 $Y=1.35
+ $X2=3.75 $Y2=1.515
r63 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.75 $Y=1.35 $X2=3.75
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A1 3 7 11 15 17 18 19 20 21 26 35
r47 34 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.73 $Y=1.515
+ $X2=5.745 $Y2=1.515
r48 32 34 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=5.455 $Y=1.515
+ $X2=5.73 $Y2=1.515
r49 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.515 $X2=5.455 $Y2=1.515
r50 30 32 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.275 $Y=1.515
+ $X2=5.455 $Y2=1.515
r51 29 33 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.115 $Y=1.565
+ $X2=5.455 $Y2=1.565
r52 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.115
+ $Y=1.515 $X2=5.115 $Y2=1.515
r53 26 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.185 $Y=1.515
+ $X2=5.275 $Y2=1.515
r54 26 28 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.185 $Y=1.515
+ $X2=5.115 $Y2=1.515
r55 20 21 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.565 $X2=6
+ $Y2=1.565
r56 20 33 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.455 $Y2=1.565
r57 19 29 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.115 $Y2=1.565
r58 18 19 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r59 17 28 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.76 $Y=1.515
+ $X2=5.115 $Y2=1.515
r60 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=1.515
r61 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=0.74
r62 9 34 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.68
+ $X2=5.73 $Y2=1.515
r63 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.73 $Y=1.68 $X2=5.73
+ $Y2=2.4
r64 5 30 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.68
+ $X2=5.275 $Y2=1.515
r65 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.275 $Y=1.68
+ $X2=5.275 $Y2=2.4
r66 1 17 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.685 $Y=1.35
+ $X2=4.76 $Y2=1.515
r67 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.685 $Y=1.35
+ $X2=4.685 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A_27_368# 1 2 3 12 16 17 18 20 27
c31 27 0 1.72955e-19 $X=2.08 $Y=2.455
c32 12 0 1.94533e-19 $X=0.28 $Y=2.115
r33 21 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.375
+ $X2=1.18 $Y2=2.375
r34 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=2.375
+ $X2=2.08 $Y2=2.375
r35 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.915 $Y=2.375
+ $X2=1.265 $Y2=2.375
r36 18 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.46 $X2=1.18
+ $Y2=2.375
r37 18 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.18 $Y=2.46
+ $X2=1.18 $Y2=2.905
r38 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=1.18 $Y2=2.905
r39 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=0.365 $Y2=2.99
r40 12 15 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=2.115 $X2=0.24
+ $Y2=2.815
r41 10 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.365 $Y2=2.99
r42 10 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=2.905 $X2=0.24
+ $Y2=2.815
r43 3 27 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.455
r44 2 25 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.455
r45 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r46 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%Y 1 2 3 4 15 19 20 21 25 27 32 33 34 35 45
+ 46
r86 45 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=1.985
+ $X2=3.09 $Y2=1.82
r87 34 45 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.09 $Y=2.035 $X2=3.09
+ $Y2=1.985
r88 34 35 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=3.09 $Y=2.12
+ $X2=3.09 $Y2=2.405
r89 29 46 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.01 $Y=1.18 $X2=3.01
+ $Y2=1.82
r90 28 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.095
+ $X2=1.71 $Y2=1.095
r91 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.925 $Y=1.095
+ $X2=3.01 $Y2=1.18
r92 27 28 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=2.925 $Y=1.095
+ $X2=1.875 $Y2=1.095
r93 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.01 $X2=1.71
+ $Y2=1.095
r94 23 25 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.71 $Y=1.01
+ $X2=1.71 $Y2=0.775
r95 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=2.035
r96 21 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=3.09 $Y2=2.035
r97 21 22 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=0.895 $Y2=2.035
r98 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=1.71 $Y2=1.095
r99 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=0.875 $Y2=1.095
r100 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.875 $Y2=1.095
r101 13 15 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.775
r102 4 45 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.84 $X2=3.09 $Y2=1.985
r103 3 32 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.115
r104 2 25 182 $w=1.7e-07 $l=4.99074e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.775
r105 1 15 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%VPWR 1 2 3 12 16 18 20 24 26 34 39 45 48 52
c64 12 0 1.87992e-19 $X=1.63 $Y=2.805
r65 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r66 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r67 45 46 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 43 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r69 43 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r70 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r71 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=3.33 $X2=5
+ $Y2=3.33
r72 40 42 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 39 51 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=6.055 $Y2=3.33
r74 39 42 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r76 37 38 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 35 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.59 $Y2=3.33
r78 35 37 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=3.33 $X2=5
+ $Y2=3.33
r80 34 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 29 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r84 28 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.59 $Y2=3.33
r87 26 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r88 24 38 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r89 24 46 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.68 $Y2=3.33
r90 20 23 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.995 $Y=2.115
+ $X2=5.995 $Y2=2.815
r91 18 51 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.995 $Y=3.245
+ $X2=6.055 $Y2=3.33
r92 18 23 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.995 $Y=3.245
+ $X2=5.995 $Y2=2.815
r93 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=3.33
r94 14 16 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=2.455
r95 10 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=3.33
r96 10 12 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=2.805
r97 3 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.84 $X2=5.955 $Y2=2.815
r98 3 20 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.84 $X2=5.955 $Y2=2.115
r99 2 16 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.84 $X2=5 $Y2=2.455
r100 1 12 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A_499_368# 1 2 3 12 14 15 18 22 26 28
r34 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.44 $Y=2.905
+ $X2=4.44 $Y2=2.455
r35 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=3.54 $Y2=2.99
r36 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.275 $Y=2.99
+ $X2=4.44 $Y2=2.905
r37 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.275 $Y=2.99
+ $X2=3.625 $Y2=2.99
r38 18 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.54 $Y=2.115 $X2=3.54
+ $Y2=2.815
r39 16 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.905
+ $X2=3.54 $Y2=2.99
r40 16 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=2.905 $X2=3.54
+ $Y2=2.815
r41 14 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=3.54 $Y2=2.99
r42 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=2.725 $Y2=2.99
r43 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.6 $Y=2.905
+ $X2=2.725 $Y2=2.99
r44 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.6 $Y=2.905 $X2=2.6
+ $Y2=2.455
r45 3 26 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.84 $X2=4.44 $Y2=2.455
r46 2 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.84 $X2=3.54 $Y2=2.815
r47 2 18 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.84 $X2=3.54 $Y2=2.115
r48 1 12 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=2.64 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A_771_368# 1 2 9 11 13 16
r26 11 18 2.63384 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.502 $Y=2.12
+ $X2=5.502 $Y2=2.035
r27 11 13 23.9089 $w=3.33e-07 $l=6.95e-07 $layer=LI1_cond $X=5.502 $Y=2.12
+ $X2=5.502 $Y2=2.815
r28 10 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.035
+ $X2=3.95 $Y2=2.035
r29 9 18 5.17472 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=5.502 $Y2=2.035
r30 9 10 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=4.075 $Y2=2.035
r31 2 18 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.84 $X2=5.5 $Y2=2.035
r32 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.84 $X2=5.5 $Y2=2.815
r33 1 16 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=3.855
+ $Y=1.84 $X2=3.99 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%A_27_74# 1 2 3 4 5 6 21 23 24 27 29 34 35 36
+ 38 39 40 43 45 49 51 53 56
r91 53 55 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.47 $Y=0.515
+ $X2=3.47 $Y2=0.755
r92 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.96 $Y=1.01
+ $X2=5.96 $Y2=0.515
r93 46 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=1.095
+ $X2=4.47 $Y2=1.095
r94 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.795 $Y=1.095
+ $X2=5.96 $Y2=1.01
r95 45 46 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.795 $Y=1.095
+ $X2=4.635 $Y2=1.095
r96 41 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=1.01 $X2=4.47
+ $Y2=1.095
r97 41 43 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.47 $Y=1.01
+ $X2=4.47 $Y2=0.515
r98 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=1.095
+ $X2=4.47 $Y2=1.095
r99 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.305 $Y=1.095
+ $X2=3.635 $Y2=1.095
r100 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.47 $Y=1.01
+ $X2=3.635 $Y2=1.095
r101 37 55 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=0.84
+ $X2=3.47 $Y2=0.755
r102 37 38 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.47 $Y=0.84
+ $X2=3.47 $Y2=1.01
r103 35 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0.755
+ $X2=3.47 $Y2=0.755
r104 35 36 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.305 $Y=0.755
+ $X2=2.375 $Y2=0.755
r105 32 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.21 $Y=0.67
+ $X2=2.375 $Y2=0.755
r106 32 34 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.21 $Y=0.67
+ $X2=2.21 $Y2=0.595
r107 31 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.21 $Y=0.425
+ $X2=2.21 $Y2=0.595
r108 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r109 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=2.21 $Y2=0.425
r110 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=1.375 $Y2=0.34
r111 25 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.34
r112 25 27 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.66
r113 23 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r114 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r115 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r116 19 21 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.24 $Y2=0.515
r117 6 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.37 $X2=5.96 $Y2=0.515
r118 5 43 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.37 $X2=4.47 $Y2=0.515
r119 4 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.33
+ $Y=0.37 $X2=3.47 $Y2=0.515
r120 3 34 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.37
+ $X2=2.21 $Y2=0.595
r121 2 27 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.66
r122 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_2%VGND 1 2 3 12 15 16 17 37 38 43 46 50 56
r66 55 56 11.2541 $w=8.88e-07 $l=9.5e-08 $layer=LI1_cond $X=5.53 $Y=0.36
+ $X2=5.625 $Y2=0.36
r67 52 55 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=5.52 $Y=0.36 $X2=5.53
+ $Y2=0.36
r68 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r69 49 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r70 48 52 6.57978 $w=8.88e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=0.36
+ $X2=5.52 $Y2=0.36
r71 48 50 13.1732 $w=8.88e-07 $l=2.35e-07 $layer=LI1_cond $X=5.04 $Y=0.36
+ $X2=4.805 $Y2=0.36
r72 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r73 45 46 12.5119 $w=5.83e-07 $l=2.85e-07 $layer=LI1_cond $X=2.84 $Y=0.207
+ $X2=3.125 $Y2=0.207
r74 41 45 4.08916 $w=5.83e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=0.207 $X2=2.84
+ $Y2=0.207
r75 41 43 8.42273 $w=5.83e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=2.555 $Y2=0.207
r76 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r77 38 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r78 37 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6 $Y=0 $X2=5.625
+ $Y2=0
r79 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r80 34 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r81 33 50 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.805
+ $Y2=0
r82 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r83 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r84 29 46 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.125
+ $Y2=0
r85 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r86 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r87 25 43 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.555
+ $Y2=0
r88 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r89 22 26 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r90 21 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r91 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r92 17 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r93 17 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r94 15 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.6
+ $Y2=0
r95 15 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.97
+ $Y2=0
r96 14 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.135 $Y=0 $X2=4.56
+ $Y2=0
r97 14 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=0 $X2=3.97
+ $Y2=0
r98 10 16 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=0.085
+ $X2=3.97 $Y2=0
r99 10 12 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.97 $Y=0.085
+ $X2=3.97 $Y2=0.635
r100 3 55 91 $w=1.7e-07 $l=8.94874e-07 $layer=licon1_NDIFF $count=2 $X=4.76
+ $Y=0.37 $X2=5.53 $Y2=0.64
r101 2 12 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=3.825
+ $Y=0.37 $X2=3.97 $Y2=0.635
r102 1 45 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.37 $X2=2.84 $Y2=0.335
.ends


* File: sky130_fd_sc_ms__or3b_2.pxi.spice
* Created: Wed Sep  2 12:28:37 2020
* 
x_PM_SKY130_FD_SC_MS__OR3B_2%C_N N_C_N_c_70_n N_C_N_M1002_g N_C_N_M1005_g C_N
+ N_C_N_c_72_n PM_SKY130_FD_SC_MS__OR3B_2%C_N
x_PM_SKY130_FD_SC_MS__OR3B_2%A_190_260# N_A_190_260#_M1007_d
+ N_A_190_260#_M1000_d N_A_190_260#_M1009_d N_A_190_260#_M1010_g
+ N_A_190_260#_M1004_g N_A_190_260#_c_97_n N_A_190_260#_M1011_g
+ N_A_190_260#_M1008_g N_A_190_260#_c_100_n N_A_190_260#_c_101_n
+ N_A_190_260#_c_102_n N_A_190_260#_c_103_n N_A_190_260#_c_104_n
+ N_A_190_260#_c_105_n N_A_190_260#_c_106_n N_A_190_260#_c_111_n
+ N_A_190_260#_c_107_n N_A_190_260#_c_108_n
+ PM_SKY130_FD_SC_MS__OR3B_2%A_190_260#
x_PM_SKY130_FD_SC_MS__OR3B_2%A N_A_M1001_g N_A_M1007_g A A N_A_c_210_n
+ N_A_c_211_n PM_SKY130_FD_SC_MS__OR3B_2%A
x_PM_SKY130_FD_SC_MS__OR3B_2%B N_B_M1003_g N_B_M1006_g B N_B_c_254_n N_B_c_255_n
+ PM_SKY130_FD_SC_MS__OR3B_2%B
x_PM_SKY130_FD_SC_MS__OR3B_2%A_27_368# N_A_27_368#_M1005_s N_A_27_368#_M1002_s
+ N_A_27_368#_M1009_g N_A_27_368#_M1000_g N_A_27_368#_c_296_n
+ N_A_27_368#_c_320_n N_A_27_368#_c_323_n N_A_27_368#_c_324_n
+ N_A_27_368#_c_344_n N_A_27_368#_c_297_n N_A_27_368#_c_298_n
+ N_A_27_368#_c_303_n N_A_27_368#_c_299_n N_A_27_368#_c_304_n
+ PM_SKY130_FD_SC_MS__OR3B_2%A_27_368#
x_PM_SKY130_FD_SC_MS__OR3B_2%VPWR N_VPWR_M1002_d N_VPWR_M1011_s N_VPWR_c_391_n
+ N_VPWR_c_392_n N_VPWR_c_393_n VPWR N_VPWR_c_394_n N_VPWR_c_390_n
+ N_VPWR_c_396_n N_VPWR_c_397_n PM_SKY130_FD_SC_MS__OR3B_2%VPWR
x_PM_SKY130_FD_SC_MS__OR3B_2%X N_X_M1004_d N_X_M1010_d N_X_c_429_n N_X_c_430_n
+ N_X_c_431_n X X PM_SKY130_FD_SC_MS__OR3B_2%X
x_PM_SKY130_FD_SC_MS__OR3B_2%VGND N_VGND_M1005_d N_VGND_M1008_s N_VGND_M1006_d
+ N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n VGND N_VGND_c_478_n
+ N_VGND_c_479_n N_VGND_c_480_n PM_SKY130_FD_SC_MS__OR3B_2%VGND
cc_1 VNB N_C_N_c_70_n 0.0646212f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.78
cc_2 VNB N_C_N_M1005_g 0.029568f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_3 VNB N_C_N_c_72_n 0.00652172f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A_190_260#_M1010_g 0.0113917f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_5 VNB N_A_190_260#_M1004_g 0.0217342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_190_260#_c_97_n 0.0363841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_190_260#_M1011_g 0.00171409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_190_260#_M1008_g 0.0236017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_190_260#_c_100_n 0.00908278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_190_260#_c_101_n 0.0089459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_190_260#_c_102_n 0.00897658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_190_260#_c_103_n 0.00328996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_190_260#_c_104_n 0.00951425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_190_260#_c_105_n 0.0272219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_190_260#_c_106_n 0.00761269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_190_260#_c_107_n 0.0226504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_190_260#_c_108_n 0.0149819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_M1007_g 0.0271057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_c_210_n 0.026818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_211_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_21 VNB N_B_M1006_g 0.0258186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_254_n 0.0266192f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_23 VNB N_B_c_255_n 0.0016559f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_24 VNB N_A_27_368#_M1000_g 0.0311299f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_25 VNB N_A_27_368#_c_296_n 0.00523497f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_26 VNB N_A_27_368#_c_297_n 0.00167078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_368#_c_298_n 0.0289629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_368#_c_299_n 0.0293174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_390_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_429_n 0.00273546f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_X_c_430_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_32 VNB N_X_c_431_n 0.00422231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_470_n 0.0111927f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_34 VNB N_VGND_c_471_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_472_n 0.0166983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_473_n 0.018099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_474_n 0.024548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_475_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_476_n 0.0205837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_477_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_478_n 0.020559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_479_n 0.247561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_480_n 0.00980973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_C_N_c_70_n 0.03071f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.78
cc_45 VPB N_C_N_c_72_n 0.00761845f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_46 VPB N_A_190_260#_M1010_g 0.0239191f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_47 VPB N_A_190_260#_M1011_g 0.0247794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_190_260#_c_111_n 0.033624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_190_260#_c_107_n 0.0300171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_M1001_g 0.0224314f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_51 VPB N_A_c_210_n 0.00576827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_c_211_n 0.00191357f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_53 VPB N_B_M1003_g 0.0208876f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_54 VPB N_B_c_254_n 0.00561656f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_55 VPB N_B_c_255_n 0.00274372f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_56 VPB N_A_27_368#_c_296_n 0.00316182f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_57 VPB N_A_27_368#_c_297_n 0.00106862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_27_368#_c_298_n 0.00945897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_27_368#_c_303_n 0.0344781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_368#_c_304_n 0.0241186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_391_n 0.0163583f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_62 VPB N_VPWR_c_392_n 0.0206218f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_63 VPB N_VPWR_c_393_n 0.0148008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_394_n 0.0552717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_390_n 0.0872715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_396_n 0.0274712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_397_n 0.00834123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_429_n 0.00152096f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_69 VPB X 0.00598134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_C_N_c_70_n N_A_190_260#_M1010_g 0.0361765f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_71 N_C_N_M1005_g N_A_190_260#_M1004_g 0.0195624f $X=0.565 $Y=0.835 $X2=0
+ $Y2=0
cc_72 N_C_N_c_70_n N_A_190_260#_c_100_n 0.00597962f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_73 N_C_N_c_70_n N_A_27_368#_c_296_n 0.00963071f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_74 N_C_N_M1005_g N_A_27_368#_c_296_n 0.00652595f $X=0.565 $Y=0.835 $X2=0
+ $Y2=0
cc_75 N_C_N_c_72_n N_A_27_368#_c_296_n 0.0355099f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_76 N_C_N_c_70_n N_A_27_368#_c_303_n 0.0333294f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_77 N_C_N_c_72_n N_A_27_368#_c_303_n 0.0258519f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_78 N_C_N_c_70_n N_A_27_368#_c_299_n 0.00470761f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_79 N_C_N_M1005_g N_A_27_368#_c_299_n 0.0242901f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_80 N_C_N_c_72_n N_A_27_368#_c_299_n 0.0214092f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_81 N_C_N_c_70_n N_VPWR_c_391_n 0.00339971f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_82 N_C_N_c_70_n N_VPWR_c_390_n 0.00555093f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_83 N_C_N_c_70_n N_VPWR_c_396_n 0.0046462f $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_84 N_C_N_c_70_n N_X_c_429_n 5.81161e-19 $X=0.505 $Y=1.78 $X2=0 $Y2=0
cc_85 N_C_N_M1005_g N_X_c_430_n 5.95409e-19 $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_86 N_C_N_M1005_g N_X_c_431_n 2.34935e-19 $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_87 N_C_N_M1005_g N_VGND_c_470_n 0.00417177f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_88 N_C_N_M1005_g N_VGND_c_474_n 0.00366404f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_89 N_C_N_M1005_g N_VGND_c_479_n 0.00487769f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_90 N_A_190_260#_M1011_g N_A_M1001_g 0.0241087f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_190_260#_c_97_n N_A_M1007_g 0.00119833f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_92 N_A_190_260#_M1008_g N_A_M1007_g 0.0147478f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_190_260#_c_101_n N_A_M1007_g 0.0162422f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_94 N_A_190_260#_c_102_n N_A_M1007_g 0.00325729f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_95 N_A_190_260#_c_103_n N_A_M1007_g 0.00299701f $X=2.515 $Y=0.615 $X2=0 $Y2=0
cc_96 N_A_190_260#_c_97_n N_A_c_210_n 0.0147986f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_97 N_A_190_260#_M1011_g N_A_c_210_n 0.00167705f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_190_260#_c_101_n N_A_c_210_n 0.00125903f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_99 N_A_190_260#_c_102_n N_A_c_210_n 0.00172393f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_100 N_A_190_260#_c_97_n N_A_c_211_n 3.15084e-19 $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_101 N_A_190_260#_M1011_g N_A_c_211_n 0.00396351f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_190_260#_c_101_n N_A_c_211_n 0.0256551f $X=2.35 $Y=1.095 $X2=0 $Y2=0
cc_103 N_A_190_260#_c_102_n N_A_c_211_n 0.0216131f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_104 N_A_190_260#_c_111_n N_B_M1003_g 0.00229611f $X=3.4 $Y=2.375 $X2=0 $Y2=0
cc_105 N_A_190_260#_c_103_n N_B_M1006_g 0.00798791f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_106 N_A_190_260#_c_104_n N_B_M1006_g 0.0116271f $X=3.35 $Y=1.095 $X2=0 $Y2=0
cc_107 N_A_190_260#_c_105_n N_B_M1006_g 6.07993e-19 $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_108 N_A_190_260#_c_106_n N_B_M1006_g 0.00171282f $X=2.515 $Y=1.095 $X2=0
+ $Y2=0
cc_109 N_A_190_260#_c_104_n N_B_c_254_n 2.7493e-19 $X=3.35 $Y=1.095 $X2=0 $Y2=0
cc_110 N_A_190_260#_c_106_n N_B_c_254_n 0.00108976f $X=2.515 $Y=1.095 $X2=0
+ $Y2=0
cc_111 N_A_190_260#_c_104_n N_B_c_255_n 0.0121392f $X=3.35 $Y=1.095 $X2=0 $Y2=0
cc_112 N_A_190_260#_c_106_n N_B_c_255_n 0.0140411f $X=2.515 $Y=1.095 $X2=0 $Y2=0
cc_113 N_A_190_260#_c_103_n N_A_27_368#_M1000_g 6.0898e-19 $X=2.515 $Y=0.615
+ $X2=0 $Y2=0
cc_114 N_A_190_260#_c_104_n N_A_27_368#_M1000_g 0.0116271f $X=3.35 $Y=1.095
+ $X2=0 $Y2=0
cc_115 N_A_190_260#_c_105_n N_A_27_368#_M1000_g 0.00816329f $X=3.515 $Y=0.615
+ $X2=0 $Y2=0
cc_116 N_A_190_260#_c_107_n N_A_27_368#_M1000_g 0.00391901f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_117 N_A_190_260#_c_108_n N_A_27_368#_M1000_g 0.00221813f $X=3.552 $Y=1.095
+ $X2=0 $Y2=0
cc_118 N_A_190_260#_M1004_g N_A_27_368#_c_296_n 0.00123682f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_119 N_A_190_260#_c_100_n N_A_27_368#_c_296_n 0.00532417f $X=1.05 $Y=1.375
+ $X2=0 $Y2=0
cc_120 N_A_190_260#_M1010_g N_A_27_368#_c_320_n 0.0170047f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_121 N_A_190_260#_M1011_g N_A_27_368#_c_320_n 0.0145159f $X=1.49 $Y=2.4 $X2=0
+ $Y2=0
cc_122 N_A_190_260#_c_111_n N_A_27_368#_c_320_n 0.00500344f $X=3.4 $Y=2.375
+ $X2=0 $Y2=0
cc_123 N_A_190_260#_c_111_n N_A_27_368#_c_323_n 7.83251e-19 $X=3.4 $Y=2.375
+ $X2=0 $Y2=0
cc_124 N_A_190_260#_M1009_d N_A_27_368#_c_324_n 0.00290398f $X=3.265 $Y=1.84
+ $X2=0 $Y2=0
cc_125 N_A_190_260#_c_111_n N_A_27_368#_c_324_n 0.0106128f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_126 N_A_190_260#_c_107_n N_A_27_368#_c_324_n 0.0140565f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_127 N_A_190_260#_M1009_d N_A_27_368#_c_297_n 0.00118548f $X=3.265 $Y=1.84
+ $X2=0 $Y2=0
cc_128 N_A_190_260#_c_104_n N_A_27_368#_c_297_n 0.0205962f $X=3.35 $Y=1.095
+ $X2=0 $Y2=0
cc_129 N_A_190_260#_c_107_n N_A_27_368#_c_297_n 0.0458135f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_130 N_A_190_260#_c_108_n N_A_27_368#_c_297_n 0.0055933f $X=3.552 $Y=1.095
+ $X2=0 $Y2=0
cc_131 N_A_190_260#_c_104_n N_A_27_368#_c_298_n 9.6679e-19 $X=3.35 $Y=1.095
+ $X2=0 $Y2=0
cc_132 N_A_190_260#_c_111_n N_A_27_368#_c_298_n 4.2865e-19 $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_133 N_A_190_260#_c_107_n N_A_27_368#_c_298_n 0.00840771f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_134 N_A_190_260#_c_108_n N_A_27_368#_c_298_n 3.08066e-19 $X=3.552 $Y=1.095
+ $X2=0 $Y2=0
cc_135 N_A_190_260#_M1010_g N_A_27_368#_c_303_n 0.00715311f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_136 N_A_190_260#_M1004_g N_A_27_368#_c_299_n 0.00203846f $X=1.075 $Y=0.74
+ $X2=0 $Y2=0
cc_137 N_A_190_260#_c_111_n N_A_27_368#_c_304_n 0.0131052f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_138 N_A_190_260#_c_107_n N_A_27_368#_c_304_n 0.00463021f $X=3.495 $Y=2.29
+ $X2=0 $Y2=0
cc_139 N_A_190_260#_M1010_g N_VPWR_c_391_n 0.012355f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_190_260#_M1011_g N_VPWR_c_391_n 0.00130014f $X=1.49 $Y=2.4 $X2=0
+ $Y2=0
cc_141 N_A_190_260#_M1010_g N_VPWR_c_392_n 0.00460063f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_190_260#_M1011_g N_VPWR_c_392_n 0.00553757f $X=1.49 $Y=2.4 $X2=0
+ $Y2=0
cc_143 N_A_190_260#_M1011_g N_VPWR_c_393_n 0.00612791f $X=1.49 $Y=2.4 $X2=0
+ $Y2=0
cc_144 N_A_190_260#_c_111_n N_VPWR_c_394_n 0.0153256f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_145 N_A_190_260#_M1010_g N_VPWR_c_390_n 0.0046086f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_190_260#_M1011_g N_VPWR_c_390_n 0.00560227f $X=1.49 $Y=2.4 $X2=0
+ $Y2=0
cc_147 N_A_190_260#_c_111_n N_VPWR_c_390_n 0.0175815f $X=3.4 $Y=2.375 $X2=0
+ $Y2=0
cc_148 N_A_190_260#_M1010_g N_X_c_429_n 0.0149133f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_190_260#_M1004_g N_X_c_429_n 0.00382206f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_190_260#_c_97_n N_X_c_429_n 0.00859318f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_151 N_A_190_260#_M1008_g N_X_c_429_n 0.00127735f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_190_260#_c_100_n N_X_c_429_n 0.00275812f $X=1.05 $Y=1.375 $X2=0 $Y2=0
cc_153 N_A_190_260#_c_102_n N_X_c_429_n 0.0321078f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_154 N_A_190_260#_M1004_g N_X_c_430_n 0.00881022f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_190_260#_M1008_g N_X_c_430_n 0.0135262f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_190_260#_M1004_g N_X_c_431_n 0.00618144f $X=1.075 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_190_260#_c_97_n N_X_c_431_n 0.00432913f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_158 N_A_190_260#_M1008_g N_X_c_431_n 0.00405854f $X=1.505 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_190_260#_c_102_n N_X_c_431_n 0.00957189f $X=1.795 $Y=1.095 $X2=0
+ $Y2=0
cc_160 N_A_190_260#_c_97_n X 0.00338917f $X=1.4 $Y=1.375 $X2=0 $Y2=0
cc_161 N_A_190_260#_M1011_g X 0.0155763f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_190_260#_c_102_n X 0.0286568f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_163 N_A_190_260#_c_101_n N_VGND_M1008_s 0.00464866f $X=2.35 $Y=1.095 $X2=0
+ $Y2=0
cc_164 N_A_190_260#_c_102_n N_VGND_M1008_s 0.002869f $X=1.795 $Y=1.095 $X2=0
+ $Y2=0
cc_165 N_A_190_260#_c_104_n N_VGND_M1006_d 0.00358162f $X=3.35 $Y=1.095 $X2=0
+ $Y2=0
cc_166 N_A_190_260#_M1004_g N_VGND_c_470_n 0.00490645f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_190_260#_M1004_g N_VGND_c_471_n 0.00434272f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_190_260#_M1008_g N_VGND_c_471_n 0.00434272f $X=1.505 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_190_260#_c_97_n N_VGND_c_472_n 4.47758e-19 $X=1.4 $Y=1.375 $X2=0
+ $Y2=0
cc_170 N_A_190_260#_M1008_g N_VGND_c_472_n 0.00820727f $X=1.505 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_190_260#_c_101_n N_VGND_c_472_n 0.0196678f $X=2.35 $Y=1.095 $X2=0
+ $Y2=0
cc_172 N_A_190_260#_c_102_n N_VGND_c_472_n 0.0112912f $X=1.795 $Y=1.095 $X2=0
+ $Y2=0
cc_173 N_A_190_260#_c_103_n N_VGND_c_472_n 0.00138617f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_174 N_A_190_260#_c_103_n N_VGND_c_473_n 0.0154242f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_175 N_A_190_260#_c_104_n N_VGND_c_473_n 0.0248957f $X=3.35 $Y=1.095 $X2=0
+ $Y2=0
cc_176 N_A_190_260#_c_105_n N_VGND_c_473_n 0.01589f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_177 N_A_190_260#_c_103_n N_VGND_c_476_n 0.0103491f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_178 N_A_190_260#_c_105_n N_VGND_c_478_n 0.0127299f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_179 N_A_190_260#_M1004_g N_VGND_c_479_n 0.00825283f $X=1.075 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_A_190_260#_M1008_g N_VGND_c_479_n 0.00825059f $X=1.505 $Y=0.74 $X2=0
+ $Y2=0
cc_181 N_A_190_260#_c_103_n N_VGND_c_479_n 0.0113354f $X=2.515 $Y=0.615 $X2=0
+ $Y2=0
cc_182 N_A_190_260#_c_105_n N_VGND_c_479_n 0.0139328f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_183 N_A_M1001_g N_B_M1003_g 0.0696191f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_184 N_A_c_211_n N_B_M1003_g 0.00146529f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A_M1007_g N_B_M1006_g 0.021941f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_186 N_A_c_210_n N_B_c_254_n 0.0201104f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_187 N_A_c_211_n N_B_c_254_n 0.00114936f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_188 N_A_M1001_g N_B_c_255_n 5.64277e-19 $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_189 N_A_c_210_n N_B_c_255_n 0.00114936f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A_c_211_n N_B_c_255_n 0.0276387f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A_M1001_g N_A_27_368#_c_320_n 0.0141605f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_192 N_A_c_210_n N_A_27_368#_c_320_n 3.56046e-19 $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A_c_211_n N_A_27_368#_c_320_n 0.0211204f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A_M1001_g N_A_27_368#_c_323_n 0.0036f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_195 N_A_c_211_n N_A_27_368#_c_323_n 0.00217881f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A_M1001_g N_A_27_368#_c_344_n 0.00103411f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_197 N_A_c_211_n N_A_27_368#_c_344_n 0.0140387f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A_c_211_n N_VPWR_M1011_s 0.00395846f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A_M1001_g N_VPWR_c_393_n 0.00551792f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_200 N_A_M1001_g N_VPWR_c_394_n 0.0059286f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_201 N_A_M1001_g N_VPWR_c_390_n 0.00610055f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_202 N_A_M1001_g X 0.00110362f $X=2.215 $Y=2.34 $X2=0 $Y2=0
cc_203 N_A_c_211_n X 0.0268279f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_204 N_A_M1007_g N_VGND_c_472_n 0.00658658f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_205 N_A_M1007_g N_VGND_c_476_n 0.00507111f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_206 N_A_M1007_g N_VGND_c_479_n 0.00514438f $X=2.23 $Y=0.79 $X2=0 $Y2=0
cc_207 N_B_M1006_g N_A_27_368#_M1000_g 0.0240664f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_208 N_B_M1003_g N_A_27_368#_c_320_n 0.00852694f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_209 N_B_M1003_g N_A_27_368#_c_323_n 0.0056859f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_210 N_B_M1003_g N_A_27_368#_c_324_n 0.00821682f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_211 N_B_c_254_n N_A_27_368#_c_324_n 5.39698e-19 $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_212 N_B_c_255_n N_A_27_368#_c_324_n 0.0132765f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_213 N_B_M1003_g N_A_27_368#_c_344_n 0.00375255f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_214 N_B_c_255_n N_A_27_368#_c_344_n 0.0093022f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_215 N_B_M1003_g N_A_27_368#_c_297_n 0.00112952f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_216 N_B_c_254_n N_A_27_368#_c_297_n 0.00121489f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_217 N_B_c_255_n N_A_27_368#_c_297_n 0.0248917f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_218 N_B_M1003_g N_A_27_368#_c_298_n 0.0447628f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_219 N_B_c_254_n N_A_27_368#_c_298_n 0.017083f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_220 N_B_c_255_n N_A_27_368#_c_298_n 0.00192255f $X=2.68 $Y=1.515 $X2=0 $Y2=0
cc_221 N_B_M1003_g N_VPWR_c_394_n 0.0059286f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_222 N_B_M1003_g N_VPWR_c_390_n 0.00610055f $X=2.635 $Y=2.34 $X2=0 $Y2=0
cc_223 N_B_M1006_g N_VGND_c_473_n 0.00564618f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_224 N_B_M1006_g N_VGND_c_476_n 0.00485498f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_225 N_B_M1006_g N_VGND_c_479_n 0.00514438f $X=2.73 $Y=0.79 $X2=0 $Y2=0
cc_226 N_A_27_368#_c_296_n N_VPWR_M1002_d 0.00115589f $X=0.69 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_27_368#_c_320_n N_VPWR_M1002_d 0.00569107f $X=2.475 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_228 N_A_27_368#_c_303_n N_VPWR_M1002_d 0.00581669f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_229 N_A_27_368#_c_320_n N_VPWR_M1011_s 0.0156629f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_230 N_A_27_368#_c_320_n N_VPWR_c_391_n 0.011474f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_231 N_A_27_368#_c_303_n N_VPWR_c_391_n 0.0127735f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_232 N_A_27_368#_c_320_n N_VPWR_c_393_n 0.0342973f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_233 N_A_27_368#_c_304_n N_VPWR_c_394_n 0.00567889f $X=3.25 $Y=1.725 $X2=0
+ $Y2=0
cc_234 N_A_27_368#_c_320_n N_VPWR_c_390_n 0.0419266f $X=2.475 $Y=2.405 $X2=0
+ $Y2=0
cc_235 N_A_27_368#_c_303_n N_VPWR_c_390_n 0.0178704f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_236 N_A_27_368#_c_304_n N_VPWR_c_390_n 0.00610055f $X=3.25 $Y=1.725 $X2=0
+ $Y2=0
cc_237 N_A_27_368#_c_303_n N_VPWR_c_396_n 0.006683f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_238 N_A_27_368#_c_320_n N_X_M1010_d 0.00479747f $X=2.475 $Y=2.405 $X2=0 $Y2=0
cc_239 N_A_27_368#_c_296_n N_X_c_429_n 0.0403904f $X=0.69 $Y=1.95 $X2=0 $Y2=0
cc_240 N_A_27_368#_c_320_n N_X_c_429_n 0.00877235f $X=2.475 $Y=2.405 $X2=0 $Y2=0
cc_241 N_A_27_368#_c_303_n N_X_c_429_n 0.0115375f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_242 N_A_27_368#_c_299_n N_X_c_430_n 0.00520473f $X=0.35 $Y=0.835 $X2=0 $Y2=0
cc_243 N_A_27_368#_c_299_n N_X_c_431_n 0.00935177f $X=0.35 $Y=0.835 $X2=0 $Y2=0
cc_244 N_A_27_368#_c_320_n X 0.0331049f $X=2.475 $Y=2.405 $X2=0 $Y2=0
cc_245 N_A_27_368#_c_320_n A_461_368# 0.0068255f $X=2.475 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_246 N_A_27_368#_c_323_n A_461_368# 0.00220282f $X=2.56 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_27_368#_c_344_n A_461_368# 0.00205147f $X=2.645 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_248 N_A_27_368#_c_324_n A_545_368# 0.0169445f $X=3.085 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_249 N_A_27_368#_c_299_n N_VGND_M1005_d 0.00517204f $X=0.35 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_250 N_A_27_368#_c_299_n N_VGND_c_470_n 0.0189052f $X=0.35 $Y=0.835 $X2=0
+ $Y2=0
cc_251 N_A_27_368#_M1000_g N_VGND_c_473_n 0.00564618f $X=3.3 $Y=0.79 $X2=0 $Y2=0
cc_252 N_A_27_368#_c_299_n N_VGND_c_474_n 0.0101249f $X=0.35 $Y=0.835 $X2=0
+ $Y2=0
cc_253 N_A_27_368#_M1000_g N_VGND_c_478_n 0.00485498f $X=3.3 $Y=0.79 $X2=0 $Y2=0
cc_254 N_A_27_368#_M1000_g N_VGND_c_479_n 0.00514438f $X=3.3 $Y=0.79 $X2=0 $Y2=0
cc_255 N_A_27_368#_c_299_n N_VGND_c_479_n 0.0134471f $X=0.35 $Y=0.835 $X2=0
+ $Y2=0
cc_256 N_VPWR_M1011_s X 0.00524448f $X=1.58 $Y=1.84 $X2=0 $Y2=0
cc_257 N_X_c_430_n N_VGND_c_470_n 0.0164567f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_258 N_X_c_430_n N_VGND_c_471_n 0.0144922f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_259 N_X_c_430_n N_VGND_c_472_n 0.0169789f $X=1.29 $Y=0.515 $X2=0 $Y2=0
cc_260 N_X_c_430_n N_VGND_c_479_n 0.0118826f $X=1.29 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__inv_8.pex.spice
* Created: Fri Aug 28 17:38:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__INV_8%A 3 5 7 8 10 13 17 21 25 29 33 37 41 45 49 53
+ 55 57 61 63 64 65 82
c143 13 0 1.53462e-19 $X=0.955 $Y=2.4
r144 81 82 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.085
+ $Y=1.515 $X2=2.085 $Y2=1.515
r145 79 81 24.3708 $w=3.56e-07 $l=1.8e-07 $layer=POLY_cond $X=1.905 $Y=1.44
+ $X2=2.085 $Y2=1.44
r146 74 75 2.0309 $w=3.56e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.44
+ $X2=0.955 $Y2=1.44
r147 72 74 29.1096 $w=3.56e-07 $l=2.15e-07 $layer=POLY_cond $X=0.725 $Y=1.44
+ $X2=0.94 $Y2=1.44
r148 72 73 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.515 $X2=0.725 $Y2=1.515
r149 70 72 29.1096 $w=3.56e-07 $l=2.15e-07 $layer=POLY_cond $X=0.51 $Y=1.44
+ $X2=0.725 $Y2=1.44
r150 69 70 0.676966 $w=3.56e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.44
+ $X2=0.51 $Y2=1.44
r151 65 82 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.085 $Y2=1.565
r152 64 65 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r153 64 73 12.7305 $w=4.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.725 $Y2=1.565
r154 63 73 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.725 $Y2=1.565
r155 59 90 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=3.755 $Y=1.68
+ $X2=3.755 $Y2=1.44
r156 59 61 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.755 $Y=1.68
+ $X2=3.755 $Y2=2.4
r157 55 90 3.38483 $w=3.56e-07 $l=2.5e-08 $layer=POLY_cond $X=3.73 $Y=1.44
+ $X2=3.755 $Y2=1.44
r158 55 88 57.5421 $w=3.56e-07 $l=4.25e-07 $layer=POLY_cond $X=3.73 $Y=1.44
+ $X2=3.305 $Y2=1.44
r159 55 57 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.73 $Y=1.35
+ $X2=3.73 $Y2=0.74
r160 51 88 0.676966 $w=3.56e-07 $l=5e-09 $layer=POLY_cond $X=3.3 $Y=1.44
+ $X2=3.305 $Y2=1.44
r161 51 86 67.0197 $w=3.56e-07 $l=4.95e-07 $layer=POLY_cond $X=3.3 $Y=1.44
+ $X2=2.805 $Y2=1.44
r162 51 53 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.3 $Y=1.35 $X2=3.3
+ $Y2=0.74
r163 47 88 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=3.305 $Y=1.68
+ $X2=3.305 $Y2=1.44
r164 47 49 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.305 $Y=1.68
+ $X2=3.305 $Y2=2.4
r165 43 86 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=2.805 $Y=1.68
+ $X2=2.805 $Y2=1.44
r166 43 45 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.805 $Y=1.68
+ $X2=2.805 $Y2=2.4
r167 39 86 10.1545 $w=3.56e-07 $l=7.5e-08 $layer=POLY_cond $X=2.73 $Y=1.44
+ $X2=2.805 $Y2=1.44
r168 39 84 50.7725 $w=3.56e-07 $l=3.75e-07 $layer=POLY_cond $X=2.73 $Y=1.44
+ $X2=2.355 $Y2=1.44
r169 39 41 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.73 $Y=1.35
+ $X2=2.73 $Y2=0.74
r170 35 84 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=2.355 $Y=1.68
+ $X2=2.355 $Y2=1.44
r171 35 37 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.355 $Y=1.68
+ $X2=2.355 $Y2=2.4
r172 31 84 7.44663 $w=3.56e-07 $l=5.5e-08 $layer=POLY_cond $X=2.3 $Y=1.44
+ $X2=2.355 $Y2=1.44
r173 31 81 29.1096 $w=3.56e-07 $l=2.15e-07 $layer=POLY_cond $X=2.3 $Y=1.44
+ $X2=2.085 $Y2=1.44
r174 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.3
+ $Y2=0.74
r175 27 79 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=1.44
r176 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=2.4
r177 23 79 14.2163 $w=3.56e-07 $l=1.05e-07 $layer=POLY_cond $X=1.8 $Y=1.44
+ $X2=1.905 $Y2=1.44
r178 23 77 46.7107 $w=3.56e-07 $l=3.45e-07 $layer=POLY_cond $X=1.8 $Y=1.44
+ $X2=1.455 $Y2=1.44
r179 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.8 $Y=1.35 $X2=1.8
+ $Y2=0.74
r180 19 77 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.44
r181 19 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r182 15 77 11.5084 $w=3.56e-07 $l=8.5e-08 $layer=POLY_cond $X=1.37 $Y=1.44
+ $X2=1.455 $Y2=1.44
r183 15 75 56.1882 $w=3.56e-07 $l=4.15e-07 $layer=POLY_cond $X=1.37 $Y=1.44
+ $X2=0.955 $Y2=1.44
r184 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.37 $Y=1.35
+ $X2=1.37 $Y2=0.74
r185 11 75 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.44
r186 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r187 8 74 23.0368 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.94 $Y=1.2 $X2=0.94
+ $Y2=1.44
r188 8 10 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.94 $Y=1.2 $X2=0.94
+ $Y2=0.74
r189 5 70 23.0368 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.51 $Y=1.2 $X2=0.51
+ $Y2=1.44
r190 5 7 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.51 $Y=1.2 $X2=0.51
+ $Y2=0.74
r191 1 69 18.7059 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.44
r192 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__INV_8%VPWR 1 2 3 4 5 16 18 24 28 32 36 38 43 44 45
+ 47 52 61 69 72 76
r67 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r68 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r69 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 64 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r72 61 75 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.092 $Y2=3.33
r73 61 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.6 $Y2=3.33
r74 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 57 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.17 $Y2=3.33
r77 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r81 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 52 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.17 $Y2=3.33
r83 52 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r85 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 48 66 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r88 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 47 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r90 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 45 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 45 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 43 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.03 $Y2=3.33
r96 42 63 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.6 $Y2=3.33
r97 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.03 $Y2=3.33
r98 38 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.03 $Y=1.985
+ $X2=4.03 $Y2=2.815
r99 36 75 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.092 $Y2=3.33
r100 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.03 $Y2=2.815
r101 32 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.03 $Y=1.985
+ $X2=3.03 $Y2=2.815
r102 30 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r103 30 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.815
r104 26 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r105 26 28 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.455
r106 22 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r107 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.455
r108 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r109 16 66 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r110 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r111 5 41 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.84 $X2=4.03 $Y2=2.815
r112 5 38 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=3.845
+ $Y=1.84 $X2=4.03 $Y2=1.985
r113 4 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.84 $X2=3.03 $Y2=2.815
r114 4 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.84 $X2=3.03 $Y2=1.985
r115 3 28 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.84 $X2=2.13 $Y2=2.455
r116 2 24 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.455
r117 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r118 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__INV_8%Y 1 2 3 4 5 6 7 8 27 29 31 33 34 35 39 43 45
+ 47 51 54 57 59 63 67 73 75 76 80 81
c130 31 0 1.53462e-19 $X=0.73 $Y=2.815
r131 79 81 9.59355 $w=4.78e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=1.38
+ $X2=4.08 $Y2=1.38
r132 79 80 1.71002 $w=4.8e-07 $l=1.73e-07 $layer=LI1_cond $X=3.695 $Y=1.38
+ $X2=3.522 $Y2=1.38
r133 67 69 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.53 $Y=1.985
+ $X2=3.53 $Y2=2.815
r134 65 80 4.64884 $w=3.3e-07 $l=2.43967e-07 $layer=LI1_cond $X=3.53 $Y=1.62
+ $X2=3.522 $Y2=1.38
r135 65 67 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.53 $Y=1.62
+ $X2=3.53 $Y2=1.985
r136 61 80 4.64884 $w=2.6e-07 $l=2.60154e-07 $layer=LI1_cond $X=3.48 $Y=1.14
+ $X2=3.522 $Y2=1.38
r137 61 63 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=3.48 $Y=1.14
+ $X2=3.48 $Y2=0.515
r138 60 76 2.29025 $w=4.8e-07 $l=5.0892e-07 $layer=LI1_cond $X=2.68 $Y=1.38
+ $X2=2.35 $Y2=1.01
r139 59 80 1.71002 $w=4.8e-07 $l=1.72e-07 $layer=LI1_cond $X=3.35 $Y=1.38
+ $X2=3.522 $Y2=1.38
r140 59 60 16.6953 $w=4.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.35 $Y=1.38
+ $X2=2.68 $Y2=1.38
r141 55 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.035
r142 55 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.4
r143 54 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.95
+ $X2=2.58 $Y2=2.035
r144 53 76 3.88572 $w=1.7e-07 $l=7.15821e-07 $layer=LI1_cond $X=2.58 $Y=1.62
+ $X2=2.35 $Y2=1.01
r145 53 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.58 $Y=1.62
+ $X2=2.58 $Y2=1.95
r146 49 76 3.88572 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.35 $Y2=1.01
r147 49 51 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.515 $Y2=0.515
r148 48 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.035
+ $X2=1.68 $Y2=2.035
r149 47 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=2.035
+ $X2=2.58 $Y2=2.035
r150 47 48 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.495 $Y=2.035
+ $X2=1.845 $Y2=2.035
r151 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.095
+ $X2=1.585 $Y2=1.095
r152 45 76 2.29025 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=2.35 $Y2=1.01
r153 45 46 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=1.67 $Y2=1.095
r154 41 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.12
+ $X2=1.68 $Y2=2.035
r155 41 43 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.68 $Y=2.12
+ $X2=1.68 $Y2=2.815
r156 37 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=1.01
+ $X2=1.585 $Y2=1.095
r157 37 39 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.585 $Y=1.01
+ $X2=1.585 $Y2=0.515
r158 36 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=2.035
+ $X2=0.69 $Y2=2.035
r159 35 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=1.68 $Y2=2.035
r160 35 36 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=0.815 $Y2=2.035
r161 33 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=1.095
+ $X2=1.585 $Y2=1.095
r162 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.5 $Y=1.095
+ $X2=0.81 $Y2=1.095
r163 29 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.12
+ $X2=0.69 $Y2=2.035
r164 29 31 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.69 $Y=2.12
+ $X2=0.69 $Y2=2.815
r165 25 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.685 $Y=1.01
+ $X2=0.81 $Y2=1.095
r166 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.685 $Y=1.01
+ $X2=0.685 $Y2=0.515
r167 8 69 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.84 $X2=3.53 $Y2=2.815
r168 8 67 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.84 $X2=3.53 $Y2=1.985
r169 7 78 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.84 $X2=2.58 $Y2=1.985
r170 7 57 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=1.84 $X2=2.58 $Y2=2.4
r171 6 75 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.115
r172 6 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.815
r173 5 72 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.115
r174 5 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r175 4 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.375
+ $Y=0.37 $X2=3.515 $Y2=0.515
r176 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.375
+ $Y=0.37 $X2=2.515 $Y2=0.515
r177 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.515
r178 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__INV_8%VGND 1 2 3 4 5 16 18 22 26 30 32 34 37 38 40
+ 41 42 44 56 64 68
r67 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r68 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r69 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 59 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r71 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r72 56 67 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=4.05
+ $Y2=0
r73 56 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.78 $Y=0 $X2=3.6
+ $Y2=0
r74 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r75 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r77 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r78 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.155
+ $Y2=0
r79 49 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.68
+ $Y2=0
r80 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r81 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r82 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r83 45 61 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r84 45 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.72
+ $Y2=0
r85 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.155
+ $Y2=0
r86 44 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r87 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r88 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r89 40 54 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.64
+ $Y2=0
r90 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.015
+ $Y2=0
r91 39 58 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.6
+ $Y2=0
r92 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.015
+ $Y2=0
r93 37 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r94 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.015
+ $Y2=0
r95 36 54 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.64
+ $Y2=0
r96 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.015
+ $Y2=0
r97 32 67 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=4.05 $Y2=0
r98 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0.515
r99 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0
r100 28 30 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.495
r101 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0
r102 24 26 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.015 $Y=0.085
+ $X2=2.015 $Y2=0.675
r103 20 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r104 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.675
r105 16 61 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r106 16 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.515
r107 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.805
+ $Y=0.37 $X2=3.945 $Y2=0.515
r108 4 30 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.37 $X2=3.015 $Y2=0.495
r109 3 26 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.37 $X2=2.015 $Y2=0.675
r110 2 22 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.675
r111 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__mux2_4.spice
* Created: Wed Sep  2 12:11:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux2_4.pex.spice"
.subckt sky130_fd_sc_ms__mux2_4  VNB VPB S A0 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_S_M1002_g N_A_27_368#_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.4 A=0.096 P=1.58 MULT=1
MM1006 N_X_M1006_d N_A_193_241#_M1006_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.157545 PD=1.06 PS=1.24406 NRD=6.48 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1006_d N_A_193_241#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1628 PD=1.06 PS=1.18 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1021 N_X_M1021_d N_A_193_241#_M1021_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1628 PD=1.02 PS=1.18 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75001.8
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1021_d N_A_193_241#_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.249804 PD=1.02 PS=1.56043 NRD=0 NRS=27.156 M=1 R=4.93333
+ SA=75002.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_709_119#_M1001_d N_S_M1001_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.216046 PD=0.99 PS=1.34957 NRD=0 NRS=73.116 M=1 R=4.26667
+ SA=75002.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1024 N_A_709_119#_M1001_d N_S_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1568 PD=0.99 PS=1.13 NRD=13.116 NRS=13.116 M=1 R=4.26667
+ SA=75003.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_937_119#_M1003_d N_A_27_368#_M1003_g N_VGND_M1024_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1568 PD=0.92 PS=1.13 NRD=0 NRS=26.244 M=1 R=4.26667
+ SA=75003.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 N_A_937_119#_M1003_d N_A_27_368#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.3692 PD=0.92 PS=2.64 NRD=0 NRS=97.848 M=1 R=4.26667
+ SA=75004.2 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1017 N_A_937_119#_M1017_d N_A0_M1017_g N_A_193_241#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.096 AS=0.4992 PD=0.94 PS=2.84 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_937_119#_M1017_d N_A0_M1022_g N_A_193_241#_M1022_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.096 AS=0.1056 PD=0.94 PS=0.97 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75001.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1014 N_A_193_241#_M1022_s N_A1_M1014_g N_A_709_119#_M1014_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1056 AS=0.0992 PD=0.97 PS=0.95 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_193_241#_M1025_d N_A1_M1025_g N_A_709_119#_M1014_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2112 AS=0.0992 PD=1.94 PS=0.95 NRD=7.488 NRS=5.616 M=1 R=4.26667
+ SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_S_M1009_g N_A_27_368#_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.191226 AS=0.28 PD=1.40566 PS=2.56 NRD=17.7103 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90004.6 A=0.18 P=2.36 MULT=1
MM1000 N_X_M1000_d N_A_193_241#_M1000_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1.12
+ AD=0.27395 AS=0.214174 PD=1.75 PS=1.57434 NRD=33.3324 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90004 A=0.2016 P=2.6 MULT=1
MM1004 N_X_M1000_d N_A_193_241#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.27395 AS=0.273225 PD=1.75 PS=1.745 NRD=14.9326 NRS=14.9326 M=1 R=6.22222
+ SA=90001.3 SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1019 N_X_M1019_d N_A_193_241#_M1019_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.258725 AS=0.273225 PD=1.645 PS=1.745 NRD=2.6201 NRS=33.2339 M=1 R=6.22222
+ SA=90001.9 SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1020 N_X_M1019_d N_A_193_241#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.258725 AS=0.276949 PD=1.645 PS=1.84377 NRD=2.6201 NRS=33.8052 M=1
+ R=6.22222 SA=90002.5 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1010 N_A_725_391#_M1010_d N_S_M1010_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.247276 PD=1.27 PS=1.64623 NRD=0 NRS=37.8634 M=1 R=5.55556
+ SA=90003.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1013 N_A_725_391#_M1010_d N_S_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.23885 PD=1.27 PS=1.57 NRD=0 NRS=16.7253 M=1 R=5.55556 SA=90003.6
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1015 N_A_939_391#_M1015_d N_A_27_368#_M1015_g N_VPWR_M1013_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.23885 PD=1.27 PS=1.57 NRD=0 NRS=16.7253 M=1 R=5.55556
+ SA=90004.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1018 N_A_939_391#_M1015_d N_A_27_368#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.4027 PD=1.27 PS=2.99 NRD=0 NRS=16.7253 M=1 R=5.55556
+ SA=90004.7 SB=90000.3 A=0.18 P=2.36 MULT=1
MM1011 N_A_725_391#_M1011_d N_A0_M1011_g N_A_193_241#_M1011_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.315 PD=1.27 PS=2.63 NRD=0 NRS=2.9353 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1016 N_A_725_391#_M1011_d N_A0_M1016_g N_A_193_241#_M1016_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.14 PD=1.27 PS=1.28 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_A_939_391#_M1005_d N_A1_M1005_g N_A_193_241#_M1016_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.14 PD=1.27 PS=1.28 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1008 N_A_939_391#_M1005_d N_A1_M1008_g N_A_193_241#_M1008_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.33 PD=1.27 PS=2.66 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX26_noxref VNB VPB NWDIODE A=17.0422 P=22.14
*
.include "sky130_fd_sc_ms__mux2_4.pxi.spice"
*
.ends
*
*

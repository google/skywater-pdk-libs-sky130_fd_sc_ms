* File: sky130_fd_sc_ms__o2111a_2.spice
* Created: Fri Aug 28 17:51:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2111a_2.pex.spice"
.subckt sky130_fd_sc_ms__o2111a_2  VNB VPB A1 A2 B1 C1 D1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D1	D1
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_54_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2627 PD=1.16 PS=2.19 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1003 N_A_54_74#_M1003_d N_A2_M1003_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=11.34 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1013 A_369_74# N_B1_M1013_g N_A_54_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=16.212 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1005 A_461_74# N_C1_M1005_g A_369_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1147 PD=1.16 PS=1.05 NRD=25.128 NRS=16.212 M=1 R=4.93333 SA=75001.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1008 N_A_239_368#_M1008_d N_D1_M1008_g A_461_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_239_368#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_239_368#_M1009_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.222 AS=0.1036 PD=2.08 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 A_155_368# N_A1_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90003.8
+ A=0.18 P=2.36 MULT=1
MM1011 N_A_239_368#_M1011_d N_A2_M1011_g A_155_368# VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.12 PD=1.39 PS=1.24 NRD=22.6353 NRS=12.7853 M=1 R=5.55556
+ SA=90000.6 SB=90003.4 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_B1_M1010_g N_A_239_368#_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.23 AS=0.195 PD=1.46 PS=1.39 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90001.2
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1002 N_A_239_368#_M1002_d N_C1_M1002_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.23 PD=1.32 PS=1.46 NRD=0 NRS=26.5753 M=1 R=5.55556 SA=90001.8
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_D1_M1000_g N_A_239_368#_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.391509 AS=0.16 PD=1.81132 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90002.3 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1000_d N_A_239_368#_M1001_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.438491 AS=0.1512 PD=2.02868 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90003 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1012_d N_A_239_368#_M1012_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__o2111a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sdfrtp_1.spice
* Created: Fri Aug 28 18:12:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfrtp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfrtp_1  VNB VPB SCE D SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1034 N_VGND_M1034_d N_SCE_M1034_g N_A_27_88#_M1034_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 noxref_25 N_A_27_88#_M1008_g N_noxref_24_M1008_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_303_464#_M1009_d N_D_M1009_g noxref_25 VNB NLOWVT L=0.15 W=0.42
+ AD=0.13125 AS=0.0504 PD=1.045 PS=0.66 NRD=98.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1025 noxref_26 N_SCE_M1025_g N_A_303_464#_M1009_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.13125 PD=0.66 PS=1.045 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 N_noxref_24_M1015_d N_SCD_M1015_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0651 AS=0.0504 PD=0.73 PS=0.66 NRD=2.856 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_RESET_B_M1036_g N_noxref_24_M1015_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0651 PD=1.41 PS=0.73 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_CLK_M1029_g N_A_835_93#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.16425 AS=0.28265 PD=1.27 PS=2.43 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75000.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1032 N_A_1037_387#_M1032_d N_A_835_93#_M1032_g N_VGND_M1029_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1961 AS=0.16425 PD=2.01 PS=1.27 NRD=0 NRS=10.536 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_1234_119#_M1035_d N_A_835_93#_M1035_g N_A_303_464#_M1035_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1001 A_1320_119# N_A_1037_387#_M1001_g N_A_1234_119#_M1035_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.04935 AS=0.0588 PD=0.655 PS=0.7 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1020 A_1397_119# N_A_1367_93#_M1020_g A_1320_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.04935 PD=0.66 PS=0.655 NRD=18.564 NRS=17.856 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_RESET_B_M1012_g A_1397_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.211634 AS=0.0504 PD=1.27189 PS=0.66 NRD=128.244 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_1367_93#_M1033_d N_A_1234_119#_M1033_g N_VGND_M1012_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.322491 PD=0.92 PS=1.93811 NRD=0 NRS=84.156 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1006 N_A_1745_74#_M1006_d N_A_1037_387#_M1006_g N_A_1367_93#_M1033_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.282989 AS=0.0896 PD=1.96226 PS=0.92 NRD=132.18 NRS=0
+ M=1 R=4.26667 SA=75002.1 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1004 A_1972_74# N_A_835_93#_M1004_g N_A_1745_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.185711 PD=0.63 PS=1.28774 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75003 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_1997_272#_M1003_g A_1972_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1038 A_2135_74# N_RESET_B_M1038_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.06405 PD=0.63 PS=0.725 NRD=14.28 NRS=7.14 M=1 R=2.8 SA=75003.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_1997_272#_M1022_d N_A_1745_74#_M1022_g A_2135_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_A_2402_424#_M1027_d N_A_1745_74#_M1027_g N_VGND_M1027_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.1595 PD=1.67 PS=1.68 NRD=0 NRS=1.08 M=1
+ R=3.66667 SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1007 N_Q_M1007_d N_A_2402_424#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_SCE_M1005_g N_A_27_88#_M1005_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.1792 PD=0.96 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90003.3 A=0.1152 P=1.64 MULT=1
MM1002 A_219_464# N_SCE_M1002_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90002.8 A=0.1152 P=1.64 MULT=1
MM1013 N_A_303_464#_M1013_d N_D_M1013_g A_219_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.3136 AS=0.0768 PD=1.62 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.1
+ SB=90002.4 A=0.1152 P=1.64 MULT=1
MM1016 A_535_464# N_A_27_88#_M1016_g N_A_303_464#_M1013_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.3136 PD=0.91 PS=1.62 NRD=24.625 NRS=0 M=1 R=3.55556
+ SA=90002.3 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1019 N_VPWR_M1019_d N_SCD_M1019_g A_535_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1248 AS=0.0864 PD=1.03 PS=0.91 NRD=0 NRS=24.625 M=1 R=3.55556 SA=90002.7
+ SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1023 N_A_303_464#_M1023_d N_RESET_B_M1023_g N_VPWR_M1019_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.1248 PD=1.84 PS=1.03 NRD=0 NRS=35.3812 M=1 R=3.55556
+ SA=90003.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1018 N_VPWR_M1018_d N_CLK_M1018_g N_A_835_93#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1030 N_A_1037_387#_M1030_d N_A_835_93#_M1030_g N_VPWR_M1018_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_1234_119#_M1000_d N_A_1037_387#_M1000_g N_A_303_464#_M1000_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.07 AS=0.1176 PD=0.765 PS=1.4 NRD=23.443 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1017 A_1346_461# N_A_835_93#_M1017_g N_A_1234_119#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.07 PD=0.66 PS=0.765 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1028 N_VPWR_M1028_d N_A_1367_93#_M1028_g A_1346_461# VPB PSHORT L=0.18 W=0.42
+ AD=0.129587 AS=0.0504 PD=1.11 PS=0.66 NRD=118.909 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1010 N_A_1234_119#_M1010_d N_RESET_B_M1010_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.129587 PD=1.4 PS=1.11 NRD=0 NRS=118.909 M=1 R=2.33333
+ SA=90001.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1026 N_A_1367_93#_M1026_d N_A_1234_119#_M1026_g N_VPWR_M1026_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1031 N_A_1745_74#_M1031_d N_A_835_93#_M1031_g N_A_1367_93#_M1026_d VPB PSHORT
+ L=0.18 W=1 AD=0.296954 AS=0.135 PD=2.52113 PS=1.27 NRD=37.43 NRS=0 M=1
+ R=5.55556 SA=90000.6 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1014 A_1996_508# N_A_1037_387#_M1014_g N_A_1745_74#_M1031_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.124721 PD=0.66 PS=1.05887 NRD=30.4759 NRS=46.886 M=1
+ R=2.33333 SA=90000.9 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1037 N_VPWR_M1037_d N_A_1997_272#_M1037_g A_1996_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.08295 AS=0.0504 PD=0.815 PS=0.66 NRD=14.0658 NRS=30.4759 M=1 R=2.33333
+ SA=90001.3 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1021 N_A_1997_272#_M1021_d N_RESET_B_M1021_g N_VPWR_M1037_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.08295 PD=0.69 PS=0.815 NRD=0 NRS=39.8531 M=1 R=2.33333
+ SA=90001.9 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_1745_74#_M1024_g N_A_1997_272#_M1021_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1029 AS=0.0567 PD=0.83 PS=0.69 NRD=37.5088 NRS=0 M=1
+ R=2.33333 SA=90002.3 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1039 N_A_2402_424#_M1039_d N_A_1745_74#_M1039_g N_VPWR_M1024_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.2058 PD=2.24 PS=1.66 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90001.6 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1011 N_Q_M1011_d N_A_2402_424#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.4373 P=31.76
c_154 VNB 0 1.61901e-19 $X=0 $Y=0
c_2103 A_1346_461# 0 1.83551e-19 $X=6.73 $Y=2.305
c_2105 A_1996_508# 0 1.04043e-19 $X=9.98 $Y=2.54
*
.include "sky130_fd_sc_ms__sdfrtp_1.pxi.spice"
*
.ends
*
*

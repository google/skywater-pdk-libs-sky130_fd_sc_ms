* File: sky130_fd_sc_ms__sdfbbn_1.pex.spice
* Created: Wed Sep  2 12:29:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%SCD 2 5 9 11 12 15 16
c32 5 0 8.66027e-20 $X=0.505 $Y=2.64
r33 15 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.37
+ $X2=0.407 $Y2=1.205
r34 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.37 $X2=0.385 $Y2=1.37
r35 12 16 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.385 $Y2=1.54
r36 9 17 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.52 $Y=0.805 $X2=0.52
+ $Y2=1.205
r37 5 11 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=0.505 $Y=2.64
+ $X2=0.505 $Y2=1.875
r38 2 11 42.8297 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.407 $Y=1.688
+ $X2=0.407 $Y2=1.875
r39 1 15 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.392
+ $X2=0.407 $Y2=1.37
r40 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.407 $Y=1.392
+ $X2=0.407 $Y2=1.688
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%D 1 3 8 10 11 17
c59 11 0 1.09459e-19 $X=1.68 $Y=1.665
r60 15 17 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.45 $Y=1.645 $X2=1.65
+ $Y2=1.645
r61 13 15 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=1.42 $Y=1.645 $X2=1.45
+ $Y2=1.645
r62 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.645 $X2=1.65 $Y2=1.645
r63 6 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.48
+ $X2=1.45 $Y2=1.645
r64 6 8 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.45 $Y=1.48 $X2=1.45
+ $Y2=0.805
r65 4 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.81
+ $X2=1.42 $Y2=1.645
r66 4 10 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.42 $Y=1.81
+ $X2=1.42 $Y2=2.115
r67 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.405 $Y=2.205
+ $X2=1.405 $Y2=2.115
r68 1 3 116.483 $w=1.8e-07 $l=4.35e-07 $layer=POLY_cond $X=1.405 $Y=2.205
+ $X2=1.405 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_353_93# 1 2 7 9 10 12 14 16 19 23 26 29
+ 37 40 43 44
c90 23 0 5.47294e-20 $X=2.13 $Y=2.125
c91 19 0 1.66897e-19 $X=2.13 $Y=1.165
r92 43 44 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=2.465
+ $X2=3.07 $Y2=2.3
r93 39 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.895 $Y=1.645
+ $X2=2.975 $Y2=1.645
r94 36 39 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.675 $Y=1.645
+ $X2=2.895 $Y2=1.645
r95 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.645 $X2=2.675 $Y2=1.645
r96 31 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=1.81
+ $X2=2.975 $Y2=1.645
r97 31 44 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.975 $Y=1.81
+ $X2=2.975 $Y2=2.3
r98 27 39 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=1.48
+ $X2=2.895 $Y2=1.645
r99 27 29 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.895 $Y=1.48
+ $X2=2.895 $Y2=0.815
r100 25 37 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=2.205 $Y=1.645
+ $X2=2.675 $Y2=1.645
r101 25 26 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=1.645
+ $X2=2.13 $Y2=1.645
r102 17 19 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.84 $Y=1.165
+ $X2=2.13 $Y2=1.165
r103 16 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=2.05
+ $X2=2.13 $Y2=2.125
r104 15 26 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=1.645
r105 15 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=2.05
r106 14 26 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.48
+ $X2=2.13 $Y2=1.645
r107 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.24
+ $X2=2.13 $Y2=1.165
r108 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.24
+ $X2=2.13 $Y2=1.48
r109 10 23 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.855 $Y=2.125
+ $X2=2.13 $Y2=2.125
r110 10 12 117.822 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=1.855 $Y=2.2
+ $X2=1.855 $Y2=2.64
r111 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.09
+ $X2=1.84 $Y2=1.165
r112 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.84 $Y=1.09 $X2=1.84
+ $Y2=0.805
r113 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.95
+ $Y=2.32 $X2=3.085 $Y2=2.465
r114 1 29 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.595 $X2=2.895 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%SCE 4 7 9 10 14 15 16 17 19 21 24 25 28 30
+ 33
c103 33 0 8.1544e-20 $X=0.97 $Y=1.37
c104 4 0 2.95072e-20 $X=0.91 $Y=0.805
r105 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.97
+ $Y=1.37 $X2=0.97 $Y2=1.37
r106 30 34 4.10594 $w=6.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.54
+ $X2=0.97 $Y2=1.54
r107 24 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.97 $Y=1.71
+ $X2=0.97 $Y2=1.37
r108 24 25 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.71
+ $X2=0.97 $Y2=1.875
r109 23 33 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.205
+ $X2=0.97 $Y2=1.37
r110 21 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.155 $Y=2.05
+ $X2=3.155 $Y2=2.125
r111 20 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.155 $Y=1.24
+ $X2=3.155 $Y2=2.05
r112 17 28 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.86 $Y=2.125
+ $X2=3.155 $Y2=2.125
r113 17 19 117.822 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=2.86 $Y=2.2
+ $X2=2.86 $Y2=2.64
r114 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.08 $Y=1.165
+ $X2=3.155 $Y2=1.24
r115 15 16 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.08 $Y=1.165
+ $X2=2.755 $Y2=1.165
r116 12 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.68 $Y=1.09
+ $X2=2.755 $Y2=1.165
r117 12 14 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.68 $Y=1.09
+ $X2=2.68 $Y2=0.805
r118 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.68 $Y=0.255
+ $X2=2.68 $Y2=0.805
r119 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.605 $Y=0.18
+ $X2=2.68 $Y2=0.255
r120 9 10 830.681 $w=1.5e-07 $l=1.62e-06 $layer=POLY_cond $X=2.605 $Y=0.18
+ $X2=0.985 $Y2=0.18
r121 7 25 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=0.985 $Y=2.64
+ $X2=0.985 $Y2=1.875
r122 4 23 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.91 $Y=0.805 $X2=0.91
+ $Y2=1.205
r123 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.985 $Y2=0.18
r124 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.91 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%CLK_N 3 7 9 13 16
c42 7 0 1.13863e-19 $X=3.87 $Y=2.4
c43 3 0 1.60531e-19 $X=3.67 $Y=0.78
r44 15 16 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=3.67 $Y=1.515 $X2=3.87
+ $Y2=1.515
r45 12 15 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.635 $Y=1.515
+ $X2=3.67 $Y2=1.515
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.635
+ $Y=1.515 $X2=3.635 $Y2=1.515
r47 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.635 $Y=1.665
+ $X2=3.635 $Y2=1.515
r48 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.87 $Y=1.68
+ $X2=3.87 $Y2=1.515
r49 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.87 $Y=1.68 $X2=3.87
+ $Y2=2.4
r50 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.35
+ $X2=3.67 $Y2=1.515
r51 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.67 $Y=1.35 $X2=3.67
+ $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_977_243# 1 2 3 12 13 14 16 20 24 28 30 31
+ 37 40 42 43 46 48 49 53 57 58 61 62 68 69 71 74 78
c201 61 0 7.4272e-20 $X=5.05 $Y=2.13
c202 58 0 1.73041e-20 $X=9.365 $Y=1.795
c203 57 0 1.73394e-19 $X=9.365 $Y=1.795
c204 31 0 1.49471e-19 $X=5.05 $Y=1.755
c205 28 0 1.99515e-19 $X=9.44 $Y=2.54
c206 20 0 8.96875e-20 $X=5.68 $Y=0.805
c207 14 0 1.01056e-19 $X=5.33 $Y=2.295
r208 76 78 3.904 $w=2.5e-07 $l=8e-08 $layer=LI1_cond $X=8.662 $Y=2.395 $X2=8.662
+ $Y2=2.475
r209 75 76 8.784 $w=2.5e-07 $l=1.8e-07 $layer=LI1_cond $X=8.662 $Y=2.215
+ $X2=8.662 $Y2=2.395
r210 71 73 10.5575 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.925 $Y=0.855
+ $X2=7.925 $Y2=1.08
r211 67 69 8.89604 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=7.335 $Y=2.862
+ $X2=7.505 $Y2=2.862
r212 67 68 15.404 $w=4.23e-07 $l=4.1e-07 $layer=LI1_cond $X=7.335 $Y=2.862
+ $X2=6.925 $Y2=2.862
r213 61 64 3.47907 $w=2.63e-07 $l=8e-08 $layer=LI1_cond $X=5.082 $Y=2.13
+ $X2=5.082 $Y2=2.21
r214 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=2.13 $X2=5.05 $Y2=2.13
r215 58 82 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.365 $Y=1.795
+ $X2=9.365 $Y2=1.96
r216 58 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.365 $Y=1.795
+ $X2=9.365 $Y2=1.63
r217 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.365
+ $Y=1.795 $X2=9.365 $Y2=1.795
r218 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.365 $Y=2.13
+ $X2=9.365 $Y2=1.795
r219 54 75 2.99516 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.83 $Y=2.215
+ $X2=8.662 $Y2=2.215
r220 53 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.2 $Y=2.215
+ $X2=9.365 $Y2=2.13
r221 53 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.2 $Y=2.215
+ $X2=8.83 $Y2=2.215
r222 50 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=2.395
+ $X2=7.845 $Y2=2.395
r223 49 76 2.99516 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=8.495 $Y=2.395
+ $X2=8.662 $Y2=2.395
r224 49 50 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=8.495 $Y=2.395
+ $X2=7.93 $Y2=2.395
r225 47 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=2.48
+ $X2=7.845 $Y2=2.395
r226 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.845 $Y=2.48
+ $X2=7.845 $Y2=2.65
r227 46 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=2.31
+ $X2=7.845 $Y2=2.395
r228 46 73 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=7.845 $Y=2.31
+ $X2=7.845 $Y2=1.08
r229 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.76 $Y=2.735
+ $X2=7.845 $Y2=2.65
r230 43 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.76 $Y=2.735
+ $X2=7.505 $Y2=2.735
r231 42 68 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=5.61 $Y=2.99
+ $X2=6.925 $Y2=2.99
r232 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.525 $Y=2.905
+ $X2=5.61 $Y2=2.99
r233 39 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.525 $Y=2.295
+ $X2=5.525 $Y2=2.905
r234 38 64 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.215 $Y=2.21
+ $X2=5.082 $Y2=2.21
r235 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.44 $Y=2.21
+ $X2=5.525 $Y2=2.295
r236 37 38 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.44 $Y=2.21
+ $X2=5.215 $Y2=2.21
r237 33 62 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.05 $Y=2.145
+ $X2=5.05 $Y2=2.13
r238 30 62 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.05 $Y=1.92
+ $X2=5.05 $Y2=2.13
r239 30 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.92
+ $X2=5.05 $Y2=1.755
r240 28 82 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=9.44 $Y=2.54
+ $X2=9.44 $Y2=1.96
r241 24 81 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.305 $Y=0.87
+ $X2=9.305 $Y2=1.63
r242 18 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.68 $Y=1.215
+ $X2=5.68 $Y2=0.805
r243 14 33 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.33 $Y=2.22
+ $X2=5.05 $Y2=2.22
r244 14 16 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=5.33 $Y=2.295
+ $X2=5.33 $Y2=2.695
r245 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=1.29
+ $X2=5.68 $Y2=1.215
r246 12 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.605 $Y=1.29
+ $X2=5.035 $Y2=1.29
r247 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.96 $Y=1.365
+ $X2=5.035 $Y2=1.29
r248 10 31 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.96 $Y=1.365
+ $X2=4.96 $Y2=1.755
r249 3 78 300 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_PDIFF $count=2 $X=8.525
+ $Y=2.12 $X2=8.66 $Y2=2.475
r250 2 67 600 $w=1.7e-07 $l=8.00125e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=2.12 $X2=7.335 $Y2=2.78
r251 1 71 182 $w=1.7e-07 $l=3.60555e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.595 $X2=7.925 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_867_82# 1 2 9 13 17 21 23 26 28 31 36 38
+ 39 45 46 47 50 51 57 58 61 68 78 79
c221 79 0 1.01056e-19 $X=5.755 $Y=1.727
c222 68 0 3.86106e-20 $X=9.905 $Y=1.775
c223 26 0 1.13863e-19 $X=4.58 $Y=2.04
c224 23 0 1.60531e-19 $X=4.61 $Y=1.045
c225 21 0 3.18534e-20 $X=10.745 $Y=0.805
c226 13 0 2.29882e-20 $X=6.47 $Y=0.805
r227 68 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.905 $Y=1.775
+ $X2=9.905 $Y2=1.94
r228 61 63 20.6118 $w=3.04e-07 $l=1.3e-07 $layer=POLY_cond $X=5.59 $Y=1.74
+ $X2=5.72 $Y2=1.74
r229 58 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.905
+ $Y=1.775 $X2=9.905 $Y2=1.775
r230 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r231 54 79 8.65129 $w=3.53e-07 $l=2.35e-07 $layer=LI1_cond $X=5.52 $Y=1.727
+ $X2=5.755 $Y2=1.727
r232 54 78 6.8759 $w=3.53e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.727
+ $X2=5.405 $Y2=1.727
r233 54 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.74 $X2=5.59 $Y2=1.74
r234 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r235 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r236 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r237 50 51 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=5.665 $Y2=1.665
r238 49 58 3.67446 $w=3.43e-07 $l=1.1e-07 $layer=LI1_cond $X=9.897 $Y=1.555
+ $X2=9.897 $Y2=1.665
r239 47 79 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=6.38 $Y=1.675
+ $X2=5.755 $Y2=1.675
r240 46 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.545 $Y=1.635
+ $X2=6.545 $Y2=1.47
r241 45 47 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.545 $Y=1.635
+ $X2=6.38 $Y2=1.635
r242 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.545
+ $Y=1.635 $X2=6.545 $Y2=1.635
r243 41 43 16.9064 $w=2.67e-07 $l=3.7e-07 $layer=LI1_cond $X=4.61 $Y=1.635
+ $X2=4.61 $Y2=2.005
r244 39 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.245
r245 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.835
+ $Y=1.41 $X2=10.835 $Y2=1.41
r246 36 49 6.87075 $w=2.95e-07 $l=2.35654e-07 $layer=LI1_cond $X=10.07 $Y=1.407
+ $X2=9.897 $Y2=1.555
r247 36 38 29.8854 $w=2.93e-07 $l=7.65e-07 $layer=LI1_cond $X=10.07 $Y=1.407
+ $X2=10.835 $Y2=1.407
r248 33 41 3.37873 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.79 $Y=1.635
+ $X2=4.61 $Y2=1.635
r249 33 78 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.79 $Y=1.635
+ $X2=5.405 $Y2=1.635
r250 31 41 5.1848 $w=2.67e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.7 $Y=1.55
+ $X2=4.61 $Y2=1.635
r251 30 31 23.4141 $w=1.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.7 $Y=1.17 $X2=4.7
+ $Y2=1.55
r252 26 43 2.41973 $w=4e-07 $l=4.7697e-08 $layer=LI1_cond $X=4.58 $Y=2.04
+ $X2=4.61 $Y2=2.005
r253 26 28 22.3286 $w=3.98e-07 $l=7.75e-07 $layer=LI1_cond $X=4.58 $Y=2.04
+ $X2=4.58 $Y2=2.815
r254 23 30 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.61 $Y=1.045
+ $X2=4.7 $Y2=1.17
r255 23 25 2.928 $w=2.5e-07 $l=6e-08 $layer=LI1_cond $X=4.61 $Y=1.045 $X2=4.55
+ $Y2=1.045
r256 21 73 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.745 $Y=0.805
+ $X2=10.745 $Y2=1.245
r257 17 71 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=9.83 $Y=2.54 $X2=9.83
+ $Y2=1.94
r258 13 65 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=6.47 $Y=0.805
+ $X2=6.47 $Y2=1.47
r259 7 63 15.0262 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.72 $Y=1.905
+ $X2=5.72 $Y2=1.74
r260 7 9 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=5.72 $Y=1.905
+ $X2=5.72 $Y2=2.695
r261 2 43 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.84 $X2=4.545 $Y2=2.005
r262 2 28 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.84 $X2=4.545 $Y2=2.815
r263 1 25 182 $w=1.7e-07 $l=6.94226e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.41 $X2=4.55 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_1162_497# 1 2 7 8 11 13 15 17 20 22 24 25
+ 29 30 31
c90 25 0 8.96875e-20 $X=6.42 $Y=1.215
c91 8 0 2.87426e-20 $X=7.25 $Y=1.33
r92 31 33 19.511 $w=2.72e-07 $l=4.35e-07 $layer=LI1_cond $X=6.03 $Y=2.055
+ $X2=6.03 $Y2=2.49
r93 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.085
+ $Y=1.42 $X2=7.085 $Y2=1.42
r94 27 29 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=7.085 $Y=1.97
+ $X2=7.085 $Y2=1.42
r95 26 29 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.085 $Y=1.3
+ $X2=7.085 $Y2=1.42
r96 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.92 $Y=1.215
+ $X2=7.085 $Y2=1.3
r97 24 25 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.92 $Y=1.215 $X2=6.42
+ $Y2=1.215
r98 23 31 3.48705 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=2.055
+ $X2=6.03 $Y2=2.055
r99 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.92 $Y=2.055
+ $X2=7.085 $Y2=1.97
r100 22 23 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.92 $Y=2.055
+ $X2=6.195 $Y2=2.055
r101 18 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.295 $Y=1.13
+ $X2=6.42 $Y2=1.215
r102 18 20 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=6.295 $Y=1.13
+ $X2=6.295 $Y2=0.815
r103 16 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.085 $Y=1.405
+ $X2=7.085 $Y2=1.42
r104 13 17 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=7.61 $Y=1.255
+ $X2=7.58 $Y2=1.33
r105 13 15 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.61 $Y=1.255
+ $X2=7.61 $Y2=0.87
r106 9 17 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.565 $Y=1.405
+ $X2=7.58 $Y2=1.33
r107 9 11 441.185 $w=1.8e-07 $l=1.135e-06 $layer=POLY_cond $X=7.565 $Y=1.405
+ $X2=7.565 $Y2=2.54
r108 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.25 $Y=1.33
+ $X2=7.085 $Y2=1.405
r109 7 17 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=7.475 $Y=1.33
+ $X2=7.58 $Y2=1.33
r110 7 8 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.475 $Y=1.33
+ $X2=7.25 $Y2=1.33
r111 2 33 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=2.485 $X2=6.03 $Y2=2.49
r112 1 20 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=6.115
+ $Y=0.595 $X2=6.255 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_1579_258# 1 2 9 13 15 17 18 20 22 25 26
+ 27 28 31 32 33 34 37 40 42 44 46 50 52 56 63
c192 56 0 9.562e-20 $X=12.365 $Y=1.215
c193 46 0 1.37209e-19 $X=8.265 $Y=1.375
c194 42 0 7.63376e-20 $X=13.78 $Y=1.915
c195 20 0 2.82259e-19 $X=12.47 $Y=2.46
c196 13 0 4.35224e-20 $X=8.14 $Y=0.87
c197 9 0 3.27703e-19 $X=7.985 $Y=2.54
r198 65 67 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=7.985 $Y=1.455
+ $X2=8.14 $Y2=1.455
r199 62 63 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=13.695 $Y=1.215
+ $X2=13.82 $Y2=1.215
r200 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.365
+ $Y=1.385 $X2=12.365 $Y2=1.385
r201 56 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.365 $Y=1.215
+ $X2=12.365 $Y2=1.385
r202 52 54 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.835 $Y=0.45
+ $X2=10.835 $Y2=0.665
r203 50 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=8.265 $Y=1.455
+ $X2=8.14 $Y2=1.455
r204 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.265
+ $Y=1.455 $X2=8.265 $Y2=1.455
r205 46 49 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.265 $Y=1.375
+ $X2=8.265 $Y2=1.455
r206 42 44 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=13.78 $Y=1.915
+ $X2=13.87 $Y2=1.915
r207 38 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.82 $Y=1.13
+ $X2=13.82 $Y2=1.215
r208 38 40 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=13.82 $Y=1.13
+ $X2=13.82 $Y2=0.9
r209 37 42 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.695 $Y=1.79
+ $X2=13.78 $Y2=1.915
r210 36 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.695 $Y=1.3
+ $X2=13.695 $Y2=1.215
r211 36 37 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=13.695 $Y=1.3
+ $X2=13.695 $Y2=1.79
r212 35 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.53 $Y=1.215
+ $X2=12.365 $Y2=1.215
r213 34 62 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=13.61 $Y=1.215
+ $X2=13.695 $Y2=1.215
r214 34 35 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=13.61 $Y=1.215
+ $X2=12.53 $Y2=1.215
r215 32 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.2 $Y=1.215
+ $X2=12.365 $Y2=1.215
r216 32 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=12.2 $Y=1.215
+ $X2=11.68 $Y2=1.215
r217 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.595 $Y=1.13
+ $X2=11.68 $Y2=1.215
r218 30 31 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.595 $Y=0.75
+ $X2=11.595 $Y2=1.13
r219 29 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.665
+ $X2=10.835 $Y2=0.665
r220 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.51 $Y=0.665
+ $X2=11.595 $Y2=0.75
r221 28 29 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.51 $Y=0.665
+ $X2=10.92 $Y2=0.665
r222 26 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.45
+ $X2=10.835 $Y2=0.45
r223 26 27 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=10.75 $Y=0.45
+ $X2=9.555 $Y2=0.45
r224 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.47 $Y=0.535
+ $X2=9.555 $Y2=0.45
r225 24 25 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.47 $Y=0.535
+ $X2=9.47 $Y2=1.29
r226 23 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.43 $Y=1.375
+ $X2=8.265 $Y2=1.375
r227 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.385 $Y=1.375
+ $X2=9.47 $Y2=1.29
r228 22 23 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=9.385 $Y=1.375
+ $X2=8.43 $Y2=1.375
r229 18 60 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=12.47 $Y=1.55
+ $X2=12.38 $Y2=1.385
r230 18 20 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=12.47 $Y=1.55
+ $X2=12.47 $Y2=2.46
r231 15 60 38.7084 $w=3.43e-07 $l=1.94808e-07 $layer=POLY_cond $X=12.315 $Y=1.22
+ $X2=12.38 $Y2=1.385
r232 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.315 $Y=1.22
+ $X2=12.315 $Y2=0.74
r233 11 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.14 $Y=1.29
+ $X2=8.14 $Y2=1.455
r234 11 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=8.14 $Y=1.29
+ $X2=8.14 $Y2=0.87
r235 7 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.985 $Y=1.62
+ $X2=7.985 $Y2=1.455
r236 7 9 357.613 $w=1.8e-07 $l=9.2e-07 $layer=POLY_cond $X=7.985 $Y=1.62
+ $X2=7.985 $Y2=2.54
r237 2 44 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=13.6
+ $Y=1.73 $X2=13.87 $Y2=1.875
r238 1 40 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=13.675
+ $Y=0.69 $X2=13.82 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%SET_B 1 3 6 10 14 16 17 20 22 25 30 31
c135 25 0 1.37209e-19 $X=8.745 $Y=1.82
c136 22 0 1.50853e-19 $X=11.76 $Y=2.035
c137 20 0 1.79798e-19 $X=8.4 $Y=2.035
c138 16 0 4.36058e-20 $X=11.615 $Y=2.035
c139 10 0 9.77748e-20 $X=11.85 $Y=2.46
c140 6 0 1.76028e-19 $X=8.745 $Y=0.87
r141 31 37 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=11.795 $Y=1.635
+ $X2=11.795 $Y2=2.035
r142 30 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.795 $Y=1.635
+ $X2=11.795 $Y2=1.8
r143 30 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.795 $Y=1.635
+ $X2=11.795 $Y2=1.47
r144 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.795
+ $Y=1.635 $X2=11.795 $Y2=1.635
r145 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.825
+ $Y=1.795 $X2=8.825 $Y2=1.795
r146 25 27 14.4419 $w=2.67e-07 $l=8e-08 $layer=POLY_cond $X=8.745 $Y=1.82
+ $X2=8.825 $Y2=1.82
r147 22 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=2.035
+ $X2=11.76 $Y2=2.035
r148 20 28 17.4579 $w=2.97e-07 $l=4.25e-07 $layer=LI1_cond $X=8.4 $Y=1.885
+ $X2=8.825 $Y2=1.885
r149 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r150 17 19 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=2.035
+ $X2=8.4 $Y2=2.035
r151 16 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=2.035
+ $X2=11.76 $Y2=2.035
r152 16 17 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=11.615 $Y=2.035
+ $X2=8.545 $Y2=2.035
r153 14 32 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=11.885 $Y=0.74
+ $X2=11.885 $Y2=1.47
r154 10 33 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=11.85 $Y=2.46
+ $X2=11.85 $Y2=1.8
r155 4 25 16.2448 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.745 $Y=1.63
+ $X2=8.745 $Y2=1.82
r156 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.745 $Y=1.63
+ $X2=8.745 $Y2=0.87
r157 1 25 55.9625 $w=2.67e-07 $l=3.937e-07 $layer=POLY_cond $X=8.435 $Y=2.01
+ $X2=8.745 $Y2=1.82
r158 1 3 141.922 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=8.435 $Y=2.01
+ $X2=8.435 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_662_82# 1 2 10 13 15 16 20 22 23 25 27 31
+ 32 33 34 36 40 42 47 48 52 54 56 59 61 67 68
c186 68 0 1.27434e-19 $X=4.335 $Y=1.505
c187 67 0 1.49471e-19 $X=4.335 $Y=1.505
c188 40 0 4.28297e-20 $X=6.04 $Y=0.18
c189 34 0 3.8609e-20 $X=10.365 $Y=2.27
c190 32 0 1.94296e-19 $X=10.28 $Y=1.295
c191 13 0 7.4272e-20 $X=4.32 $Y=2.4
r192 68 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.505
+ $X2=4.335 $Y2=1.67
r193 68 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.505
+ $X2=4.335 $Y2=1.34
r194 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.335
+ $Y=1.505 $X2=4.335 $Y2=1.505
r195 64 67 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.055 $Y=1.505
+ $X2=4.335 $Y2=1.505
r196 60 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=1.67
+ $X2=4.055 $Y2=1.505
r197 60 61 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.055 $Y=1.67
+ $X2=4.055 $Y2=1.95
r198 59 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=1.34
+ $X2=4.055 $Y2=1.505
r199 58 59 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.055 $Y=1.17
+ $X2=4.055 $Y2=1.34
r200 57 63 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.73 $Y=2.035
+ $X2=3.605 $Y2=2.035
r201 56 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.97 $Y=2.035
+ $X2=4.055 $Y2=1.95
r202 56 57 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.97 $Y=2.035
+ $X2=3.73 $Y2=2.035
r203 52 63 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=2.12
+ $X2=3.605 $Y2=2.035
r204 52 54 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.605 $Y=2.12
+ $X2=3.605 $Y2=2.815
r205 48 58 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.97 $Y=1.045
+ $X2=4.055 $Y2=1.17
r206 48 50 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=3.97 $Y=1.045
+ $X2=3.455 $Y2=1.045
r207 41 42 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.067 $Y=1.09
+ $X2=6.067 $Y2=1.24
r208 38 47 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.355 $Y=1.37
+ $X2=10.355 $Y2=2.18
r209 34 47 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.365 $Y=2.27
+ $X2=10.365 $Y2=2.18
r210 34 36 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=10.365 $Y=2.27
+ $X2=10.365 $Y2=2.75
r211 32 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.28 $Y=1.295
+ $X2=10.355 $Y2=1.37
r212 32 33 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=10.28 $Y=1.295
+ $X2=9.77 $Y2=1.295
r213 29 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.695 $Y=1.22
+ $X2=9.77 $Y2=1.295
r214 29 31 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.695 $Y=1.22
+ $X2=9.695 $Y2=0.87
r215 28 31 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=9.695 $Y=0.255
+ $X2=9.695 $Y2=0.87
r216 25 43 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=6.255 $Y=2.115
+ $X2=6.095 $Y2=2.115
r217 25 27 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.255 $Y=2.19
+ $X2=6.255 $Y2=2.585
r218 24 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.115 $Y=0.18
+ $X2=6.04 $Y2=0.18
r219 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.62 $Y=0.18
+ $X2=9.695 $Y2=0.255
r220 23 24 1797.24 $w=1.5e-07 $l=3.505e-06 $layer=POLY_cond $X=9.62 $Y=0.18
+ $X2=6.115 $Y2=0.18
r221 22 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.095 $Y=2.04
+ $X2=6.095 $Y2=2.115
r222 22 42 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.095 $Y=2.04
+ $X2=6.095 $Y2=1.24
r223 20 41 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.04 $Y=0.805
+ $X2=6.04 $Y2=1.09
r224 17 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.04 $Y=0.255
+ $X2=6.04 $Y2=0.18
r225 17 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.04 $Y=0.255
+ $X2=6.04 $Y2=0.805
r226 15 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.965 $Y=0.18
+ $X2=6.04 $Y2=0.18
r227 15 16 835.809 $w=1.5e-07 $l=1.63e-06 $layer=POLY_cond $X=5.965 $Y=0.18
+ $X2=4.335 $Y2=0.18
r228 13 72 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=4.32 $Y=2.4
+ $X2=4.32 $Y2=1.67
r229 10 71 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.26 $Y=0.78
+ $X2=4.26 $Y2=1.34
r230 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.26 $Y=0.255
+ $X2=4.335 $Y2=0.18
r231 7 10 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.26 $Y=0.255
+ $X2=4.26 $Y2=0.78
r232 2 63 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.645 $Y2=2.115
r233 2 54 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.645 $Y2=2.815
r234 1 50 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.31
+ $Y=0.41 $X2=3.455 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_2133_410# 1 2 3 12 14 18 22 26 28 32 36
+ 38 41 45 46 48 50 51 52 55 56 57 59 60 61 65 68 69 71 78 80 82 90
c239 50 0 1.31405e-19 $X=13.115 $Y=2.38
c240 26 0 1.65234e-19 $X=14.785 $Y=0.74
r241 89 90 28.3072 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=14.785 $Y=1.465
+ $X2=14.935 $Y2=1.465
r242 79 89 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=14.77 $Y=1.465
+ $X2=14.785 $Y2=1.465
r243 79 86 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=14.77 $Y=1.465
+ $X2=14.75 $Y2=1.465
r244 78 81 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=14.742 $Y=1.465
+ $X2=14.742 $Y2=1.63
r245 78 80 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=14.742 $Y=1.465
+ $X2=14.742 $Y2=1.3
r246 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.77
+ $Y=1.465 $X2=14.77 $Y2=1.465
r247 71 73 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=12.63 $Y=0.775
+ $X2=12.63 $Y2=0.875
r248 67 69 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=2.805
+ $X2=11.79 $Y2=2.805
r249 67 68 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=2.805
+ $X2=11.46 $Y2=2.805
r250 65 81 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=14.635 $Y=2.21
+ $X2=14.635 $Y2=1.63
r251 62 80 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=14.635 $Y=1.02
+ $X2=14.635 $Y2=1.3
r252 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.55 $Y=0.935
+ $X2=14.635 $Y2=1.02
r253 60 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.55 $Y=0.935
+ $X2=14.245 $Y2=0.935
r254 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.16 $Y=0.85
+ $X2=14.245 $Y2=0.935
r255 58 59 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=14.16 $Y=0.5
+ $X2=14.16 $Y2=0.85
r256 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.075 $Y=0.415
+ $X2=14.16 $Y2=0.5
r257 56 57 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=14.075 $Y=0.415
+ $X2=13.565 $Y2=0.415
r258 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.48 $Y=0.5
+ $X2=13.565 $Y2=0.415
r259 54 55 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.48 $Y=0.5
+ $X2=13.48 $Y2=0.79
r260 53 76 4.65971 $w=1.7e-07 $l=1.98997e-07 $layer=LI1_cond $X=13.28 $Y=2.295
+ $X2=13.115 $Y2=2.22
r261 52 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.55 $Y=2.295
+ $X2=14.635 $Y2=2.21
r262 52 53 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=14.55 $Y=2.295
+ $X2=13.28 $Y2=2.295
r263 50 76 3.10647 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=13.115 $Y=2.38
+ $X2=13.115 $Y2=2.22
r264 50 51 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=13.115 $Y=2.38
+ $X2=13.115 $Y2=2.63
r265 49 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.795 $Y=0.875
+ $X2=12.63 $Y2=0.875
r266 48 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.395 $Y=0.875
+ $X2=13.48 $Y2=0.79
r267 48 49 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=13.395 $Y=0.875
+ $X2=12.795 $Y2=0.875
r268 46 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.95 $Y=2.715
+ $X2=13.115 $Y2=2.63
r269 46 69 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=12.95 $Y=2.715
+ $X2=11.79 $Y2=2.715
r270 45 68 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=10.995 $Y=2.715
+ $X2=11.46 $Y2=2.715
r271 42 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.83 $Y=2.215
+ $X2=10.83 $Y2=2.38
r272 42 82 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.83 $Y=2.215
+ $X2=10.83 $Y2=2.125
r273 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.83
+ $Y=2.215 $X2=10.83 $Y2=2.215
r274 39 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.83 $Y=2.63
+ $X2=10.995 $Y2=2.715
r275 39 41 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=10.83 $Y=2.63
+ $X2=10.83 $Y2=2.215
r276 34 38 30.0832 $w=1.65e-07 $l=1.42302e-07 $layer=POLY_cond $X=15.775 $Y=1.3
+ $X2=15.76 $Y2=1.435
r277 34 36 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=15.775 $Y=1.3
+ $X2=15.775 $Y2=0.645
r278 30 38 30.0832 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=15.76 $Y=1.57
+ $X2=15.76 $Y2=1.435
r279 30 32 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=15.76 $Y=1.57
+ $X2=15.76 $Y2=2.34
r280 28 38 1.40033 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=15.67 $Y=1.435
+ $X2=15.76 $Y2=1.435
r281 28 90 163.298 $w=2.7e-07 $l=7.35e-07 $layer=POLY_cond $X=15.67 $Y=1.435
+ $X2=14.935 $Y2=1.435
r282 24 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.785 $Y=1.3
+ $X2=14.785 $Y2=1.465
r283 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.785 $Y=1.3
+ $X2=14.785 $Y2=0.74
r284 20 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.75 $Y=1.63
+ $X2=14.75 $Y2=1.465
r285 20 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=14.75 $Y=1.63
+ $X2=14.75 $Y2=2.4
r286 16 18 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=11.285 $Y=2.05
+ $X2=11.285 $Y2=0.805
r287 15 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.995 $Y=2.125
+ $X2=10.83 $Y2=2.125
r288 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.21 $Y=2.125
+ $X2=11.285 $Y2=2.05
r289 14 15 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=11.21 $Y=2.125
+ $X2=10.995 $Y2=2.125
r290 12 85 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=10.755 $Y=2.75
+ $X2=10.755 $Y2=2.38
r291 3 76 300 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=2 $X=12.98
+ $Y=1.96 $X2=13.115 $Y2=2.225
r292 2 67 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=11.48
+ $Y=1.96 $X2=11.625 $Y2=2.805
r293 1 71 182 $w=1.7e-07 $l=5.11102e-07 $layer=licon1_NDIFF $count=1 $X=12.39
+ $Y=0.37 $X2=12.63 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_1954_119# 1 2 9 13 16 21 24 25 26 27 30
+ 32 33 34 36 37 39 40 45 48 49 50
c153 50 0 9.77748e-20 $X=11.255 $Y=1.81
c154 49 0 1.86341e-19 $X=10.58 $Y=0.897
c155 48 0 1.23089e-20 $X=10.415 $Y=0.87
c156 45 0 1.99515e-19 $X=10.325 $Y=2.195
c157 40 0 7.63376e-20 $X=13.275 $Y=1.635
c158 26 0 1.94296e-19 $X=10.41 $Y=1.81
c159 24 0 3.8609e-20 $X=10.325 $Y=2.11
c160 16 0 9.562e-20 $X=12.875 $Y=1.635
r161 48 49 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=0.897
+ $X2=10.58 $Y2=0.897
r162 43 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.055 $Y=2.195
+ $X2=10.325 $Y2=2.195
r163 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.275
+ $Y=1.635 $X2=13.275 $Y2=1.635
r164 37 39 13.5824 $w=4.18e-07 $l=4.95e-07 $layer=LI1_cond $X=12.78 $Y=1.68
+ $X2=13.275 $Y2=1.68
r165 35 37 7.86469 $w=3.2e-07 $l=2.48898e-07 $layer=LI1_cond $X=12.695 $Y=1.89
+ $X2=12.78 $Y2=1.68
r166 35 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=12.695 $Y=1.89
+ $X2=12.695 $Y2=2.29
r167 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.61 $Y=2.375
+ $X2=12.695 $Y2=2.29
r168 33 34 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=12.61 $Y=2.375
+ $X2=11.34 $Y2=2.375
r169 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.255 $Y=2.29
+ $X2=11.34 $Y2=2.375
r170 31 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=1.895
+ $X2=11.255 $Y2=1.81
r171 31 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.255 $Y=1.895
+ $X2=11.255 $Y2=2.29
r172 30 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=1.725
+ $X2=11.255 $Y2=1.81
r173 29 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.255 $Y=1.09
+ $X2=11.255 $Y2=1.725
r174 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.17 $Y=1.005
+ $X2=11.255 $Y2=1.09
r175 27 49 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.17 $Y=1.005
+ $X2=10.58 $Y2=1.005
r176 25 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.17 $Y=1.81
+ $X2=11.255 $Y2=1.81
r177 25 26 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=11.17 $Y=1.81
+ $X2=10.41 $Y2=1.81
r178 24 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.325 $Y=2.11
+ $X2=10.325 $Y2=2.195
r179 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.325 $Y=1.895
+ $X2=10.41 $Y2=1.81
r180 23 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.325 $Y=1.895
+ $X2=10.325 $Y2=2.11
r181 21 43 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=10.055 $Y=2.815
+ $X2=10.055 $Y2=2.28
r182 15 40 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=12.98 $Y=1.635
+ $X2=13.275 $Y2=1.635
r183 15 16 3.90195 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=12.98 $Y=1.635
+ $X2=12.875 $Y2=1.635
r184 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.89 $Y=1.8
+ $X2=12.875 $Y2=1.635
r185 11 13 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=12.89 $Y=1.8
+ $X2=12.89 $Y2=2.46
r186 7 16 34.7346 $w=1.65e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.845 $Y=1.47
+ $X2=12.875 $Y2=1.635
r187 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=12.845 $Y=1.47
+ $X2=12.845 $Y2=0.74
r188 2 43 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=9.92
+ $Y=2.12 $X2=10.055 $Y2=2.275
r189 2 21 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=9.92
+ $Y=2.12 $X2=10.055 $Y2=2.815
r190 1 48 91 $w=1.7e-07 $l=7.70325e-07 $layer=licon1_NDIFF $count=2 $X=9.77
+ $Y=0.595 $X2=10.415 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%RESET_B 1 3 4 6 7 8 10 11 18
c54 11 0 1.65234e-19 $X=14.16 $Y=1.295
r55 16 18 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=14.23 $Y=1.385
+ $X2=14.26 $Y2=1.385
r56 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.23
+ $Y=1.385 $X2=14.23 $Y2=1.385
r57 13 16 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=14.035 $Y=1.385
+ $X2=14.23 $Y2=1.385
r58 11 17 3.40065 $w=3.03e-07 $l=9e-08 $layer=LI1_cond $X=14.227 $Y=1.295
+ $X2=14.227 $Y2=1.385
r59 9 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.26 $Y=1.55
+ $X2=14.26 $Y2=1.385
r60 9 10 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=14.26 $Y=1.55
+ $X2=14.26 $Y2=2.095
r61 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.185 $Y=2.17
+ $X2=14.26 $Y2=2.095
r62 7 8 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=14.185 $Y=2.17
+ $X2=14.03 $Y2=2.17
r63 4 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.035 $Y=1.22
+ $X2=14.035 $Y2=1.385
r64 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=14.035 $Y=1.22
+ $X2=14.035 $Y2=0.9
r65 1 8 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=13.94 $Y=2.245
+ $X2=14.03 $Y2=2.17
r66 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=13.94 $Y=2.245
+ $X2=13.94 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_3078_384# 1 2 9 13 16 20 24 25 27 29
c53 25 0 1.99629e-19 $X=16.225 $Y=1.385
r54 25 30 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=16.225 $Y=1.385
+ $X2=16.225 $Y2=1.55
r55 25 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=16.225 $Y=1.385
+ $X2=16.225 $Y2=1.22
r56 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.225
+ $Y=1.385 $X2=16.225 $Y2=1.385
r57 22 27 0.533013 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=15.725 $Y=1.385
+ $X2=15.587 $Y2=1.385
r58 22 24 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=15.725 $Y=1.385
+ $X2=16.225 $Y2=1.385
r59 18 27 6.22203 $w=2.62e-07 $l=1.70895e-07 $layer=LI1_cond $X=15.575 $Y=1.55
+ $X2=15.587 $Y2=1.385
r60 18 20 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=15.575 $Y=1.55
+ $X2=15.575 $Y2=2.065
r61 14 27 6.22203 $w=2.62e-07 $l=1.65e-07 $layer=LI1_cond $X=15.587 $Y=1.22
+ $X2=15.587 $Y2=1.385
r62 14 16 24.0965 $w=2.73e-07 $l=5.75e-07 $layer=LI1_cond $X=15.587 $Y=1.22
+ $X2=15.587 $Y2=0.645
r63 13 29 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=16.285 $Y=0.74
+ $X2=16.285 $Y2=1.22
r64 9 30 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=16.295 $Y=2.4
+ $X2=16.295 $Y2=1.55
r65 2 20 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=15.39
+ $Y=1.92 $X2=15.535 $Y2=2.065
r66 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=15.415
+ $Y=0.37 $X2=15.56 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_27_464# 1 2 9 11 12 14 15 16 19
c49 16 0 8.66027e-20 $X=1.235 $Y=2.99
r50 17 19 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.08 $Y2=2.465
r51 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.915 $Y=2.99
+ $X2=2.08 $Y2=2.905
r52 15 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.915 $Y=2.99
+ $X2=1.235 $Y2=2.99
r53 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.905
+ $X2=1.235 $Y2=2.99
r54 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.15 $Y=2.215
+ $X2=1.15 $Y2=2.905
r55 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.13
+ $X2=1.15 $Y2=2.215
r56 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=2.13
+ $X2=0.395 $Y2=2.13
r57 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.255 $Y=2.215
+ $X2=0.395 $Y2=2.13
r58 7 9 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.255 $Y=2.215
+ $X2=0.255 $Y2=2.465
r59 2 19 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=2.32 $X2=2.08 $Y2=2.465
r60 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 43 47 51
+ 55 59 63 68 69 71 74 78 79 80 82 87 95 107 115 119 132 133 136 139 142 145 148
+ 151 158
c190 41 0 1.27434e-19 $X=4.095 $Y=2.455
c191 6 0 1.73394e-19 $X=9.07 $Y=2.12
c192 5 0 1.79798e-19 $X=8.075 $Y=2.12
r193 159 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r194 158 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r195 158 159 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r196 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r197 151 154 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.16 $Y=3.055
+ $X2=12.16 $Y2=3.33
r198 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r199 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r200 143 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r201 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r202 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r203 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r205 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.56 $Y2=3.33
r206 130 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=14.64 $Y2=3.33
r207 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r208 127 158 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=14.69 $Y=3.33
+ $X2=14.345 $Y2=3.33
r209 127 129 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=14.69 $Y=3.33
+ $X2=15.6 $Y2=3.33
r210 126 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r211 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r212 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r213 123 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r214 122 125 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r215 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r216 120 154 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.16 $Y2=3.33
r217 120 122 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.72 $Y2=3.33
r218 119 158 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=14 $Y=3.33
+ $X2=14.345 $Y2=3.33
r219 119 125 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=14 $Y=3.33
+ $X2=13.68 $Y2=3.33
r220 118 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r221 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r222 115 154 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.995 $Y=3.33
+ $X2=12.16 $Y2=3.33
r223 115 117 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.995 $Y=3.33
+ $X2=11.76 $Y2=3.33
r224 114 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r225 114 149 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.36 $Y2=3.33
r226 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r227 111 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.38 $Y=3.33
+ $X2=9.215 $Y2=3.33
r228 111 113 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=9.38 $Y=3.33
+ $X2=10.8 $Y2=3.33
r229 110 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r230 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r231 107 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.05 $Y=3.33
+ $X2=9.215 $Y2=3.33
r232 107 109 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.05 $Y=3.33
+ $X2=8.88 $Y2=3.33
r233 105 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r234 103 106 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r235 103 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r236 102 105 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r237 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r238 100 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.145 $Y2=3.33
r239 100 102 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.52 $Y2=3.33
r240 99 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r241 99 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r242 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r243 96 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=2.595 $Y2=3.33
r244 96 98 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=3.6 $Y2=3.33
r245 95 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=4.055 $Y2=3.33
r246 95 98 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=3.6 $Y2=3.33
r247 94 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r248 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r249 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r250 91 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r251 90 93 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r252 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r253 88 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r254 88 90 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r255 87 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.595 $Y2=3.33
r256 87 93 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.16 $Y2=3.33
r257 85 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r258 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r259 82 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r260 82 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r261 80 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r262 80 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r263 78 129 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=15.905 $Y=3.33
+ $X2=15.6 $Y2=3.33
r264 78 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.905 $Y=3.33
+ $X2=16.03 $Y2=3.33
r265 77 132 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=16.56 $Y2=3.33
r266 77 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=16.03 $Y2=3.33
r267 75 117 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=11.76 $Y2=3.33
r268 74 113 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=10.9 $Y=3.33
+ $X2=10.8 $Y2=3.33
r269 73 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=3.33
+ $X2=11.23 $Y2=3.33
r270 73 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=3.33
+ $X2=10.9 $Y2=3.33
r271 71 73 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=11.065 $Y=3.055
+ $X2=11.065 $Y2=3.33
r272 68 105 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.92 $Y2=3.33
r273 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.21 $Y2=3.33
r274 67 109 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.88 $Y2=3.33
r275 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.21 $Y2=3.33
r276 63 66 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=16.03 $Y=2.065
+ $X2=16.03 $Y2=2.815
r277 61 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.03 $Y=3.245
+ $X2=16.03 $Y2=3.33
r278 61 66 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.03 $Y=3.245
+ $X2=16.03 $Y2=2.815
r279 57 158 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=14.345 $Y=3.245
+ $X2=14.345 $Y2=3.33
r280 57 59 9.7073 $w=6.88e-07 $l=5.6e-07 $layer=LI1_cond $X=14.345 $Y=3.245
+ $X2=14.345 $Y2=2.685
r281 53 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.215 $Y=3.245
+ $X2=9.215 $Y2=3.33
r282 53 55 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=9.215 $Y=3.245
+ $X2=9.215 $Y2=2.635
r283 49 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=3.33
r284 49 51 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=2.815
r285 45 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=3.33
r286 45 47 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=2.695
r287 44 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=3.33
+ $X2=4.055 $Y2=3.33
r288 43 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=5.145 $Y2=3.33
r289 43 44 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=4.18 $Y2=3.33
r290 39 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=3.245
+ $X2=4.055 $Y2=3.33
r291 39 41 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.055 $Y=3.245
+ $X2=4.055 $Y2=2.455
r292 35 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=3.33
r293 35 37 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=2.465
r294 31 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r295 31 33 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.47
r296 10 66 600 $w=1.7e-07 $l=9.98962e-07 $layer=licon1_PDIFF $count=1 $X=15.85
+ $Y=1.92 $X2=16.07 $Y2=2.815
r297 10 63 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=15.85
+ $Y=1.92 $X2=16.07 $Y2=2.065
r298 9 59 300 $w=1.7e-07 $l=6.52457e-07 $layer=licon1_PDIFF $count=2 $X=14.03
+ $Y=2.32 $X2=14.525 $Y2=2.685
r299 8 151 600 $w=1.7e-07 $l=1.19997e-06 $layer=licon1_PDIFF $count=1 $X=11.94
+ $Y=1.96 $X2=12.16 $Y2=3.055
r300 7 71 600 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_PDIFF $count=1 $X=10.845
+ $Y=2.54 $X2=11.065 $Y2=3.055
r301 6 55 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=2.12 $X2=9.215 $Y2=2.635
r302 5 51 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=8.075
+ $Y=2.12 $X2=8.21 $Y2=2.815
r303 4 47 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=2.485 $X2=5.105 $Y2=2.695
r304 3 41 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.96
+ $Y=1.84 $X2=4.095 $Y2=2.455
r305 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=2.32 $X2=2.635 $Y2=2.465
r306 1 33 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.32 $X2=0.73 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_197_119# 1 2 3 4 13 15 17 21 23 24 26 27
+ 30 31 32 34 35 36 38 39 40 42 43 44 48 49 51 52 54 56 60 61 65 66
c223 61 0 1.93711e-19 $X=1.57 $Y=0.95
c224 54 0 4.35224e-20 $X=7.505 $Y=2.31
c225 52 0 2.87426e-20 $X=6.925 $Y=0.875
c226 49 0 1.51675e-19 $X=7.42 $Y=2.395
c227 44 0 4.28297e-20 $X=5.97 $Y=0.34
c228 39 0 2.29882e-20 $X=5.8 $Y=1.29
c229 13 0 2.95072e-20 $X=1.485 $Y=0.95
r230 66 69 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=6.53 $Y=2.395
+ $X2=6.53 $Y2=2.52
r231 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.57 $Y=0.95
+ $X2=1.57 $Y2=1.225
r232 56 58 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.125 $Y=0.805
+ $X2=1.125 $Y2=0.95
r233 53 54 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=7.505 $Y=0.96
+ $X2=7.505 $Y2=2.31
r234 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.42 $Y=0.875
+ $X2=7.505 $Y2=0.96
r235 51 52 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.42 $Y=0.875
+ $X2=6.925 $Y2=0.875
r236 50 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=2.395
+ $X2=6.53 $Y2=2.395
r237 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.42 $Y=2.395
+ $X2=7.505 $Y2=2.31
r238 49 50 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.42 $Y=2.395
+ $X2=6.695 $Y2=2.395
r239 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.76 $Y=0.79
+ $X2=6.925 $Y2=0.875
r240 46 48 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.76 $Y=0.79
+ $X2=6.76 $Y2=0.765
r241 45 48 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.76 $Y=0.425
+ $X2=6.76 $Y2=0.765
r242 43 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.595 $Y=0.34
+ $X2=6.76 $Y2=0.425
r243 43 44 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.595 $Y=0.34
+ $X2=5.97 $Y2=0.34
r244 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.885 $Y=0.425
+ $X2=5.97 $Y2=0.34
r245 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.885 $Y=0.425
+ $X2=5.885 $Y2=1.205
r246 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.8 $Y=1.29
+ $X2=5.885 $Y2=1.205
r247 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.8 $Y=1.29
+ $X2=5.13 $Y2=1.29
r248 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.045 $Y=1.205
+ $X2=5.13 $Y2=1.29
r249 37 38 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.045 $Y=0.75
+ $X2=5.045 $Y2=1.205
r250 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.96 $Y=0.665
+ $X2=5.045 $Y2=0.75
r251 35 36 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=4.96 $Y=0.665
+ $X2=3.4 $Y2=0.665
r252 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.315 $Y=0.58
+ $X2=3.4 $Y2=0.665
r253 33 34 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.315 $Y=0.425
+ $X2=3.315 $Y2=0.58
r254 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.23 $Y=0.34
+ $X2=3.315 $Y2=0.425
r255 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.23 $Y=0.34
+ $X2=2.56 $Y2=0.34
r256 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.425
+ $X2=2.56 $Y2=0.34
r257 29 30 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.475 $Y=0.425
+ $X2=2.475 $Y2=1.14
r258 28 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.225
+ $X2=2.07 $Y2=1.225
r259 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.39 $Y=1.225
+ $X2=2.475 $Y2=1.14
r260 27 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.39 $Y=1.225
+ $X2=2.155 $Y2=1.225
r261 25 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.31
+ $X2=2.07 $Y2=1.225
r262 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=1.31
+ $X2=2.07 $Y2=1.98
r263 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=2.065
+ $X2=2.07 $Y2=1.98
r264 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.985 $Y=2.065
+ $X2=1.715 $Y2=2.065
r265 22 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=1.225
+ $X2=1.57 $Y2=1.225
r266 21 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.225
+ $X2=2.07 $Y2=1.225
r267 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.985 $Y=1.225
+ $X2=1.655 $Y2=1.225
r268 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.715 $Y2=2.065
r269 19 60 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.63 $Y2=2.3
r270 15 60 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.59 $Y=2.425
+ $X2=1.59 $Y2=2.3
r271 15 17 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=2.425
+ $X2=1.59 $Y2=2.515
r272 14 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0.95
+ $X2=1.125 $Y2=0.95
r273 13 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=0.95
+ $X2=1.57 $Y2=0.95
r274 13 14 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.485 $Y=0.95
+ $X2=1.29 $Y2=0.95
r275 4 69 600 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=2.265 $X2=6.53 $Y2=2.52
r276 3 17 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.32 $X2=1.63 $Y2=2.515
r277 2 48 182 $w=1.7e-07 $l=2.87706e-07 $layer=licon1_NDIFF $count=1 $X=6.545
+ $Y=0.595 $X2=6.76 $Y2=0.765
r278 1 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.595 $X2=1.125 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%Q_N 1 2 9 13 14 15 16 23 33
r35 21 35 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=15.082 $Y=2.012
+ $X2=15.082 $Y2=1.985
r36 21 23 0.688472 $w=3.83e-07 $l=2.3e-08 $layer=LI1_cond $X=15.082 $Y=2.012
+ $X2=15.082 $Y2=2.035
r37 16 30 1.19734 $w=3.83e-07 $l=4e-08 $layer=LI1_cond $X=15.082 $Y=2.775
+ $X2=15.082 $Y2=2.815
r38 15 16 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=15.082 $Y=2.405
+ $X2=15.082 $Y2=2.775
r39 14 35 0.119734 $w=3.83e-07 $l=4e-09 $layer=LI1_cond $X=15.082 $Y=1.981
+ $X2=15.082 $Y2=1.985
r40 14 33 8.4692 $w=3.83e-07 $l=1.61e-07 $layer=LI1_cond $X=15.082 $Y=1.981
+ $X2=15.082 $Y2=1.82
r41 14 15 10.1475 $w=3.83e-07 $l=3.39e-07 $layer=LI1_cond $X=15.082 $Y=2.066
+ $X2=15.082 $Y2=2.405
r42 14 23 0.927941 $w=3.83e-07 $l=3.1e-08 $layer=LI1_cond $X=15.082 $Y=2.066
+ $X2=15.082 $Y2=2.035
r43 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.19 $Y=1.13
+ $X2=15.19 $Y2=1.82
r44 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=15.095 $Y=0.95
+ $X2=15.095 $Y2=1.13
r45 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=15.095 $Y=0.95
+ $X2=15.095 $Y2=0.515
r46 2 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.84
+ $Y=1.84 $X2=14.975 $Y2=1.985
r47 2 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.84
+ $Y=1.84 $X2=14.975 $Y2=2.815
r48 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.86
+ $Y=0.37 $X2=15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%Q 1 2 9 13 14 15 16 23 32
c24 14 0 1.99629e-19 $X=16.475 $Y=1.95
r25 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=16.535 $Y=2
+ $X2=16.535 $Y2=2.035
r26 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=16.535 $Y=2.405
+ $X2=16.535 $Y2=2.775
r27 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=16.535 $Y=1.975
+ $X2=16.535 $Y2=2
r28 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=16.535 $Y=1.975
+ $X2=16.535 $Y2=1.82
r29 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=16.535 $Y=2.06
+ $X2=16.535 $Y2=2.405
r30 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=16.535 $Y=2.06
+ $X2=16.535 $Y2=2.035
r31 13 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=16.63 $Y=1.05
+ $X2=16.63 $Y2=1.82
r32 7 13 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=16.525 $Y=0.86
+ $X2=16.525 $Y2=1.05
r33 7 9 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=16.525 $Y=0.86
+ $X2=16.525 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=16.385
+ $Y=1.84 $X2=16.52 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=16.385
+ $Y=1.84 $X2=16.52 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=16.36
+ $Y=0.37 $X2=16.5 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%VGND 1 2 3 4 5 6 7 8 25 27 31 35 39 43 47
+ 51 52 59 60 61 63 71 76 81 96 108 109 115 119 125 128 131
c171 109 0 3.18534e-20 $X=16.56 $Y=0
r172 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r173 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r174 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r175 119 122 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.965 $Y=0
+ $X2=3.965 $Y2=0.325
r176 119 120 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r177 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r178 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r179 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r180 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.56 $Y2=0
r181 106 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=14.64 $Y2=0
r182 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r183 103 131 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=14.735 $Y=0
+ $X2=14.575 $Y2=0
r184 103 105 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=14.735 $Y=0
+ $X2=15.6 $Y2=0
r185 102 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r186 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r187 99 102 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=14.16 $Y2=0
r188 98 101 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=14.16 $Y2=0
r189 98 99 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r190 96 131 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=14.415 $Y=0
+ $X2=14.575 $Y2=0
r191 96 101 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.415 $Y=0
+ $X2=14.16 $Y2=0
r192 95 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r193 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r194 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r195 92 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r196 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r197 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r198 89 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.96 $Y2=0
r199 89 91 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.36 $Y2=0
r200 85 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r201 84 87 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r202 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r203 82 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=0
+ $X2=5.465 $Y2=0
r204 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.63 $Y=0 $X2=6
+ $Y2=0
r205 81 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.96 $Y2=0
r206 81 87 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.4
+ $Y2=0
r207 80 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r208 80 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.08 $Y2=0
r209 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r210 77 119 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=0
+ $X2=3.965 $Y2=0
r211 77 79 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=4.13 $Y=0 $X2=5.04
+ $Y2=0
r212 76 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.465
+ $Y2=0
r213 76 79 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.04
+ $Y2=0
r214 75 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r215 75 116 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=2.16 $Y2=0
r216 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r217 72 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0
+ $X2=2.055 $Y2=0
r218 72 74 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.22 $Y=0 $X2=3.6
+ $Y2=0
r219 71 119 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.965
+ $Y2=0
r220 71 74 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.6
+ $Y2=0
r221 70 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r222 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r223 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r224 67 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r225 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r226 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r227 64 112 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0
+ $X2=0.235 $Y2=0
r228 64 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r229 63 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0
+ $X2=2.055 $Y2=0
r230 63 69 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r231 61 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r232 61 85 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=6
+ $Y2=0
r233 61 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r234 59 105 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=15.905 $Y=0
+ $X2=15.6 $Y2=0
r235 59 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.905 $Y=0
+ $X2=16.03 $Y2=0
r236 58 108 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.155 $Y=0
+ $X2=16.56 $Y2=0
r237 58 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.155 $Y=0
+ $X2=16.03 $Y2=0
r238 54 98 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=11.755 $Y=0
+ $X2=11.76 $Y2=0
r239 52 94 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=11.415 $Y=0
+ $X2=11.28 $Y2=0
r240 51 56 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.585 $Y2=0.325
r241 51 54 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.755 $Y2=0
r242 51 52 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.415 $Y2=0
r243 47 49 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=16.03 $Y=0.515
+ $X2=16.03 $Y2=0.885
r244 45 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.03 $Y=0.085
+ $X2=16.03 $Y2=0
r245 45 47 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.03 $Y=0.085
+ $X2=16.03 $Y2=0.515
r246 41 131 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=14.575 $Y=0.085
+ $X2=14.575 $Y2=0
r247 41 43 15.486 $w=3.18e-07 $l=4.3e-07 $layer=LI1_cond $X=14.575 $Y=0.085
+ $X2=14.575 $Y2=0.515
r248 37 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0
r249 37 39 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0.845
r250 33 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.465 $Y2=0
r251 33 35 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.465 $Y2=0.805
r252 29 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r253 29 31 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.77
r254 25 112 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.235 $Y2=0
r255 25 27 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.305 $Y2=0.805
r256 8 49 182 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_NDIFF $count=1 $X=15.85
+ $Y=0.37 $X2=16.07 $Y2=0.885
r257 8 47 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=15.85
+ $Y=0.37 $X2=16.07 $Y2=0.515
r258 7 43 182 $w=1.7e-07 $l=5.04975e-07 $layer=licon1_NDIFF $count=1 $X=14.11
+ $Y=0.69 $X2=14.535 $Y2=0.515
r259 6 56 182 $w=1.7e-07 $l=3.65582e-07 $layer=licon1_NDIFF $count=1 $X=11.36
+ $Y=0.595 $X2=11.585 $Y2=0.325
r260 5 39 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.82
+ $Y=0.595 $X2=8.96 $Y2=0.845
r261 4 35 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.595 $X2=5.465 $Y2=0.805
r262 3 122 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.41 $X2=3.965 $Y2=0.325
r263 2 31 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.595 $X2=2.055 $Y2=0.77
r264 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_1434_78# 1 2 7 11 13
r29 13 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.315 $Y=0.34
+ $X2=7.315 $Y2=0.535
r30 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.425 $Y=0.425
+ $X2=8.425 $Y2=0.855
r31 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.48 $Y=0.34
+ $X2=7.315 $Y2=0.34
r32 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.26 $Y=0.34
+ $X2=8.425 $Y2=0.425
r33 7 8 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=8.26 $Y=0.34 $X2=7.48
+ $Y2=0.34
r34 2 11 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.595 $X2=8.425 $Y2=0.855
r35 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=7.17
+ $Y=0.39 $X2=7.315 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_1%A_2392_74# 1 2 9 11 12 13
r31 13 16 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=13.1 $Y=0.34
+ $X2=13.1 $Y2=0.455
r32 11 13 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.975 $Y=0.34
+ $X2=13.1 $Y2=0.34
r33 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=12.975 $Y=0.34
+ $X2=12.265 $Y2=0.34
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.1 $Y=0.425
+ $X2=12.265 $Y2=0.34
r35 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=12.1 $Y=0.425 $X2=12.1
+ $Y2=0.495
r36 2 16 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.14 $Y2=0.455
r37 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=11.96
+ $Y=0.37 $X2=12.1 $Y2=0.495
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_343_368# A3 a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 a_230_94# B1 a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VPWR A1 a_259_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 VGND A1 a_230_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VGND A3 a_230_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_259_368# A2 a_343_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 X a_84_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_84_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 a_230_94# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 X a_84_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_1 A B C VGND VNB VPB VPWR X
M1000 a_601_384# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=7.15e+11p ps=5.61e+06u
M1001 VPWR a_84_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1002 VGND a_84_74# X VNB nlowvt w=740000u l=150000u
+  ad=5.466e+11p pd=4.39e+06u as=2.081e+11p ps=2.05e+06u
M1003 a_84_74# C a_601_384# VPB pshort w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 a_84_74# B a_223_120# VNB nlowvt w=640000u l=150000u
+  ad=4.177e+11p pd=4.01e+06u as=1.536e+11p ps=1.76e+06u
M1005 a_595_136# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1006 a_229_384# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND C a_403_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1008 a_84_74# C a_595_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_409_384# B a_84_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1010 a_84_74# B a_229_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_223_120# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C a_409_384# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_403_136# B a_84_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

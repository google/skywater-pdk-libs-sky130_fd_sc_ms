* File: sky130_fd_sc_ms__dlrtn_2.pex.spice
* Created: Wed Sep  2 12:05:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRTN_2%D 3 7 9 16
r30 14 16 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.6 $Y=1.615
+ $X2=0.675 $Y2=1.615
r31 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.615 $X2=0.6 $Y2=1.615
r32 11 14 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.495 $Y=1.615
+ $X2=0.6 $Y2=1.615
r33 9 15 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.615 $X2=0.6
+ $Y2=1.615
r34 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=1.78
+ $X2=0.675 $Y2=1.615
r35 5 7 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.675 $Y=1.78
+ $X2=0.675 $Y2=2.39
r36 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=1.615
r37 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%GATE_N 3 7 9 12
c39 12 0 1.5038e-19 $X=1.17 $Y=1.615
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.78
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.45
r42 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r43 7 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.225 $Y=2.39
+ $X2=1.225 $Y2=1.78
r44 3 14 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.085 $Y=0.86
+ $X2=1.085 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%A_232_98# 1 2 7 11 15 19 23 25 26 31 32 34
+ 35 38 39 42 43 48
c119 42 0 1.5038e-19 $X=1.45 $Y=2.115
r120 52 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.8 $Y=2.195
+ $X2=3.815 $Y2=2.195
r121 47 48 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.74 $Y=1.505
+ $X2=1.74 $Y2=1.415
r122 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.505 $X2=1.74 $Y2=1.505
r123 42 43 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=2.115
+ $X2=1.48 $Y2=1.95
r124 39 54 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=4.16 $Y=2.195
+ $X2=3.815 $Y2=2.195
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.16
+ $Y=2.195 $X2=4.16 $Y2=2.195
r126 36 38 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.16 $Y=2.52
+ $X2=4.16 $Y2=2.195
r127 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.995 $Y=2.605
+ $X2=4.16 $Y2=2.52
r128 34 35 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=3.995 $Y=2.605
+ $X2=1.675 $Y2=2.605
r129 32 46 9.11389 $w=2.71e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.675 $Y2=1.505
r130 32 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.59 $Y2=1.95
r131 31 35 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=1.48 $Y=2.52
+ $X2=1.675 $Y2=2.605
r132 30 42 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.48 $Y=2.145
+ $X2=1.48 $Y2=2.115
r133 30 31 11.0812 $w=3.88e-07 $l=3.75e-07 $layer=LI1_cond $X=1.48 $Y=2.145
+ $X2=1.48 $Y2=2.52
r134 26 46 18.9077 $w=2.71e-07 $l=4.2e-07 $layer=LI1_cond $X=1.675 $Y=1.085
+ $X2=1.675 $Y2=1.505
r135 26 28 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.505 $Y=1.085
+ $X2=1.3 $Y2=1.085
r136 21 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=2.36
+ $X2=3.815 $Y2=2.195
r137 21 23 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.815 $Y=2.36
+ $X2=3.815 $Y2=2.73
r138 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=2.03
+ $X2=3.8 $Y2=2.195
r139 17 19 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=3.8 $Y=2.03
+ $X2=3.8 $Y2=0.69
r140 13 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.235 $Y2=1.415
r141 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.25 $Y2=0.78
r142 9 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.235 $Y=1.49
+ $X2=2.235 $Y2=1.415
r143 9 11 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.235 $Y=1.49
+ $X2=2.235 $Y2=2.38
r144 8 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.415
+ $X2=1.74 $Y2=1.415
r145 7 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.145 $Y=1.415
+ $X2=2.235 $Y2=1.415
r146 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.145 $Y=1.415
+ $X2=1.905 $Y2=1.415
r147 2 42 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.315
+ $Y=1.97 $X2=1.45 $Y2=2.115
r148 1 28 182 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.3 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%A_27_136# 1 2 7 9 11 13 15 19 24 25 28 31 33
+ 34
c77 7 0 5.22992e-20 $X=2.855 $Y=1.59
r78 33 34 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.355 $Y=2.115
+ $X2=0.355 $Y2=1.95
r79 31 34 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.18 $Y=1.25 $X2=0.18
+ $Y2=1.95
r80 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.425 $X2=2.78 $Y2=1.425
r81 26 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.78 $Y=0.75
+ $X2=2.78 $Y2=1.425
r82 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.615 $Y=0.665
+ $X2=2.78 $Y2=0.75
r83 24 25 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=2.615 $Y=0.665
+ $X2=0.445 $Y2=0.665
r84 17 31 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=1.25
r85 17 19 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=0.955
r86 16 25 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.445 $Y2=0.665
r87 16 19 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.27 $Y2=0.955
r88 13 15 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.41 $Y=1.11 $X2=3.41
+ $Y2=0.69
r89 12 29 42.3736 $w=2.73e-07 $l=3.11769e-07 $layer=POLY_cond $X=2.945 $Y=1.185
+ $X2=2.78 $Y2=1.425
r90 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.335 $Y=1.185
+ $X2=3.41 $Y2=1.11
r91 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.335 $Y=1.185
+ $X2=2.945 $Y2=1.185
r92 7 29 34.7287 $w=2.73e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.855 $Y=1.59
+ $X2=2.78 $Y2=1.425
r93 7 9 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=2.855 $Y=1.59
+ $X2=2.855 $Y2=2.46
r94 2 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.305
+ $Y=1.97 $X2=0.45 $Y2=2.115
r95 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%A_373_82# 1 2 9 13 17 22 23 24 26 27 32 34
+ 35
c95 32 0 5.22992e-20 $X=2.16 $Y=1.045
c96 9 0 1.94055e-19 $X=3.275 $Y=2.46
r97 34 37 6.33844 $w=3.98e-07 $l=2.2e-07 $layer=LI1_cond $X=2.045 $Y=1.925
+ $X2=2.045 $Y2=2.145
r98 34 35 6.34273 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=1.925
+ $X2=2.045 $Y2=1.84
r99 30 32 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.02 $Y=1.045
+ $X2=2.16 $Y2=1.045
r100 27 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.355
+ $X2=4.25 $Y2=1.19
r101 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=1.355 $X2=4.25 $Y2=1.355
r102 24 26 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.485 $Y=1.355
+ $X2=4.25 $Y2=1.355
r103 23 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.32 $Y=1.635
+ $X2=3.32 $Y2=1.8
r104 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.635 $X2=3.32 $Y2=1.635
r105 20 22 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.32 $Y=1.84
+ $X2=3.32 $Y2=1.635
r106 19 24 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.32 $Y=1.52
+ $X2=3.485 $Y2=1.355
r107 19 22 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.32 $Y=1.52
+ $X2=3.32 $Y2=1.635
r108 18 34 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.245 $Y=1.925
+ $X2=2.045 $Y2=1.925
r109 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.155 $Y=1.925
+ $X2=3.32 $Y2=1.84
r110 17 18 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=3.155 $Y=1.925
+ $X2=2.245 $Y2=1.925
r111 15 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.045
r112 15 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.84
r113 13 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.275 $Y=0.58
+ $X2=4.275 $Y2=1.19
r114 9 41 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.275 $Y=2.46
+ $X2=3.275 $Y2=1.8
r115 2 37 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.96 $X2=2.01 $Y2=2.145
r116 1 30 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.41 $X2=2.02 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%A_913_406# 1 2 9 13 15 17 21 25 27 31 35 38
+ 39 40 43 47 53 55 57 58 59 65 69 71
c137 59 0 3.65537e-20 $X=5.795 $Y=1.72
c138 55 0 7.11433e-20 $X=6.505 $Y=1.805
r139 66 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.68 $Y=1.485
+ $X2=6.68 $Y2=1.395
r140 65 67 14.5672 $w=2.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.675 $Y=1.485
+ $X2=6.675 $Y2=1.805
r141 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.68
+ $Y=1.485 $X2=6.68 $Y2=1.485
r142 62 63 5.33075 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=2.195
+ $X2=5.795 $Y2=2.36
r143 61 62 5.02353 $w=4.98e-07 $l=2.1e-07 $layer=LI1_cond $X=5.795 $Y=1.985
+ $X2=5.795 $Y2=2.195
r144 58 61 4.30588 $w=4.98e-07 $l=1.8e-07 $layer=LI1_cond $X=5.795 $Y=1.805
+ $X2=5.795 $Y2=1.985
r145 58 59 7.60339 $w=4.98e-07 $l=8.5e-08 $layer=LI1_cond $X=5.795 $Y=1.805
+ $X2=5.795 $Y2=1.72
r146 57 59 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.63 $Y=1.13
+ $X2=5.63 $Y2=1.72
r147 56 58 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.045 $Y=1.805
+ $X2=5.795 $Y2=1.805
r148 55 67 3.40055 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.505 $Y=1.805
+ $X2=6.675 $Y2=1.805
r149 55 56 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.505 $Y=1.805
+ $X2=6.045 $Y2=1.805
r150 53 63 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.88 $Y=2.815
+ $X2=5.88 $Y2=2.36
r151 45 57 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=5.512 $Y=0.928
+ $X2=5.512 $Y2=1.13
r152 45 47 11.7521 $w=4.03e-07 $l=4.13e-07 $layer=LI1_cond $X=5.512 $Y=0.928
+ $X2=5.512 $Y2=0.515
r153 43 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.73 $Y=2.195
+ $X2=4.73 $Y2=2.36
r154 43 69 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.73 $Y=2.195
+ $X2=4.73 $Y2=2.03
r155 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.73
+ $Y=2.195 $X2=4.73 $Y2=2.195
r156 40 62 3.16914 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=5.545 $Y=2.195
+ $X2=5.795 $Y2=2.195
r157 40 42 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=5.545 $Y=2.195
+ $X2=4.73 $Y2=2.195
r158 33 39 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=7.585 $Y=1.32
+ $X2=7.595 $Y2=1.395
r159 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.585 $Y=1.32
+ $X2=7.585 $Y2=0.74
r160 29 39 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.47
+ $X2=7.595 $Y2=1.395
r161 29 31 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=7.595 $Y=1.47
+ $X2=7.595 $Y2=2.4
r162 28 38 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.235 $Y=1.395
+ $X2=7.145 $Y2=1.395
r163 27 39 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=1.395
+ $X2=7.595 $Y2=1.395
r164 27 28 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.505 $Y=1.395
+ $X2=7.235 $Y2=1.395
r165 23 38 10.9219 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=7.155 $Y=1.32
+ $X2=7.145 $Y2=1.395
r166 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.155 $Y=1.32
+ $X2=7.155 $Y2=0.74
r167 19 38 10.9219 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=7.145 $Y=1.47
+ $X2=7.145 $Y2=1.395
r168 19 21 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=7.145 $Y=1.47
+ $X2=7.145 $Y2=2.4
r169 18 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=1.395
+ $X2=6.68 $Y2=1.395
r170 17 38 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.055 $Y=1.395
+ $X2=7.145 $Y2=1.395
r171 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.055 $Y=1.395
+ $X2=6.845 $Y2=1.395
r172 15 37 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.715 $Y=1.77
+ $X2=4.715 $Y2=1.68
r173 15 69 101.065 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=4.715 $Y=1.77
+ $X2=4.715 $Y2=2.03
r174 13 37 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=4.7 $Y=0.58 $X2=4.7
+ $Y2=1.68
r175 9 70 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.655 $Y=2.73
+ $X2=4.655 $Y2=2.36
r176 2 61 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.84 $X2=5.88 $Y2=1.985
r177 2 53 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.84 $X2=5.88 $Y2=2.815
r178 1 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.33
+ $Y=0.37 $X2=5.475 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%A_673_392# 1 2 9 13 15 16 17 22 23 24 27 29
+ 30 34 36
c100 24 0 1.94055e-19 $X=3.825 $Y=1.775
c101 15 0 1.01066e-19 $X=5.555 $Y=1.515
c102 9 0 7.11433e-20 $X=5.645 $Y=2.4
r103 34 36 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=5.172 $Y=1.515
+ $X2=5.172 $Y2=1.35
r104 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.21
+ $Y=1.515 $X2=5.21 $Y2=1.515
r105 31 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.055 $Y=1.02
+ $X2=5.055 $Y2=1.35
r106 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.97 $Y=0.935
+ $X2=5.055 $Y2=1.02
r107 29 30 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.97 $Y=0.935
+ $X2=4.225 $Y2=0.935
r108 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.06 $Y=0.85
+ $X2=4.225 $Y2=0.935
r109 25 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.06 $Y=0.85
+ $X2=4.06 $Y2=0.58
r110 23 34 7.3984 $w=4.03e-07 $l=2.6e-07 $layer=LI1_cond $X=5.172 $Y=1.775
+ $X2=5.172 $Y2=1.515
r111 23 24 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=4.97 $Y=1.775
+ $X2=3.825 $Y2=1.775
r112 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.74 $Y=1.86
+ $X2=3.825 $Y2=1.775
r113 21 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.74 $Y=1.86
+ $X2=3.74 $Y2=2.18
r114 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=2.265
+ $X2=3.74 $Y2=2.18
r115 17 19 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.655 $Y=2.265
+ $X2=3.5 $Y2=2.265
r116 15 35 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=5.555 $Y=1.515
+ $X2=5.21 $Y2=1.515
r117 15 16 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.555 $Y=1.515
+ $X2=5.555 $Y2=1.35
r118 11 16 34.7346 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=5.69 $Y=1.35
+ $X2=5.555 $Y2=1.35
r119 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.69 $Y=1.35
+ $X2=5.69 $Y2=0.74
r120 7 16 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=5.645 $Y=1.68
+ $X2=5.555 $Y2=1.35
r121 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.645 $Y=1.68
+ $X2=5.645 $Y2=2.4
r122 2 19 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=1.96 $X2=3.5 $Y2=2.265
r123 1 27 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.37 $X2=4.06 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%RESET_B 3 6 8 11 12 13
c37 13 0 3.65537e-20 $X=6.14 $Y=1.22
r38 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.385
+ $X2=6.14 $Y2=1.55
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.385
+ $X2=6.14 $Y2=1.22
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.14
+ $Y=1.385 $X2=6.14 $Y2=1.385
r41 8 12 4.3606 $w=3.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6 $Y=1.365 $X2=6.14
+ $Y2=1.365
r42 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.105 $Y=2.4
+ $X2=6.105 $Y2=1.55
r43 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.08 $Y=0.74 $X2=6.08
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%VPWR 1 2 3 4 5 18 22 26 28 30 35 36 37 43 55
+ 60 66 71 74 76 80
r83 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r84 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r85 73 74 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.38 $Y=3.022
+ $X2=5.545 $Y2=3.022
r86 69 73 5.18047 $w=7.83e-07 $l=3.4e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=5.38 $Y2=3.022
r87 69 71 13.7794 $w=7.83e-07 $l=3.25e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=4.715 $Y2=3.022
r88 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r89 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r91 64 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r93 61 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.485 $Y2=3.33
r94 61 63 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 60 79 4.82984 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.932 $Y2=3.33
r96 60 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 59 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r98 59 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r99 58 74 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6 $Y=3.33 $X2=5.545
+ $Y2=3.33
r100 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r101 55 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=3.33
+ $X2=6.485 $Y2=3.33
r102 55 58 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.32 $Y=3.33 $X2=6
+ $Y2=3.33
r103 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 53 71 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.715 $Y2=3.33
r105 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r106 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r107 51 53 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=4.56 $Y2=3.33
r108 49 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r111 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r112 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r113 43 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r114 43 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 41 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r116 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 37 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 37 67 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 35 40 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.95 $Y2=3.33
r121 34 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.95 $Y2=3.33
r123 30 33 28.1332 $w=3.38e-07 $l=8.3e-07 $layer=LI1_cond $X=7.875 $Y=1.985
+ $X2=7.875 $Y2=2.815
r124 28 79 3.02131 $w=3.4e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.875 $Y=3.245
+ $X2=7.932 $Y2=3.33
r125 28 33 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=7.875 $Y=3.245
+ $X2=7.875 $Y2=2.815
r126 24 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=3.33
r127 24 26 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=2.225
r128 20 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r129 20 22 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.025
r130 16 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=3.33
r131 16 18 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=2.115
r132 5 33 400 $w=1.7e-07 $l=1.06577e-06 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.84 $X2=7.875 $Y2=2.815
r133 5 30 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.84 $X2=7.875 $Y2=1.985
r134 4 26 300 $w=1.7e-07 $l=5.09779e-07 $layer=licon1_PDIFF $count=2 $X=6.195
+ $Y=1.84 $X2=6.485 $Y2=2.225
r135 3 73 300 $w=1.7e-07 $l=7.60164e-07 $layer=licon1_PDIFF $count=2 $X=4.745
+ $Y=2.52 $X2=5.38 $Y2=2.795
r136 2 22 600 $w=1.7e-07 $l=1.16984e-06 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.96 $X2=2.545 $Y2=3.025
r137 1 18 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.765
+ $Y=1.97 $X2=0.95 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%Q 1 2 9 13 14 15 16 29 30
r35 29 30 10.7408 $w=6.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.19 $Y=1.985
+ $X2=7.19 $Y2=1.82
r36 16 26 0.693379 $w=6.88e-07 $l=4e-08 $layer=LI1_cond $X=7.19 $Y=2.775
+ $X2=7.19 $Y2=2.815
r37 15 16 6.41375 $w=6.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.19 $Y=2.405
+ $X2=7.19 $Y2=2.775
r38 15 20 4.16027 $w=6.88e-07 $l=2.4e-07 $layer=LI1_cond $X=7.19 $Y=2.405
+ $X2=7.19 $Y2=2.165
r39 14 20 2.25348 $w=6.88e-07 $l=1.3e-07 $layer=LI1_cond $X=7.19 $Y=2.035
+ $X2=7.19 $Y2=2.165
r40 14 29 0.866723 $w=6.88e-07 $l=5e-08 $layer=LI1_cond $X=7.19 $Y=2.035
+ $X2=7.19 $Y2=1.985
r41 13 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.45 $Y=1.47
+ $X2=7.45 $Y2=1.82
r42 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.305
+ $X2=7.37 $Y2=1.47
r43 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7.37 $Y=1.305 $X2=7.37
+ $Y2=0.515
r44 2 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.235
+ $Y=1.84 $X2=7.37 $Y2=1.985
r45 2 26 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.235
+ $Y=1.84 $X2=7.37 $Y2=2.815
r46 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.23
+ $Y=0.37 $X2=7.37 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_2%VGND 1 2 3 4 5 18 22 24 26 28 30 43 51 56 63
+ 70 74 76 79 83
c75 18 0 1.01066e-19 $X=4.915 $Y=0.515
r76 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r77 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r78 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r79 72 74 9.36575 $w=4.93e-07 $l=1.6e-07 $layer=LI1_cond $X=3.12 $Y=0.162
+ $X2=3.28 $Y2=0.162
r80 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r81 69 72 0.120816 $w=4.93e-07 $l=5e-09 $layer=LI1_cond $X=3.115 $Y=0.162
+ $X2=3.12 $Y2=0.162
r82 69 70 23.2596 $w=4.93e-07 $l=7.35e-07 $layer=LI1_cond $X=3.115 $Y=0.162
+ $X2=2.38 $Y2=0.162
r83 63 66 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r84 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r85 60 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r86 60 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r87 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r88 57 79 15.5458 $w=1.7e-07 $l=4.53e-07 $layer=LI1_cond $X=7.035 $Y=0 $X2=6.582
+ $Y2=0
r89 57 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.035 $Y=0 $X2=7.44
+ $Y2=0
r90 56 82 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=0 $X2=7.932
+ $Y2=0
r91 56 59 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=0 $X2=7.44
+ $Y2=0
r92 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r93 55 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r94 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r95 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.915
+ $Y2=0
r96 52 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=6
+ $Y2=0
r97 51 79 15.5458 $w=1.7e-07 $l=4.52e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.582
+ $Y2=0
r98 51 54 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6
+ $Y2=0
r99 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r100 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r101 47 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r102 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r103 46 74 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.28
+ $Y2=0
r104 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r105 43 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.915
+ $Y2=0
r106 43 49 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r107 42 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r108 41 70 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.38
+ $Y2=0
r109 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r111 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r112 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r113 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r114 36 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r115 36 38 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r116 33 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r117 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 30 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r119 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r120 28 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r121 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r122 24 82 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.932 $Y2=0
r123 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.515
r124 20 79 3.35974 $w=9.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.582 $Y=0.085
+ $X2=6.582 $Y2=0
r125 20 22 5.79669 $w=9.03e-07 $l=4.3e-07 $layer=LI1_cond $X=6.582 $Y=0.085
+ $X2=6.582 $Y2=0.515
r126 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0
r127 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0.515
r128 5 26 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.66
+ $Y=0.37 $X2=7.87 $Y2=0.515
r129 4 22 45.5 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=4 $X=6.155
+ $Y=0.37 $X2=6.87 $Y2=0.515
r130 3 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.37 $X2=4.915 $Y2=0.515
r131 2 69 91 $w=1.7e-07 $l=8.31414e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.41 $X2=3.115 $Y2=0.325
r132 1 66 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends


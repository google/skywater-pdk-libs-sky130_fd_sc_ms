* File: sky130_fd_sc_ms__a2bb2oi_2.spice
* Created: Wed Sep  2 11:54:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2bb2oi_2.pex.spice"
.subckt sky130_fd_sc_ms__a2bb2oi_2  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1011 N_A_212_102#_M1011_d N_A1_N_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.104 AS=0.1696 PD=0.965 PS=1.81 NRD=3.744 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A2_N_M1007_g N_A_212_102#_M1011_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.113206 AS=0.104 PD=1.00174 PS=0.965 NRD=11.244 NRS=4.68 M=1
+ R=4.26667 SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_Y_M1002_d N_A_212_102#_M1002_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1002_d N_A_212_102#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g N_A_615_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1000_d N_B2_M1006_g N_A_615_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_615_74#_M1006_s N_B1_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_A_615_74#_M1014_d N_B1_M1014_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 A_212_392# N_A1_N_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1 AD=0.105
+ AS=0.26 PD=1.21 PS=2.52 NRD=9.8303 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90000.6
+ A=0.18 P=2.36 MULT=1
MM1015 N_A_212_102#_M1015_d N_A2_N_M1015_g A_212_392# VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_A_212_102#_M1003_g N_A_424_368#_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1003_d N_A_212_102#_M1004_g N_A_424_368#_M1004_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90002 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_B2_M1008_g N_A_424_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1008_d N_B2_M1009_g N_A_424_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1010_d N_B1_M1010_g N_A_424_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1010_d N_B1_M1013_g N_A_424_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_58 VNB 0 1.56524e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a2bb2oi_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a21boi_1.pxi.spice
* Created: Wed Sep  2 11:50:57 2020
* 
x_PM_SKY130_FD_SC_MS__A21BOI_1%B1_N N_B1_N_c_60_n N_B1_N_M1007_g N_B1_N_c_61_n
+ N_B1_N_c_62_n N_B1_N_M1001_g B1_N B1_N B1_N N_B1_N_c_63_n N_B1_N_c_64_n
+ PM_SKY130_FD_SC_MS__A21BOI_1%B1_N
x_PM_SKY130_FD_SC_MS__A21BOI_1%A_29_424# N_A_29_424#_M1001_s N_A_29_424#_M1007_s
+ N_A_29_424#_M1002_g N_A_29_424#_c_107_n N_A_29_424#_M1005_g
+ N_A_29_424#_c_116_n N_A_29_424#_c_117_n N_A_29_424#_c_118_n
+ N_A_29_424#_c_108_n N_A_29_424#_c_109_n N_A_29_424#_c_110_n
+ N_A_29_424#_c_111_n N_A_29_424#_c_112_n N_A_29_424#_c_113_n
+ N_A_29_424#_c_114_n PM_SKY130_FD_SC_MS__A21BOI_1%A_29_424#
x_PM_SKY130_FD_SC_MS__A21BOI_1%A1 N_A1_M1004_g N_A1_M1000_g A1 N_A1_c_181_n
+ N_A1_c_182_n PM_SKY130_FD_SC_MS__A21BOI_1%A1
x_PM_SKY130_FD_SC_MS__A21BOI_1%A2 N_A2_M1006_g N_A2_M1003_g A2 A2 N_A2_c_223_n
+ N_A2_c_224_n PM_SKY130_FD_SC_MS__A21BOI_1%A2
x_PM_SKY130_FD_SC_MS__A21BOI_1%VPWR N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_c_251_n
+ N_VPWR_c_252_n N_VPWR_c_253_n N_VPWR_c_254_n VPWR N_VPWR_c_255_n
+ N_VPWR_c_256_n N_VPWR_c_250_n N_VPWR_c_258_n PM_SKY130_FD_SC_MS__A21BOI_1%VPWR
x_PM_SKY130_FD_SC_MS__A21BOI_1%Y N_Y_M1005_d N_Y_M1002_s N_Y_c_291_n N_Y_c_288_n
+ N_Y_c_289_n N_Y_c_290_n Y Y Y N_Y_c_294_n PM_SKY130_FD_SC_MS__A21BOI_1%Y
x_PM_SKY130_FD_SC_MS__A21BOI_1%A_351_368# N_A_351_368#_M1002_d
+ N_A_351_368#_M1003_d N_A_351_368#_c_341_n N_A_351_368#_c_337_n
+ N_A_351_368#_c_338_n N_A_351_368#_c_339_n
+ PM_SKY130_FD_SC_MS__A21BOI_1%A_351_368#
x_PM_SKY130_FD_SC_MS__A21BOI_1%VGND N_VGND_M1001_d N_VGND_M1006_d N_VGND_c_364_n
+ N_VGND_c_365_n VGND N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n
+ N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n PM_SKY130_FD_SC_MS__A21BOI_1%VGND
cc_1 VNB N_B1_N_c_60_n 0.0621915f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.695
cc_2 VNB N_B1_N_c_61_n 0.0296109f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.26
cc_3 VNB N_B1_N_c_62_n 0.0169054f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.185
cc_4 VNB N_B1_N_c_63_n 0.125025f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=0.42
cc_5 VNB N_B1_N_c_64_n 0.00504936f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=0.42
cc_6 VNB N_A_29_424#_M1002_g 0.00667008f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.835
cc_7 VNB N_A_29_424#_c_107_n 0.0192839f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_8 VNB N_A_29_424#_c_108_n 0.00600215f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.44
cc_9 VNB N_A_29_424#_c_109_n 5.48582e-19 $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=0.42
cc_10 VNB N_A_29_424#_c_110_n 0.0031525f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=0.555
cc_11 VNB N_A_29_424#_c_111_n 0.0108997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_29_424#_c_112_n 0.00221045f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.44
cc_13 VNB N_A_29_424#_c_113_n 0.00329669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_29_424#_c_114_n 0.0431674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1000_g 0.0249694f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.185
cc_16 VNB N_A1_c_181_n 0.0259698f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A1_c_182_n 0.0041984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_M1003_g 0.00909003f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.26
cc_19 VNB A2 0.0455343f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.835
cc_20 VNB N_A2_c_223_n 0.0339369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_224_n 0.0215298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_250_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_288_n 0.00343427f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_24 VNB N_Y_c_289_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_290_n 0.00446143f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.185
cc_26 VNB N_VGND_c_364_n 0.0125231f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.835
cc_27 VNB N_VGND_c_365_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_28 VNB N_VGND_c_366_n 0.032726f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.42
cc_29 VNB N_VGND_c_367_n 0.029505f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.44
cc_30 VNB N_VGND_c_368_n 0.0148721f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=0.925
cc_31 VNB N_VGND_c_369_n 0.232561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_370_n 0.00962017f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.44
cc_33 VNB N_VGND_c_371_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_B1_N_c_60_n 0.00313824f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.695
cc_35 VPB N_B1_N_M1007_g 0.0505523f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_36 VPB N_A_29_424#_M1002_g 0.0258932f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.835
cc_37 VPB N_A_29_424#_c_116_n 0.0431662f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.185
cc_38 VPB N_A_29_424#_c_117_n 0.00982697f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=0.42
cc_39 VPB N_A_29_424#_c_118_n 0.0100261f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=0.42
cc_40 VPB N_A_29_424#_c_110_n 0.00313134f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=0.555
cc_41 VPB N_A1_M1004_g 0.02134f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_42 VPB N_A1_c_181_n 0.00559054f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB N_A1_c_182_n 0.00203881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A2_M1003_g 0.0311153f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.26
cc_45 VPB N_VPWR_c_251_n 0.020139f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.835
cc_46 VPB N_VPWR_c_252_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_253_n 0.0355956f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.185
cc_48 VPB N_VPWR_c_254_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=0.42
cc_49 VPB N_VPWR_c_255_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_256_n 0.0264269f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=1.44
cc_51 VPB N_VPWR_c_250_n 0.0789553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_258_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_Y_c_291_n 0.00146579f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.185
cc_54 VPB N_Y_c_288_n 3.48972e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_55 VPB Y 0.0175722f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=0.42
cc_56 VPB N_Y_c_294_n 0.0110082f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=1.44
cc_57 VPB N_A_351_368#_c_337_n 0.0314181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_351_368#_c_338_n 0.00242978f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.185
cc_59 VPB N_A_351_368#_c_339_n 0.0187294f $X=-0.19 $Y=1.66 $X2=0.285 $Y2=0.42
cc_60 N_B1_N_c_62_n N_A_29_424#_c_107_n 0.00907454f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_61 N_B1_N_M1007_g N_A_29_424#_c_116_n 0.0221138f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_62 N_B1_N_M1007_g N_A_29_424#_c_117_n 0.0177373f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_63 N_B1_N_c_61_n N_A_29_424#_c_117_n 0.00459448f $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_64 N_B1_N_c_64_n N_A_29_424#_c_117_n 0.0010324f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_65 N_B1_N_c_60_n N_A_29_424#_c_118_n 0.00222095f $X=0.495 $Y=1.695 $X2=0
+ $Y2=0
cc_66 N_B1_N_M1007_g N_A_29_424#_c_118_n 0.0043353f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_67 N_B1_N_c_64_n N_A_29_424#_c_118_n 0.0278594f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_68 N_B1_N_c_62_n N_A_29_424#_c_108_n 0.00467438f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_69 N_B1_N_c_63_n N_A_29_424#_c_108_n 0.0050246f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_70 N_B1_N_c_64_n N_A_29_424#_c_108_n 0.0403141f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_71 N_B1_N_c_61_n N_A_29_424#_c_109_n 0.00401161f $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_72 N_B1_N_c_62_n N_A_29_424#_c_109_n 0.0041311f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_73 N_B1_N_c_63_n N_A_29_424#_c_109_n 0.0011876f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_74 N_B1_N_c_64_n N_A_29_424#_c_109_n 0.00829248f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_75 N_B1_N_c_60_n N_A_29_424#_c_110_n 0.00731867f $X=0.495 $Y=1.695 $X2=0
+ $Y2=0
cc_76 N_B1_N_c_64_n N_A_29_424#_c_110_n 0.00271322f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_77 N_B1_N_c_61_n N_A_29_424#_c_111_n 0.0106117f $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_78 N_B1_N_c_61_n N_A_29_424#_c_112_n 0.00407965f $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_79 N_B1_N_c_62_n N_A_29_424#_c_112_n 0.00246642f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_80 N_B1_N_c_60_n N_A_29_424#_c_113_n 0.00557769f $X=0.495 $Y=1.695 $X2=0
+ $Y2=0
cc_81 N_B1_N_c_61_n N_A_29_424#_c_113_n 0.0090613f $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_82 N_B1_N_c_64_n N_A_29_424#_c_113_n 0.0179229f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_83 N_B1_N_c_61_n N_A_29_424#_c_114_n 0.00751861f $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_84 N_B1_N_M1007_g N_VPWR_c_251_n 0.00804508f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_85 N_B1_N_M1007_g N_VPWR_c_255_n 0.005209f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_86 N_B1_N_M1007_g N_VPWR_c_250_n 0.00991105f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_87 N_B1_N_c_61_n N_Y_c_288_n 4.43758e-19 $X=0.925 $Y=1.26 $X2=0 $Y2=0
cc_88 N_B1_N_c_62_n N_Y_c_290_n 4.02742e-19 $X=1 $Y=1.185 $X2=0 $Y2=0
cc_89 N_B1_N_M1007_g N_Y_c_294_n 0.0038131f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_90 N_B1_N_c_62_n N_VGND_c_364_n 0.00587808f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_91 N_B1_N_c_63_n N_VGND_c_364_n 0.00352148f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_92 N_B1_N_c_64_n N_VGND_c_364_n 0.00819751f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_93 N_B1_N_c_62_n N_VGND_c_366_n 0.0043356f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_94 N_B1_N_c_63_n N_VGND_c_366_n 0.00613683f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_95 N_B1_N_c_64_n N_VGND_c_366_n 0.0223605f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_96 N_B1_N_c_62_n N_VGND_c_369_n 0.00487769f $X=1 $Y=1.185 $X2=0 $Y2=0
cc_97 N_B1_N_c_63_n N_VGND_c_369_n 0.00385956f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_98 N_B1_N_c_64_n N_VGND_c_369_n 0.012558f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_99 N_A_29_424#_M1002_g N_A1_M1004_g 0.0307168f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_29_424#_c_107_n N_A1_M1000_g 0.018275f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A_29_424#_c_114_n N_A1_c_181_n 0.0203918f $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_102 N_A_29_424#_c_114_n N_A1_c_182_n 3.91289e-19 $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A_29_424#_M1002_g N_VPWR_c_251_n 0.00326547f $X=1.665 $Y=2.4 $X2=0
+ $Y2=0
cc_104 N_A_29_424#_c_116_n N_VPWR_c_251_n 0.0293161f $X=0.27 $Y=2.265 $X2=0
+ $Y2=0
cc_105 N_A_29_424#_c_117_n N_VPWR_c_251_n 0.0221455f $X=0.745 $Y=1.86 $X2=0
+ $Y2=0
cc_106 N_A_29_424#_M1002_g N_VPWR_c_252_n 7.62978e-19 $X=1.665 $Y=2.4 $X2=0
+ $Y2=0
cc_107 N_A_29_424#_M1002_g N_VPWR_c_253_n 0.005209f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_29_424#_c_116_n N_VPWR_c_255_n 0.014549f $X=0.27 $Y=2.265 $X2=0 $Y2=0
cc_109 N_A_29_424#_M1002_g N_VPWR_c_250_n 0.00988607f $X=1.665 $Y=2.4 $X2=0
+ $Y2=0
cc_110 N_A_29_424#_c_116_n N_VPWR_c_250_n 0.0119743f $X=0.27 $Y=2.265 $X2=0
+ $Y2=0
cc_111 N_A_29_424#_M1002_g N_Y_c_291_n 0.0190155f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_29_424#_c_111_n N_Y_c_291_n 7.13932e-19 $X=1.45 $Y=1.385 $X2=0 $Y2=0
cc_113 N_A_29_424#_c_114_n N_Y_c_291_n 0.00172466f $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_114 N_A_29_424#_M1002_g N_Y_c_288_n 0.00806386f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A_29_424#_c_107_n N_Y_c_288_n 0.00110635f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_116 N_A_29_424#_c_111_n N_Y_c_288_n 0.0249855f $X=1.45 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A_29_424#_c_114_n N_Y_c_288_n 0.00778846f $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_118 N_A_29_424#_c_107_n N_Y_c_289_n 3.97481e-19 $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_119 N_A_29_424#_c_107_n N_Y_c_290_n 0.00699147f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A_29_424#_M1002_g Y 0.00148248f $X=1.665 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_29_424#_c_116_n N_Y_c_294_n 0.00497542f $X=0.27 $Y=2.265 $X2=0 $Y2=0
cc_122 N_A_29_424#_c_117_n N_Y_c_294_n 0.0101435f $X=0.745 $Y=1.86 $X2=0 $Y2=0
cc_123 N_A_29_424#_c_110_n N_Y_c_294_n 0.00270822f $X=0.83 $Y=1.775 $X2=0 $Y2=0
cc_124 N_A_29_424#_c_111_n N_Y_c_294_n 0.0309215f $X=1.45 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A_29_424#_c_114_n N_Y_c_294_n 0.00559096f $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_29_424#_M1002_g N_A_351_368#_c_338_n 0.0143327f $X=1.665 $Y=2.4 $X2=0
+ $Y2=0
cc_127 N_A_29_424#_c_107_n N_VGND_c_364_n 0.0146184f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_128 N_A_29_424#_c_108_n N_VGND_c_364_n 0.0200379f $X=0.785 $Y=0.795 $X2=0
+ $Y2=0
cc_129 N_A_29_424#_c_111_n N_VGND_c_364_n 0.03064f $X=1.45 $Y=1.385 $X2=0 $Y2=0
cc_130 N_A_29_424#_c_114_n N_VGND_c_364_n 0.00684864f $X=1.68 $Y=1.385 $X2=0
+ $Y2=0
cc_131 N_A_29_424#_c_108_n N_VGND_c_366_n 0.00808397f $X=0.785 $Y=0.795 $X2=0
+ $Y2=0
cc_132 N_A_29_424#_c_107_n N_VGND_c_367_n 0.00383152f $X=1.68 $Y=1.22 $X2=0
+ $Y2=0
cc_133 N_A_29_424#_c_107_n N_VGND_c_369_n 0.00757637f $X=1.68 $Y=1.22 $X2=0
+ $Y2=0
cc_134 N_A_29_424#_c_108_n N_VGND_c_369_n 0.01059f $X=0.785 $Y=0.795 $X2=0 $Y2=0
cc_135 N_A1_M1004_g N_A2_M1003_g 0.0306283f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A1_c_182_n N_A2_M1003_g 0.00215789f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A1_M1000_g A2 6.65781e-19 $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A1_c_181_n A2 6.91666e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_c_182_n A2 0.0131385f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A1_c_181_n N_A2_c_223_n 0.0210016f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A1_c_182_n N_A2_c_223_n 0.00114066f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_A2_c_224_n 0.0399035f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1004_g N_VPWR_c_252_n 0.00995413f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A1_M1004_g N_VPWR_c_253_n 0.0050621f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A1_M1004_g N_VPWR_c_250_n 0.00998985f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A1_M1004_g N_Y_c_291_n 0.00338828f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A1_c_182_n N_Y_c_291_n 0.00491347f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_Y_c_288_n 2.25762e-19 $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A1_M1000_g N_Y_c_288_n 0.00174323f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A1_c_181_n N_Y_c_288_n 0.00204642f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A1_c_182_n N_Y_c_288_n 0.0271535f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A1_M1000_g N_Y_c_289_n 0.0130209f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1000_g N_Y_c_290_n 0.00480013f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_c_181_n N_Y_c_290_n 0.00315033f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A1_c_182_n N_Y_c_290_n 0.00106339f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A1_M1004_g N_A_351_368#_c_341_n 0.0161289f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A1_c_181_n N_A_351_368#_c_341_n 3.28371e-19 $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_158 N_A1_c_182_n N_A_351_368#_c_341_n 0.0113544f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A1_M1004_g N_A_351_368#_c_338_n 0.00110512f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A1_c_181_n N_A_351_368#_c_338_n 9.49345e-19 $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_161 N_A1_M1004_g N_A_351_368#_c_339_n 0.00120755f $X=2.115 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A1_M1000_g N_VGND_c_364_n 7.01115e-19 $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A1_M1000_g N_VGND_c_365_n 0.00253715f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_M1000_g N_VGND_c_367_n 0.00434272f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1000_g N_VGND_c_369_n 0.00821825f $X=2.11 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A2_M1003_g N_VPWR_c_252_n 0.0128939f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A2_M1003_g N_VPWR_c_256_n 0.0050621f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VPWR_c_250_n 0.0100324f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_169 A2 N_Y_c_288_n 0.00489165f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_c_224_n N_Y_c_289_n 0.00281399f $X=2.67 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A2_M1003_g N_A_351_368#_c_341_n 0.0149451f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_172 A2 N_A_351_368#_c_341_n 0.00440887f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A2_M1003_g N_A_351_368#_c_337_n 0.00101635f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A2_M1003_g N_A_351_368#_c_339_n 0.00845189f $X=2.595 $Y=2.4 $X2=0 $Y2=0
cc_175 A2 N_A_351_368#_c_339_n 0.0201859f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A2_c_223_n N_A_351_368#_c_339_n 0.00330217f $X=2.67 $Y=1.385 $X2=0
+ $Y2=0
cc_177 A2 N_VGND_c_365_n 0.0259407f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A2_c_223_n N_VGND_c_365_n 0.0011179f $X=2.67 $Y=1.385 $X2=0 $Y2=0
cc_179 N_A2_c_224_n N_VGND_c_365_n 0.0176088f $X=2.67 $Y=1.22 $X2=0 $Y2=0
cc_180 N_A2_c_224_n N_VGND_c_367_n 0.00383152f $X=2.67 $Y=1.22 $X2=0 $Y2=0
cc_181 N_A2_c_224_n N_VGND_c_369_n 0.00757998f $X=2.67 $Y=1.22 $X2=0 $Y2=0
cc_182 N_VPWR_c_251_n Y 0.062468f $X=0.72 $Y=2.28 $X2=0 $Y2=0
cc_183 N_VPWR_c_253_n Y 0.019544f $X=2.19 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_250_n Y 0.0161768f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_251_n N_Y_c_294_n 0.00186751f $X=0.72 $Y=2.28 $X2=0 $Y2=0
cc_186 N_VPWR_M1004_d N_A_351_368#_c_341_n 0.00820977f $X=2.205 $Y=1.84 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_252_n N_A_351_368#_c_341_n 0.0171814f $X=2.355 $Y=2.485 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_252_n N_A_351_368#_c_337_n 0.0225402f $X=2.355 $Y=2.485 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_256_n N_A_351_368#_c_337_n 0.0130739f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_250_n N_A_351_368#_c_337_n 0.0108215f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_252_n N_A_351_368#_c_338_n 0.0225402f $X=2.355 $Y=2.485 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_253_n N_A_351_368#_c_338_n 0.0129872f $X=2.19 $Y=3.33 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_250_n N_A_351_368#_c_338_n 0.0106816f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_Y_c_291_n N_A_351_368#_M1002_d 0.00136368f $X=1.705 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_195 N_Y_c_291_n N_A_351_368#_c_338_n 0.00817739f $X=1.705 $Y=1.805 $X2=0
+ $Y2=0
cc_196 Y N_A_351_368#_c_338_n 0.0249923f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_197 N_Y_c_289_n N_VGND_c_364_n 0.00662748f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_198 N_Y_c_290_n N_VGND_c_364_n 0.00229541f $X=1.882 $Y=1.18 $X2=0 $Y2=0
cc_199 N_Y_c_289_n N_VGND_c_365_n 0.0178888f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_200 N_Y_c_289_n N_VGND_c_367_n 0.0109942f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_201 N_Y_c_289_n N_VGND_c_369_n 0.00904371f $X=1.895 $Y=0.515 $X2=0 $Y2=0

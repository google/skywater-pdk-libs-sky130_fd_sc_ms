* File: sky130_fd_sc_ms__o21a_2.spice
* Created: Wed Sep  2 12:21:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21a_2.pex.spice"
.subckt sky130_fd_sc_ms__o21a_2  VNB VPB A1 A2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_54_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1702 AS=0.2627 PD=1.2 PS=2.19 NRD=12.156 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1005 N_A_54_74#_M1005_d N_A2_M1005_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.1702 PD=1.065 PS=1.2 NRD=7.296 NRS=17.016 M=1 R=4.93333
+ SA=75000.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1009 N_A_247_368#_M1009_d N_B1_M1009_g N_A_54_74#_M1005_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.12025 PD=2.19 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.4 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 N_X_M1003_d N_A_247_368#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1003_d N_A_247_368#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 A_163_368# N_A1_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90002.4
+ A=0.18 P=2.36 MULT=1
MM1001 N_A_247_368#_M1001_d N_A2_M1001_g A_163_368# VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.12 PD=1.39 PS=1.24 NRD=22.6353 NRS=12.7853 M=1 R=5.55556
+ SA=90000.6 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_A_247_368#_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.261509 AS=0.195 PD=1.53774 PS=1.39 NRD=36.7602 NRS=0 M=1 R=5.55556
+ SA=90001.2 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1002 N_X_M1002_d N_A_247_368#_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.292891 PD=1.39 PS=1.72226 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.7 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1004 N_X_M1002_d N_A_247_368#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o21a_2.pxi.spice"
*
.ends
*
*

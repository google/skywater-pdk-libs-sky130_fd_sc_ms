* File: sky130_fd_sc_ms__ha_4.pex.spice
* Created: Wed Sep  2 12:10:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__HA_4%A_435_99# 1 2 3 10 12 13 14 15 17 20 24 28 32
+ 36 40 44 48 52 56 58 61 65 69 72 74 75 80 84 87 100
c188 74 0 1.09796e-19 $X=5.965 $Y=1.82
c189 10 0 1.8401e-19 $X=2.25 $Y=1.34
r190 100 101 11.2969 $w=3.2e-07 $l=7.5e-08 $layer=POLY_cond $X=7.515 $Y=1.485
+ $X2=7.59 $Y2=1.485
r191 99 100 53.4719 $w=3.2e-07 $l=3.55e-07 $layer=POLY_cond $X=7.16 $Y=1.485
+ $X2=7.515 $Y2=1.485
r192 98 99 14.3094 $w=3.2e-07 $l=9.5e-08 $layer=POLY_cond $X=7.065 $Y=1.485
+ $X2=7.16 $Y2=1.485
r193 95 96 17.3219 $w=3.2e-07 $l=1.15e-07 $layer=POLY_cond $X=6.615 $Y=1.485
+ $X2=6.73 $Y2=1.485
r194 94 95 47.4469 $w=3.2e-07 $l=3.15e-07 $layer=POLY_cond $X=6.3 $Y=1.485
+ $X2=6.615 $Y2=1.485
r195 84 86 0.122819 $w=2.98e-07 $l=3e-09 $layer=LI1_cond $X=4.07 $Y=1.907
+ $X2=4.07 $Y2=1.91
r196 83 84 13.7966 $w=2.98e-07 $l=3.37e-07 $layer=LI1_cond $X=4.07 $Y=1.57
+ $X2=4.07 $Y2=1.907
r197 81 98 41.4219 $w=3.2e-07 $l=2.75e-07 $layer=POLY_cond $X=6.79 $Y=1.485
+ $X2=7.065 $Y2=1.485
r198 81 96 9.0375 $w=3.2e-07 $l=6e-08 $layer=POLY_cond $X=6.79 $Y=1.485 $X2=6.73
+ $Y2=1.485
r199 80 81 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=1.485 $X2=6.79 $Y2=1.485
r200 78 94 28.6187 $w=3.2e-07 $l=1.9e-07 $layer=POLY_cond $X=6.11 $Y=1.485
+ $X2=6.3 $Y2=1.485
r201 78 92 15.8156 $w=3.2e-07 $l=1.05e-07 $layer=POLY_cond $X=6.11 $Y=1.485
+ $X2=6.005 $Y2=1.485
r202 77 80 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.11 $Y=1.485
+ $X2=6.79 $Y2=1.485
r203 77 78 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.485 $X2=6.11 $Y2=1.485
r204 75 77 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=6.05 $Y=1.485
+ $X2=6.11 $Y2=1.485
r205 73 75 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.965 $Y=1.65
+ $X2=6.05 $Y2=1.485
r206 73 74 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.965 $Y=1.65
+ $X2=5.965 $Y2=1.82
r207 72 87 8.29065 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.12 $Y=1.985
+ $X2=4.955 $Y2=1.985
r208 69 74 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.88 $Y=1.985
+ $X2=5.965 $Y2=1.82
r209 69 72 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.88 $Y=1.985
+ $X2=5.12 $Y2=1.985
r210 68 84 3.87205 $w=1.75e-07 $l=1.6e-07 $layer=LI1_cond $X=4.23 $Y=1.907
+ $X2=4.07 $Y2=1.907
r211 68 87 45.9481 $w=1.73e-07 $l=7.25e-07 $layer=LI1_cond $X=4.23 $Y=1.907
+ $X2=4.955 $Y2=1.907
r212 63 83 6.24057 $w=3.3e-07 $l=1.86145e-07 $layer=LI1_cond $X=4.115 $Y=1.405
+ $X2=4.07 $Y2=1.57
r213 63 65 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=4.115 $Y=1.405
+ $X2=4.115 $Y2=0.74
r214 61 91 10.2408 $w=3.53e-07 $l=7.5e-08 $layer=POLY_cond $X=3.24 $Y=1.537
+ $X2=3.315 $Y2=1.537
r215 61 89 51.204 $w=3.53e-07 $l=3.75e-07 $layer=POLY_cond $X=3.24 $Y=1.537
+ $X2=2.865 $Y2=1.537
r216 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.57 $X2=3.24 $Y2=1.57
r217 58 83 0.0845041 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=3.9 $Y=1.57
+ $X2=4.07 $Y2=1.57
r218 58 60 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=3.9 $Y=1.57
+ $X2=3.24 $Y2=1.57
r219 54 101 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.59 $Y=1.32
+ $X2=7.59 $Y2=1.485
r220 54 56 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.59 $Y=1.32
+ $X2=7.59 $Y2=0.74
r221 50 100 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.515 $Y=1.65
+ $X2=7.515 $Y2=1.485
r222 50 52 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.515 $Y=1.65
+ $X2=7.515 $Y2=2.4
r223 46 99 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.16 $Y=1.32
+ $X2=7.16 $Y2=1.485
r224 46 48 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.16 $Y=1.32
+ $X2=7.16 $Y2=0.74
r225 42 98 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.065 $Y=1.65
+ $X2=7.065 $Y2=1.485
r226 42 44 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.065 $Y=1.65
+ $X2=7.065 $Y2=2.4
r227 38 96 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.73 $Y=1.32
+ $X2=6.73 $Y2=1.485
r228 38 40 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.73 $Y=1.32
+ $X2=6.73 $Y2=0.74
r229 34 95 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.615 $Y=1.65
+ $X2=6.615 $Y2=1.485
r230 34 36 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.615 $Y=1.65
+ $X2=6.615 $Y2=2.4
r231 30 94 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.3 $Y=1.32
+ $X2=6.3 $Y2=1.485
r232 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.3 $Y=1.32 $X2=6.3
+ $Y2=0.74
r233 26 92 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.005 $Y=1.65
+ $X2=6.005 $Y2=1.485
r234 26 28 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.005 $Y=1.65
+ $X2=6.005 $Y2=2.4
r235 22 91 18.5072 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=3.315 $Y=1.735
+ $X2=3.315 $Y2=1.537
r236 22 24 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.315 $Y=1.735
+ $X2=3.315 $Y2=2.315
r237 18 89 18.5072 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=2.865 $Y=1.735
+ $X2=2.865 $Y2=1.537
r238 18 20 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.865 $Y=1.735
+ $X2=2.865 $Y2=2.315
r239 15 89 19.7989 $w=3.53e-07 $l=2.59565e-07 $layer=POLY_cond $X=2.72 $Y=1.34
+ $X2=2.865 $Y2=1.537
r240 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.72 $Y=1.34
+ $X2=2.72 $Y2=0.945
r241 13 15 26.5307 $w=3.53e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.645 $Y=1.415
+ $X2=2.72 $Y2=1.34
r242 13 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.645 $Y=1.415
+ $X2=2.325 $Y2=1.415
r243 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.325 $Y2=1.415
r244 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.25 $Y2=0.945
r245 3 72 600 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=2.05 $X2=5.12 $Y2=1.985
r246 2 86 600 $w=1.7e-07 $l=2.17371e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.895 $X2=4.065 $Y2=1.91
r247 1 65 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.975
+ $Y=0.595 $X2=4.115 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%B 3 5 7 10 12 14 15 16 18 19 20 24 27 29 31 35
+ 39 41 42 43 44
c123 44 0 1.898e-19 $X=2.16 $Y=1.665
c124 39 0 6.08632e-20 $X=4.37 $Y=2.47
c125 12 0 7.39997e-20 $X=1.845 $Y=1.88
c126 5 0 3.95329e-20 $X=1.395 $Y=1.88
c127 3 0 1.44963e-19 $X=1.36 $Y=0.945
r128 52 53 6.3726 $w=4.16e-07 $l=5.5e-08 $layer=POLY_cond $X=1.79 $Y=1.667
+ $X2=1.845 $Y2=1.667
r129 50 52 6.95192 $w=4.16e-07 $l=6e-08 $layer=POLY_cond $X=1.73 $Y=1.667
+ $X2=1.79 $Y2=1.667
r130 48 50 38.8149 $w=4.16e-07 $l=3.35e-07 $layer=POLY_cond $X=1.395 $Y=1.667
+ $X2=1.73 $Y2=1.667
r131 47 48 4.05529 $w=4.16e-07 $l=3.5e-08 $layer=POLY_cond $X=1.36 $Y=1.667
+ $X2=1.395 $Y2=1.667
r132 43 44 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.62
+ $X2=2.16 $Y2=1.62
r133 43 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.62 $X2=1.73 $Y2=1.62
r134 37 39 235.169 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=4.37 $Y=3.075
+ $X2=4.37 $Y2=2.47
r135 33 35 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.33 $Y=1.53
+ $X2=4.33 $Y2=0.915
r136 32 41 6.66866 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.975 $Y=1.605
+ $X2=3.825 $Y2=1.605
r137 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.255 $Y=1.605
+ $X2=4.33 $Y2=1.53
r138 31 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.255 $Y=1.605
+ $X2=3.975 $Y2=1.605
r139 30 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=3.15
+ $X2=3.765 $Y2=3.15
r140 29 37 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.28 $Y=3.15
+ $X2=4.37 $Y2=3.075
r141 29 30 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.28 $Y=3.15
+ $X2=3.855 $Y2=3.15
r142 25 41 18.8402 $w=1.65e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.9 $Y=1.53
+ $X2=3.825 $Y2=1.605
r143 25 27 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.9 $Y=1.53
+ $X2=3.9 $Y2=0.915
r144 22 42 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=3.075
+ $X2=3.765 $Y2=3.15
r145 22 24 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=3.765 $Y=3.075
+ $X2=3.765 $Y2=2.315
r146 21 41 18.8402 $w=1.65e-07 $l=1.00623e-07 $layer=POLY_cond $X=3.765 $Y=1.68
+ $X2=3.825 $Y2=1.605
r147 21 24 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=3.765 $Y=1.68
+ $X2=3.765 $Y2=2.315
r148 19 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.675 $Y=3.15
+ $X2=3.765 $Y2=3.15
r149 19 20 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=3.675 $Y=3.15
+ $X2=2.43 $Y2=3.15
r150 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.355 $Y=3.075
+ $X2=2.43 $Y2=3.15
r151 17 18 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=2.355 $Y=1.88
+ $X2=2.355 $Y2=3.075
r152 16 53 31.2225 $w=4.16e-07 $l=1.77381e-07 $layer=POLY_cond $X=1.935 $Y=1.805
+ $X2=1.845 $Y2=1.667
r153 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.28 $Y=1.805
+ $X2=2.355 $Y2=1.88
r154 15 16 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.28 $Y=1.805
+ $X2=1.935 $Y2=1.805
r155 12 53 22.3993 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=1.845 $Y=1.88
+ $X2=1.845 $Y2=1.667
r156 12 14 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.845 $Y=1.88
+ $X2=1.845 $Y2=2.46
r157 8 52 26.8236 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=1.79 $Y=1.455
+ $X2=1.79 $Y2=1.667
r158 8 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.79 $Y=1.455
+ $X2=1.79 $Y2=0.945
r159 5 48 22.3993 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=1.395 $Y=1.88
+ $X2=1.395 $Y2=1.667
r160 5 7 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.395 $Y=1.88
+ $X2=1.395 $Y2=2.46
r161 1 47 26.8236 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=1.36 $Y=1.455
+ $X2=1.36 $Y2=1.667
r162 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.36 $Y=1.455
+ $X2=1.36 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%A 3 7 12 13 15 16 17 20 25 26 28 30 33 35 36 37
+ 38 39 47
c113 47 0 1.898e-19 $X=0.93 $Y=1.665
c114 28 0 1.39181e-20 $X=5.33 $Y=1.31
c115 13 0 5.44618e-20 $X=0.945 $Y=1.875
c116 3 0 2.18257e-19 $X=0.495 $Y=2.46
r117 47 48 2.12647 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=0.93 $Y=1.665
+ $X2=0.945 $Y2=1.665
r118 45 47 29.0618 $w=3.4e-07 $l=2.05e-07 $layer=POLY_cond $X=0.725 $Y=1.665
+ $X2=0.93 $Y2=1.665
r119 38 39 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.62
+ $X2=1.2 $Y2=1.62
r120 38 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.62 $X2=0.725 $Y2=1.62
r121 37 38 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.62
+ $X2=0.72 $Y2=1.62
r122 31 36 33.9972 $w=1.65e-07 $l=3.62215e-07 $layer=POLY_cond $X=5.345 $Y=1.63
+ $X2=5.255 $Y2=1.31
r123 31 33 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=5.345 $Y=1.63
+ $X2=5.345 $Y2=2.26
r124 28 36 33.9972 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=5.33 $Y=1.31
+ $X2=5.255 $Y2=1.31
r125 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.33 $Y=1.31
+ $X2=5.33 $Y2=0.915
r126 27 35 3.5291 $w=3.2e-07 $l=1.84932e-07 $layer=POLY_cond $X=4.91 $Y=1.47
+ $X2=4.73 $Y2=1.46
r127 26 36 3.5291 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=5.255 $Y=1.47
+ $X2=5.255 $Y2=1.31
r128 26 27 62.2124 $w=3.2e-07 $l=3.45e-07 $layer=POLY_cond $X=5.255 $Y=1.47
+ $X2=4.91 $Y2=1.47
r129 23 35 33.9972 $w=1.65e-07 $l=1.93649e-07 $layer=POLY_cond $X=4.83 $Y=1.31
+ $X2=4.73 $Y2=1.46
r130 23 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.83 $Y=1.31
+ $X2=4.83 $Y2=0.915
r131 22 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.83 $Y2=0.915
r132 18 35 33.9972 $w=1.65e-07 $l=2.10238e-07 $layer=POLY_cond $X=4.82 $Y=1.63
+ $X2=4.73 $Y2=1.46
r133 18 20 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=4.82 $Y=1.63
+ $X2=4.82 $Y2=2.47
r134 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.755 $Y=0.18
+ $X2=4.83 $Y2=0.255
r135 16 17 1922.87 $w=1.5e-07 $l=3.75e-06 $layer=POLY_cond $X=4.755 $Y=0.18
+ $X2=1.005 $Y2=0.18
r136 13 48 17.6285 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.945 $Y=1.875
+ $X2=0.945 $Y2=1.665
r137 13 15 156.65 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=0.945 $Y=1.875
+ $X2=0.945 $Y2=2.46
r138 10 47 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.93 $Y=1.455
+ $X2=0.93 $Y2=1.665
r139 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.93 $Y=1.455
+ $X2=0.93 $Y2=0.945
r140 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=0.255
+ $X2=1.005 $Y2=0.18
r141 9 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.93 $Y=0.255
+ $X2=0.93 $Y2=0.945
r142 5 7 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.495 $Y=1.455
+ $X2=0.495 $Y2=0.945
r143 1 45 32.6059 $w=3.4e-07 $l=2.3e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.725 $Y2=1.665
r144 1 5 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.495 $Y2=1.455
r145 1 3 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=0.495 $Y=1.785
+ $X2=0.495 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%A_297_392# 1 2 3 12 16 20 24 28 32 34 35 38 42
+ 46 50 53 54 56 58 61 62 67 68 71 72 73 76 78
c200 71 0 5.44618e-20 $X=1.62 $Y=2.12
c201 61 0 5.29972e-20 $X=7.81 $Y=2.32
c202 53 0 1.00633e-19 $X=2.585 $Y=1.905
c203 35 0 9.40988e-20 $X=9.025 $Y=1.485
c204 12 0 1.7493e-19 $X=7.965 $Y=2.4
r205 88 89 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=8.865 $Y=1.485
+ $X2=8.95 $Y2=1.485
r206 87 88 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.45 $Y=1.485
+ $X2=8.865 $Y2=1.485
r207 86 87 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.415 $Y=1.485
+ $X2=8.45 $Y2=1.485
r208 82 84 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=7.965 $Y=1.485
+ $X2=8.02 $Y2=1.485
r209 78 80 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.985 $Y=2.25
+ $X2=3.985 $Y2=2.405
r210 76 77 7.52055 $w=2.92e-07 $l=1.8e-07 $layer=LI1_cond $X=3.09 $Y=2.07
+ $X2=3.09 $Y2=2.25
r211 74 76 2.29795 $w=2.92e-07 $l=5.5e-08 $layer=LI1_cond $X=3.09 $Y=2.015
+ $X2=3.09 $Y2=2.07
r212 67 68 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.56
+ $Y=1.485 $X2=9.56 $Y2=1.485
r213 65 86 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=8.04 $Y=1.485
+ $X2=8.415 $Y2=1.485
r214 65 84 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.04 $Y=1.485
+ $X2=8.02 $Y2=1.485
r215 64 67 53.0822 $w=3.28e-07 $l=1.52e-06 $layer=LI1_cond $X=8.04 $Y=1.485
+ $X2=9.56 $Y2=1.485
r216 64 65 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.04
+ $Y=1.485 $X2=8.04 $Y2=1.485
r217 62 64 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.895 $Y=1.485
+ $X2=8.04 $Y2=1.485
r218 60 62 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.81 $Y=1.65
+ $X2=7.895 $Y2=1.485
r219 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.81 $Y=1.65
+ $X2=7.81 $Y2=2.32
r220 59 80 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.405
+ $X2=3.985 $Y2=2.405
r221 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.725 $Y=2.405
+ $X2=7.81 $Y2=2.32
r222 58 59 238.455 $w=1.68e-07 $l=3.655e-06 $layer=LI1_cond $X=7.725 $Y=2.405
+ $X2=4.07 $Y2=2.405
r223 57 77 3.90229 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.25
+ $X2=3.09 $Y2=2.25
r224 56 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=2.25
+ $X2=3.985 $Y2=2.25
r225 56 57 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.9 $Y=2.25
+ $X2=3.255 $Y2=2.25
r226 55 73 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.015
+ $X2=2.585 $Y2=2.015
r227 54 74 2.3974 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=2.015
+ $X2=3.09 $Y2=2.015
r228 54 55 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.925 $Y=2.015
+ $X2=2.67 $Y2=2.015
r229 53 73 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.585 $Y=1.905
+ $X2=2.585 $Y2=2.015
r230 53 72 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.585 $Y=1.905
+ $X2=2.585 $Y2=1.285
r231 48 72 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.12
+ $X2=2.505 $Y2=1.285
r232 48 50 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.505 $Y=1.12
+ $X2=2.505 $Y2=0.77
r233 47 71 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.735 $Y=2.04
+ $X2=1.595 $Y2=2.04
r234 46 73 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=2.5 $Y=2.04
+ $X2=2.585 $Y2=2.015
r235 46 47 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.5 $Y=2.04
+ $X2=1.735 $Y2=2.04
r236 40 68 34.7346 $w=1.65e-07 $l=1.65997e-07 $layer=POLY_cond $X=9.575 $Y=1.65
+ $X2=9.577 $Y2=1.485
r237 40 42 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=9.575 $Y=1.65
+ $X2=9.575 $Y2=2.4
r238 36 68 34.7346 $w=1.65e-07 $l=1.9775e-07 $layer=POLY_cond $X=9.505 $Y=1.32
+ $X2=9.577 $Y2=1.485
r239 36 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.505 $Y=1.32
+ $X2=9.505 $Y2=0.74
r240 35 89 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.025 $Y=1.485
+ $X2=8.95 $Y2=1.485
r241 34 68 3.90195 $w=3.3e-07 $l=1.47e-07 $layer=POLY_cond $X=9.43 $Y=1.485
+ $X2=9.577 $Y2=1.485
r242 34 35 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=9.43 $Y=1.485
+ $X2=9.025 $Y2=1.485
r243 30 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.95 $Y=1.32
+ $X2=8.95 $Y2=1.485
r244 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.95 $Y=1.32
+ $X2=8.95 $Y2=0.74
r245 26 88 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.865 $Y=1.65
+ $X2=8.865 $Y2=1.485
r246 26 28 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.865 $Y=1.65
+ $X2=8.865 $Y2=2.4
r247 22 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.45 $Y=1.32
+ $X2=8.45 $Y2=1.485
r248 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.45 $Y=1.32
+ $X2=8.45 $Y2=0.74
r249 18 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.415 $Y=1.65
+ $X2=8.415 $Y2=1.485
r250 18 20 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.415 $Y=1.65
+ $X2=8.415 $Y2=2.4
r251 14 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.02 $Y=1.32
+ $X2=8.02 $Y2=1.485
r252 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.02 $Y=1.32
+ $X2=8.02 $Y2=0.74
r253 10 82 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.965 $Y=1.65
+ $X2=7.965 $Y2=1.485
r254 10 12 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.965 $Y=1.65
+ $X2=7.965 $Y2=2.4
r255 3 76 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.895 $X2=3.09 $Y2=2.07
r256 2 71 300 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.96 $X2=1.62 $Y2=2.12
r257 1 50 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.625 $X2=2.505 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%A_27_392# 1 2 3 10 12 14 16 19 20 21 24
c41 21 0 1.01045e-19 $X=1.255 $Y=2.99
c42 16 0 3.95329e-20 $X=1.13 $Y=2.125
c43 12 0 1.17212e-19 $X=0.27 $Y=2.8
r44 22 24 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=2.38
r45 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=2.07 $Y2=2.905
r46 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=1.255 $Y2=2.99
r47 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.13 $Y=2.905
+ $X2=1.255 $Y2=2.99
r48 17 19 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.13 $Y=2.905 $X2=1.13
+ $Y2=2.815
r49 16 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=2.125
+ $X2=1.13 $Y2=2.04
r50 16 19 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=1.13 $Y=2.125
+ $X2=1.13 $Y2=2.815
r51 15 27 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.385 $Y=2.04
+ $X2=0.245 $Y2=2.04
r52 14 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=2.04
+ $X2=1.13 $Y2=2.04
r53 14 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.005 $Y=2.04
+ $X2=0.385 $Y2=2.04
r54 10 27 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.125
+ $X2=0.245 $Y2=2.04
r55 10 12 27.7821 $w=2.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.245 $Y=2.125
+ $X2=0.245 $Y2=2.8
r56 3 24 300 $w=1.7e-07 $l=4.82804e-07 $layer=licon1_PDIFF $count=2 $X=1.935
+ $Y=1.96 $X2=2.07 $Y2=2.38
r57 2 29 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.96 $X2=1.17 $Y2=2.12
r58 2 19 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.96 $X2=1.17 $Y2=2.815
r59 1 27 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.27 $Y2=2.12
r60 1 12 400 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.27 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 44 48 52 56
+ 60 62 64 67 68 70 71 73 74 75 77 82 90 95 110 115 118 121 124 127 131
c151 34 0 7.39997e-20 $X=2.64 $Y=2.57
c152 2 0 1.00633e-19 $X=2.505 $Y=1.895
r153 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r154 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r155 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r157 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r158 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r159 113 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r160 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 110 130 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.857 $Y2=3.33
r162 110 112 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r164 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r165 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r166 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r167 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r168 103 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r169 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r170 100 127 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=5.717 $Y2=3.33
r171 100 102 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=6.48 $Y2=3.33
r172 99 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r173 99 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r174 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 96 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.54 $Y2=3.33
r176 96 98 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r177 95 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.595 $Y2=3.33
r178 95 98 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r179 94 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r180 94 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r181 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r182 91 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r183 91 93 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=3.12 $Y2=3.33
r184 90 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.54 $Y2=3.33
r185 90 93 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r186 89 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r187 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r188 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r189 86 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r190 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r191 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r192 83 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.68 $Y2=3.33
r193 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 82 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.64 $Y2=3.33
r195 82 88 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.16 $Y2=3.33
r196 80 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r197 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r198 77 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.68 $Y2=3.33
r199 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r200 75 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r201 75 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 73 108 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=8.475 $Y=3.33
+ $X2=8.4 $Y2=3.33
r203 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.475 $Y=3.33
+ $X2=8.64 $Y2=3.33
r204 72 112 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=9.36 $Y2=3.33
r205 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=8.64 $Y2=3.33
r206 70 105 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.44 $Y2=3.33
r207 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=3.33
+ $X2=7.74 $Y2=3.33
r208 69 108 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=7.74 $Y2=3.33
r210 67 102 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.48 $Y2=3.33
r211 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.84 $Y2=3.33
r212 66 105 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.005 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=3.33
+ $X2=6.84 $Y2=3.33
r214 62 130 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.857 $Y2=3.33
r215 62 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.415
r216 58 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.64 $Y=3.245
+ $X2=8.64 $Y2=3.33
r217 58 60 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.64 $Y=3.245
+ $X2=8.64 $Y2=2.405
r218 54 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.74 $Y=3.245
+ $X2=7.74 $Y2=3.33
r219 54 56 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.74 $Y=3.245
+ $X2=7.74 $Y2=2.78
r220 50 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=3.245
+ $X2=6.84 $Y2=3.33
r221 50 52 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.84 $Y=3.245
+ $X2=6.84 $Y2=2.78
r222 46 127 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.717 $Y=3.245
+ $X2=5.717 $Y2=3.33
r223 46 48 13.1437 $w=4.53e-07 $l=5e-07 $layer=LI1_cond $X=5.717 $Y=3.245
+ $X2=5.717 $Y2=2.745
r224 45 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=4.595 $Y2=3.33
r225 44 127 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.717 $Y2=3.33
r226 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=4.76 $Y2=3.33
r227 40 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=3.33
r228 40 42 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=2.745
r229 36 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=3.33
r230 36 38 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=2.59
r231 32 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=3.245
+ $X2=2.64 $Y2=3.33
r232 32 34 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.64 $Y=3.245
+ $X2=2.64 $Y2=2.57
r233 28 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=3.33
r234 28 30 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=2.46
r235 9 64 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=2.415
r236 8 60 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=8.505
+ $Y=1.84 $X2=8.64 $Y2=2.405
r237 7 56 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=7.605
+ $Y=1.84 $X2=7.74 $Y2=2.78
r238 6 52 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=6.705
+ $Y=1.84 $X2=6.84 $Y2=2.78
r239 5 48 600 $w=1.7e-07 $l=1.03558e-06 $layer=licon1_PDIFF $count=1 $X=5.435
+ $Y=1.84 $X2=5.715 $Y2=2.745
r240 4 42 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=2.05 $X2=4.595 $Y2=2.745
r241 3 38 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.895 $X2=3.54 $Y2=2.59
r242 2 34 600 $w=1.7e-07 $l=7.39425e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.895 $X2=2.64 $Y2=2.57
r243 1 30 300 $w=1.7e-07 $l=5.63471e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.96 $X2=0.72 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%COUT 1 2 3 4 13 17 19 21 25 28 29 30 34
c51 28 0 9.9062e-20 $X=7.44 $Y=1.295
r52 30 34 3.3396 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=7.382 $Y=1.985
+ $X2=7.382 $Y2=1.82
r53 29 34 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=7.382 $Y=1.665
+ $X2=7.382 $Y2=1.82
r54 28 29 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=7.382 $Y=1.295
+ $X2=7.382 $Y2=1.665
r55 25 28 5.51168 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.382 $Y=1.13
+ $X2=7.382 $Y2=1.295
r56 25 27 2.96505 $w=3.45e-07 $l=1.25e-07 $layer=LI1_cond $X=7.382 $Y=1.13
+ $X2=7.382 $Y2=1.005
r57 22 24 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.6 $Y=1.005
+ $X2=6.475 $Y2=1.005
r58 21 27 4.07991 $w=2.5e-07 $l=1.72e-07 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=7.382 $Y2=1.005
r59 21 22 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=6.6 $Y2=1.005
r60 17 24 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=0.88
+ $X2=6.475 $Y2=1.005
r61 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=6.475 $Y=0.88
+ $X2=6.475 $Y2=0.515
r62 13 30 3.48128 $w=3.3e-07 $l=1.72e-07 $layer=LI1_cond $X=7.21 $Y=1.985
+ $X2=7.382 $Y2=1.985
r63 13 15 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=7.21 $Y=1.985
+ $X2=6.385 $Y2=1.985
r64 4 30 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.155
+ $Y=1.84 $X2=7.29 $Y2=1.985
r65 3 15 600 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=1 $X=6.095
+ $Y=1.84 $X2=6.385 $Y2=1.985
r66 2 27 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.235
+ $Y=0.37 $X2=7.375 $Y2=0.965
r67 1 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.375
+ $Y=0.37 $X2=6.515 $Y2=0.965
r68 1 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.375
+ $Y=0.37 $X2=6.515 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%SUM 1 2 3 4 13 15 19 21 22 25 29 31 33 36 40 41
+ 43 44 45 50
c89 13 0 1.7493e-19 $X=8.19 $Y=2.15
r90 50 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=2.035
+ $X2=9.84 $Y2=2.035
r91 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r92 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.025 $Y=2.035
+ $X2=8.88 $Y2=2.035
r93 44 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=9.84 $Y2=2.035
r94 44 45 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=9.025 $Y2=2.035
r95 41 48 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=9.075 $Y=1.985
+ $X2=8.88 $Y2=1.985
r96 41 43 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=1.985
+ $X2=9.24 $Y2=1.985
r97 37 48 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=8.305 $Y=1.985
+ $X2=8.88 $Y2=1.985
r98 37 39 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=8.305 $Y=1.985
+ $X2=8.19 $Y2=1.985
r99 36 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.91 $Y=1.82
+ $X2=9.91 $Y2=1.985
r100 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.91 $Y=1.15
+ $X2=9.91 $Y2=1.82
r101 34 43 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.405 $Y=1.985
+ $X2=9.24 $Y2=1.985
r102 33 54 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.825 $Y=1.985
+ $X2=9.91 $Y2=1.985
r103 33 34 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.825 $Y=1.985
+ $X2=9.405 $Y2=1.985
r104 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.4 $Y=1.065
+ $X2=9.235 $Y2=1.065
r105 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.825 $Y=1.065
+ $X2=9.91 $Y2=1.15
r106 31 32 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.825 $Y=1.065
+ $X2=9.4 $Y2=1.065
r107 27 43 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.24 $Y=2.15
+ $X2=9.24 $Y2=1.985
r108 27 29 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=9.24 $Y=2.15
+ $X2=9.24 $Y2=2.43
r109 23 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.235 $Y=0.98
+ $X2=9.235 $Y2=1.065
r110 23 25 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.235 $Y=0.98
+ $X2=9.235 $Y2=0.515
r111 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.07 $Y=1.065
+ $X2=9.235 $Y2=1.065
r112 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.07 $Y=1.065
+ $X2=8.4 $Y2=1.065
r113 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.275 $Y=0.98
+ $X2=8.4 $Y2=1.065
r114 17 19 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.275 $Y=0.98
+ $X2=8.275 $Y2=0.515
r115 13 39 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=2.15
+ $X2=8.19 $Y2=1.985
r116 13 15 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=8.19 $Y=2.15
+ $X2=8.19 $Y2=2.43
r117 4 43 600 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_PDIFF $count=1 $X=8.955
+ $Y=1.84 $X2=9.24 $Y2=1.985
r118 4 29 300 $w=1.7e-07 $l=7.18505e-07 $layer=licon1_PDIFF $count=2 $X=8.955
+ $Y=1.84 $X2=9.24 $Y2=2.43
r119 3 39 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.055
+ $Y=1.84 $X2=8.19 $Y2=1.985
r120 3 15 300 $w=1.7e-07 $l=6.54026e-07 $layer=licon1_PDIFF $count=2 $X=8.055
+ $Y=1.84 $X2=8.19 $Y2=2.43
r121 2 25 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.025
+ $Y=0.37 $X2=9.235 $Y2=0.515
r122 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.095
+ $Y=0.37 $X2=8.235 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%A_27_125# 1 2 3 4 15 17 18 21 23 28 29 30 33 35
c66 23 0 1.8401e-19 $X=1.84 $Y=1.2
c67 21 0 1.44963e-19 $X=1.145 $Y=0.77
r68 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.005 $Y=0.435
+ $X2=3.005 $Y2=0.77
r69 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.84 $Y=0.35
+ $X2=3.005 $Y2=0.435
r70 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=0.35
+ $X2=2.17 $Y2=0.35
r71 26 28 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.005 $Y=1.115
+ $X2=2.005 $Y2=0.77
r72 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.005 $Y=0.435
+ $X2=2.17 $Y2=0.35
r73 25 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.005 $Y=0.435
+ $X2=2.005 $Y2=0.77
r74 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.23 $Y=1.2
+ $X2=1.105 $Y2=1.2
r75 23 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.84 $Y=1.2
+ $X2=2.005 $Y2=1.115
r76 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.84 $Y=1.2 $X2=1.23
+ $Y2=1.2
r77 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=1.115
+ $X2=1.105 $Y2=1.2
r78 19 21 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=1.105 $Y=1.115
+ $X2=1.105 $Y2=0.77
r79 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.98 $Y=1.2
+ $X2=1.105 $Y2=1.2
r80 17 18 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.98 $Y=1.2
+ $X2=0.365 $Y2=1.2
r81 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.115
+ $X2=0.365 $Y2=1.2
r82 13 15 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.115
+ $X2=0.24 $Y2=0.77
r83 4 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.795
+ $Y=0.625 $X2=3.005 $Y2=0.77
r84 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.625 $X2=2.005 $Y2=0.77
r85 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.625 $X2=1.145 $Y2=0.77
r86 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%VGND 1 2 3 4 5 6 7 8 27 31 35 37 41 45 49 53 55
+ 57 60 61 63 64 66 67 69 70 71 80 87 99 104 107 110 114
c126 49 0 9.40988e-20 $X=7.805 $Y=0.53
r127 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r128 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r129 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r130 102 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r131 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r132 99 113 4.36388 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=9.58 $Y=0 $X2=9.83
+ $Y2=0
r133 99 101 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.58 $Y=0 $X2=9.36
+ $Y2=0
r134 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r135 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r136 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r137 95 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r138 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r139 92 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.11 $Y=0
+ $X2=6.945 $Y2=0
r140 92 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.44
+ $Y2=0
r141 91 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r142 91 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r143 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r144 88 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.17 $Y=0
+ $X2=6.045 $Y2=0
r145 88 90 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.48
+ $Y2=0
r146 87 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=0
+ $X2=6.945 $Y2=0
r147 87 90 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.78 $Y=0 $X2=6.48
+ $Y2=0
r148 85 86 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r149 83 86 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=4.56 $Y2=0
r150 82 85 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=4.56
+ $Y2=0
r151 82 83 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r152 80 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.95 $Y=0
+ $X2=5.115 $Y2=0
r153 80 85 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.95 $Y=0 $X2=4.56
+ $Y2=0
r154 79 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r155 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r156 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r157 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r158 71 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r159 71 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r160 71 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r161 69 97 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.57 $Y=0 $X2=8.4
+ $Y2=0
r162 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=0 $X2=8.735
+ $Y2=0
r163 68 101 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.9 $Y=0 $X2=9.36
+ $Y2=0
r164 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.9 $Y=0 $X2=8.735
+ $Y2=0
r165 66 94 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.44
+ $Y2=0
r166 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.805
+ $Y2=0
r167 65 97 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.97 $Y=0 $X2=8.4
+ $Y2=0
r168 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.97 $Y=0 $X2=7.805
+ $Y2=0
r169 63 78 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.2
+ $Y2=0
r170 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.535
+ $Y2=0
r171 62 82 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.68
+ $Y2=0
r172 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.535
+ $Y2=0
r173 60 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r174 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r175 59 78 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r176 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r177 55 113 3.19436 $w=3.05e-07 $l=1.33918e-07 $layer=LI1_cond $X=9.732 $Y=0.085
+ $X2=9.83 $Y2=0
r178 55 57 21.1596 $w=3.03e-07 $l=5.6e-07 $layer=LI1_cond $X=9.732 $Y=0.085
+ $X2=9.732 $Y2=0.645
r179 51 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0
r180 51 53 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.735 $Y=0.085
+ $X2=8.735 $Y2=0.58
r181 47 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.805 $Y=0.085
+ $X2=7.805 $Y2=0
r182 47 49 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.805 $Y=0.085
+ $X2=7.805 $Y2=0.53
r183 43 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.945 $Y=0.085
+ $X2=6.945 $Y2=0
r184 43 45 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.945 $Y=0.085
+ $X2=6.945 $Y2=0.53
r185 39 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=0.085
+ $X2=6.045 $Y2=0
r186 39 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.045 $Y=0.085
+ $X2=6.045 $Y2=0.515
r187 38 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.28 $Y=0
+ $X2=5.115 $Y2=0
r188 37 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.92 $Y=0
+ $X2=6.045 $Y2=0
r189 37 38 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=5.28
+ $Y2=0
r190 33 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0
r191 33 35 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.115 $Y=0.085
+ $X2=5.115 $Y2=0.74
r192 29 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0.085
+ $X2=1.535 $Y2=0
r193 29 31 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=1.535 $Y=0.085
+ $X2=1.535 $Y2=0.775
r194 25 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r195 25 27 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.775
r196 8 57 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.58
+ $Y=0.37 $X2=9.72 $Y2=0.645
r197 7 53 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=8.525
+ $Y=0.37 $X2=8.735 $Y2=0.58
r198 6 49 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=7.665
+ $Y=0.37 $X2=7.805 $Y2=0.53
r199 5 45 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.37 $X2=6.945 $Y2=0.53
r200 4 41 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.95
+ $Y=0.37 $X2=6.085 $Y2=0.515
r201 3 35 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.905
+ $Y=0.595 $X2=5.115 $Y2=0.74
r202 2 31 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.625 $X2=1.575 $Y2=0.775
r203 1 27 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.625 $X2=0.71 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__HA_4%A_707_119# 1 2 3 12 14 15 19 20 21 24
c52 21 0 6.08632e-20 $X=4.78 $Y=1.51
c53 14 0 1.39181e-20 $X=4.45 $Y=0.4
r54 22 24 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.585 $Y=1.425
+ $X2=5.585 $Y2=0.74
r55 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.46 $Y=1.51
+ $X2=5.585 $Y2=1.425
r56 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.46 $Y=1.51
+ $X2=4.78 $Y2=1.51
r57 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.615 $Y=1.425
+ $X2=4.78 $Y2=1.51
r58 17 19 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.615 $Y=1.425
+ $X2=4.615 $Y2=0.74
r59 16 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.615 $Y=0.485
+ $X2=4.615 $Y2=0.74
r60 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.45 $Y=0.4
+ $X2=4.615 $Y2=0.485
r61 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.45 $Y=0.4 $X2=3.78
+ $Y2=0.4
r62 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.65 $Y=0.485
+ $X2=3.78 $Y2=0.4
r63 10 12 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=3.65 $Y=0.485
+ $X2=3.65 $Y2=0.73
r64 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.405
+ $Y=0.595 $X2=5.545 $Y2=0.74
r65 2 19 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.405
+ $Y=0.595 $X2=4.615 $Y2=0.74
r66 1 12 91 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=2 $X=3.535
+ $Y=0.595 $X2=3.685 $Y2=0.73
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_643_74# a_219_424# a_571_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR a_219_424# a_363_74# VPB pshort w=840000u l=180000u
+  ad=1.4754e+12p pd=1.132e+07u as=2.352e+11p ps=2.24e+06u
M1002 VPWR RESET_B a_817_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1003 a_817_48# a_643_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Q a_817_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 a_762_508# a_363_74# a_643_74# VPB pshort w=420000u l=180000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1006 a_219_424# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=4.2675e+11p pd=2.84e+06u as=0p ps=0u
M1007 a_219_424# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=9.349e+11p ps=8.16e+06u
M1008 VPWR D a_27_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 VGND RESET_B a_1045_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1010 a_769_74# a_219_424# a_643_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.907e+11p ps=2.24e+06u
M1011 VGND a_817_48# a_769_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_219_424# a_363_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.2225e+11p ps=2.64e+06u
M1013 VPWR a_817_48# a_762_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q a_817_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1015 a_1045_74# a_643_74# a_817_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 a_571_392# a_27_424# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND D a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 a_565_74# a_27_424# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_643_74# a_363_74# a_565_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a22oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 1.350000 1.875000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.755000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.350000 1.335000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.624600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.010000 1.570000 1.180000 ;
        RECT 0.605000 1.180000 0.835000 1.950000 ;
        RECT 0.605000 1.950000 1.015000 2.120000 ;
        RECT 0.845000 2.120000 1.015000 2.735000 ;
        RECT 1.130000 0.350000 1.570000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.315000  2.290000 0.645000 2.905000 ;
      RECT 0.315000  2.905000 1.545000 3.075000 ;
      RECT 0.340000  0.085000 0.670000 0.840000 ;
      RECT 1.215000  1.950000 2.565000 2.120000 ;
      RECT 1.215000  2.120000 1.545000 2.905000 ;
      RECT 1.715000  2.290000 2.065000 3.245000 ;
      RECT 2.210000  0.085000 2.540000 1.130000 ;
      RECT 2.235000  2.120000 2.565000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_ms__a22oi_1
END LIBRARY

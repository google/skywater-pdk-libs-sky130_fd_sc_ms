* File: sky130_fd_sc_ms__and3b_4.spice
* Created: Fri Aug 28 17:13:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and3b_4.pex.spice"
.subckt sky130_fd_sc_ms__and3b_4  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_N_M1018_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1888 AS=0.1824 PD=1.87 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_239_98#_M1002_d N_A_27_74#_M1002_g N_A_301_368#_M1002_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1013 N_A_239_98#_M1013_d N_A_27_74#_M1013_g N_A_301_368#_M1002_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1010 N_A_239_98#_M1013_d N_B_M1010_g N_A_498_98#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1011 N_A_239_98#_M1011_d N_B_M1011_g N_A_498_98#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_498_98#_M1003_d N_C_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1009 N_A_498_98#_M1003_d N_C_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.12007 PD=0.92 PS=1.02029 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75000.6 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1009_s N_A_301_368#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13883 AS=0.1295 PD=1.17971 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_301_368#_M1007_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1295 PD=1.04 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1007_d N_A_301_368#_M1008_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1036 PD=1.04 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_301_368#_M1012_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.185 AS=0.28 PD=1.37 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90005.3 A=0.18 P=2.36 MULT=1
MM1016 N_A_301_368#_M1016_d N_A_27_74#_M1016_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90000.7 SB=90004.8 A=0.18 P=2.36 MULT=1
MM1020 N_A_301_368#_M1016_d N_A_27_74#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90001.2 SB=90004.3 A=0.18 P=2.36 MULT=1
MM1015 N_A_301_368#_M1015_d N_B_M1015_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90001.7
+ SB=90003.8 A=0.18 P=2.36 MULT=1
MM1019 N_A_301_368#_M1015_d N_B_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.215 PD=1.27 PS=1.43 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.2
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1005 N_A_301_368#_M1005_d N_C_M1005_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.215 PD=1.27 PS=1.43 NRD=0 NRS=20.685 M=1 R=5.55556 SA=90002.8
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1006 N_A_301_368#_M1005_d N_C_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.209717 PD=1.27 PS=1.43868 NRD=0 NRS=16.0752 M=1 R=5.55556
+ SA=90003.2 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1006_s N_A_301_368#_M1001_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.234883 AS=0.1512 PD=1.61132 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90003.4 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_301_368#_M1014_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.9
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1014_d N_A_301_368#_M1017_g N_X_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90004.4
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_301_368#_M1021_g N_X_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90004.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ms__and3b_4.pxi.spice"
*
.ends
*
*

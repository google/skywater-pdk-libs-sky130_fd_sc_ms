* File: sky130_fd_sc_ms__dlxtn_2.spice
* Created: Wed Sep  2 12:06:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlxtn_2.pex.spice"
.subckt sky130_fd_sc_ms__dlxtn_2  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_D_M1016_g N_A_27_120#_M1016_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.161184 AS=0.15675 PD=1.20233 PS=1.67 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1004 N_A_232_82#_M1004_d N_GATE_N_M1004_g N_VGND_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_232_82#_M1008_g N_A_369_392#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.25707 AS=0.2109 PD=1.55507 PS=2.05 NRD=66.48 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 A_658_79# N_A_27_120#_M1003_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.22233 PD=0.88 PS=1.34493 NRD=12.18 NRS=3.744 M=1 R=4.26667
+ SA=75001.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_672_392#_M1002_d N_A_232_82#_M1002_g A_658_79# VNB NLOWVT L=0.15
+ W=0.64 AD=0.169238 AS=0.0768 PD=1.52755 PS=0.88 NRD=24.372 NRS=12.18 M=1
+ R=4.26667 SA=75001.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1013 A_875_139# N_A_369_392#_M1013_g N_A_672_392#_M1002_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.111062 PD=0.66 PS=1.00245 NRD=18.564 NRS=38.568 M=1
+ R=2.8 SA=75001.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_842_405#_M1006_g A_875_139# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_A_842_405#_M1011_d N_A_672_392#_M1011_g N_VGND_M1006_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Q_M1000_d N_A_842_405#_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2109 PD=1.08 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_Q_M1000_d N_A_842_405#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2294 PD=1.08 PS=2.1 NRD=8.916 NRS=4.044 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_A_27_120#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1017 N_A_232_82#_M1017_d N_GATE_N_M1017_g N_VPWR_M1001_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1554 PD=2.24 PS=1.21 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1018 N_VPWR_M1018_d N_A_232_82#_M1018_g N_A_369_392#_M1018_s VPB PSHORT L=0.18
+ W=0.84 AD=0.22034 AS=0.2352 PD=1.44717 PS=2.24 NRD=48.5999 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1009 A_588_392# N_A_27_120#_M1009_g N_VPWR_M1018_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.26231 PD=1.24 PS=1.72283 NRD=12.7853 NRS=18.6953 M=1 R=5.55556
+ SA=90000.7 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1012 N_A_672_392#_M1012_d N_A_369_392#_M1012_g A_588_392# VPB PSHORT L=0.18
+ W=1 AD=0.270335 AS=0.12 PD=2.01408 PS=1.24 NRD=5.8903 NRS=12.7853 M=1
+ R=5.55556 SA=90001.2 SB=90001 A=0.18 P=2.36 MULT=1
MM1015 A_794_503# N_A_232_82#_M1015_g N_A_672_392#_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.11354 PD=0.66 PS=0.845915 NRD=30.4759 NRS=56.2829 M=1
+ R=2.33333 SA=90001.7 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_842_405#_M1007_g A_794_503# VPB PSHORT L=0.18 W=0.42
+ AD=0.129055 AS=0.0504 PD=0.998182 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333
+ SA=90002.1 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1014 N_A_842_405#_M1014_d N_A_672_392#_M1014_g N_VPWR_M1007_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.344145 PD=2.8 PS=2.66182 NRD=0 NRS=0 M=1
+ R=6.22222 SA=90001.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_842_405#_M1005_g N_Q_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1764 PD=2.8 PS=1.435 NRD=0 NRS=2.6201 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1019_d N_A_842_405#_M1019_g N_Q_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1764 PD=2.8 PS=1.435 NRD=0 NRS=3.5066 M=1 R=6.22222 SA=90000.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.1255 P=18.93
c_78 VNB 0 1.98766e-19 $X=0 $Y=0
c_950 A_658_79# 0 3.15497e-20 $X=3.29 $Y=0.395
*
.include "sky130_fd_sc_ms__dlxtn_2.pxi.spice"
*
.ends
*
*

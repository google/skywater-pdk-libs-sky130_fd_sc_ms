# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__xnor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.916200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575000 1.180000 0.865000 1.225000 ;
        RECT 0.575000 1.225000 3.265000 1.365000 ;
        RECT 0.575000 1.365000 0.865000 1.410000 ;
        RECT 2.975000 1.180000 3.265000 1.225000 ;
        RECT 2.975000 1.365000 3.265000 1.410000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.916200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.350000 1.675000 1.720000 ;
        RECT 1.345000 1.720000 2.775000 1.890000 ;
        RECT 2.605000 1.890000 2.775000 2.060000 ;
        RECT 2.605000 2.060000 5.195000 2.230000 ;
        RECT 3.925000 1.010000 5.195000 1.180000 ;
        RECT 3.925000 1.180000 4.255000 1.550000 ;
        RECT 5.025000 1.180000 5.195000 2.060000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.005600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.835000 1.010000 ;
        RECT 0.085000 1.010000 0.255000 2.320000 ;
        RECT 0.085000 2.320000 2.435000 2.400000 ;
        RECT 0.085000 2.400000 4.135000 2.490000 ;
        RECT 0.665000 0.255000 2.575000 0.425000 ;
        RECT 0.665000 0.425000 0.835000 0.840000 ;
        RECT 2.045000 2.060000 2.435000 2.320000 ;
        RECT 2.045000 2.490000 4.135000 2.570000 ;
        RECT 2.045000 2.570000 2.435000 2.980000 ;
        RECT 2.190000 0.425000 2.575000 0.500000 ;
        RECT 3.805000 2.570000 4.135000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.495000 0.670000 ;
      RECT 0.115000  2.660000 0.445000 3.245000 ;
      RECT 0.425000  1.180000 0.835000 1.550000 ;
      RECT 0.650000  1.820000 1.175000 2.150000 ;
      RECT 1.005000  0.635000 1.450000 1.010000 ;
      RECT 1.005000  1.010000 2.585000 1.180000 ;
      RECT 1.005000  1.180000 1.175000 1.820000 ;
      RECT 1.230000  2.660000 1.875000 3.245000 ;
      RECT 1.680000  0.595000 2.010000 0.670000 ;
      RECT 1.680000  0.670000 5.165000 0.840000 ;
      RECT 1.915000  1.180000 2.585000 1.550000 ;
      RECT 2.640000  2.740000 2.970000 3.245000 ;
      RECT 2.755000  0.350000 3.085000 0.670000 ;
      RECT 2.755000  0.840000 3.085000 1.010000 ;
      RECT 3.005000  1.180000 3.355000 1.550000 ;
      RECT 3.025000  1.550000 3.355000 1.720000 ;
      RECT 3.025000  1.720000 4.675000 1.890000 ;
      RECT 3.260000  2.740000 3.600000 2.905000 ;
      RECT 3.260000  2.905000 4.635000 3.075000 ;
      RECT 3.265000  0.085000 3.600000 0.500000 ;
      RECT 3.780000  0.490000 4.110000 0.670000 ;
      RECT 4.305000  2.400000 4.635000 2.905000 ;
      RECT 4.310000  0.085000 4.655000 0.500000 ;
      RECT 4.445000  1.350000 4.855000 1.680000 ;
      RECT 4.445000  1.680000 4.675000 1.720000 ;
      RECT 4.805000  2.400000 5.135000 3.245000 ;
      RECT 4.835000  0.490000 5.165000 0.670000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  1.210000 0.805000 1.380000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  1.210000 3.205000 1.380000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_ms__xnor2_2
END LIBRARY

* File: sky130_fd_sc_ms__and3b_2.spice
* Created: Fri Aug 28 17:12:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and3b_2.pex.spice"
.subckt sky130_fd_sc_ms__and3b_2  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_N_M1009_g N_A_27_88#_M1009_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.16225 AS=0.15675 PD=1.69 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1008 A_376_74# N_A_27_88#_M1008_g N_A_284_368#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1006 A_454_74# N_B_M1006_g A_376_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g A_454_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.2 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1004 N_X_M1004_d N_A_284_368#_M1004_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=22.692 M=1 R=4.93333 SA=75001.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1004_d N_A_284_368#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_88#_M1005_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2436 AS=0.2352 PD=2.26 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1002 N_VPWR_M1002_d N_A_27_88#_M1002_g N_A_284_368#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.195 AS=0.28 PD=1.39 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_284_368#_M1001_d N_B_M1001_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.195 PD=1.27 PS=1.39 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90000.8
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_C_M1003_g N_A_284_368#_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.18566 AS=0.135 PD=1.39623 PS=1.27 NRD=16.7253 NRS=0 M=1 R=5.55556
+ SA=90001.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1007_d N_A_284_368#_M1007_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.20794 PD=1.405 PS=1.56377 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1007_d N_A_284_368#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.3136 PD=1.405 PS=2.8 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__and3b_2.pxi.spice"
*
.ends
*
*

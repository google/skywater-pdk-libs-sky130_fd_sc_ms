* File: sky130_fd_sc_ms__a22oi_4.pxi.spice
* Created: Fri Aug 28 17:03:35 2020
* 
x_PM_SKY130_FD_SC_MS__A22OI_4%B2 N_B2_c_125_n N_B2_M1003_g N_B2_M1005_g
+ N_B2_M1010_g N_B2_M1004_g N_B2_M1014_g N_B2_M1006_g N_B2_M1028_g N_B2_M1007_g
+ B2 B2 B2 N_B2_c_129_n N_B2_c_124_n PM_SKY130_FD_SC_MS__A22OI_4%B2
x_PM_SKY130_FD_SC_MS__A22OI_4%B1 N_B1_M1001_g N_B1_M1008_g N_B1_M1002_g
+ N_B1_M1011_g N_B1_M1024_g N_B1_M1016_g N_B1_M1025_g N_B1_M1019_g B1 B1
+ N_B1_c_206_n PM_SKY130_FD_SC_MS__A22OI_4%B1
x_PM_SKY130_FD_SC_MS__A22OI_4%A1 N_A1_M1018_g N_A1_c_295_n N_A1_c_296_n
+ N_A1_M1009_g N_A1_M1020_g N_A1_M1017_g N_A1_M1022_g N_A1_M1027_g N_A1_M1031_g
+ N_A1_M1030_g A1 A1 A1 N_A1_c_302_n PM_SKY130_FD_SC_MS__A22OI_4%A1
x_PM_SKY130_FD_SC_MS__A22OI_4%A2 N_A2_M1000_g N_A2_M1012_g N_A2_M1021_g
+ N_A2_M1013_g N_A2_M1023_g N_A2_M1015_g N_A2_M1026_g N_A2_M1029_g A2 A2 A2
+ N_A2_c_387_n N_A2_c_388_n PM_SKY130_FD_SC_MS__A22OI_4%A2
x_PM_SKY130_FD_SC_MS__A22OI_4%A_45_368# N_A_45_368#_M1003_s N_A_45_368#_M1004_s
+ N_A_45_368#_M1007_s N_A_45_368#_M1011_s N_A_45_368#_M1019_s
+ N_A_45_368#_M1020_d N_A_45_368#_M1031_d N_A_45_368#_M1021_d
+ N_A_45_368#_M1026_d N_A_45_368#_c_462_n N_A_45_368#_c_463_n
+ N_A_45_368#_c_464_n N_A_45_368#_c_480_n N_A_45_368#_c_465_n
+ N_A_45_368#_c_486_n N_A_45_368#_c_466_n N_A_45_368#_c_495_n
+ N_A_45_368#_c_467_n N_A_45_368#_c_468_n N_A_45_368#_c_502_n
+ N_A_45_368#_c_509_n N_A_45_368#_c_469_n N_A_45_368#_c_515_n
+ N_A_45_368#_c_470_n N_A_45_368#_c_526_n N_A_45_368#_c_471_n
+ N_A_45_368#_c_532_n N_A_45_368#_c_472_n N_A_45_368#_c_473_n
+ N_A_45_368#_c_474_n N_A_45_368#_c_475_n N_A_45_368#_c_476_n
+ N_A_45_368#_c_521_n N_A_45_368#_c_524_n N_A_45_368#_c_539_n
+ PM_SKY130_FD_SC_MS__A22OI_4%A_45_368#
x_PM_SKY130_FD_SC_MS__A22OI_4%Y N_Y_M1001_s N_Y_M1024_s N_Y_M1009_s N_Y_M1027_s
+ N_Y_M1003_d N_Y_M1006_d N_Y_M1008_d N_Y_M1016_d N_Y_c_606_n N_Y_c_609_n
+ N_Y_c_610_n N_Y_c_669_n N_Y_c_614_n N_Y_c_621_n N_Y_c_672_n N_Y_c_600_n
+ N_Y_c_601_n N_Y_c_632_n N_Y_c_605_n N_Y_c_602_n N_Y_c_616_n N_Y_c_645_n
+ N_Y_c_678_n N_Y_c_603_n N_Y_c_604_n Y Y PM_SKY130_FD_SC_MS__A22OI_4%Y
x_PM_SKY130_FD_SC_MS__A22OI_4%VPWR N_VPWR_M1018_s N_VPWR_M1022_s N_VPWR_M1000_s
+ N_VPWR_M1023_s N_VPWR_c_700_n N_VPWR_c_701_n N_VPWR_c_702_n N_VPWR_c_703_n
+ N_VPWR_c_704_n N_VPWR_c_705_n N_VPWR_c_706_n N_VPWR_c_707_n VPWR
+ N_VPWR_c_708_n N_VPWR_c_709_n N_VPWR_c_710_n N_VPWR_c_699_n N_VPWR_c_712_n
+ N_VPWR_c_713_n PM_SKY130_FD_SC_MS__A22OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A22OI_4%A_48_74# N_A_48_74#_M1005_s N_A_48_74#_M1010_s
+ N_A_48_74#_M1028_s N_A_48_74#_M1002_d N_A_48_74#_M1025_d N_A_48_74#_c_799_n
+ N_A_48_74#_c_800_n N_A_48_74#_c_801_n N_A_48_74#_c_802_n N_A_48_74#_c_803_n
+ N_A_48_74#_c_804_n N_A_48_74#_c_805_n N_A_48_74#_c_806_n N_A_48_74#_c_807_n
+ N_A_48_74#_c_808_n PM_SKY130_FD_SC_MS__A22OI_4%A_48_74#
x_PM_SKY130_FD_SC_MS__A22OI_4%VGND N_VGND_M1005_d N_VGND_M1014_d N_VGND_M1012_d
+ N_VGND_M1015_d N_VGND_c_865_n N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n
+ N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n VGND
+ N_VGND_c_873_n N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n
+ N_VGND_c_878_n PM_SKY130_FD_SC_MS__A22OI_4%VGND
x_PM_SKY130_FD_SC_MS__A22OI_4%A_840_74# N_A_840_74#_M1009_d N_A_840_74#_M1017_d
+ N_A_840_74#_M1030_d N_A_840_74#_M1013_s N_A_840_74#_M1029_s
+ N_A_840_74#_c_959_n N_A_840_74#_c_960_n N_A_840_74#_c_961_n
+ N_A_840_74#_c_962_n N_A_840_74#_c_963_n N_A_840_74#_c_964_n
+ N_A_840_74#_c_965_n N_A_840_74#_c_966_n N_A_840_74#_c_967_n
+ PM_SKY130_FD_SC_MS__A22OI_4%A_840_74#
cc_1 VNB N_B2_M1005_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.74
cc_2 VNB N_B2_M1010_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.74
cc_3 VNB N_B2_M1014_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_4 VNB N_B2_M1028_g 0.0229726f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_5 VNB N_B2_c_124_n 0.0816419f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.56
cc_6 VNB N_B1_M1001_g 0.0213573f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_7 VNB N_B1_M1002_g 0.0206638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_M1024_g 0.0206542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_M1025_g 0.0248723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB B1 0.0014908f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_11 VNB N_B1_c_206_n 0.081918f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.515
cc_12 VNB N_A1_M1018_g 4.92955e-19 $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_13 VNB N_A1_c_295_n 0.0108754f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.74
cc_14 VNB N_A1_c_296_n 0.0109186f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.74
cc_15 VNB N_A1_M1009_g 0.0269428f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.74
cc_16 VNB N_A1_M1017_g 0.0234062f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_17 VNB N_A1_M1027_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_18 VNB N_A1_M1030_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_19 VNB A1 0.00163664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_302_n 0.0620733f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_21 VNB N_A2_M1012_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_M1013_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1015_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_M1029_g 0.0326336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_c_387_n 0.00356131f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.56
cc_26 VNB N_A2_c_388_n 0.080392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_600_n 0.00224682f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.56
cc_28 VNB N_Y_c_601_n 0.00229069f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.56
cc_29 VNB N_Y_c_602_n 0.0229782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_603_n 0.00510981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_604_n 0.00826357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_699_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_48_74#_c_799_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.74
cc_34 VNB N_A_48_74#_c_800_n 0.00367897f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.68
cc_35 VNB N_A_48_74#_c_801_n 0.0120073f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.4
cc_36 VNB N_A_48_74#_c_802_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_37 VNB N_A_48_74#_c_803_n 0.0102323f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_38 VNB N_A_48_74#_c_804_n 0.00299433f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_39 VNB N_A_48_74#_c_805_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_40 VNB N_A_48_74#_c_806_n 0.00938494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_48_74#_c_807_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.56
cc_42 VNB N_A_48_74#_c_808_n 0.00164253f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.56
cc_43 VNB N_VGND_c_865_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_866_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_867_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_868_n 0.00497771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_869_n 0.108097f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.4
cc_48 VNB N_VGND_c_870_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_871_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_50 VNB N_VGND_c_872_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_51 VNB N_VGND_c_873_n 0.0200958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_874_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_53 VNB N_VGND_c_875_n 0.0231293f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_54 VNB N_VGND_c_876_n 0.445534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_877_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_878_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_840_74#_c_959_n 0.00754101f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.35
cc_58 VNB N_A_840_74#_c_960_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.68
cc_59 VNB N_A_840_74#_c_961_n 0.00257879f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_60 VNB N_A_840_74#_c_962_n 0.00230622f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_61 VNB N_A_840_74#_c_963_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.68
cc_62 VNB N_A_840_74#_c_964_n 0.0166385f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=2.4
cc_63 VNB N_A_840_74#_c_965_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_64 VNB N_A_840_74#_c_966_n 0.00646965f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.56
cc_65 VNB N_A_840_74#_c_967_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_66 VPB N_B2_c_125_n 0.0194702f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.77
cc_67 VPB N_B2_M1004_g 0.0196336f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_68 VPB N_B2_M1006_g 0.0196343f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.4
cc_69 VPB N_B2_M1007_g 0.0203472f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=2.4
cc_70 VPB N_B2_c_129_n 0.00755402f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_71 VPB N_B2_c_124_n 0.020257f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.56
cc_72 VPB N_B1_M1008_g 0.0197821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_B1_M1011_g 0.0196326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_B1_M1016_g 0.0199999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_B1_M1019_g 0.02059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB B1 0.00615807f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_77 VPB N_B1_c_206_n 0.0121998f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_78 VPB N_A1_M1018_g 0.0223262f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_79 VPB N_A1_M1020_g 0.0198939f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_80 VPB N_A1_M1022_g 0.0227028f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.4
cc_81 VPB N_A1_M1031_g 0.0239636f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=2.4
cc_82 VPB A1 0.00976728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A1_c_302_n 0.0167577f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_84 VPB N_A2_M1000_g 0.0202433f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_85 VPB N_A2_M1021_g 0.0198928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A2_M1023_g 0.0198921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A2_M1026_g 0.0281481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A2_c_387_n 0.0103635f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=1.56
cc_89 VPB N_A2_c_388_n 0.012272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_45_368#_c_462_n 0.0454702f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=2.4
cc_91 VPB N_A_45_368#_c_463_n 0.00227131f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_92 VPB N_A_45_368#_c_464_n 0.00933537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_45_368#_c_465_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.56
cc_94 VPB N_A_45_368#_c_466_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.56
cc_95 VPB N_A_45_368#_c_467_n 0.00440264f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_96 VPB N_A_45_368#_c_468_n 0.00275273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_45_368#_c_469_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_45_368#_c_470_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_45_368#_c_471_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_45_368#_c_472_n 0.0168839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_45_368#_c_473_n 0.0345796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_45_368#_c_474_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_45_368#_c_475_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_45_368#_c_476_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_Y_c_605_n 0.00250628f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_106 VPB N_VPWR_c_700_n 0.00335558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_701_n 0.0094781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_702_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_703_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_704_n 0.0993924f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=2.4
cc_111 VPB N_VPWR_c_705_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_706_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_113 VPB N_VPWR_c_707_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_114 VPB N_VPWR_c_708_n 0.0175706f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.56
cc_115 VPB N_VPWR_c_709_n 0.0175706f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.515
cc_116 VPB N_VPWR_c_710_n 0.0212096f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_117 VPB N_VPWR_c_699_n 0.0905491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_712_n 0.0088221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_713_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 N_B2_M1028_g N_B1_M1001_g 0.0189918f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B2_M1007_g N_B1_M1008_g 0.0328829f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B2_M1007_g B1 7.28948e-19 $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B2_c_129_n B1 0.0227445f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_124 N_B2_c_124_n B1 0.00140489f $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_125 N_B2_c_129_n N_B1_c_206_n 6.87613e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_126 N_B2_c_124_n N_B1_c_206_n 0.0197381f $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_127 N_B2_c_125_n N_A_45_368#_c_462_n 0.00181594f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_128 N_B2_c_125_n N_A_45_368#_c_463_n 0.0149887f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_129 N_B2_M1004_g N_A_45_368#_c_463_n 0.0116345f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_130 N_B2_c_125_n N_A_45_368#_c_480_n 6.24073e-19 $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_131 N_B2_M1004_g N_A_45_368#_c_480_n 0.00970901f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_132 N_B2_M1006_g N_A_45_368#_c_480_n 0.00951061f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_133 N_B2_M1007_g N_A_45_368#_c_480_n 5.73047e-19 $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_134 N_B2_M1006_g N_A_45_368#_c_465_n 0.0116345f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_135 N_B2_M1007_g N_A_45_368#_c_465_n 0.0116345f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_136 N_B2_M1006_g N_A_45_368#_c_486_n 5.73047e-19 $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_137 N_B2_M1007_g N_A_45_368#_c_486_n 0.00949909f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_138 N_B2_M1004_g N_A_45_368#_c_474_n 0.00194226f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_139 N_B2_M1006_g N_A_45_368#_c_474_n 0.00194226f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B2_M1007_g N_A_45_368#_c_475_n 0.001916f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_141 N_B2_c_125_n N_Y_c_606_n 0.0025567f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_142 N_B2_c_129_n N_Y_c_606_n 0.0189743f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B2_c_124_n N_Y_c_606_n 5.54777e-19 $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_144 N_B2_c_125_n N_Y_c_609_n 0.00936614f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_145 N_B2_M1004_g N_Y_c_610_n 0.0142562f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_146 N_B2_M1006_g N_Y_c_610_n 0.0142562f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_147 N_B2_c_129_n N_Y_c_610_n 0.0478981f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B2_c_124_n N_Y_c_610_n 4.89356e-19 $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_149 N_B2_M1007_g N_Y_c_614_n 0.0159441f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_150 N_B2_c_129_n N_Y_c_614_n 0.0108884f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_151 N_B2_c_129_n N_Y_c_616_n 0.0143992f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_152 N_B2_c_124_n N_Y_c_616_n 5.51948e-19 $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_153 N_B2_c_125_n N_VPWR_c_704_n 0.00333926f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_154 N_B2_M1004_g N_VPWR_c_704_n 0.00333896f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_155 N_B2_M1006_g N_VPWR_c_704_n 0.00333896f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_156 N_B2_M1007_g N_VPWR_c_704_n 0.00333896f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_157 N_B2_c_125_n N_VPWR_c_699_n 0.00426649f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_158 N_B2_M1004_g N_VPWR_c_699_n 0.00422685f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_159 N_B2_M1006_g N_VPWR_c_699_n 0.00422685f $X=1.475 $Y=2.4 $X2=0 $Y2=0
cc_160 N_B2_M1007_g N_VPWR_c_699_n 0.00422796f $X=1.925 $Y=2.4 $X2=0 $Y2=0
cc_161 N_B2_M1005_g N_A_48_74#_c_799_n 0.00159319f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_162 N_B2_M1005_g N_A_48_74#_c_800_n 0.0167076f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_163 N_B2_M1010_g N_A_48_74#_c_800_n 0.01115f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B2_c_129_n N_A_48_74#_c_800_n 0.0342156f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_165 N_B2_c_124_n N_A_48_74#_c_800_n 0.00286877f $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_166 N_B2_M1005_g N_A_48_74#_c_802_n 6.58468e-19 $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_167 N_B2_M1010_g N_A_48_74#_c_802_n 0.00918302f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B2_M1014_g N_A_48_74#_c_802_n 3.97481e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B2_M1014_g N_A_48_74#_c_803_n 0.0130453f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B2_M1028_g N_A_48_74#_c_803_n 0.0128967f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B2_c_129_n N_A_48_74#_c_803_n 0.0483191f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_172 N_B2_c_124_n N_A_48_74#_c_803_n 0.00527888f $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_173 N_B2_M1028_g N_A_48_74#_c_805_n 9.48753e-19 $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B2_M1010_g N_A_48_74#_c_807_n 0.00157732f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B2_c_129_n N_A_48_74#_c_807_n 0.0213626f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_176 N_B2_c_124_n N_A_48_74#_c_807_n 0.00244789f $X=1.87 $Y=1.56 $X2=0 $Y2=0
cc_177 N_B2_M1005_g N_VGND_c_865_n 0.0128874f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_178 N_B2_M1010_g N_VGND_c_865_n 0.00204878f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B2_M1010_g N_VGND_c_866_n 5.19194e-19 $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B2_M1014_g N_VGND_c_866_n 0.0108127f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B2_M1028_g N_VGND_c_866_n 0.0100301f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B2_M1028_g N_VGND_c_869_n 0.00383152f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B2_M1005_g N_VGND_c_873_n 0.00383152f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_184 N_B2_M1010_g N_VGND_c_874_n 0.00434272f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_185 N_B2_M1014_g N_VGND_c_874_n 0.00383152f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B2_M1005_g N_VGND_c_876_n 0.00761455f $X=0.58 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B2_M1010_g N_VGND_c_876_n 0.00820284f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B2_M1014_g N_VGND_c_876_n 0.0075754f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B2_M1028_g N_VGND_c_876_n 0.00757637f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B1_M1019_g N_A1_M1018_g 0.0125409f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_191 N_B1_c_206_n N_A1_c_296_n 0.0125409f $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_192 N_B1_c_206_n N_A1_M1009_g 0.0020658f $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_193 N_B1_c_206_n A1 8.7484e-19 $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_194 N_B1_M1008_g N_A_45_368#_c_486_n 0.00949909f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_195 N_B1_M1011_g N_A_45_368#_c_486_n 5.73047e-19 $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_196 N_B1_M1008_g N_A_45_368#_c_466_n 0.0116345f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_197 N_B1_M1011_g N_A_45_368#_c_466_n 0.0116345f $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_198 N_B1_M1008_g N_A_45_368#_c_495_n 5.73047e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_199 N_B1_M1011_g N_A_45_368#_c_495_n 0.00951061f $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_200 N_B1_M1016_g N_A_45_368#_c_495_n 0.00951061f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_201 N_B1_M1019_g N_A_45_368#_c_495_n 5.73047e-19 $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_202 N_B1_M1016_g N_A_45_368#_c_467_n 0.0115958f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_203 N_B1_M1019_g N_A_45_368#_c_467_n 0.0132535f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_204 N_B1_M1019_g N_A_45_368#_c_468_n 0.00410764f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_205 N_B1_M1016_g N_A_45_368#_c_502_n 6.01317e-19 $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_206 N_B1_M1019_g N_A_45_368#_c_502_n 0.010544f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_207 N_B1_M1008_g N_A_45_368#_c_475_n 0.001916f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_208 N_B1_M1011_g N_A_45_368#_c_476_n 0.00194226f $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_209 N_B1_M1016_g N_A_45_368#_c_476_n 0.00194226f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_210 N_B1_M1008_g N_Y_c_614_n 0.0142175f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_211 B1 N_Y_c_614_n 0.0161329f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_212 N_B1_c_206_n N_Y_c_614_n 7.35521e-19 $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_213 N_B1_M1001_g N_Y_c_621_n 0.00525476f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B1_M1002_g N_Y_c_621_n 0.00642147f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B1_M1024_g N_Y_c_621_n 5.71377e-19 $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B1_M1002_g N_Y_c_600_n 0.00900535f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B1_M1024_g N_Y_c_600_n 0.00841735f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_218 B1 N_Y_c_600_n 0.0396537f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B1_c_206_n N_Y_c_600_n 0.00272949f $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_220 N_B1_M1001_g N_Y_c_601_n 0.00413664f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B1_M1002_g N_Y_c_601_n 0.00277633f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_222 B1 N_Y_c_601_n 0.027784f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_223 N_B1_c_206_n N_Y_c_601_n 0.00277132f $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_224 N_B1_M1011_g N_Y_c_632_n 0.0142175f $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_225 N_B1_M1016_g N_Y_c_632_n 0.0169129f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_226 B1 N_Y_c_632_n 0.0391986f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B1_c_206_n N_Y_c_632_n 4.84419e-19 $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_228 N_B1_M1016_g N_Y_c_605_n 0.00447513f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B1_M1019_g N_Y_c_605_n 0.00400958f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_230 B1 N_Y_c_605_n 0.0200227f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B1_c_206_n N_Y_c_605_n 0.00951622f $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_232 N_B1_M1002_g N_Y_c_602_n 5.1907e-19 $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B1_M1024_g N_Y_c_602_n 0.0093565f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B1_M1025_g N_Y_c_602_n 0.0241822f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_235 B1 N_Y_c_602_n 0.0195623f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B1_c_206_n N_Y_c_602_n 0.0319577f $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_237 B1 N_Y_c_645_n 0.0143992f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B1_c_206_n N_Y_c_645_n 5.4904e-19 $X=3.59 $Y=1.5 $X2=0 $Y2=0
cc_239 N_B1_M1019_g N_VPWR_c_700_n 3.91772e-19 $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_240 N_B1_M1008_g N_VPWR_c_704_n 0.00333896f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B1_M1011_g N_VPWR_c_704_n 0.00333896f $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_242 N_B1_M1016_g N_VPWR_c_704_n 0.00333896f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_243 N_B1_M1019_g N_VPWR_c_704_n 0.00333896f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_244 N_B1_M1008_g N_VPWR_c_699_n 0.00422796f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B1_M1011_g N_VPWR_c_699_n 0.00422685f $X=2.825 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B1_M1016_g N_VPWR_c_699_n 0.00422685f $X=3.275 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B1_M1019_g N_VPWR_c_699_n 0.00422796f $X=3.725 $Y=2.4 $X2=0 $Y2=0
cc_248 N_B1_M1001_g N_A_48_74#_c_803_n 5.7448e-19 $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B1_M1001_g N_A_48_74#_c_804_n 0.0119575f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B1_M1002_g N_A_48_74#_c_804_n 0.00942802f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B1_M1024_g N_A_48_74#_c_806_n 0.0135458f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B1_M1025_g N_A_48_74#_c_806_n 0.013953f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B1_M1002_g N_A_48_74#_c_808_n 2.84754e-19 $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B1_M1024_g N_A_48_74#_c_808_n 2.84754e-19 $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B1_M1001_g N_VGND_c_869_n 0.00278271f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B1_M1002_g N_VGND_c_869_n 0.00278271f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B1_M1024_g N_VGND_c_869_n 0.00278271f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B1_M1025_g N_VGND_c_869_n 0.00278271f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_259 N_B1_M1001_g N_VGND_c_876_n 0.00353526f $X=2.3 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B1_M1002_g N_VGND_c_876_n 0.00353428f $X=2.73 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B1_M1024_g N_VGND_c_876_n 0.00353428f $X=3.16 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B1_M1025_g N_VGND_c_876_n 0.00358427f $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_263 N_B1_M1025_g N_A_840_74#_c_966_n 5.02354e-19 $X=3.59 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A1_M1031_g N_A2_M1000_g 0.0149277f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A1_M1030_g N_A2_M1012_g 0.019323f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A1_M1031_g N_A2_c_387_n 9.87744e-19 $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_267 A1 N_A2_c_387_n 0.0274602f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_268 N_A1_c_302_n N_A2_c_387_n 0.0108039f $X=5.755 $Y=1.515 $X2=0 $Y2=0
cc_269 N_A1_c_302_n N_A2_c_388_n 0.0216032f $X=5.755 $Y=1.515 $X2=0 $Y2=0
cc_270 N_A1_M1018_g N_A_45_368#_c_467_n 0.00101073f $X=4.175 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A1_M1018_g N_A_45_368#_c_468_n 4.97677e-19 $X=4.175 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A1_M1018_g N_A_45_368#_c_509_n 0.0171838f $X=4.175 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A1_c_295_n N_A_45_368#_c_509_n 0.00268172f $X=4.465 $Y=1.575 $X2=0
+ $Y2=0
cc_274 N_A1_M1020_g N_A_45_368#_c_509_n 0.0142562f $X=4.625 $Y=2.4 $X2=0 $Y2=0
cc_275 A1 N_A_45_368#_c_509_n 0.0203648f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A1_M1022_g N_A_45_368#_c_469_n 0.0121815f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A1_M1031_g N_A_45_368#_c_469_n 8.40609e-19 $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A1_M1022_g N_A_45_368#_c_515_n 0.0140172f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A1_M1031_g N_A_45_368#_c_515_n 0.0185678f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_280 A1 N_A_45_368#_c_515_n 0.0452959f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_281 N_A1_c_302_n N_A_45_368#_c_515_n 0.00172308f $X=5.755 $Y=1.515 $X2=0
+ $Y2=0
cc_282 N_A1_M1022_g N_A_45_368#_c_470_n 8.40609e-19 $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A1_M1031_g N_A_45_368#_c_470_n 0.0124458f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A1_M1022_g N_A_45_368#_c_521_n 8.84614e-19 $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_285 A1 N_A_45_368#_c_521_n 0.0189743f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_286 N_A1_c_302_n N_A_45_368#_c_521_n 5.48413e-19 $X=5.755 $Y=1.515 $X2=0
+ $Y2=0
cc_287 N_A1_M1031_g N_A_45_368#_c_524_n 0.00196977f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_288 N_A1_c_296_n N_Y_c_605_n 7.92155e-19 $X=4.265 $Y=1.575 $X2=0 $Y2=0
cc_289 N_A1_c_296_n N_Y_c_602_n 0.00605014f $X=4.265 $Y=1.575 $X2=0 $Y2=0
cc_290 N_A1_M1009_g N_Y_c_602_n 0.0102495f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_291 A1 N_Y_c_602_n 0.0118787f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_292 N_A1_c_302_n N_Y_c_602_n 7.30532e-19 $X=5.755 $Y=1.515 $X2=0 $Y2=0
cc_293 N_A1_M1017_g N_Y_c_603_n 3.85913e-19 $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A1_M1027_g N_Y_c_603_n 0.00304036f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A1_M1030_g N_Y_c_603_n 0.0054657f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A1_c_302_n N_Y_c_603_n 0.00304816f $X=5.755 $Y=1.515 $X2=0 $Y2=0
cc_297 N_A1_c_296_n N_Y_c_604_n 0.00825396f $X=4.265 $Y=1.575 $X2=0 $Y2=0
cc_298 N_A1_M1009_g N_Y_c_604_n 0.0156902f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A1_M1017_g N_Y_c_604_n 0.0123927f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A1_M1027_g N_Y_c_604_n 0.0106768f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_301 A1 N_Y_c_604_n 0.0766192f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_302 N_A1_c_302_n N_Y_c_604_n 0.00514547f $X=5.755 $Y=1.515 $X2=0 $Y2=0
cc_303 N_A1_M1018_g N_VPWR_c_700_n 0.012709f $X=4.175 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A1_M1020_g N_VPWR_c_700_n 0.013449f $X=4.625 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A1_M1022_g N_VPWR_c_700_n 5.60473e-19 $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A1_M1022_g N_VPWR_c_701_n 0.007417f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_307 N_A1_M1031_g N_VPWR_c_701_n 0.007417f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_308 N_A1_M1031_g N_VPWR_c_702_n 5.56271e-19 $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_309 N_A1_M1018_g N_VPWR_c_704_n 0.00460063f $X=4.175 $Y=2.4 $X2=0 $Y2=0
cc_310 N_A1_M1020_g N_VPWR_c_708_n 0.00460063f $X=4.625 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A1_M1022_g N_VPWR_c_708_n 0.005209f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A1_M1031_g N_VPWR_c_709_n 0.005209f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A1_M1018_g N_VPWR_c_699_n 0.00908665f $X=4.175 $Y=2.4 $X2=0 $Y2=0
cc_314 N_A1_M1020_g N_VPWR_c_699_n 0.00908554f $X=4.625 $Y=2.4 $X2=0 $Y2=0
cc_315 N_A1_M1022_g N_VPWR_c_699_n 0.00983498f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A1_M1031_g N_VPWR_c_699_n 0.00983609f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_317 N_A1_M1009_g N_A_48_74#_c_806_n 0.0032792f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A1_M1030_g N_VGND_c_867_n 6.37019e-19 $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A1_M1009_g N_VGND_c_869_n 0.00291649f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A1_M1017_g N_VGND_c_869_n 0.00291649f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A1_M1027_g N_VGND_c_869_n 0.00291649f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A1_M1030_g N_VGND_c_869_n 0.00291649f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A1_M1009_g N_VGND_c_876_n 0.0036412f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A1_M1017_g N_VGND_c_876_n 0.00359121f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A1_M1027_g N_VGND_c_876_n 0.00359121f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A1_M1030_g N_VGND_c_876_n 0.00359219f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A1_M1009_g N_A_840_74#_c_959_n 0.00920696f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A1_M1017_g N_A_840_74#_c_959_n 0.0106927f $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_M1027_g N_A_840_74#_c_959_n 0.0105443f $X=5.4 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1030_g N_A_840_74#_c_959_n 0.014175f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1030_g N_A_840_74#_c_962_n 0.0017668f $X=5.83 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1009_g N_A_840_74#_c_966_n 0.00296395f $X=4.54 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1017_g N_A_840_74#_c_966_n 3.85913e-19 $X=4.97 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A2_M1000_g N_A_45_368#_c_470_n 3.25185e-19 $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A2_M1000_g N_A_45_368#_c_526_n 0.0142562f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A2_M1021_g N_A_45_368#_c_526_n 0.0142562f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_337 N_A2_c_387_n N_A_45_368#_c_526_n 0.0478981f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_338 N_A2_c_388_n N_A_45_368#_c_526_n 4.87946e-19 $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_339 N_A2_M1021_g N_A_45_368#_c_471_n 3.19438e-19 $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_340 N_A2_M1023_g N_A_45_368#_c_471_n 3.19438e-19 $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_341 N_A2_M1023_g N_A_45_368#_c_532_n 0.0142562f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_342 N_A2_M1026_g N_A_45_368#_c_532_n 0.0196896f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A2_c_387_n N_A_45_368#_c_532_n 0.0326319f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_344 N_A2_c_388_n N_A_45_368#_c_532_n 4.90767e-19 $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_345 N_A2_M1026_g N_A_45_368#_c_472_n 8.13654e-19 $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_346 N_A2_M1026_g N_A_45_368#_c_473_n 0.00147311f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_347 N_A2_c_387_n N_A_45_368#_c_524_n 0.0148344f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_348 N_A2_c_387_n N_A_45_368#_c_539_n 0.0143992f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_349 N_A2_c_388_n N_A_45_368#_c_539_n 5.53363e-19 $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_350 N_A2_M1000_g N_VPWR_c_702_n 0.013449f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A2_M1021_g N_VPWR_c_702_n 0.0133668f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A2_M1023_g N_VPWR_c_702_n 5.41206e-19 $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_353 N_A2_M1021_g N_VPWR_c_703_n 5.41206e-19 $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_354 N_A2_M1023_g N_VPWR_c_703_n 0.0133668f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_355 N_A2_M1026_g N_VPWR_c_703_n 0.0164749f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_356 N_A2_M1021_g N_VPWR_c_706_n 0.00460063f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A2_M1023_g N_VPWR_c_706_n 0.00460063f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_358 N_A2_M1000_g N_VPWR_c_709_n 0.00460063f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A2_M1026_g N_VPWR_c_710_n 0.00460063f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A2_M1000_g N_VPWR_c_699_n 0.00908665f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A2_M1021_g N_VPWR_c_699_n 0.00908554f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A2_M1023_g N_VPWR_c_699_n 0.00908554f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_363 N_A2_M1026_g N_VPWR_c_699_n 0.00912597f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_364 N_A2_M1012_g N_VGND_c_867_n 0.00977449f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_365 N_A2_M1013_g N_VGND_c_867_n 0.00192252f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A2_M1013_g N_VGND_c_868_n 5.20618e-19 $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A2_M1015_g N_VGND_c_868_n 0.00985915f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A2_M1029_g N_VGND_c_868_n 0.00328502f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A2_M1012_g N_VGND_c_869_n 0.00383152f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A2_M1013_g N_VGND_c_871_n 0.00434272f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A2_M1015_g N_VGND_c_871_n 0.00383152f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A2_M1029_g N_VGND_c_875_n 0.00434272f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A2_M1012_g N_VGND_c_876_n 0.00757637f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A2_M1013_g N_VGND_c_876_n 0.00820284f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A2_M1015_g N_VGND_c_876_n 0.0075754f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A2_M1029_g N_VGND_c_876_n 0.00824275f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A2_M1012_g N_A_840_74#_c_961_n 0.0128967f $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A2_M1013_g N_A_840_74#_c_961_n 0.0111034f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A2_c_387_n N_A_840_74#_c_961_n 0.0456932f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_380 N_A2_c_388_n N_A_840_74#_c_961_n 0.00388668f $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_381 N_A2_c_387_n N_A_840_74#_c_962_n 0.0152645f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_382 N_A2_c_388_n N_A_840_74#_c_962_n 4.08598e-19 $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_383 N_A2_M1012_g N_A_840_74#_c_963_n 7.09663e-19 $X=6.26 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A2_M1013_g N_A_840_74#_c_963_n 0.00918302f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A2_M1015_g N_A_840_74#_c_963_n 3.97481e-19 $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A2_M1015_g N_A_840_74#_c_964_n 0.0130918f $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A2_M1029_g N_A_840_74#_c_964_n 0.0180198f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A2_c_387_n N_A_840_74#_c_964_n 0.0358403f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_389 N_A2_c_388_n N_A_840_74#_c_964_n 0.00324916f $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_390 N_A2_M1015_g N_A_840_74#_c_965_n 7.07591e-19 $X=7.12 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A2_M1029_g N_A_840_74#_c_965_n 0.0100626f $X=7.55 $Y=0.74 $X2=0 $Y2=0
cc_392 N_A2_M1013_g N_A_840_74#_c_967_n 0.00157732f $X=6.69 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A2_c_387_n N_A_840_74#_c_967_n 0.0213626f $X=7.3 $Y=1.515 $X2=0 $Y2=0
cc_394 N_A2_c_388_n N_A_840_74#_c_967_n 0.00244789f $X=7.555 $Y=1.515 $X2=0
+ $Y2=0
cc_395 N_A_45_368#_c_463_n N_Y_M1003_d 0.00165831f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_396 N_A_45_368#_c_465_n N_Y_M1006_d 0.00165831f $X=1.985 $Y=2.99 $X2=0 $Y2=0
cc_397 N_A_45_368#_c_466_n N_Y_M1008_d 0.00165831f $X=2.885 $Y=2.99 $X2=0 $Y2=0
cc_398 N_A_45_368#_c_467_n N_Y_M1016_d 0.00165831f $X=3.785 $Y=2.99 $X2=0 $Y2=0
cc_399 N_A_45_368#_c_463_n N_Y_c_609_n 0.0139027f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_400 N_A_45_368#_M1004_s N_Y_c_610_n 0.00314376f $X=1.115 $Y=1.84 $X2=0 $Y2=0
cc_401 N_A_45_368#_c_480_n N_Y_c_610_n 0.0170259f $X=1.25 $Y=2.375 $X2=0 $Y2=0
cc_402 N_A_45_368#_c_465_n N_Y_c_669_n 0.0118736f $X=1.985 $Y=2.99 $X2=0 $Y2=0
cc_403 N_A_45_368#_M1007_s N_Y_c_614_n 0.00749611f $X=2.015 $Y=1.84 $X2=0 $Y2=0
cc_404 N_A_45_368#_c_486_n N_Y_c_614_n 0.0170259f $X=2.15 $Y=2.375 $X2=0 $Y2=0
cc_405 N_A_45_368#_c_466_n N_Y_c_672_n 0.0118736f $X=2.885 $Y=2.99 $X2=0 $Y2=0
cc_406 N_A_45_368#_M1011_s N_Y_c_632_n 0.00314376f $X=2.915 $Y=1.84 $X2=0 $Y2=0
cc_407 N_A_45_368#_c_495_n N_Y_c_632_n 0.0170259f $X=3.05 $Y=2.375 $X2=0 $Y2=0
cc_408 N_A_45_368#_c_468_n N_Y_c_605_n 0.00542049f $X=3.91 $Y=2.12 $X2=0 $Y2=0
cc_409 N_A_45_368#_c_468_n N_Y_c_602_n 0.0154538f $X=3.91 $Y=2.12 $X2=0 $Y2=0
cc_410 N_A_45_368#_c_509_n N_Y_c_602_n 0.00514862f $X=4.765 $Y=2.035 $X2=0 $Y2=0
cc_411 N_A_45_368#_c_467_n N_Y_c_678_n 0.0118736f $X=3.785 $Y=2.99 $X2=0 $Y2=0
cc_412 N_A_45_368#_c_509_n N_VPWR_M1018_s 0.00442649f $X=4.765 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_413 N_A_45_368#_c_515_n N_VPWR_M1022_s 0.00888936f $X=5.815 $Y=2.035 $X2=0
+ $Y2=0
cc_414 N_A_45_368#_c_526_n N_VPWR_M1000_s 0.00314376f $X=6.795 $Y=2.035 $X2=0
+ $Y2=0
cc_415 N_A_45_368#_c_532_n N_VPWR_M1023_s 0.00314376f $X=7.695 $Y=2.035 $X2=0
+ $Y2=0
cc_416 N_A_45_368#_c_467_n N_VPWR_c_700_n 0.0103602f $X=3.785 $Y=2.99 $X2=0
+ $Y2=0
cc_417 N_A_45_368#_c_509_n N_VPWR_c_700_n 0.0170259f $X=4.765 $Y=2.035 $X2=0
+ $Y2=0
cc_418 N_A_45_368#_c_469_n N_VPWR_c_700_n 0.0234083f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_419 N_A_45_368#_c_469_n N_VPWR_c_701_n 0.0256432f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_420 N_A_45_368#_c_515_n N_VPWR_c_701_n 0.0314044f $X=5.815 $Y=2.035 $X2=0
+ $Y2=0
cc_421 N_A_45_368#_c_470_n N_VPWR_c_701_n 0.0256432f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_45_368#_c_470_n N_VPWR_c_702_n 0.0234083f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_45_368#_c_526_n N_VPWR_c_702_n 0.0170259f $X=6.795 $Y=2.035 $X2=0
+ $Y2=0
cc_424 N_A_45_368#_c_471_n N_VPWR_c_702_n 0.0233699f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_45_368#_c_471_n N_VPWR_c_703_n 0.0233699f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A_45_368#_c_532_n N_VPWR_c_703_n 0.0170259f $X=7.695 $Y=2.035 $X2=0
+ $Y2=0
cc_427 N_A_45_368#_c_473_n N_VPWR_c_703_n 0.0234083f $X=7.78 $Y=2.4 $X2=0 $Y2=0
cc_428 N_A_45_368#_c_463_n N_VPWR_c_704_n 0.0408559f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_429 N_A_45_368#_c_464_n N_VPWR_c_704_n 0.0179217f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_430 N_A_45_368#_c_465_n N_VPWR_c_704_n 0.0357927f $X=1.985 $Y=2.99 $X2=0
+ $Y2=0
cc_431 N_A_45_368#_c_466_n N_VPWR_c_704_n 0.0357927f $X=2.885 $Y=2.99 $X2=0
+ $Y2=0
cc_432 N_A_45_368#_c_467_n N_VPWR_c_704_n 0.0536089f $X=3.785 $Y=2.99 $X2=0
+ $Y2=0
cc_433 N_A_45_368#_c_474_n N_VPWR_c_704_n 0.0234458f $X=1.25 $Y=2.99 $X2=0 $Y2=0
cc_434 N_A_45_368#_c_475_n N_VPWR_c_704_n 0.0234458f $X=2.15 $Y=2.99 $X2=0 $Y2=0
cc_435 N_A_45_368#_c_476_n N_VPWR_c_704_n 0.0234458f $X=3.05 $Y=2.99 $X2=0 $Y2=0
cc_436 N_A_45_368#_c_471_n N_VPWR_c_706_n 0.00749631f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_437 N_A_45_368#_c_469_n N_VPWR_c_708_n 0.0109793f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_438 N_A_45_368#_c_470_n N_VPWR_c_709_n 0.0109793f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_439 N_A_45_368#_c_473_n N_VPWR_c_710_n 0.011066f $X=7.78 $Y=2.4 $X2=0 $Y2=0
cc_440 N_A_45_368#_c_463_n N_VPWR_c_699_n 0.0229294f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_441 N_A_45_368#_c_464_n N_VPWR_c_699_n 0.00971942f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_442 N_A_45_368#_c_465_n N_VPWR_c_699_n 0.0200586f $X=1.985 $Y=2.99 $X2=0
+ $Y2=0
cc_443 N_A_45_368#_c_466_n N_VPWR_c_699_n 0.0200586f $X=2.885 $Y=2.99 $X2=0
+ $Y2=0
cc_444 N_A_45_368#_c_467_n N_VPWR_c_699_n 0.0296408f $X=3.785 $Y=2.99 $X2=0
+ $Y2=0
cc_445 N_A_45_368#_c_469_n N_VPWR_c_699_n 0.00901959f $X=4.85 $Y=2.415 $X2=0
+ $Y2=0
cc_446 N_A_45_368#_c_470_n N_VPWR_c_699_n 0.00901959f $X=5.98 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_45_368#_c_471_n N_VPWR_c_699_n 0.0062048f $X=6.88 $Y=2.465 $X2=0
+ $Y2=0
cc_448 N_A_45_368#_c_473_n N_VPWR_c_699_n 0.00915947f $X=7.78 $Y=2.4 $X2=0 $Y2=0
cc_449 N_A_45_368#_c_474_n N_VPWR_c_699_n 0.0125551f $X=1.25 $Y=2.99 $X2=0 $Y2=0
cc_450 N_A_45_368#_c_475_n N_VPWR_c_699_n 0.0125551f $X=2.15 $Y=2.99 $X2=0 $Y2=0
cc_451 N_A_45_368#_c_476_n N_VPWR_c_699_n 0.0125551f $X=3.05 $Y=2.99 $X2=0 $Y2=0
cc_452 N_A_45_368#_c_462_n N_A_48_74#_c_801_n 0.00864987f $X=0.35 $Y=1.985 $X2=0
+ $Y2=0
cc_453 N_A_45_368#_c_472_n N_A_840_74#_c_964_n 0.00868683f $X=7.82 $Y=2.12 $X2=0
+ $Y2=0
cc_454 N_Y_c_600_n N_A_48_74#_M1002_d 0.00176461f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_455 N_Y_c_602_n N_A_48_74#_M1025_d 0.00386132f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_456 N_Y_c_601_n N_A_48_74#_c_803_n 0.00997012f $X=2.68 $Y=1.095 $X2=0 $Y2=0
cc_457 N_Y_M1001_s N_A_48_74#_c_804_n 0.00176461f $X=2.375 $Y=0.37 $X2=0 $Y2=0
cc_458 N_Y_c_621_n N_A_48_74#_c_804_n 0.0157965f $X=2.515 $Y=0.76 $X2=0 $Y2=0
cc_459 N_Y_c_600_n N_A_48_74#_c_804_n 0.0030313f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_460 N_Y_M1024_s N_A_48_74#_c_806_n 0.00180346f $X=3.235 $Y=0.37 $X2=0 $Y2=0
cc_461 N_Y_c_600_n N_A_48_74#_c_806_n 0.00436902f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_462 N_Y_c_602_n N_A_48_74#_c_806_n 0.0472031f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_463 N_Y_c_600_n N_A_48_74#_c_808_n 0.0133411f $X=3.21 $Y=1.095 $X2=0 $Y2=0
cc_464 N_Y_c_602_n N_VGND_c_876_n 0.00898375f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_465 N_Y_c_604_n N_A_840_74#_M1009_d 0.00344035f $X=5.45 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_466 N_Y_c_604_n N_A_840_74#_M1017_d 0.00209854f $X=5.45 $Y=0.95 $X2=0 $Y2=0
cc_467 N_Y_M1009_s N_A_840_74#_c_959_n 0.00212678f $X=4.615 $Y=0.37 $X2=0 $Y2=0
cc_468 N_Y_M1027_s N_A_840_74#_c_959_n 0.00179007f $X=5.475 $Y=0.37 $X2=0 $Y2=0
cc_469 N_Y_c_603_n N_A_840_74#_c_959_n 0.016201f $X=5.615 $Y=0.95 $X2=0 $Y2=0
cc_470 N_Y_c_604_n N_A_840_74#_c_959_n 0.0379865f $X=5.45 $Y=0.95 $X2=0 $Y2=0
cc_471 N_Y_c_603_n N_A_840_74#_c_962_n 0.00561736f $X=5.615 $Y=0.95 $X2=0 $Y2=0
cc_472 N_Y_c_602_n N_A_840_74#_c_966_n 0.0030156f $X=4.195 $Y=0.99 $X2=0 $Y2=0
cc_473 N_Y_c_604_n N_A_840_74#_c_966_n 0.0182263f $X=5.45 $Y=0.95 $X2=0 $Y2=0
cc_474 N_A_48_74#_c_800_n N_VGND_M1005_d 0.00176461f $X=1.06 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_475 N_A_48_74#_c_803_n N_VGND_M1014_d 0.00176461f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_476 N_A_48_74#_c_799_n N_VGND_c_865_n 0.0175587f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_477 N_A_48_74#_c_800_n N_VGND_c_865_n 0.0152916f $X=1.06 $Y=1.095 $X2=0 $Y2=0
cc_478 N_A_48_74#_c_802_n N_VGND_c_865_n 0.0175587f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_479 N_A_48_74#_c_802_n N_VGND_c_866_n 0.0182902f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_480 N_A_48_74#_c_803_n N_VGND_c_866_n 0.0170777f $X=2 $Y=1.095 $X2=0 $Y2=0
cc_481 N_A_48_74#_c_805_n N_VGND_c_866_n 0.0112234f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_482 N_A_48_74#_c_804_n N_VGND_c_869_n 0.0435462f $X=2.86 $Y=0.34 $X2=0 $Y2=0
cc_483 N_A_48_74#_c_805_n N_VGND_c_869_n 0.0121867f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_484 N_A_48_74#_c_806_n N_VGND_c_869_n 0.0626962f $X=3.805 $Y=0.515 $X2=0
+ $Y2=0
cc_485 N_A_48_74#_c_808_n N_VGND_c_869_n 0.0119073f $X=2.945 $Y=0.34 $X2=0 $Y2=0
cc_486 N_A_48_74#_c_799_n N_VGND_c_873_n 0.011066f $X=0.365 $Y=0.515 $X2=0 $Y2=0
cc_487 N_A_48_74#_c_802_n N_VGND_c_874_n 0.0109942f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_488 N_A_48_74#_c_799_n N_VGND_c_876_n 0.00915947f $X=0.365 $Y=0.515 $X2=0
+ $Y2=0
cc_489 N_A_48_74#_c_802_n N_VGND_c_876_n 0.00904371f $X=1.225 $Y=0.515 $X2=0
+ $Y2=0
cc_490 N_A_48_74#_c_804_n N_VGND_c_876_n 0.0245733f $X=2.86 $Y=0.34 $X2=0 $Y2=0
cc_491 N_A_48_74#_c_805_n N_VGND_c_876_n 0.00660921f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_492 N_A_48_74#_c_806_n N_VGND_c_876_n 0.0345365f $X=3.805 $Y=0.515 $X2=0
+ $Y2=0
cc_493 N_A_48_74#_c_808_n N_VGND_c_876_n 0.00650586f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_494 N_A_48_74#_c_806_n N_A_840_74#_c_966_n 0.0214676f $X=3.805 $Y=0.515 $X2=0
+ $Y2=0
cc_495 N_VGND_c_867_n N_A_840_74#_c_960_n 0.00947603f $X=6.475 $Y=0.595 $X2=0
+ $Y2=0
cc_496 N_VGND_c_869_n N_A_840_74#_c_960_n 0.00758556f $X=6.31 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_876_n N_A_840_74#_c_960_n 0.00627867f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_498 N_VGND_M1012_d N_A_840_74#_c_961_n 0.00176461f $X=6.335 $Y=0.37 $X2=0
+ $Y2=0
cc_499 N_VGND_c_867_n N_A_840_74#_c_961_n 0.0153337f $X=6.475 $Y=0.595 $X2=0
+ $Y2=0
cc_500 N_VGND_c_867_n N_A_840_74#_c_963_n 0.0175587f $X=6.475 $Y=0.595 $X2=0
+ $Y2=0
cc_501 N_VGND_c_868_n N_A_840_74#_c_963_n 0.0175587f $X=7.335 $Y=0.595 $X2=0
+ $Y2=0
cc_502 N_VGND_c_871_n N_A_840_74#_c_963_n 0.0109942f $X=7.17 $Y=0 $X2=0 $Y2=0
cc_503 N_VGND_c_876_n N_A_840_74#_c_963_n 0.00904371f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_504 N_VGND_M1015_d N_A_840_74#_c_964_n 0.00176461f $X=7.195 $Y=0.37 $X2=0
+ $Y2=0
cc_505 N_VGND_c_868_n N_A_840_74#_c_964_n 0.0153337f $X=7.335 $Y=0.595 $X2=0
+ $Y2=0
cc_506 N_VGND_c_868_n N_A_840_74#_c_965_n 0.0182902f $X=7.335 $Y=0.595 $X2=0
+ $Y2=0
cc_507 N_VGND_c_875_n N_A_840_74#_c_965_n 0.0145639f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_876_n N_A_840_74#_c_965_n 0.0119984f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_869_n N_A_840_74#_c_966_n 0.0731929f $X=6.31 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_876_n N_A_840_74#_c_966_n 0.0615691f $X=7.92 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dlrbp_2.spice
* Created: Fri Aug 28 17:27:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrbp_2.pex.spice"
.subckt sky130_fd_sc_ms__dlrbp_2  VNB VPB D GATE RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_D_M1015_g N_A_27_112#_M1015_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1013 N_A_230_74#_M1013_d N_GATE_M1013_g N_VGND_M1015_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_230_74#_M1002_g N_A_363_82#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.201864 AS=0.2109 PD=1.51754 PS=2.05 NRD=35.316 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 A_569_80# N_A_27_112#_M1004_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.174586 PD=0.85 PS=1.31246 NRD=9.372 NRS=16.872 M=1 R=4.26667
+ SA=75000.8 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_641_80#_M1023_d N_A_363_82#_M1023_g A_569_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.162536 AS=0.0672 PD=1.38868 PS=0.85 NRD=21.552 NRS=9.372 M=1
+ R=4.26667 SA=75001.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1003 A_773_124# N_A_230_74#_M1003_g N_A_641_80#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.106664 PD=0.66 PS=0.911321 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_821_98#_M1018_g A_773_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 A_1049_74# N_A_641_80#_M1016_g N_A_821_98#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_1049_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0888 PD=1.13 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1024 N_Q_M1024_d N_A_821_98#_M1024_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1443 PD=1.02 PS=1.13 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_Q_M1024_d N_A_821_98#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_821_98#_M1006_g N_A_1449_368#_M1006_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1011 N_Q_N_M1011_d N_A_1449_368#_M1011_g N_VGND_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.157545 PD=1.02 PS=1.24406 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1019 N_Q_N_M1011_d N_A_1449_368#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_112#_M1000_s VPB PSHORT L=0.18 W=0.84
+ AD=0.21525 AS=0.2352 PD=1.49 PS=2.24 NRD=47.1815 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1017 N_A_230_74#_M1017_d N_GATE_M1017_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2772 AS=0.21525 PD=2.34 PS=1.49 NRD=0 NRS=47.1815 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1001_d N_A_230_74#_M1001_g N_A_363_82#_M1001_s VPB PSHORT L=0.18
+ W=0.84 AD=0.172565 AS=0.2352 PD=1.26913 PS=2.24 NRD=23.443 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1010 A_569_392# N_A_27_112#_M1010_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.205435 PD=1.24 PS=1.51087 NRD=12.7853 NRS=2.9353 M=1 R=5.55556
+ SA=90000.7 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1014 N_A_641_80#_M1014_d N_A_230_74#_M1014_g A_569_392# VPB PSHORT L=0.18 W=1
+ AD=0.219366 AS=0.12 PD=1.90845 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1020 A_760_508# N_A_363_82#_M1020_g N_A_641_80#_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09975 AS=0.0921338 PD=0.895 PS=0.801549 NRD=85.5965 NRS=39.8531
+ M=1 R=2.33333 SA=90001.5 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_821_98#_M1007_g A_760_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.114164 AS=0.09975 PD=0.927273 PS=0.895 NRD=70.3487 NRS=85.5965 M=1
+ R=2.33333 SA=90002.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1027 N_A_821_98#_M1027_d N_A_641_80#_M1027_g N_VPWR_M1007_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.304436 PD=1.44 PS=2.47273 NRD=7.8997 NRS=26.3783 M=1
+ R=6.22222 SA=90001.2 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1026 N_VPWR_M1026_d N_RESET_B_M1026_g N_A_821_98#_M1027_d VPB PSHORT L=0.18
+ W=1.12 AD=0.196 AS=0.1792 PD=1.47 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90001.7 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1021 N_Q_M1021_d N_A_821_98#_M1021_g N_VPWR_M1026_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196 PD=1.39 PS=1.47 NRD=0 NRS=4.3931 M=1 R=6.22222 SA=90002.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1022 N_Q_M1021_d N_A_821_98#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1012_d N_A_821_98#_M1012_g N_A_1449_368#_M1012_s VPB PSHORT
+ L=0.18 W=1 AD=0.188679 AS=0.28 PD=1.40566 PS=2.56 NRD=8.8453 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1005 N_Q_N_M1005_d N_A_1449_368#_M1005_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.211321 PD=1.39 PS=1.57434 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.7 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1008 N_Q_N_M1005_d N_A_1449_368#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ms__dlrbp_2.pxi.spice"
*
.ends
*
*

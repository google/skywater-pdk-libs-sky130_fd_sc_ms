* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_231_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_465_368# C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_159_368# B1 a_465_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_159_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_159_74# A2 a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR A1 a_159_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 VPWR A3 a_159_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND A3 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__o2111a_1.spice
* Created: Fri Aug 28 17:51:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2111a_1.pex.spice"
.subckt sky130_fd_sc_ms__o2111a_1  VNB VPB D1 C1 B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_82_48#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.2035 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 A_321_74# N_D1_M1011_g N_A_82_48#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.259 PD=0.95 PS=2.18 NRD=8.1 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1000 A_393_74# N_C1_M1000_g A_321_74# VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.0777 PD=0.98 PS=0.95 NRD=10.536 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1001 N_A_471_74#_M1001_d N_B1_M1001_g A_393_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.0888 PD=1.1 PS=0.98 NRD=8.1 NRS=10.536 M=1 R=4.93333 SA=75001
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_471_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1332 PD=1.13 PS=1.1 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75001.5
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_A_471_74#_M1009_d N_A1_M1009_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1443 PD=2.05 PS=1.13 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_82_48#_M1003_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2593 AS=0.3136 PD=1.79429 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1008 N_A_82_48#_M1008_d N_D1_M1008_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.194475 PD=1.16 PS=1.34571 NRD=0 NRS=29.8849 M=1 R=4.66667
+ SA=90000.8 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1005_d N_C1_M1005_g N_A_82_48#_M1008_d VPB PSHORT L=0.18 W=0.84
+ AD=0.2415 AS=0.1344 PD=1.415 PS=1.16 NRD=35.1645 NRS=10.5395 M=1 R=4.66667
+ SA=90001.3 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1002 N_A_82_48#_M1002_d N_B1_M1002_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=0.84
+ AD=0.156587 AS=0.2415 PD=1.23717 PS=1.415 NRD=18.7544 NRS=34.0022 M=1
+ R=4.66667 SA=90002.1 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1010 A_603_381# N_A2_M1010_g N_A_82_48#_M1002_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.186413 PD=1.24 PS=1.47283 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90002.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_603_381# VPB PSHORT L=0.18 W=1 AD=0.27
+ AS=0.12 PD=2.54 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90002.6 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o2111a_1.pxi.spice"
*
.ends
*
*

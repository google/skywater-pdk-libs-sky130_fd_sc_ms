* File: sky130_fd_sc_ms__xnor2_4.spice
* Created: Fri Aug 28 18:17:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xnor2_4.pex.spice"
.subckt sky130_fd_sc_ms__xnor2_4  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1019 N_A_27_74#_M1019_d N_A_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1028 N_A_27_74#_M1028_d N_A_M1028_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.7
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1022 N_A_27_74#_M1028_d N_B_M1022_g N_A_119_368#_M1022_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1026 N_A_27_74#_M1026_d N_B_M1026_g N_A_119_368#_M1022_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_A_511_74#_M1010_d N_A_119_368#_M1010_g N_Y_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.2 SB=75005.9 A=0.111 P=1.78 MULT=1
MM1014 N_A_511_74#_M1014_d N_A_119_368#_M1014_g N_Y_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.16465 AS=0.1295 PD=1.185 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75005.4 A=0.111 P=1.78 MULT=1
MM1017 N_A_511_74#_M1014_d N_A_119_368#_M1017_g N_Y_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.16465 AS=0.1036 PD=1.185 PS=1.02 NRD=15.396 NRS=0 M=1 R=4.93333
+ SA=75001.3 SB=75004.8 A=0.111 P=1.78 MULT=1
MM1029 N_A_511_74#_M1029_d N_A_119_368#_M1029_g N_Y_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.7 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1002 N_A_511_74#_M1029_d N_A_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1889 PD=1.09 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75002.2
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_511_74#_M1009_d N_A_M1009_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75002.8
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1021 N_A_511_74#_M1009_d N_A_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75003.3
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1023 N_A_511_74#_M1023_d N_A_M1023_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75003.8
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g N_A_511_74#_M1023_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.205 AS=0.1036 PD=1.395 PS=1.02 NRD=36 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1001_d N_B_M1015_g N_A_511_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.205 AS=0.1036 PD=1.395 PS=1.02 NRD=36 NRS=0 M=1 R=4.93333 SA=75004.9
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_B_M1016_g N_A_511_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1889 AS=0.1036 PD=1.36 PS=1.02 NRD=32.472 NRS=0 M=1 R=4.93333 SA=75005.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1016_d N_B_M1024_g N_A_511_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1889 AS=0.2109 PD=1.36 PS=2.05 NRD=32.472 NRS=0 M=1 R=4.93333 SA=75005.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_119_368#_M1012_d N_A_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1013 N_A_119_368#_M1012_d N_A_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1134 PD=1.11 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.6
+ SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1018 N_A_119_368#_M1018_d N_B_M1018_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1134 PD=1.11 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667 SA=90001.1
+ SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1020 N_A_119_368#_M1018_d N_B_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.237214 PD=1.11 PS=1.54714 NRD=0 NRS=53.3279 M=1 R=4.66667
+ SA=90001.5 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1025 N_Y_M1025_d N_A_119_368#_M1025_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.316286 PD=1.39 PS=2.06286 NRD=0 NRS=39.991 M=1 R=6.22222
+ SA=90001.7 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1027 N_Y_M1025_d N_A_119_368#_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.47695 PD=1.39 PS=3.44 NRD=0 NRS=65.2267 M=1 R=6.22222
+ SA=90002.1 SB=90000.3 A=0.2016 P=2.6 MULT=1
MM1000 N_A_950_368#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.283862 PD=2.8 PS=1.8 NRD=0 NRS=34.8887 M=1 R=6.22222 SA=90000.2
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1004 N_A_950_368#_M1004_d N_A_M1004_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.283862 PD=1.39 PS=1.8 NRD=0 NRS=34.8887 M=1 R=6.22222
+ SA=90000.8 SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1006 N_A_950_368#_M1004_d N_A_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.280475 PD=1.39 PS=1.795 NRD=0 NRS=34.3568 M=1 R=6.22222
+ SA=90001.3 SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1007 N_A_950_368#_M1007_d N_A_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.280475 PD=1.39 PS=1.795 NRD=0 NRS=34.3568 M=1 R=6.22222
+ SA=90001.9 SB=90002 A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_A_950_368#_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1003_d N_B_M1005_g N_A_950_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.8
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_B_M1008_g N_A_950_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1008_d N_B_M1011_g N_A_950_368#_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX30_noxref VNB VPB NWDIODE A=17.67 P=22.72
c_79 VNB 0 1.57454e-19 $X=0 $Y=0
c_143 VPB 0 3.00577e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__xnor2_4.pxi.spice"
*
.ends
*
*

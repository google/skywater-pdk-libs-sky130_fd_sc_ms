* File: sky130_fd_sc_ms__conb_1.pxi.spice
* Created: Wed Sep  2 12:02:02 2020
* 
x_PM_SKY130_FD_SC_MS__CONB_1%HI HI HI HI HI HI N_HI_R0_pos N_HI_c_24_n
+ N_HI_c_25_n HI PM_SKY130_FD_SC_MS__CONB_1%HI
x_PM_SKY130_FD_SC_MS__CONB_1%VPWR N_VPWR_c_44_n N_VPWR_c_42_n N_VPWR_c_46_n
+ N_VPWR_c_47_n VPWR N_VPWR_R0_neg N_VPWR_c_48_n N_VPWR_c_43_n
+ PM_SKY130_FD_SC_MS__CONB_1%VPWR
x_PM_SKY130_FD_SC_MS__CONB_1%VGND N_VGND_c_61_n N_VGND_c_62_n N_VGND_c_63_n
+ N_VGND_c_64_n N_VGND_c_65_n VGND N_VGND_R1_pos N_VGND_c_66_n
+ PM_SKY130_FD_SC_MS__CONB_1%VGND
x_PM_SKY130_FD_SC_MS__CONB_1%LO LO LO LO LO LO N_LO_R1_neg N_LO_c_79_n LO
+ PM_SKY130_FD_SC_MS__CONB_1%LO
cc_1 VNB N_HI_c_24_n 0.144349f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=0.34
cc_2 VNB N_HI_c_25_n 0.0234388f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=0.34
cc_3 VNB HI 0.0301052f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.925
cc_4 VNB N_VPWR_c_42_n 0.0163332f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_5 VNB N_VPWR_c_43_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.925
cc_6 VNB N_VGND_c_61_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_VGND_c_62_n 0.163296f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_VGND_c_63_n 0.0104949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_64_n 0.0224837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_65_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_66_n 0.115863f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.927
cc_12 VNB LO 0.0252697f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_13 VNB N_LO_c_79_n 0.0163328f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=0.34
cc_14 VPB HI 0.0257382f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.925
cc_15 VPB N_VPWR_c_44_n 0.00177638f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_16 VPB N_VPWR_c_42_n 0.185307f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_17 VPB N_VPWR_c_46_n 0.0104949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_47_n 0.00497896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_48_n 0.0224837f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.925
cc_20 VPB N_VPWR_c_43_n 0.0516935f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.925
cc_21 VPB LO 0.0303528f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_22 VPB LO 0.0234388f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_23 VPB N_LO_c_79_n 0.166357f $X=-0.19 $Y=1.66 $X2=0.45 $Y2=0.34
cc_24 HI N_VPWR_c_44_n 0.00914229f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_25 HI N_VPWR_c_42_n 0.0617789f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_26 N_HI_c_24_n N_VGND_c_61_n 0.00301226f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_27 N_HI_c_25_n N_VGND_c_61_n 0.03748f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_28 N_HI_c_24_n N_VGND_c_62_n 0.0875407f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_29 N_HI_c_25_n N_VGND_c_62_n 0.00229804f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_30 HI N_VGND_c_62_n 0.00205142f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_31 N_HI_c_24_n N_VGND_c_64_n 0.0106827f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_32 N_HI_c_25_n N_VGND_c_64_n 0.0359088f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_33 N_HI_c_24_n N_VGND_c_66_n 0.0139097f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_34 N_HI_c_25_n N_VGND_c_66_n 0.0181672f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_35 N_HI_c_24_n LO 0.00132481f $X=0.45 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_36 HI LO 0.0323696f $X=0.24 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_37 HI N_LO_c_79_n 0.00249655f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_38 N_VPWR_c_42_n LO 0.00313643f $X=0.45 $Y=2.605 $X2=-0.19 $Y2=-0.245
cc_39 N_VPWR_c_44_n LO 0.03748f $X=0.45 $Y=2.605 $X2=0 $Y2=0
cc_40 N_VPWR_c_42_n LO 0.00229804f $X=0.45 $Y=2.605 $X2=0 $Y2=0
cc_41 N_VPWR_c_48_n LO 0.0359018f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_42 N_VPWR_c_43_n LO 0.0181658f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_43 N_VPWR_c_44_n N_LO_c_79_n 0.00301226f $X=0.45 $Y=2.605 $X2=0 $Y2=0
cc_44 N_VPWR_c_42_n N_LO_c_79_n 0.114704f $X=0.45 $Y=2.605 $X2=0 $Y2=0
cc_45 N_VPWR_c_48_n N_LO_c_79_n 0.0106827f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_46 N_VPWR_c_43_n N_LO_c_79_n 0.0139097f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_47 N_VGND_c_61_n LO 0.00829579f $X=0.99 $Y=0.32 $X2=-0.19 $Y2=-0.245
cc_48 N_VGND_c_62_n LO 0.0379897f $X=0.99 $Y=0.32 $X2=-0.19 $Y2=-0.245

* File: sky130_fd_sc_ms__einvn_8.pex.spice
* Created: Fri Aug 28 17:33:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EINVN_8%TE_B 1 3 6 8 10 12 13 15 17 18 20 22 23 25
+ 27 28 30 32 33 35 37 38 40 42 43 45 47 48 49 50 51 52 53 54 55 62
c172 55 0 1.9459e-20 $X=0.24 $Y=1.295
c173 40 0 2.46858e-19 $X=4.415 $Y=1.725
r174 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r175 55 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.465
r176 45 47 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.965 $Y=1.725
+ $X2=4.965 $Y2=2.4
r177 44 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.505 $Y=1.65
+ $X2=4.415 $Y2=1.65
r178 43 45 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.875 $Y=1.65
+ $X2=4.965 $Y2=1.725
r179 43 44 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.875 $Y=1.65
+ $X2=4.505 $Y2=1.65
r180 40 54 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.415 $Y=1.725
+ $X2=4.415 $Y2=1.65
r181 40 42 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.415 $Y=1.725
+ $X2=4.415 $Y2=2.4
r182 39 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.055 $Y=1.65
+ $X2=3.965 $Y2=1.65
r183 38 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=4.415 $Y2=1.65
r184 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=4.055 $Y2=1.65
r185 35 53 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.965 $Y=1.725
+ $X2=3.965 $Y2=1.65
r186 35 37 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.965 $Y=1.725
+ $X2=3.965 $Y2=2.4
r187 34 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.555 $Y=1.65
+ $X2=3.465 $Y2=1.65
r188 33 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.875 $Y=1.65
+ $X2=3.965 $Y2=1.65
r189 33 34 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.875 $Y=1.65
+ $X2=3.555 $Y2=1.65
r190 30 52 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.465 $Y=1.725
+ $X2=3.465 $Y2=1.65
r191 30 32 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.465 $Y=1.725
+ $X2=3.465 $Y2=2.4
r192 29 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.105 $Y=1.65
+ $X2=3.015 $Y2=1.65
r193 28 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.375 $Y=1.65
+ $X2=3.465 $Y2=1.65
r194 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.375 $Y=1.65
+ $X2=3.105 $Y2=1.65
r195 25 51 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=1.725
+ $X2=3.015 $Y2=1.65
r196 25 27 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.015 $Y=1.725
+ $X2=3.015 $Y2=2.4
r197 24 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.605 $Y=1.65
+ $X2=2.515 $Y2=1.65
r198 23 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.925 $Y=1.65
+ $X2=3.015 $Y2=1.65
r199 23 24 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.925 $Y=1.65
+ $X2=2.605 $Y2=1.65
r200 20 50 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.515 $Y=1.725
+ $X2=2.515 $Y2=1.65
r201 20 22 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.515 $Y=1.725
+ $X2=2.515 $Y2=2.4
r202 19 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.155 $Y=1.65
+ $X2=2.065 $Y2=1.65
r203 18 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.425 $Y=1.65
+ $X2=2.515 $Y2=1.65
r204 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.425 $Y=1.65
+ $X2=2.155 $Y2=1.65
r205 15 49 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.065 $Y=1.725
+ $X2=2.065 $Y2=1.65
r206 15 17 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.065 $Y=1.725
+ $X2=2.065 $Y2=2.4
r207 14 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.655 $Y=1.65
+ $X2=1.565 $Y2=1.65
r208 13 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.975 $Y=1.65
+ $X2=2.065 $Y2=1.65
r209 13 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.975 $Y=1.65
+ $X2=1.655 $Y2=1.65
r210 10 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.565 $Y=1.725
+ $X2=1.565 $Y2=1.65
r211 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.565 $Y=1.725
+ $X2=1.565 $Y2=2.4
r212 8 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.475 $Y=1.65
+ $X2=1.565 $Y2=1.65
r213 8 62 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.475 $Y=1.65
+ $X2=0.645 $Y2=1.65
r214 4 62 36.463 $w=4.25e-07 $l=9e-08 $layer=POLY_cond $X=0.555 $Y=1.512
+ $X2=0.645 $Y2=1.512
r215 4 58 37.295 $w=4.25e-07 $l=2.85e-07 $layer=POLY_cond $X=0.555 $Y=1.512
+ $X2=0.27 $Y2=1.512
r216 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.555 $Y2=0.74
r217 1 4 22.9127 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=0.555 $Y=1.725
+ $X2=0.555 $Y2=1.512
r218 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=0.555 $Y=1.725
+ $X2=0.555 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%A_126_74# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 27 29 31 32 34 36 37 39 41 42 44 46 48 49 50 51 52 53 54 57 63 64 69
c154 64 0 3.46022e-20 $X=1.19 $Y=0.49
c155 42 0 1.72182e-19 $X=4.9 $Y=1.26
c156 8 0 1.9459e-20 $X=1.355 $Y=1.26
r157 69 72 6.39005 $w=7.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=1.17
+ $X2=0.985 $Y2=1.335
r158 69 71 0.778307 $w=7.38e-07 $l=4e-08 $layer=LI1_cond $X=0.985 $Y=1.17
+ $X2=0.985 $Y2=1.13
r159 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.17 $X2=1.19 $Y2=1.17
r160 67 71 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.02 $Y=0.515
+ $X2=1.02 $Y2=1.13
r161 64 70 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=1.19 $Y=0.49
+ $X2=1.19 $Y2=1.17
r162 63 67 0.446298 $w=6.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.02 $Y=0.49
+ $X2=1.02 $Y2=0.515
r163 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=0.49 $X2=1.19 $Y2=0.49
r164 57 59 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=2.815
r165 57 72 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=1.335
r166 47 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.19 $Y=1.185
+ $X2=1.19 $Y2=1.17
r167 44 46 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.975 $Y=1.185
+ $X2=4.975 $Y2=0.74
r168 43 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.62 $Y=1.26
+ $X2=4.545 $Y2=1.26
r169 42 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.9 $Y=1.26
+ $X2=4.975 $Y2=1.185
r170 42 43 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.9 $Y=1.26
+ $X2=4.62 $Y2=1.26
r171 39 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=1.185
+ $X2=4.545 $Y2=1.26
r172 39 41 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.545 $Y=1.185
+ $X2=4.545 $Y2=0.74
r173 38 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.19 $Y=1.26
+ $X2=4.115 $Y2=1.26
r174 37 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.47 $Y=1.26
+ $X2=4.545 $Y2=1.26
r175 37 38 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.47 $Y=1.26
+ $X2=4.19 $Y2=1.26
r176 34 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.115 $Y=1.185
+ $X2=4.115 $Y2=1.26
r177 34 36 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.115 $Y=1.185
+ $X2=4.115 $Y2=0.74
r178 33 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=1.26
+ $X2=3.615 $Y2=1.26
r179 32 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=1.26
+ $X2=4.115 $Y2=1.26
r180 32 33 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.04 $Y=1.26
+ $X2=3.69 $Y2=1.26
r181 29 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.615 $Y=1.185
+ $X2=3.615 $Y2=1.26
r182 29 31 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.615 $Y=1.185
+ $X2=3.615 $Y2=0.74
r183 28 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.26 $Y=1.26
+ $X2=3.185 $Y2=1.26
r184 27 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.54 $Y=1.26
+ $X2=3.615 $Y2=1.26
r185 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.54 $Y=1.26
+ $X2=3.26 $Y2=1.26
r186 24 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.185 $Y=1.185
+ $X2=3.185 $Y2=1.26
r187 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.185 $Y=1.185
+ $X2=3.185 $Y2=0.74
r188 23 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.76 $Y=1.26
+ $X2=2.685 $Y2=1.26
r189 22 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.11 $Y=1.26
+ $X2=3.185 $Y2=1.26
r190 22 23 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.11 $Y=1.26
+ $X2=2.76 $Y2=1.26
r191 19 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.685 $Y=1.185
+ $X2=2.685 $Y2=1.26
r192 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.685 $Y=1.185
+ $X2=2.685 $Y2=0.74
r193 18 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.33 $Y=1.26
+ $X2=2.255 $Y2=1.26
r194 17 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.61 $Y=1.26
+ $X2=2.685 $Y2=1.26
r195 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.61 $Y=1.26
+ $X2=2.33 $Y2=1.26
r196 14 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.255 $Y=1.185
+ $X2=2.255 $Y2=1.26
r197 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.255 $Y=1.185
+ $X2=2.255 $Y2=0.74
r198 13 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.9 $Y=1.26
+ $X2=1.825 $Y2=1.26
r199 12 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.18 $Y=1.26
+ $X2=2.255 $Y2=1.26
r200 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.18 $Y=1.26
+ $X2=1.9 $Y2=1.26
r201 9 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.185
+ $X2=1.825 $Y2=1.26
r202 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.825 $Y=1.185
+ $X2=1.825 $Y2=0.74
r203 8 47 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.355 $Y=1.26
+ $X2=1.19 $Y2=1.185
r204 7 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.26
+ $X2=1.825 $Y2=1.26
r205 7 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.75 $Y=1.26
+ $X2=1.355 $Y2=1.26
r206 2 59 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.84 $X2=0.78 $Y2=2.815
r207 2 57 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.84 $X2=0.78 $Y2=1.985
r208 1 67 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.37 $X2=0.77 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 66 67 68 69 97
c158 97 0 1.32147e-19 $X=8.625 $Y=1.515
c159 35 0 1.56455e-19 $X=7.195 $Y=0.74
c160 11 0 1.47232e-19 $X=5.835 $Y=0.74
r161 96 97 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.515
+ $X2=8.625 $Y2=1.515
r162 94 96 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.54 $Y=1.515
+ $X2=8.615 $Y2=1.515
r163 94 95 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=8.54
+ $Y=1.515 $X2=8.54 $Y2=1.515
r164 92 94 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=8.165 $Y=1.515
+ $X2=8.54 $Y2=1.515
r165 91 92 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.055 $Y=1.515
+ $X2=8.165 $Y2=1.515
r166 90 91 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.715 $Y=1.515
+ $X2=8.055 $Y2=1.515
r167 89 90 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.625 $Y=1.515
+ $X2=7.715 $Y2=1.515
r168 88 89 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=7.265 $Y=1.515
+ $X2=7.625 $Y2=1.515
r169 87 88 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.195 $Y=1.515
+ $X2=7.265 $Y2=1.515
r170 86 87 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=6.815 $Y=1.515
+ $X2=7.195 $Y2=1.515
r171 85 86 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=6.695 $Y=1.515
+ $X2=6.815 $Y2=1.515
r172 84 85 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=6.315 $Y=1.515
+ $X2=6.695 $Y2=1.515
r173 83 84 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=6.265 $Y=1.515
+ $X2=6.315 $Y2=1.515
r174 81 83 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.16 $Y=1.515
+ $X2=6.265 $Y2=1.515
r175 81 82 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=6.16
+ $Y=1.515 $X2=6.16 $Y2=1.515
r176 79 81 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=5.865 $Y=1.515
+ $X2=6.16 $Y2=1.515
r177 78 79 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.835 $Y=1.515
+ $X2=5.865 $Y2=1.515
r178 77 78 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.415 $Y=1.515
+ $X2=5.835 $Y2=1.515
r179 75 77 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.405 $Y=1.515
+ $X2=5.415 $Y2=1.515
r180 69 95 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=8.54 $Y2=1.565
r181 68 95 3.75214 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.54 $Y2=1.565
r182 67 68 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r183 66 67 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r184 65 66 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r185 65 82 21.4408 $w=4.28e-07 $l=8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.16 $Y2=1.565
r186 61 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=1.515
r187 61 63 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=0.74
r188 57 96 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.68
+ $X2=8.615 $Y2=1.515
r189 57 59 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.615 $Y=1.68
+ $X2=8.615 $Y2=2.4
r190 53 92 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.165 $Y=1.68
+ $X2=8.165 $Y2=1.515
r191 53 55 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.165 $Y=1.68
+ $X2=8.165 $Y2=2.4
r192 49 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=1.35
+ $X2=8.055 $Y2=1.515
r193 49 51 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.055 $Y=1.35
+ $X2=8.055 $Y2=0.74
r194 45 90 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.715 $Y=1.68
+ $X2=7.715 $Y2=1.515
r195 45 47 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.715 $Y=1.68
+ $X2=7.715 $Y2=2.4
r196 41 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.625 $Y=1.35
+ $X2=7.625 $Y2=1.515
r197 41 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.625 $Y=1.35
+ $X2=7.625 $Y2=0.74
r198 37 88 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.265 $Y=1.68
+ $X2=7.265 $Y2=1.515
r199 37 39 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.265 $Y=1.68
+ $X2=7.265 $Y2=2.4
r200 33 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.35
+ $X2=7.195 $Y2=1.515
r201 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.195 $Y=1.35
+ $X2=7.195 $Y2=0.74
r202 29 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.68
+ $X2=6.815 $Y2=1.515
r203 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.815 $Y=1.68
+ $X2=6.815 $Y2=2.4
r204 25 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.515
r205 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=0.74
r206 21 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.68
+ $X2=6.315 $Y2=1.515
r207 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.315 $Y=1.68
+ $X2=6.315 $Y2=2.4
r208 17 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.515
r209 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=0.74
r210 13 79 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.865 $Y=1.68
+ $X2=5.865 $Y2=1.515
r211 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.865 $Y=1.68
+ $X2=5.865 $Y2=2.4
r212 9 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.515
r213 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=0.74
r214 5 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.515
r215 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=0.74
r216 1 77 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.68
+ $X2=5.415 $Y2=1.515
r217 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.415 $Y=1.68
+ $X2=5.415 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%VPWR 1 2 3 4 5 16 18 24 28 32 36 40 44 48 50
+ 52 62 63 69 72 75 78
r107 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r109 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 62 63 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r114 60 63 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 59 62 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 59 60 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.69 $Y2=3.33
r118 57 59 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 56 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 56 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r121 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 53 66 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r123 53 55 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 52 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=1.79 $Y2=3.33
r125 52 55 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.625 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 50 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r127 50 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 50 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r129 46 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=3.33
r130 46 48 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=2.455
r131 45 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.69 $Y2=3.33
r132 44 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.69 $Y2=3.33
r133 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=3.855 $Y2=3.33
r134 40 43 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=3.69 $Y=2.09
+ $X2=3.69 $Y2=2.815
r135 38 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=3.33
r136 38 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=2.815
r137 37 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.74 $Y2=3.33
r138 36 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.69 $Y2=3.33
r139 36 37 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=2.905 $Y2=3.33
r140 32 35 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=2.74 $Y=2.09
+ $X2=2.74 $Y2=2.815
r141 30 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=3.245
+ $X2=2.74 $Y2=3.33
r142 30 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.74 $Y=3.245
+ $X2=2.74 $Y2=2.815
r143 29 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.79 $Y2=3.33
r144 28 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=2.74 $Y2=3.33
r145 28 29 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.575 $Y=3.33
+ $X2=1.955 $Y2=3.33
r146 24 27 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=1.79 $Y=2.09
+ $X2=1.79 $Y2=2.815
r147 22 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=3.245
+ $X2=1.79 $Y2=3.33
r148 22 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.79 $Y=3.245
+ $X2=1.79 $Y2=2.815
r149 18 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r150 16 66 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r151 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r152 5 48 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=1.84 $X2=4.69 $Y2=2.455
r153 4 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=1.84 $X2=3.69 $Y2=2.815
r154 4 40 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=1.84 $X2=3.69 $Y2=2.09
r155 3 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=1.84 $X2=2.74 $Y2=2.815
r156 3 32 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=1.84 $X2=2.74 $Y2=2.09
r157 2 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.84 $X2=1.79 $Y2=2.815
r158 2 24 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.84 $X2=1.79 $Y2=2.09
r159 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r160 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%A_239_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 42
+ 46 50 54 56 58 61 62 63 66 68 72 74 78 80 84 88 89 90 98 99 100
c166 56 0 5.39614e-20 $X=5.025 $Y=2.035
c167 50 0 6.43406e-20 $X=4.025 $Y=1.75
r168 94 95 1.20266 $w=4.68e-07 $l=5e-09 $layer=LI1_cond $X=4.26 $Y=2.115
+ $X2=4.26 $Y2=2.12
r169 92 94 2.03588 $w=4.68e-07 $l=8e-08 $layer=LI1_cond $X=4.26 $Y=2.035
+ $X2=4.26 $Y2=2.115
r170 90 92 7.25282 $w=4.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.26 $Y=1.75
+ $X2=4.26 $Y2=2.035
r171 84 87 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=8.88 $Y=2.115
+ $X2=8.88 $Y2=2.815
r172 82 87 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=2.905
+ $X2=8.88 $Y2=2.815
r173 81 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=2.99
+ $X2=7.94 $Y2=2.99
r174 80 82 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.88 $Y2=2.905
r175 80 81 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.025 $Y2=2.99
r176 76 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.99
r177 76 78 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.455
r178 75 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.125 $Y=2.99
+ $X2=7.04 $Y2=2.99
r179 74 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.94 $Y2=2.99
r180 74 75 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.125 $Y2=2.99
r181 70 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=2.905
+ $X2=7.04 $Y2=2.99
r182 70 72 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.04 $Y=2.905
+ $X2=7.04 $Y2=2.455
r183 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=2.99
+ $X2=6.09 $Y2=2.99
r184 68 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=2.99
+ $X2=7.04 $Y2=2.99
r185 68 69 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.955 $Y=2.99
+ $X2=6.255 $Y2=2.99
r186 64 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=2.905
+ $X2=6.09 $Y2=2.99
r187 64 66 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.09 $Y=2.905
+ $X2=6.09 $Y2=2.455
r188 62 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.925 $Y=2.99
+ $X2=6.09 $Y2=2.99
r189 62 63 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.925 $Y=2.99
+ $X2=5.355 $Y2=2.99
r190 59 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.19 $Y=2.905
+ $X2=5.355 $Y2=2.99
r191 59 61 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.19 $Y=2.905
+ $X2=5.19 $Y2=2.815
r192 58 97 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=2.12 $X2=5.19
+ $Y2=2.035
r193 58 61 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.19 $Y=2.12
+ $X2=5.19 $Y2=2.815
r194 57 92 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.495 $Y=2.035
+ $X2=4.26 $Y2=2.035
r195 56 97 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=2.035
+ $X2=5.19 $Y2=2.035
r196 56 57 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.025 $Y=2.035
+ $X2=4.495 $Y2=2.035
r197 54 95 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.19 $Y=2.815
+ $X2=4.19 $Y2=2.12
r198 51 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.325 $Y=1.75
+ $X2=3.2 $Y2=1.75
r199 50 90 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.025 $Y=1.75
+ $X2=4.26 $Y2=1.75
r200 50 51 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.025 $Y=1.75
+ $X2=3.325 $Y2=1.75
r201 46 48 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=3.2 $Y=2.115 $X2=3.2
+ $Y2=2.815
r202 44 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.835
+ $X2=3.2 $Y2=1.75
r203 44 46 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.2 $Y=1.835
+ $X2=3.2 $Y2=2.115
r204 43 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.375 $Y=1.75
+ $X2=2.25 $Y2=1.75
r205 42 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.075 $Y=1.75
+ $X2=3.2 $Y2=1.75
r206 42 43 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.075 $Y=1.75
+ $X2=2.375 $Y2=1.75
r207 38 40 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.25 $Y=2.115
+ $X2=2.25 $Y2=2.815
r208 36 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=1.835
+ $X2=2.25 $Y2=1.75
r209 36 38 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.25 $Y=1.835
+ $X2=2.25 $Y2=2.115
r210 34 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=1.75
+ $X2=2.25 $Y2=1.75
r211 34 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.125 $Y=1.75
+ $X2=1.425 $Y2=1.75
r212 30 32 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.3 $Y=2.115 $X2=1.3
+ $Y2=2.815
r213 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.3 $Y=1.835
+ $X2=1.425 $Y2=1.75
r214 28 30 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.3 $Y=1.835
+ $X2=1.3 $Y2=2.115
r215 9 87 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.815
r216 9 84 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.115
r217 8 78 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.805
+ $Y=1.84 $X2=7.94 $Y2=2.455
r218 7 72 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.905
+ $Y=1.84 $X2=7.04 $Y2=2.455
r219 6 66 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.84 $X2=6.09 $Y2=2.455
r220 5 97 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=1.84 $X2=5.19 $Y2=2.115
r221 5 61 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=1.84 $X2=5.19 $Y2=2.815
r222 4 94 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.84 $X2=4.19 $Y2=2.115
r223 4 54 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.84 $X2=4.19 $Y2=2.815
r224 3 48 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.84 $X2=3.24 $Y2=2.815
r225 3 46 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.84 $X2=3.24 $Y2=2.115
r226 2 40 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.84 $X2=2.29 $Y2=2.815
r227 2 38 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.84 $X2=2.29 $Y2=2.115
r228 1 32 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=1.84 $X2=1.34 $Y2=2.815
r229 1 30 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=1.84 $X2=1.34 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%Z 1 2 3 4 5 6 7 8 25 26 28 31 35 39 41 43 47
+ 51 53 57 63 64 69 70 72 73 75 77 78
c112 70 0 1.47232e-19 $X=6.645 $Y=0.975
c113 63 0 1.82517e-19 $X=5.455 $Y=1.665
c114 26 0 1.1822e-19 $X=5.59 $Y=1.55
r115 68 70 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.975
+ $X2=6.645 $Y2=0.975
r116 68 69 4.83878 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.975
+ $X2=6.315 $Y2=0.975
r117 63 78 20.7941 $w=2.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.455 $Y=1.665
+ $X2=5.04 $Y2=1.665
r118 63 64 1.18299 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=5.455 $Y=1.665
+ $X2=5.59 $Y2=1.665
r119 55 57 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=8.34 $Y=1.01
+ $X2=8.34 $Y2=0.78
r120 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=2.035
+ $X2=7.49 $Y2=2.035
r121 53 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=2.035
+ $X2=8.39 $Y2=2.035
r122 53 54 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.225 $Y=2.035
+ $X2=7.655 $Y2=2.035
r123 52 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=1.095
+ $X2=7.41 $Y2=1.095
r124 51 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.175 $Y=1.095
+ $X2=8.34 $Y2=1.01
r125 51 52 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.175 $Y=1.095
+ $X2=7.495 $Y2=1.095
r126 45 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=1.01
+ $X2=7.41 $Y2=1.095
r127 45 47 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.41 $Y=1.01
+ $X2=7.41 $Y2=0.78
r128 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.59 $Y2=2.035
r129 43 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.325 $Y=2.035
+ $X2=7.49 $Y2=2.035
r130 43 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.325 $Y=2.035
+ $X2=6.755 $Y2=2.035
r131 41 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=1.095
+ $X2=7.41 $Y2=1.095
r132 41 70 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.325 $Y=1.095
+ $X2=6.645 $Y2=1.095
r133 37 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=2.12
+ $X2=6.59 $Y2=2.035
r134 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.59 $Y=2.12
+ $X2=6.59 $Y2=2.615
r135 36 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=2.035
+ $X2=5.64 $Y2=2.035
r136 35 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=6.59 $Y2=2.035
r137 35 36 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=5.725 $Y2=2.035
r138 34 62 2.99957 $w=3.6e-07 $l=1.35e-07 $layer=LI1_cond $X=5.725 $Y=0.95
+ $X2=5.59 $Y2=0.95
r139 34 69 18.8873 $w=3.58e-07 $l=5.9e-07 $layer=LI1_cond $X=5.725 $Y=0.95
+ $X2=6.315 $Y2=0.95
r140 29 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=2.12
+ $X2=5.64 $Y2=2.035
r141 29 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.64 $Y=2.12
+ $X2=5.64 $Y2=2.57
r142 28 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=1.95
+ $X2=5.64 $Y2=2.035
r143 27 64 5.35987 $w=2.2e-07 $l=1.3775e-07 $layer=LI1_cond $X=5.64 $Y=1.78
+ $X2=5.59 $Y2=1.665
r144 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.64 $Y=1.78
+ $X2=5.64 $Y2=1.95
r145 26 64 5.35987 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=5.59 $Y=1.55
+ $X2=5.59 $Y2=1.665
r146 25 62 3.99943 $w=2.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.59 $Y=1.13
+ $X2=5.59 $Y2=0.95
r147 25 26 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.59 $Y=1.13
+ $X2=5.59 $Y2=1.55
r148 8 77 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=2.035
r149 7 75 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=7.355
+ $Y=1.84 $X2=7.49 $Y2=2.035
r150 6 72 600 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=1.84 $X2=6.59 $Y2=2.035
r151 6 39 600 $w=1.7e-07 $l=8.62554e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=1.84 $X2=6.59 $Y2=2.615
r152 5 66 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.84 $X2=5.64 $Y2=1.985
r153 5 31 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=1.84 $X2=5.64 $Y2=2.57
r154 4 57 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=8.13
+ $Y=0.37 $X2=8.34 $Y2=0.78
r155 3 47 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=7.27
+ $Y=0.37 $X2=7.41 $Y2=0.78
r156 2 68 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.37 $X2=6.48 $Y2=0.91
r157 1 62 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.37 $X2=5.62 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 70 71
c108 71 0 3.46022e-20 $X=8.88 $Y=0
r109 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r111 68 71 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=8.88
+ $Y2=0
r112 67 70 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=8.88
+ $Y2=0
r113 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r114 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r115 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r116 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r117 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r118 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r119 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r120 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r121 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r122 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 50 74 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.252 $Y2=0
r124 50 52 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.72 $Y2=0
r125 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r126 48 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r127 48 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r128 46 64 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.56
+ $Y2=0
r129 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.76
+ $Y2=0
r130 45 67 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.925 $Y=0
+ $X2=5.04 $Y2=0
r131 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0 $X2=4.76
+ $Y2=0
r132 43 61 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.6
+ $Y2=0
r133 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.83
+ $Y2=0
r134 42 64 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.56
+ $Y2=0
r135 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.83
+ $Y2=0
r136 40 58 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.64
+ $Y2=0
r137 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.9
+ $Y2=0
r138 39 61 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=3.6
+ $Y2=0
r139 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=2.9
+ $Y2=0
r140 37 55 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.68 $Y2=0
r141 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2
+ $Y2=0
r142 36 58 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.125 $Y=0
+ $X2=2.64 $Y2=0
r143 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2
+ $Y2=0
r144 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0
r145 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.76 $Y=0.085
+ $X2=4.76 $Y2=0.515
r146 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0
r147 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0.515
r148 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0
r149 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.9 $Y=0.085
+ $X2=2.9 $Y2=0.515
r150 20 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r151 20 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.515
r152 16 74 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.252 $Y2=0
r153 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.34 $Y2=0.515
r154 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.62
+ $Y=0.37 $X2=4.76 $Y2=0.515
r155 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.69
+ $Y=0.37 $X2=3.83 $Y2=0.515
r156 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.76
+ $Y=0.37 $X2=2.9 $Y2=0.515
r157 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.9
+ $Y=0.37 $X2=2.04 $Y2=0.515
r158 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.195
+ $Y=0.37 $X2=0.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_8%A_293_74# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 52 55 56 60 64 66 70 72 73 74 77 83
c165 70 0 1.32147e-19 $X=8.84 $Y=0.515
c166 56 0 1.56455e-19 $X=6.815 $Y=0.427
r167 79 81 8.13695 $w=3.28e-07 $l=2.33e-07 $layer=LI1_cond $X=6.98 $Y=0.427
+ $X2=6.98 $Y2=0.66
r168 77 79 3.03826 $w=3.28e-07 $l=8.7e-08 $layer=LI1_cond $X=6.98 $Y=0.34
+ $X2=6.98 $Y2=0.427
r169 68 70 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.84 $Y=0.425
+ $X2=8.84 $Y2=0.515
r170 67 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.005 $Y=0.34
+ $X2=7.84 $Y2=0.34
r171 66 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.675 $Y=0.34
+ $X2=8.84 $Y2=0.425
r172 66 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.675 $Y=0.34
+ $X2=8.005 $Y2=0.34
r173 62 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=0.425
+ $X2=7.84 $Y2=0.34
r174 62 64 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.84 $Y=0.425
+ $X2=7.84 $Y2=0.66
r175 61 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=0.34
+ $X2=6.98 $Y2=0.34
r176 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.84 $Y2=0.34
r177 60 61 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.145 $Y2=0.34
r178 57 76 2.60071 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.275 $Y=0.427
+ $X2=5.19 $Y2=0.427
r179 57 59 25.8882 $w=3.43e-07 $l=7.75e-07 $layer=LI1_cond $X=5.275 $Y=0.427
+ $X2=6.05 $Y2=0.427
r180 56 79 0.462083 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=6.815 $Y=0.427
+ $X2=6.98 $Y2=0.427
r181 56 59 25.5542 $w=3.43e-07 $l=7.65e-07 $layer=LI1_cond $X=6.815 $Y=0.427
+ $X2=6.05 $Y2=0.427
r182 53 55 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.19 $Y=1.21
+ $X2=5.19 $Y2=0.965
r183 52 76 5.29321 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.19 $Y=0.6
+ $X2=5.19 $Y2=0.427
r184 52 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.19 $Y=0.6
+ $X2=5.19 $Y2=0.965
r185 51 74 7.02821 $w=1.7e-07 $l=1.45774e-07 $layer=LI1_cond $X=4.415 $Y=1.295
+ $X2=4.29 $Y2=1.34
r186 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.105 $Y=1.295
+ $X2=5.19 $Y2=1.21
r187 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.105 $Y=1.295
+ $X2=4.415 $Y2=1.295
r188 46 74 0.00168595 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=4.29 $Y=1.21
+ $X2=4.29 $Y2=1.34
r189 46 48 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.29 $Y=1.21
+ $X2=4.29 $Y2=0.515
r190 45 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.485 $Y=1.385
+ $X2=3.36 $Y2=1.385
r191 44 74 7.02821 $w=1.7e-07 $l=1.45774e-07 $layer=LI1_cond $X=4.165 $Y=1.385
+ $X2=4.29 $Y2=1.34
r192 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.165 $Y=1.385
+ $X2=3.485 $Y2=1.385
r193 40 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=1.3
+ $X2=3.36 $Y2=1.385
r194 40 42 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=3.36 $Y=1.3
+ $X2=3.36 $Y2=0.515
r195 39 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=1.385
+ $X2=2.43 $Y2=1.385
r196 38 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=1.385
+ $X2=3.36 $Y2=1.385
r197 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.235 $Y=1.385
+ $X2=2.555 $Y2=1.385
r198 34 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=1.3
+ $X2=2.43 $Y2=1.385
r199 34 36 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=2.43 $Y=1.3
+ $X2=2.43 $Y2=0.515
r200 32 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.305 $Y=1.385
+ $X2=2.43 $Y2=1.385
r201 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.305 $Y=1.385
+ $X2=1.695 $Y2=1.385
r202 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.61 $Y=1.3
+ $X2=1.695 $Y2=1.385
r203 28 30 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.61 $Y=1.3
+ $X2=1.61 $Y2=0.515
r204 9 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r205 8 64 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=7.7
+ $Y=0.37 $X2=7.84 $Y2=0.66
r206 7 81 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.37 $X2=6.98 $Y2=0.66
r207 6 59 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.37 $X2=6.05 $Y2=0.515
r208 5 76 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.515
r209 5 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.965
r210 4 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.19
+ $Y=0.37 $X2=4.33 $Y2=0.515
r211 3 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.26
+ $Y=0.37 $X2=3.4 $Y2=0.515
r212 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.33
+ $Y=0.37 $X2=2.47 $Y2=0.515
r213 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.465
+ $Y=0.37 $X2=1.61 $Y2=0.515
.ends


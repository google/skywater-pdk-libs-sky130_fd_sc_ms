* File: sky130_fd_sc_ms__a2bb2oi_4.pxi.spice
* Created: Fri Aug 28 17:05:14 2020
* 
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%A2_N N_A2_N_M1017_g N_A2_N_M1018_g
+ N_A2_N_c_142_n N_A2_N_c_143_n N_A2_N_c_144_n N_A2_N_M1027_g A2_N A2_N A2_N
+ N_A2_N_c_146_n PM_SKY130_FD_SC_MS__A2BB2OI_4%A2_N
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%A1_N N_A1_N_M1020_g N_A1_N_M1006_g
+ N_A1_N_M1022_g A1_N A1_N N_A1_N_c_194_n PM_SKY130_FD_SC_MS__A2BB2OI_4%A1_N
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%A_117_392# N_A_117_392#_M1027_d
+ N_A_117_392#_M1017_d N_A_117_392#_c_239_n N_A_117_392#_M1003_g
+ N_A_117_392#_c_240_n N_A_117_392#_c_241_n N_A_117_392#_M1004_g
+ N_A_117_392#_M1015_g N_A_117_392#_c_243_n N_A_117_392#_M1014_g
+ N_A_117_392#_M1021_g N_A_117_392#_c_245_n N_A_117_392#_M1028_g
+ N_A_117_392#_c_246_n N_A_117_392#_M1023_g N_A_117_392#_c_248_n
+ N_A_117_392#_M1024_g N_A_117_392#_c_250_n N_A_117_392#_c_264_n
+ N_A_117_392#_c_251_n N_A_117_392#_c_252_n N_A_117_392#_c_253_n
+ N_A_117_392#_c_254_n N_A_117_392#_c_255_n N_A_117_392#_c_256_n
+ N_A_117_392#_c_257_n N_A_117_392#_c_258_n N_A_117_392#_c_259_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_4%A_117_392#
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%B2 N_B2_M1002_g N_B2_M1001_g N_B2_M1005_g
+ N_B2_M1009_g N_B2_M1007_g N_B2_M1012_g N_B2_M1026_g N_B2_M1013_g B2 B2 B2 B2
+ N_B2_c_384_n PM_SKY130_FD_SC_MS__A2BB2OI_4%B2
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%B1 N_B1_M1000_g N_B1_M1008_g N_B1_M1011_g
+ N_B1_M1010_g N_B1_M1025_g N_B1_M1016_g N_B1_M1029_g N_B1_M1019_g B1 B1 B1 B1
+ N_B1_c_470_n PM_SKY130_FD_SC_MS__A2BB2OI_4%B1
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%A_29_392# N_A_29_392#_M1017_s
+ N_A_29_392#_M1018_s N_A_29_392#_M1022_s N_A_29_392#_c_548_n
+ N_A_29_392#_c_549_n N_A_29_392#_c_550_n N_A_29_392#_c_551_n
+ N_A_29_392#_c_562_n N_A_29_392#_c_552_n N_A_29_392#_c_553_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_4%A_29_392#
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%VPWR N_VPWR_M1020_d N_VPWR_M1002_s
+ N_VPWR_M1007_s N_VPWR_M1008_d N_VPWR_M1016_d N_VPWR_c_594_n N_VPWR_c_595_n
+ N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n
+ N_VPWR_c_601_n N_VPWR_c_602_n N_VPWR_c_603_n VPWR N_VPWR_c_604_n
+ N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_593_n N_VPWR_c_608_n N_VPWR_c_609_n
+ N_VPWR_c_610_n PM_SKY130_FD_SC_MS__A2BB2OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%A_539_368# N_A_539_368#_M1015_s
+ N_A_539_368#_M1021_s N_A_539_368#_M1024_s N_A_539_368#_M1005_d
+ N_A_539_368#_M1026_d N_A_539_368#_M1010_s N_A_539_368#_M1019_s
+ N_A_539_368#_c_697_n N_A_539_368#_c_698_n N_A_539_368#_c_699_n
+ N_A_539_368#_c_715_n N_A_539_368#_c_700_n N_A_539_368#_c_721_n
+ N_A_539_368#_c_722_n N_A_539_368#_c_731_n N_A_539_368#_c_701_n
+ N_A_539_368#_c_739_n N_A_539_368#_c_702_n N_A_539_368#_c_750_n
+ N_A_539_368#_c_703_n N_A_539_368#_c_758_n N_A_539_368#_c_704_n
+ N_A_539_368#_c_705_n N_A_539_368#_c_706_n N_A_539_368#_c_744_n
+ N_A_539_368#_c_707_n N_A_539_368#_c_767_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_4%A_539_368#
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%Y N_Y_M1003_s N_Y_M1014_s N_Y_M1001_d
+ N_Y_M1012_d N_Y_M1015_d N_Y_M1023_d N_Y_c_826_n N_Y_c_814_n N_Y_c_830_n
+ N_Y_c_872_n N_Y_c_815_n N_Y_c_822_n N_Y_c_823_n N_Y_c_816_n N_Y_c_876_n
+ N_Y_c_817_n N_Y_c_818_n N_Y_c_844_n N_Y_c_824_n N_Y_c_819_n Y Y
+ PM_SKY130_FD_SC_MS__A2BB2OI_4%Y
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%VGND N_VGND_M1027_s N_VGND_M1006_d
+ N_VGND_M1004_d N_VGND_M1028_d N_VGND_M1000_s N_VGND_M1025_s N_VGND_c_900_n
+ N_VGND_c_901_n N_VGND_c_902_n N_VGND_c_903_n N_VGND_c_904_n N_VGND_c_905_n
+ N_VGND_c_906_n N_VGND_c_907_n N_VGND_c_908_n N_VGND_c_909_n N_VGND_c_910_n
+ N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n
+ N_VGND_c_916_n VGND N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_4%VGND
x_PM_SKY130_FD_SC_MS__A2BB2OI_4%A_914_74# N_A_914_74#_M1001_s
+ N_A_914_74#_M1009_s N_A_914_74#_M1013_s N_A_914_74#_M1011_d
+ N_A_914_74#_M1029_d N_A_914_74#_c_1011_n N_A_914_74#_c_1012_n
+ N_A_914_74#_c_1013_n N_A_914_74#_c_1014_n N_A_914_74#_c_1015_n
+ N_A_914_74#_c_1016_n N_A_914_74#_c_1017_n N_A_914_74#_c_1018_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_4%A_914_74#
cc_1 VNB N_A2_N_c_142_n 0.0251068f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.26
cc_2 VNB N_A2_N_c_143_n 0.085031f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.26
cc_3 VNB N_A2_N_c_144_n 0.0173058f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=1.185
cc_4 VNB A2_N 0.00316394f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_5 VNB N_A2_N_c_146_n 0.122325f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_6 VNB N_A1_N_M1006_g 0.033515f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.46
cc_7 VNB A1_N 0.00955002f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_8 VNB N_A1_N_c_194_n 0.028665f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.29
cc_9 VNB N_A_117_392#_c_239_n 0.0169153f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.46
cc_10 VNB N_A_117_392#_c_240_n 0.00949263f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=1.185
cc_11 VNB N_A_117_392#_c_241_n 0.0157654f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=0.74
cc_12 VNB N_A_117_392#_M1015_g 0.00745612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_117_392#_c_243_n 0.0157622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_117_392#_M1021_g 0.00579105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_117_392#_c_245_n 0.0192435f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_16 VNB N_A_117_392#_c_246_n 0.0143567f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.477
cc_17 VNB N_A_117_392#_M1023_g 0.00534292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_117_392#_c_248_n 0.0242974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_117_392#_M1024_g 0.00531883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_117_392#_c_250_n 0.00832624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_117_392#_c_251_n 0.00712702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_117_392#_c_252_n 0.0111501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_117_392#_c_253_n 0.00211602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_117_392#_c_254_n 0.0073757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_117_392#_c_255_n 0.00618867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_117_392#_c_256_n 0.00167115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_117_392#_c_257_n 0.0120196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_117_392#_c_258_n 0.0218365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_117_392#_c_259_n 0.0656908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B2_M1001_g 0.0299032f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.46
cc_31 VNB N_B2_M1009_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_32 VNB N_B2_M1012_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_33 VNB N_B2_M1013_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.555
cc_34 VNB B2 0.00365188f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_35 VNB N_B2_c_384_n 0.0715777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B1_M1000_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.46
cc_37 VNB N_B1_M1011_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=1.32 $Y2=1.185
cc_38 VNB N_B1_M1025_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B1_M1029_g 0.0326336f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_40 VNB B1 0.0257216f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_41 VNB N_B1_c_470_n 0.0751108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_593_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_814_n 0.00206283f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.585
cc_44 VNB N_Y_c_815_n 0.00178621f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.555
cc_45 VNB N_Y_c_816_n 0.00312482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_817_n 0.00135831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_818_n 0.00645039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_819_n 0.0149701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB Y 0.0116167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB Y 0.00762606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_900_n 0.0176435f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.585
cc_52 VNB N_VGND_c_901_n 0.00451436f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.477
cc_53 VNB N_VGND_c_902_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.477
cc_54 VNB N_VGND_c_903_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.555
cc_55 VNB N_VGND_c_904_n 0.0138193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_905_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_906_n 0.00497771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_907_n 0.0298226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_908_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_909_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_910_n 0.00538852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_911_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_912_n 0.00601765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_913_n 0.0731998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_914_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_915_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_916_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_917_n 0.0266297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_918_n 0.484031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_919_n 0.00613324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_914_74#_c_1011_n 0.0151254f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_72 VNB N_A_914_74#_c_1012_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.585
cc_73 VNB N_A_914_74#_c_1013_n 0.00472705f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_74 VNB N_A_914_74#_c_1014_n 0.0037698f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.605
cc_75 VNB N_A_914_74#_c_1015_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=1.477
cc_76 VNB N_A_914_74#_c_1016_n 0.0126873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_914_74#_c_1017_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_78 VNB N_A_914_74#_c_1018_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_A2_N_M1017_g 0.0296314f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.46
cc_80 VPB N_A2_N_M1018_g 0.0215973f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.46
cc_81 VPB N_A2_N_c_143_n 0.0293941f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.26
cc_82 VPB A2_N 0.00261477f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_83 VPB N_A1_N_M1020_g 0.0211945f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.46
cc_84 VPB N_A1_N_M1022_g 0.0298886f $X=-0.19 $Y=1.66 $X2=1.32 $Y2=1.185
cc_85 VPB A1_N 0.00756726f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_86 VPB N_A1_N_c_194_n 0.0181778f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.29
cc_87 VPB N_A_117_392#_M1015_g 0.0267092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_117_392#_M1021_g 0.0205091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_117_392#_M1023_g 0.0202624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_117_392#_M1024_g 0.02117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_117_392#_c_264_n 0.00174737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_B2_M1002_g 0.0202491f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.46
cc_93 VPB N_B2_M1005_g 0.020498f $X=-0.19 $Y=1.66 $X2=1.32 $Y2=1.185
cc_94 VPB N_B2_M1007_g 0.0204973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_B2_M1026_g 0.0208119f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.605
cc_96 VPB B2 0.0100717f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_97 VPB N_B2_c_384_n 0.0116115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_B1_M1008_g 0.0208115f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.46
cc_99 VPB N_B1_M1010_g 0.0204973f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.84
cc_100 VPB N_B1_M1016_g 0.020498f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.585
cc_101 VPB N_B1_M1019_g 0.027583f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.555
cc_102 VPB B1 0.0213025f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_103 VPB N_B1_c_470_n 0.011923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_29_392#_c_548_n 0.0398572f $X=-0.19 $Y=1.66 $X2=1.32 $Y2=0.74
cc_105 VPB N_A_29_392#_c_549_n 0.00438754f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_106 VPB N_A_29_392#_c_550_n 0.00969936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_29_392#_c_551_n 0.00251695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_29_392#_c_552_n 0.00288429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_29_392#_c_553_n 0.0151573f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.605
cc_110 VPB N_VPWR_c_594_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_595_n 0.0810193f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.29
cc_112 VPB N_VPWR_c_596_n 0.00768638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_597_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.477
cc_114 VPB N_VPWR_c_598_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_599_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_116 VPB N_VPWR_c_600_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_601_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_602_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_603_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_604_n 0.037172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_605_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_606_n 0.0245612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_593_n 0.114962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_608_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_609_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_610_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_539_368#_c_697_n 0.0220728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_539_368#_c_698_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.477
cc_129 VPB N_A_539_368#_c_699_n 0.00767107f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.477
cc_130 VPB N_A_539_368#_c_700_n 0.00388794f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.925
cc_131 VPB N_A_539_368#_c_701_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_539_368#_c_702_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_539_368#_c_703_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_539_368#_c_704_n 0.0075508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_539_368#_c_705_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_539_368#_c_706_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_539_368#_c_707_n 0.00322238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_Y_c_822_n 0.00749758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_Y_c_823_n 0.00266104f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.925
cc_140 VPB N_Y_c_824_n 0.00116786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB Y 3.55613e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 N_A2_N_M1018_g N_A1_N_M1020_g 0.0106332f $X=0.945 $Y=2.46 $X2=0 $Y2=0
cc_143 N_A2_N_c_143_n N_A1_N_M1006_g 0.0036141f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_144 N_A2_N_c_144_n N_A1_N_M1006_g 0.0176901f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_145 N_A2_N_c_143_n A1_N 0.00445792f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_146 N_A2_N_c_142_n N_A1_N_c_194_n 0.00410217f $X=1.245 $Y=1.26 $X2=0 $Y2=0
cc_147 N_A2_N_c_143_n N_A1_N_c_194_n 0.013805f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_148 N_A2_N_M1017_g N_A_117_392#_c_264_n 0.00487324f $X=0.495 $Y=2.46 $X2=0
+ $Y2=0
cc_149 N_A2_N_M1018_g N_A_117_392#_c_264_n 0.0152803f $X=0.945 $Y=2.46 $X2=0
+ $Y2=0
cc_150 N_A2_N_c_143_n N_A_117_392#_c_264_n 0.0359645f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_151 A2_N N_A_117_392#_c_264_n 0.0329548f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_152 N_A2_N_c_142_n N_A_117_392#_c_251_n 0.0153082f $X=1.245 $Y=1.26 $X2=0
+ $Y2=0
cc_153 N_A2_N_c_143_n N_A_117_392#_c_251_n 0.0104437f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_154 N_A2_N_c_144_n N_A_117_392#_c_251_n 0.00832909f $X=1.32 $Y=1.185 $X2=0
+ $Y2=0
cc_155 N_A2_N_c_143_n N_A_117_392#_c_252_n 0.00589853f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_156 A2_N N_A_117_392#_c_252_n 0.0136491f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A2_N_c_146_n N_A_117_392#_c_252_n 0.00181472f $X=0.29 $Y=0.585 $X2=0
+ $Y2=0
cc_158 N_A2_N_c_144_n N_A_117_392#_c_253_n 8.30306e-19 $X=1.32 $Y=1.185 $X2=0
+ $Y2=0
cc_159 N_A2_N_M1017_g N_A_29_392#_c_548_n 0.013679f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_160 N_A2_N_M1018_g N_A_29_392#_c_548_n 7.38944e-19 $X=0.945 $Y=2.46 $X2=0
+ $Y2=0
cc_161 N_A2_N_c_143_n N_A_29_392#_c_548_n 0.00218185f $X=1.035 $Y=1.26 $X2=0
+ $Y2=0
cc_162 A2_N N_A_29_392#_c_548_n 0.027329f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_163 N_A2_N_M1017_g N_A_29_392#_c_549_n 0.0115958f $X=0.495 $Y=2.46 $X2=0
+ $Y2=0
cc_164 N_A2_N_M1018_g N_A_29_392#_c_549_n 0.0137017f $X=0.945 $Y=2.46 $X2=0
+ $Y2=0
cc_165 N_A2_N_M1017_g N_A_29_392#_c_550_n 0.00291744f $X=0.495 $Y=2.46 $X2=0
+ $Y2=0
cc_166 N_A2_N_c_142_n N_A_29_392#_c_551_n 0.00264727f $X=1.245 $Y=1.26 $X2=0
+ $Y2=0
cc_167 N_A2_N_c_142_n N_A_29_392#_c_562_n 2.60891e-19 $X=1.245 $Y=1.26 $X2=0
+ $Y2=0
cc_168 N_A2_N_M1017_g N_VPWR_c_604_n 0.00333896f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_169 N_A2_N_M1018_g N_VPWR_c_604_n 0.00333926f $X=0.945 $Y=2.46 $X2=0 $Y2=0
cc_170 N_A2_N_M1017_g N_VPWR_c_593_n 0.00426392f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_171 N_A2_N_M1018_g N_VPWR_c_593_n 0.00422798f $X=0.945 $Y=2.46 $X2=0 $Y2=0
cc_172 N_A2_N_c_143_n N_VGND_c_900_n 0.00192874f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_173 N_A2_N_c_144_n N_VGND_c_900_n 0.011643f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_174 A2_N N_VGND_c_900_n 0.0195009f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A2_N_c_146_n N_VGND_c_900_n 0.00569436f $X=0.29 $Y=0.585 $X2=0 $Y2=0
cc_176 N_A2_N_c_144_n N_VGND_c_901_n 4.85748e-19 $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_177 A2_N N_VGND_c_907_n 0.0105202f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_178 N_A2_N_c_146_n N_VGND_c_907_n 0.00476771f $X=0.29 $Y=0.585 $X2=0 $Y2=0
cc_179 N_A2_N_c_144_n N_VGND_c_909_n 0.00383152f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_180 N_A2_N_c_144_n N_VGND_c_918_n 0.00757637f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_181 A2_N N_VGND_c_918_n 0.0112802f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_182 N_A2_N_c_146_n N_VGND_c_918_n 0.00333647f $X=0.29 $Y=0.585 $X2=0 $Y2=0
cc_183 N_A1_N_M1006_g N_A_117_392#_c_239_n 0.0280367f $X=1.75 $Y=0.74 $X2=0
+ $Y2=0
cc_184 A1_N N_A_117_392#_c_240_n 0.00377293f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_185 A1_N N_A_117_392#_M1015_g 0.00613866f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A1_N_c_194_n N_A_117_392#_c_264_n 0.00149611f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_187 N_A1_N_c_194_n N_A_117_392#_c_251_n 0.0018193f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_188 N_A1_N_M1006_g N_A_117_392#_c_253_n 8.30306e-19 $X=1.75 $Y=0.74 $X2=0
+ $Y2=0
cc_189 A1_N N_A_117_392#_c_254_n 0.00455708f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_190 A1_N N_A_117_392#_c_256_n 0.00480329f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A1_N_c_194_n N_A_117_392#_c_256_n 0.00368739f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_192 N_A1_N_M1006_g N_A_117_392#_c_257_n 0.0145425f $X=1.75 $Y=0.74 $X2=0
+ $Y2=0
cc_193 A1_N N_A_117_392#_c_257_n 0.04954f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A1_N_c_194_n N_A_117_392#_c_257_n 0.00416999f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_195 A1_N N_A_117_392#_c_259_n 4.03225e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A1_N_c_194_n N_A_117_392#_c_259_n 9.7315e-19 $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_197 N_A1_N_M1020_g N_A_29_392#_c_549_n 0.00101073f $X=1.395 $Y=2.46 $X2=0
+ $Y2=0
cc_198 N_A1_N_M1020_g N_A_29_392#_c_551_n 4.63009e-19 $X=1.395 $Y=2.46 $X2=0
+ $Y2=0
cc_199 N_A1_N_M1020_g N_A_29_392#_c_562_n 0.0159055f $X=1.395 $Y=2.46 $X2=0
+ $Y2=0
cc_200 N_A1_N_M1022_g N_A_29_392#_c_562_n 0.0128923f $X=1.845 $Y=2.46 $X2=0
+ $Y2=0
cc_201 A1_N N_A_29_392#_c_562_n 0.0226372f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A1_N_c_194_n N_A_29_392#_c_562_n 0.00191796f $X=1.77 $Y=1.635 $X2=0
+ $Y2=0
cc_203 N_A1_N_M1022_g N_A_29_392#_c_552_n 8.84614e-19 $X=1.845 $Y=2.46 $X2=0
+ $Y2=0
cc_204 A1_N N_A_29_392#_c_552_n 0.0258724f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A1_N_M1020_g N_A_29_392#_c_553_n 6.67908e-19 $X=1.395 $Y=2.46 $X2=0
+ $Y2=0
cc_206 N_A1_N_M1022_g N_A_29_392#_c_553_n 0.0120613f $X=1.845 $Y=2.46 $X2=0
+ $Y2=0
cc_207 N_A1_N_M1020_g N_VPWR_c_594_n 0.0114961f $X=1.395 $Y=2.46 $X2=0 $Y2=0
cc_208 N_A1_N_M1022_g N_VPWR_c_594_n 0.002979f $X=1.845 $Y=2.46 $X2=0 $Y2=0
cc_209 N_A1_N_M1022_g N_VPWR_c_595_n 0.005209f $X=1.845 $Y=2.46 $X2=0 $Y2=0
cc_210 N_A1_N_M1020_g N_VPWR_c_604_n 0.00460063f $X=1.395 $Y=2.46 $X2=0 $Y2=0
cc_211 N_A1_N_M1020_g N_VPWR_c_593_n 0.00908665f $X=1.395 $Y=2.46 $X2=0 $Y2=0
cc_212 N_A1_N_M1022_g N_VPWR_c_593_n 0.00987399f $X=1.845 $Y=2.46 $X2=0 $Y2=0
cc_213 N_A1_N_M1006_g N_VGND_c_900_n 5.07446e-19 $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_N_M1006_g N_VGND_c_901_n 0.0114017f $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A1_N_M1006_g N_VGND_c_909_n 0.00383152f $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A1_N_M1006_g N_VGND_c_918_n 0.00757637f $X=1.75 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_117_392#_M1024_g N_B2_M1002_g 0.015594f $X=4.395 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_117_392#_c_248_n B2 0.00520824f $X=4.305 $Y=1.475 $X2=0 $Y2=0
cc_219 N_A_117_392#_M1024_g B2 0.00633961f $X=4.395 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_117_392#_c_248_n N_B2_c_384_n 0.015594f $X=4.305 $Y=1.475 $X2=0 $Y2=0
cc_221 N_A_117_392#_c_264_n N_A_29_392#_c_548_n 0.0268676f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_222 N_A_117_392#_M1017_d N_A_29_392#_c_549_n 0.00165831f $X=0.585 $Y=1.96
+ $X2=0 $Y2=0
cc_223 N_A_117_392#_c_264_n N_A_29_392#_c_549_n 0.0139027f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_224 N_A_117_392#_c_264_n N_A_29_392#_c_551_n 0.0069809f $X=0.72 $Y=2.105
+ $X2=0 $Y2=0
cc_225 N_A_117_392#_c_251_n N_A_29_392#_c_551_n 0.00503831f $X=1.45 $Y=1.215
+ $X2=0 $Y2=0
cc_226 N_A_117_392#_c_251_n N_A_29_392#_c_562_n 0.00383038f $X=1.45 $Y=1.215
+ $X2=0 $Y2=0
cc_227 N_A_117_392#_c_256_n N_A_29_392#_c_562_n 0.00271207f $X=1.535 $Y=1.215
+ $X2=0 $Y2=0
cc_228 N_A_117_392#_M1015_g N_VPWR_c_595_n 0.00333896f $X=3.045 $Y=2.4 $X2=0
+ $Y2=0
cc_229 N_A_117_392#_M1021_g N_VPWR_c_595_n 0.00333896f $X=3.495 $Y=2.4 $X2=0
+ $Y2=0
cc_230 N_A_117_392#_M1023_g N_VPWR_c_595_n 0.00333896f $X=3.945 $Y=2.4 $X2=0
+ $Y2=0
cc_231 N_A_117_392#_M1024_g N_VPWR_c_595_n 0.00333896f $X=4.395 $Y=2.4 $X2=0
+ $Y2=0
cc_232 N_A_117_392#_M1015_g N_VPWR_c_593_n 0.00427818f $X=3.045 $Y=2.4 $X2=0
+ $Y2=0
cc_233 N_A_117_392#_M1021_g N_VPWR_c_593_n 0.00422685f $X=3.495 $Y=2.4 $X2=0
+ $Y2=0
cc_234 N_A_117_392#_M1023_g N_VPWR_c_593_n 0.00422685f $X=3.945 $Y=2.4 $X2=0
+ $Y2=0
cc_235 N_A_117_392#_M1024_g N_VPWR_c_593_n 0.00422796f $X=4.395 $Y=2.4 $X2=0
+ $Y2=0
cc_236 N_A_117_392#_M1015_g N_A_539_368#_c_697_n 0.0160259f $X=3.045 $Y=2.4
+ $X2=0 $Y2=0
cc_237 N_A_117_392#_M1021_g N_A_539_368#_c_697_n 7.29961e-19 $X=3.495 $Y=2.4
+ $X2=0 $Y2=0
cc_238 N_A_117_392#_c_254_n N_A_539_368#_c_697_n 0.0197823f $X=2.995 $Y=1.34
+ $X2=0 $Y2=0
cc_239 N_A_117_392#_c_259_n N_A_539_368#_c_697_n 0.00729208f $X=3.585 $Y=1.385
+ $X2=0 $Y2=0
cc_240 N_A_117_392#_M1015_g N_A_539_368#_c_698_n 0.0116345f $X=3.045 $Y=2.4
+ $X2=0 $Y2=0
cc_241 N_A_117_392#_M1021_g N_A_539_368#_c_698_n 0.0116345f $X=3.495 $Y=2.4
+ $X2=0 $Y2=0
cc_242 N_A_117_392#_M1015_g N_A_539_368#_c_699_n 0.00291744f $X=3.045 $Y=2.4
+ $X2=0 $Y2=0
cc_243 N_A_117_392#_M1015_g N_A_539_368#_c_715_n 6.45773e-19 $X=3.045 $Y=2.4
+ $X2=0 $Y2=0
cc_244 N_A_117_392#_M1021_g N_A_539_368#_c_715_n 0.0139917f $X=3.495 $Y=2.4
+ $X2=0 $Y2=0
cc_245 N_A_117_392#_M1023_g N_A_539_368#_c_715_n 0.0139917f $X=3.945 $Y=2.4
+ $X2=0 $Y2=0
cc_246 N_A_117_392#_M1024_g N_A_539_368#_c_715_n 6.45773e-19 $X=4.395 $Y=2.4
+ $X2=0 $Y2=0
cc_247 N_A_117_392#_M1023_g N_A_539_368#_c_700_n 0.0116345f $X=3.945 $Y=2.4
+ $X2=0 $Y2=0
cc_248 N_A_117_392#_M1024_g N_A_539_368#_c_700_n 0.0135505f $X=4.395 $Y=2.4
+ $X2=0 $Y2=0
cc_249 N_A_117_392#_M1024_g N_A_539_368#_c_721_n 0.00244698f $X=4.395 $Y=2.4
+ $X2=0 $Y2=0
cc_250 N_A_117_392#_M1023_g N_A_539_368#_c_722_n 6.26485e-19 $X=3.945 $Y=2.4
+ $X2=0 $Y2=0
cc_251 N_A_117_392#_M1024_g N_A_539_368#_c_722_n 0.0105282f $X=4.395 $Y=2.4
+ $X2=0 $Y2=0
cc_252 N_A_117_392#_M1021_g N_A_539_368#_c_706_n 0.00194226f $X=3.495 $Y=2.4
+ $X2=0 $Y2=0
cc_253 N_A_117_392#_M1023_g N_A_539_368#_c_706_n 0.00194226f $X=3.945 $Y=2.4
+ $X2=0 $Y2=0
cc_254 N_A_117_392#_c_239_n N_Y_c_826_n 0.00273433f $X=2.22 $Y=1.22 $X2=0 $Y2=0
cc_255 N_A_117_392#_c_257_n N_Y_c_826_n 0.0176844f $X=2.575 $Y=1.34 $X2=0 $Y2=0
cc_256 N_A_117_392#_c_258_n N_Y_c_826_n 6.28576e-19 $X=2.575 $Y=1.385 $X2=0
+ $Y2=0
cc_257 N_A_117_392#_c_239_n N_Y_c_814_n 0.004978f $X=2.22 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A_117_392#_c_241_n N_Y_c_830_n 0.00947324f $X=2.65 $Y=1.22 $X2=0 $Y2=0
cc_259 N_A_117_392#_c_243_n N_Y_c_830_n 0.00947324f $X=3.08 $Y=1.22 $X2=0 $Y2=0
cc_260 N_A_117_392#_c_257_n N_Y_c_830_n 0.0442631f $X=2.575 $Y=1.34 $X2=0 $Y2=0
cc_261 N_A_117_392#_c_259_n N_Y_c_830_n 5.58069e-19 $X=3.585 $Y=1.385 $X2=0
+ $Y2=0
cc_262 N_A_117_392#_M1021_g N_Y_c_822_n 0.0152733f $X=3.495 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A_117_392#_c_246_n N_Y_c_822_n 0.0030813f $X=3.855 $Y=1.475 $X2=0 $Y2=0
cc_264 N_A_117_392#_M1023_g N_Y_c_822_n 0.0119502f $X=3.945 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A_117_392#_c_255_n N_Y_c_822_n 0.0168996f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_266 N_A_117_392#_M1015_g N_Y_c_823_n 0.00336f $X=3.045 $Y=2.4 $X2=0 $Y2=0
cc_267 N_A_117_392#_c_255_n N_Y_c_823_n 0.0145791f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_268 N_A_117_392#_c_259_n N_Y_c_823_n 0.00217549f $X=3.585 $Y=1.385 $X2=0
+ $Y2=0
cc_269 N_A_117_392#_c_245_n N_Y_c_816_n 0.0115138f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_270 N_A_117_392#_c_246_n N_Y_c_816_n 0.0105789f $X=3.855 $Y=1.475 $X2=0 $Y2=0
cc_271 N_A_117_392#_c_255_n N_Y_c_816_n 0.0132645f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_272 N_A_117_392#_c_255_n N_Y_c_844_n 0.0147027f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_273 N_A_117_392#_c_259_n N_Y_c_844_n 6.18925e-19 $X=3.585 $Y=1.385 $X2=0
+ $Y2=0
cc_274 N_A_117_392#_M1023_g N_Y_c_824_n 0.00568574f $X=3.945 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A_117_392#_M1024_g N_Y_c_824_n 0.00242454f $X=4.395 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A_117_392#_c_248_n N_Y_c_819_n 0.00780731f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_277 N_A_117_392#_c_245_n Y 0.00559274f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A_117_392#_M1021_g Y 8.65913e-19 $X=3.495 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A_117_392#_c_245_n Y 0.00168909f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_280 N_A_117_392#_M1023_g Y 0.00514907f $X=3.945 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A_117_392#_c_248_n Y 0.0124449f $X=4.305 $Y=1.475 $X2=0 $Y2=0
cc_282 N_A_117_392#_M1024_g Y 0.00131661f $X=4.395 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A_117_392#_c_250_n Y 0.00582537f $X=3.945 $Y=1.475 $X2=0 $Y2=0
cc_284 N_A_117_392#_c_255_n Y 0.0183585f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_285 N_A_117_392#_c_251_n N_VGND_c_900_n 0.0244338f $X=1.45 $Y=1.215 $X2=0
+ $Y2=0
cc_286 N_A_117_392#_c_253_n N_VGND_c_900_n 0.0225498f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_287 N_A_117_392#_c_239_n N_VGND_c_901_n 0.00242169f $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_288 N_A_117_392#_c_253_n N_VGND_c_901_n 0.0194859f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_289 N_A_117_392#_c_257_n N_VGND_c_901_n 0.0161099f $X=2.575 $Y=1.34 $X2=0
+ $Y2=0
cc_290 N_A_117_392#_c_239_n N_VGND_c_902_n 4.26297e-19 $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_291 N_A_117_392#_c_241_n N_VGND_c_902_n 0.00720343f $X=2.65 $Y=1.22 $X2=0
+ $Y2=0
cc_292 N_A_117_392#_c_243_n N_VGND_c_902_n 0.00706632f $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_293 N_A_117_392#_c_245_n N_VGND_c_902_n 4.05984e-19 $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_294 N_A_117_392#_c_243_n N_VGND_c_903_n 0.00383152f $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_295 N_A_117_392#_c_245_n N_VGND_c_903_n 0.00383152f $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_296 N_A_117_392#_c_243_n N_VGND_c_904_n 4.05984e-19 $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_297 N_A_117_392#_c_245_n N_VGND_c_904_n 0.00812981f $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_298 N_A_117_392#_c_253_n N_VGND_c_909_n 0.00749631f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_299 N_A_117_392#_c_239_n N_VGND_c_911_n 0.00434272f $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_300 N_A_117_392#_c_241_n N_VGND_c_911_n 0.00383152f $X=2.65 $Y=1.22 $X2=0
+ $Y2=0
cc_301 N_A_117_392#_c_239_n N_VGND_c_918_n 0.00820742f $X=2.22 $Y=1.22 $X2=0
+ $Y2=0
cc_302 N_A_117_392#_c_241_n N_VGND_c_918_n 0.00373475f $X=2.65 $Y=1.22 $X2=0
+ $Y2=0
cc_303 N_A_117_392#_c_243_n N_VGND_c_918_n 0.00373475f $X=3.08 $Y=1.22 $X2=0
+ $Y2=0
cc_304 N_A_117_392#_c_245_n N_VGND_c_918_n 0.00373475f $X=3.51 $Y=1.22 $X2=0
+ $Y2=0
cc_305 N_A_117_392#_c_253_n N_VGND_c_918_n 0.0062048f $X=1.535 $Y=0.515 $X2=0
+ $Y2=0
cc_306 N_B2_M1013_g N_B1_M1000_g 0.019323f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_307 N_B2_M1026_g N_B1_M1008_g 0.0164444f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_308 N_B2_M1026_g B1 2.74111e-19 $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_309 B2 B1 0.0122682f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_310 N_B2_c_384_n B1 0.00116712f $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_311 B2 N_B1_c_470_n 0.00146902f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_312 N_B2_c_384_n N_B1_c_470_n 0.0164444f $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_313 N_B2_M1002_g N_VPWR_c_595_n 0.00517089f $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_314 N_B2_M1002_g N_VPWR_c_596_n 0.00120619f $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_315 N_B2_M1005_g N_VPWR_c_596_n 0.0027763f $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_316 N_B2_M1007_g N_VPWR_c_597_n 0.002979f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_317 N_B2_M1026_g N_VPWR_c_597_n 0.0124151f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_318 N_B2_M1026_g N_VPWR_c_598_n 5.43099e-19 $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_319 N_B2_M1026_g N_VPWR_c_600_n 0.00460063f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_320 N_B2_M1005_g N_VPWR_c_605_n 0.005209f $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_321 N_B2_M1007_g N_VPWR_c_605_n 0.005209f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_322 N_B2_M1002_g N_VPWR_c_593_n 0.00977588f $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_323 N_B2_M1005_g N_VPWR_c_593_n 0.00982266f $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_324 N_B2_M1007_g N_VPWR_c_593_n 0.00982266f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_325 N_B2_M1026_g N_VPWR_c_593_n 0.00908665f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_326 N_B2_M1002_g N_A_539_368#_c_700_n 0.00347836f $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_327 N_B2_M1002_g N_A_539_368#_c_721_n 8.84614e-19 $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_328 B2 N_A_539_368#_c_721_n 0.0235495f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_329 N_B2_M1002_g N_A_539_368#_c_722_n 0.0105282f $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_330 N_B2_M1005_g N_A_539_368#_c_722_n 6.26485e-19 $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_331 N_B2_M1002_g N_A_539_368#_c_731_n 0.012931f $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_332 N_B2_M1005_g N_A_539_368#_c_731_n 0.012931f $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_333 B2 N_A_539_368#_c_731_n 0.0391869f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_334 N_B2_c_384_n N_A_539_368#_c_731_n 4.8724e-19 $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_335 N_B2_M1002_g N_A_539_368#_c_701_n 6.50516e-19 $X=4.845 $Y=2.4 $X2=0 $Y2=0
cc_336 N_B2_M1005_g N_A_539_368#_c_701_n 0.0119382f $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_337 N_B2_M1007_g N_A_539_368#_c_701_n 0.0121366f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_338 N_B2_M1026_g N_A_539_368#_c_701_n 6.74232e-19 $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_339 N_B2_M1007_g N_A_539_368#_c_739_n 0.012931f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_340 N_B2_M1026_g N_A_539_368#_c_739_n 0.0194018f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_341 B2 N_A_539_368#_c_739_n 0.0290059f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_342 N_B2_c_384_n N_A_539_368#_c_739_n 4.90062e-19 $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_343 N_B2_M1026_g N_A_539_368#_c_702_n 3.62369e-19 $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_344 N_B2_M1005_g N_A_539_368#_c_744_n 8.84614e-19 $X=5.295 $Y=2.4 $X2=0 $Y2=0
cc_345 N_B2_M1007_g N_A_539_368#_c_744_n 8.84614e-19 $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_346 B2 N_A_539_368#_c_744_n 0.0235495f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_347 N_B2_c_384_n N_A_539_368#_c_744_n 5.52655e-19 $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_348 N_B2_M1026_g N_A_539_368#_c_707_n 4.63009e-19 $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_349 N_B2_M1001_g N_Y_c_817_n 0.00262032f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_350 N_B2_c_384_n N_Y_c_817_n 0.00243719f $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_351 N_B2_M1009_g N_Y_c_818_n 0.0140439f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_352 N_B2_M1012_g N_Y_c_818_n 0.0140439f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_353 N_B2_M1013_g N_Y_c_818_n 0.0054657f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_354 N_B2_c_384_n N_Y_c_818_n 0.00465635f $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_355 B2 N_Y_c_824_n 0.00483333f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_356 N_B2_M1001_g N_Y_c_819_n 0.0159385f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_357 B2 N_Y_c_819_n 0.111129f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_358 N_B2_c_384_n N_Y_c_819_n 0.0020685f $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_359 N_B2_M1001_g Y 0.005219f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_360 B2 Y 0.0277233f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_361 N_B2_c_384_n Y 2.69051e-19 $X=6.2 $Y=1.515 $X2=0 $Y2=0
cc_362 N_B2_M1013_g N_VGND_c_905_n 6.37019e-19 $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_363 N_B2_M1001_g N_VGND_c_913_n 0.00291649f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_364 N_B2_M1009_g N_VGND_c_913_n 0.00291649f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_365 N_B2_M1012_g N_VGND_c_913_n 0.00291649f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_366 N_B2_M1013_g N_VGND_c_913_n 0.00291649f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_367 N_B2_M1001_g N_VGND_c_918_n 0.0036412f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_368 N_B2_M1009_g N_VGND_c_918_n 0.00359121f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_369 N_B2_M1012_g N_VGND_c_918_n 0.00359121f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_370 N_B2_M1013_g N_VGND_c_918_n 0.00359219f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_371 N_B2_M1001_g N_A_914_74#_c_1011_n 0.0104692f $X=4.91 $Y=0.74 $X2=0 $Y2=0
cc_372 N_B2_M1009_g N_A_914_74#_c_1011_n 0.010218f $X=5.34 $Y=0.74 $X2=0 $Y2=0
cc_373 N_B2_M1012_g N_A_914_74#_c_1011_n 0.0101492f $X=5.77 $Y=0.74 $X2=0 $Y2=0
cc_374 N_B2_M1013_g N_A_914_74#_c_1011_n 0.014175f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_375 N_B2_M1013_g N_A_914_74#_c_1014_n 0.0017668f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_376 N_B1_M1008_g N_VPWR_c_597_n 5.43099e-19 $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_377 N_B1_M1008_g N_VPWR_c_598_n 0.0124151f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_378 N_B1_M1010_g N_VPWR_c_598_n 0.002979f $X=7.095 $Y=2.4 $X2=0 $Y2=0
cc_379 N_B1_M1016_g N_VPWR_c_599_n 0.0027763f $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_380 N_B1_M1019_g N_VPWR_c_599_n 0.0027763f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_381 N_B1_M1008_g N_VPWR_c_600_n 0.00460063f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_382 N_B1_M1010_g N_VPWR_c_602_n 0.005209f $X=7.095 $Y=2.4 $X2=0 $Y2=0
cc_383 N_B1_M1016_g N_VPWR_c_602_n 0.005209f $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_384 N_B1_M1019_g N_VPWR_c_606_n 0.005209f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_385 N_B1_M1008_g N_VPWR_c_593_n 0.00908665f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_386 N_B1_M1010_g N_VPWR_c_593_n 0.00982266f $X=7.095 $Y=2.4 $X2=0 $Y2=0
cc_387 N_B1_M1016_g N_VPWR_c_593_n 0.00982266f $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_388 N_B1_M1019_g N_VPWR_c_593_n 0.00986405f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_389 N_B1_M1008_g N_A_539_368#_c_702_n 3.62369e-19 $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_390 N_B1_M1008_g N_A_539_368#_c_750_n 0.0197231f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_391 N_B1_M1010_g N_A_539_368#_c_750_n 0.012931f $X=7.095 $Y=2.4 $X2=0 $Y2=0
cc_392 B1 N_A_539_368#_c_750_n 0.0282763f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_393 N_B1_c_470_n N_A_539_368#_c_750_n 4.89356e-19 $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_394 N_B1_M1008_g N_A_539_368#_c_703_n 6.74232e-19 $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_395 N_B1_M1010_g N_A_539_368#_c_703_n 0.0121366f $X=7.095 $Y=2.4 $X2=0 $Y2=0
cc_396 N_B1_M1016_g N_A_539_368#_c_703_n 0.0119382f $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_397 N_B1_M1019_g N_A_539_368#_c_703_n 6.50516e-19 $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_398 N_B1_M1016_g N_A_539_368#_c_758_n 0.012931f $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_399 N_B1_M1019_g N_A_539_368#_c_758_n 0.012931f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_400 B1 N_A_539_368#_c_758_n 0.0391869f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_401 N_B1_c_470_n N_A_539_368#_c_758_n 4.86535e-19 $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_402 N_B1_M1019_g N_A_539_368#_c_704_n 8.84614e-19 $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_403 B1 N_A_539_368#_c_704_n 0.0264312f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_404 N_B1_M1016_g N_A_539_368#_c_705_n 6.50516e-19 $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_405 N_B1_M1019_g N_A_539_368#_c_705_n 0.0121004f $X=7.995 $Y=2.4 $X2=0 $Y2=0
cc_406 N_B1_M1008_g N_A_539_368#_c_707_n 4.63009e-19 $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_407 N_B1_M1010_g N_A_539_368#_c_767_n 8.84614e-19 $X=7.095 $Y=2.4 $X2=0 $Y2=0
cc_408 N_B1_M1016_g N_A_539_368#_c_767_n 8.84614e-19 $X=7.545 $Y=2.4 $X2=0 $Y2=0
cc_409 B1 N_A_539_368#_c_767_n 0.0235495f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_410 N_B1_c_470_n N_A_539_368#_c_767_n 5.51948e-19 $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_411 N_B1_M1000_g N_VGND_c_905_n 0.0100344f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_412 N_B1_M1011_g N_VGND_c_905_n 0.00204878f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_413 N_B1_M1011_g N_VGND_c_906_n 5.20618e-19 $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_414 N_B1_M1025_g N_VGND_c_906_n 0.0101191f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_415 N_B1_M1029_g N_VGND_c_906_n 0.00341128f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_416 N_B1_M1000_g N_VGND_c_913_n 0.00383152f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_417 N_B1_M1011_g N_VGND_c_915_n 0.00434272f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_418 N_B1_M1025_g N_VGND_c_915_n 0.00383152f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_419 N_B1_M1029_g N_VGND_c_917_n 0.00434272f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_420 N_B1_M1000_g N_VGND_c_918_n 0.00757637f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_421 N_B1_M1011_g N_VGND_c_918_n 0.00820284f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_422 N_B1_M1025_g N_VGND_c_918_n 0.0075754f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_423 N_B1_M1029_g N_VGND_c_918_n 0.00824501f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_424 N_B1_M1000_g N_A_914_74#_c_1013_n 0.0174779f $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_425 N_B1_M1011_g N_A_914_74#_c_1013_n 0.0111034f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_426 B1 N_A_914_74#_c_1013_n 0.0282658f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_427 N_B1_c_470_n N_A_914_74#_c_1013_n 0.00236025f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_428 N_B1_M1000_g N_A_914_74#_c_1015_n 6.58468e-19 $X=6.63 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B1_M1011_g N_A_914_74#_c_1015_n 0.00918302f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_430 N_B1_M1025_g N_A_914_74#_c_1015_n 3.97481e-19 $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_431 N_B1_M1025_g N_A_914_74#_c_1016_n 0.0130918f $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_432 N_B1_M1029_g N_A_914_74#_c_1016_n 0.0132972f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_433 B1 N_A_914_74#_c_1016_n 0.0748451f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_434 N_B1_c_470_n N_A_914_74#_c_1016_n 0.00496943f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_435 N_B1_M1025_g N_A_914_74#_c_1017_n 6.56397e-19 $X=7.49 $Y=0.74 $X2=0 $Y2=0
cc_436 N_B1_M1029_g N_A_914_74#_c_1017_n 0.0100626f $X=7.92 $Y=0.74 $X2=0 $Y2=0
cc_437 N_B1_M1011_g N_A_914_74#_c_1018_n 0.00157732f $X=7.06 $Y=0.74 $X2=0 $Y2=0
cc_438 B1 N_A_914_74#_c_1018_n 0.0213626f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_439 N_B1_c_470_n N_A_914_74#_c_1018_n 0.00252677f $X=7.995 $Y=1.515 $X2=0
+ $Y2=0
cc_440 N_A_29_392#_c_562_n N_VPWR_M1020_d 0.00335477f $X=1.905 $Y=2.055
+ $X2=-0.19 $Y2=1.66
cc_441 N_A_29_392#_c_549_n N_VPWR_c_594_n 0.010126f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_442 N_A_29_392#_c_562_n N_VPWR_c_594_n 0.0148589f $X=1.905 $Y=2.055 $X2=0
+ $Y2=0
cc_443 N_A_29_392#_c_553_n N_VPWR_c_594_n 0.0227494f $X=2.07 $Y=2.815 $X2=0
+ $Y2=0
cc_444 N_A_29_392#_c_553_n N_VPWR_c_595_n 0.014549f $X=2.07 $Y=2.815 $X2=0 $Y2=0
cc_445 N_A_29_392#_c_549_n N_VPWR_c_604_n 0.0530426f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_446 N_A_29_392#_c_550_n N_VPWR_c_604_n 0.0235512f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_447 N_A_29_392#_c_549_n N_VPWR_c_593_n 0.0295386f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_448 N_A_29_392#_c_550_n N_VPWR_c_593_n 0.0126924f $X=0.435 $Y=2.99 $X2=0
+ $Y2=0
cc_449 N_A_29_392#_c_553_n N_VPWR_c_593_n 0.0119743f $X=2.07 $Y=2.815 $X2=0
+ $Y2=0
cc_450 N_A_29_392#_c_552_n N_A_539_368#_c_697_n 0.00803119f $X=2.07 $Y=2.14
+ $X2=0 $Y2=0
cc_451 N_A_29_392#_c_553_n N_A_539_368#_c_697_n 0.0340606f $X=2.07 $Y=2.815
+ $X2=0 $Y2=0
cc_452 N_A_29_392#_c_553_n N_A_539_368#_c_699_n 0.00354317f $X=2.07 $Y=2.815
+ $X2=0 $Y2=0
cc_453 N_VPWR_c_595_n N_A_539_368#_c_698_n 0.0357927f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_593_n N_A_539_368#_c_698_n 0.0200586f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_455 N_VPWR_c_595_n N_A_539_368#_c_699_n 0.0235512f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_593_n N_A_539_368#_c_699_n 0.0126924f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_457 N_VPWR_c_595_n N_A_539_368#_c_700_n 0.0592384f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_596_n N_A_539_368#_c_700_n 0.0101219f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_593_n N_A_539_368#_c_700_n 0.0326137f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_460 N_VPWR_M1002_s N_A_539_368#_c_731_n 0.00314376f $X=4.935 $Y=1.84 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_596_n N_A_539_368#_c_731_n 0.0126919f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_596_n N_A_539_368#_c_701_n 0.0233699f $X=5.07 $Y=2.455 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_597_n N_A_539_368#_c_701_n 0.0234083f $X=5.97 $Y=2.455 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_605_n N_A_539_368#_c_701_n 0.0144623f $X=5.885 $Y=3.33 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_593_n N_A_539_368#_c_701_n 0.0118344f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_466 N_VPWR_M1007_s N_A_539_368#_c_739_n 0.00314376f $X=5.835 $Y=1.84 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_597_n N_A_539_368#_c_739_n 0.0148589f $X=5.97 $Y=2.455 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_597_n N_A_539_368#_c_702_n 0.022423f $X=5.97 $Y=2.455 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_598_n N_A_539_368#_c_702_n 0.022423f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_600_n N_A_539_368#_c_702_n 0.00749631f $X=6.705 $Y=3.33 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_593_n N_A_539_368#_c_702_n 0.0062048f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_472 N_VPWR_M1008_d N_A_539_368#_c_750_n 0.00314376f $X=6.735 $Y=1.84 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_598_n N_A_539_368#_c_750_n 0.0148589f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_598_n N_A_539_368#_c_703_n 0.0234083f $X=6.87 $Y=2.455 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_599_n N_A_539_368#_c_703_n 0.0233699f $X=7.77 $Y=2.455 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_602_n N_A_539_368#_c_703_n 0.0144623f $X=7.685 $Y=3.33 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_593_n N_A_539_368#_c_703_n 0.0118344f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_478 N_VPWR_M1016_d N_A_539_368#_c_758_n 0.00314376f $X=7.635 $Y=1.84 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_599_n N_A_539_368#_c_758_n 0.0126919f $X=7.77 $Y=2.455 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_599_n N_A_539_368#_c_705_n 0.0233699f $X=7.77 $Y=2.455 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_606_n N_A_539_368#_c_705_n 0.014549f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_482 N_VPWR_c_593_n N_A_539_368#_c_705_n 0.0119743f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_c_595_n N_A_539_368#_c_706_n 0.0234458f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_593_n N_A_539_368#_c_706_n 0.0125551f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_485 N_A_539_368#_c_698_n N_Y_M1015_d 0.00165831f $X=3.555 $Y=2.99 $X2=0 $Y2=0
cc_486 N_A_539_368#_c_700_n N_Y_M1023_d 0.00165831f $X=4.455 $Y=2.99 $X2=0 $Y2=0
cc_487 N_A_539_368#_c_698_n N_Y_c_872_n 0.0118736f $X=3.555 $Y=2.99 $X2=0 $Y2=0
cc_488 N_A_539_368#_M1021_s N_Y_c_822_n 0.00165831f $X=3.585 $Y=1.84 $X2=0 $Y2=0
cc_489 N_A_539_368#_c_715_n N_Y_c_822_n 0.0170259f $X=3.72 $Y=2.225 $X2=0 $Y2=0
cc_490 N_A_539_368#_c_697_n N_Y_c_823_n 0.00310493f $X=2.82 $Y=1.985 $X2=0 $Y2=0
cc_491 N_A_539_368#_c_700_n N_Y_c_876_n 0.0118736f $X=4.455 $Y=2.99 $X2=0 $Y2=0
cc_492 N_A_539_368#_c_707_n N_A_914_74#_c_1014_n 0.00609927f $X=6.42 $Y=1.985
+ $X2=0 $Y2=0
cc_493 N_Y_c_830_n N_VGND_M1004_d 0.00330219f $X=3.21 $Y=0.875 $X2=0 $Y2=0
cc_494 N_Y_c_816_n N_VGND_M1028_d 0.00668617f $X=3.965 $Y=0.875 $X2=0 $Y2=0
cc_495 N_Y_c_814_n N_VGND_c_901_n 0.0158235f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_496 N_Y_c_814_n N_VGND_c_902_n 0.0104051f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_497 N_Y_c_830_n N_VGND_c_902_n 0.0166744f $X=3.21 $Y=0.875 $X2=0 $Y2=0
cc_498 N_Y_c_815_n N_VGND_c_902_n 0.0103637f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_499 N_Y_c_815_n N_VGND_c_903_n 0.00743725f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_500 N_Y_c_815_n N_VGND_c_904_n 0.0103637f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_501 N_Y_c_816_n N_VGND_c_904_n 0.0214241f $X=3.965 $Y=0.875 $X2=0 $Y2=0
cc_502 N_Y_c_814_n N_VGND_c_911_n 0.0109081f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_503 N_Y_c_814_n N_VGND_c_918_n 0.00901008f $X=2.435 $Y=0.515 $X2=0 $Y2=0
cc_504 N_Y_c_830_n N_VGND_c_918_n 0.0122738f $X=3.21 $Y=0.875 $X2=0 $Y2=0
cc_505 N_Y_c_815_n N_VGND_c_918_n 0.00618197f $X=3.295 $Y=0.515 $X2=0 $Y2=0
cc_506 N_Y_c_816_n N_VGND_c_918_n 0.00943228f $X=3.965 $Y=0.875 $X2=0 $Y2=0
cc_507 N_Y_c_819_n N_VGND_c_918_n 0.0113458f $X=4.96 $Y=0.95 $X2=0 $Y2=0
cc_508 Y N_VGND_c_918_n 0.0119508f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_509 N_Y_c_819_n N_A_914_74#_M1001_s 0.00382948f $X=4.96 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_510 N_Y_c_818_n N_A_914_74#_M1009_s 0.00177442f $X=5.985 $Y=0.95 $X2=0 $Y2=0
cc_511 N_Y_M1001_d N_A_914_74#_c_1011_n 0.00179007f $X=4.985 $Y=0.37 $X2=0 $Y2=0
cc_512 N_Y_M1012_d N_A_914_74#_c_1011_n 0.00179007f $X=5.845 $Y=0.37 $X2=0 $Y2=0
cc_513 N_Y_c_817_n N_A_914_74#_c_1011_n 0.0628697f $X=5.14 $Y=0.95 $X2=0 $Y2=0
cc_514 N_Y_c_819_n N_A_914_74#_c_1011_n 0.0253733f $X=4.96 $Y=0.95 $X2=0 $Y2=0
cc_515 N_Y_c_818_n N_A_914_74#_c_1014_n 0.00561736f $X=5.985 $Y=0.95 $X2=0 $Y2=0
cc_516 N_VGND_c_904_n N_A_914_74#_c_1011_n 0.00868144f $X=3.725 $Y=0.525 $X2=0
+ $Y2=0
cc_517 N_VGND_c_913_n N_A_914_74#_c_1011_n 0.0729484f $X=6.68 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_918_n N_A_914_74#_c_1011_n 0.0614753f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_905_n N_A_914_74#_c_1012_n 0.00947603f $X=6.845 $Y=0.675 $X2=0
+ $Y2=0
cc_520 N_VGND_c_913_n N_A_914_74#_c_1012_n 0.00758556f $X=6.68 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_918_n N_A_914_74#_c_1012_n 0.00627867f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_M1000_s N_A_914_74#_c_1013_n 0.00176461f $X=6.705 $Y=0.37 $X2=0
+ $Y2=0
cc_523 N_VGND_c_905_n N_A_914_74#_c_1013_n 0.0152916f $X=6.845 $Y=0.675 $X2=0
+ $Y2=0
cc_524 N_VGND_c_905_n N_A_914_74#_c_1015_n 0.0175587f $X=6.845 $Y=0.675 $X2=0
+ $Y2=0
cc_525 N_VGND_c_906_n N_A_914_74#_c_1015_n 0.0175587f $X=7.705 $Y=0.675 $X2=0
+ $Y2=0
cc_526 N_VGND_c_915_n N_A_914_74#_c_1015_n 0.0109942f $X=7.54 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_918_n N_A_914_74#_c_1015_n 0.00904371f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_M1025_s N_A_914_74#_c_1016_n 0.00176461f $X=7.565 $Y=0.37 $X2=0
+ $Y2=0
cc_529 N_VGND_c_906_n N_A_914_74#_c_1016_n 0.0152916f $X=7.705 $Y=0.675 $X2=0
+ $Y2=0
cc_530 N_VGND_c_906_n N_A_914_74#_c_1017_n 0.0182902f $X=7.705 $Y=0.675 $X2=0
+ $Y2=0
cc_531 N_VGND_c_917_n N_A_914_74#_c_1017_n 0.0145639f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_918_n N_A_914_74#_c_1017_n 0.0119984f $X=8.4 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfbbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.24000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.460000 1.815000 1.790000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.370000 0.350000 17.705000 1.050000 ;
        RECT 17.395000 1.820000 17.705000 2.980000 ;
        RECT 17.535000 1.050000 17.705000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.280000 0.350000 15.610000 1.220000 ;
        RECT 15.375000 1.220000 15.610000 1.550000 ;
        RECT 15.375000 1.550000 15.715000 1.780000 ;
        RECT 15.375000 1.780000 15.625000 2.980000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.945000 1.505000 14.275000 1.835000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.125000 0.550000 2.135000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.125000 1.315000 1.795000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.524700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.790000 1.450000  9.445000 1.780000 ;
        RECT 11.955000 1.180000 12.325000 1.750000 ;
      LAYER mcon ;
        RECT  9.275000 1.580000  9.445000 1.750000 ;
        RECT 12.155000 1.580000 12.325000 1.750000 ;
      LAYER met1 ;
        RECT  9.215000 1.550000  9.505000 1.595000 ;
        RECT  9.215000 1.595000 12.385000 1.735000 ;
        RECT  9.215000 1.735000  9.505000 1.780000 ;
        RECT 12.095000 1.550000 12.385000 1.595000 ;
        RECT 12.095000 1.735000 12.385000 1.780000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.895000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 18.240000 0.085000 ;
        RECT  0.140000  0.085000  0.470000 0.955000 ;
        RECT  2.180000  0.085000  2.430000 0.950000 ;
        RECT  3.930000  0.085000  4.180000 0.490000 ;
        RECT  5.450000  0.085000  5.720000 0.670000 ;
        RECT  9.055000  0.085000  9.385000 0.940000 ;
        RECT 11.680000  0.085000 12.055000 0.430000 ;
        RECT 14.825000  0.085000 15.110000 1.130000 ;
        RECT 15.780000  0.085000 16.110000 1.130000 ;
        RECT 16.870000  0.085000 17.200000 1.050000 ;
        RECT 17.880000  0.085000 18.130000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
        RECT 16.955000 -0.085000 17.125000 0.085000 ;
        RECT 17.435000 -0.085000 17.605000 0.085000 ;
        RECT 17.915000 -0.085000 18.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 18.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 18.240000 3.415000 ;
        RECT  0.565000 2.645000  0.895000 3.245000 ;
        RECT  2.415000 2.300000  2.745000 3.245000 ;
        RECT  3.875000 2.290000  4.205000 3.245000 ;
        RECT  4.965000 2.350000  5.215000 3.245000 ;
        RECT  8.365000 2.465000  8.695000 3.245000 ;
        RECT  9.465000 2.290000  9.795000 3.245000 ;
        RECT 11.230000 2.600000 11.560000 3.245000 ;
        RECT 12.305000 2.600000 12.635000 3.245000 ;
        RECT 14.280000 2.845000 15.170000 3.245000 ;
        RECT 14.825000 1.950000 15.170000 2.845000 ;
        RECT 15.825000 1.950000 16.155000 3.245000 ;
        RECT 16.895000 1.820000 17.225000 3.245000 ;
        RECT 17.875000 1.820000 18.125000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
        RECT 16.475000 3.245000 16.645000 3.415000 ;
        RECT 16.955000 3.245000 17.125000 3.415000 ;
        RECT 17.435000 3.245000 17.605000 3.415000 ;
        RECT 17.915000 3.245000 18.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 18.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 2.305000  1.235000 2.475000 ;
      RECT  0.115000 2.475000  0.365000 2.980000 ;
      RECT  0.960000 0.625000  1.690000 0.955000 ;
      RECT  1.065000 2.475000  1.235000 2.905000 ;
      RECT  1.065000 2.905000  2.185000 3.075000 ;
      RECT  1.405000 2.300000  1.655000 2.735000 ;
      RECT  1.485000 0.955000  1.690000 1.120000 ;
      RECT  1.485000 1.120000  2.770000 1.290000 ;
      RECT  1.485000 1.960000  2.155000 2.130000 ;
      RECT  1.485000 2.130000  1.655000 2.300000 ;
      RECT  1.855000 2.300000  2.185000 2.905000 ;
      RECT  1.985000 1.290000  2.155000 1.960000 ;
      RECT  2.600000 0.255000  3.535000 0.425000 ;
      RECT  2.600000 0.425000  2.770000 1.120000 ;
      RECT  2.605000 1.480000  3.195000 1.810000 ;
      RECT  2.940000 0.595000  3.195000 1.480000 ;
      RECT  2.945000 1.810000  3.195000 2.980000 ;
      RECT  3.365000 0.425000  3.535000 0.660000 ;
      RECT  3.365000 0.660000  4.520000 0.830000 ;
      RECT  3.420000 1.000000  4.235000 1.170000 ;
      RECT  3.425000 1.950000  4.235000 2.120000 ;
      RECT  3.425000 2.120000  3.675000 2.980000 ;
      RECT  4.065000 1.170000  4.235000 1.340000 ;
      RECT  4.065000 1.340000  4.445000 1.670000 ;
      RECT  4.065000 1.670000  4.235000 1.950000 ;
      RECT  4.350000 0.255000  5.280000 0.425000 ;
      RECT  4.350000 0.425000  4.520000 0.660000 ;
      RECT  4.405000 1.840000  4.785000 2.980000 ;
      RECT  4.615000 1.180000  6.115000 1.350000 ;
      RECT  4.615000 1.350000  4.785000 1.840000 ;
      RECT  4.690000 0.595000  4.940000 1.180000 ;
      RECT  5.035000 1.830000  5.365000 2.010000 ;
      RECT  5.035000 2.010000  5.555000 2.180000 ;
      RECT  5.110000 0.425000  5.280000 0.840000 ;
      RECT  5.110000 0.840000  6.115000 1.010000 ;
      RECT  5.385000 2.180000  5.555000 2.905000 ;
      RECT  5.385000 2.905000  7.825000 3.075000 ;
      RECT  5.595000 1.350000  6.115000 1.525000 ;
      RECT  5.595000 1.525000  6.825000 1.840000 ;
      RECT  5.840000 2.040000  7.365000 2.210000 ;
      RECT  5.840000 2.210000  6.170000 2.735000 ;
      RECT  5.945000 0.265000  7.115000 0.435000 ;
      RECT  5.945000 0.435000  6.115000 0.840000 ;
      RECT  6.285000 0.605000  6.615000 1.185000 ;
      RECT  6.285000 1.185000  7.365000 1.355000 ;
      RECT  6.340000 2.380000  7.705000 2.550000 ;
      RECT  6.340000 2.550000  6.670000 2.735000 ;
      RECT  6.495000 1.840000  6.825000 1.855000 ;
      RECT  6.785000 0.435000  7.115000 0.845000 ;
      RECT  6.785000 0.845000  7.705000 1.015000 ;
      RECT  6.900000 2.730000  8.045000 2.900000 ;
      RECT  6.900000 2.900000  7.825000 2.905000 ;
      RECT  7.035000 1.355000  7.365000 2.040000 ;
      RECT  7.345000 0.265000  8.620000 0.435000 ;
      RECT  7.345000 0.435000  7.770000 0.675000 ;
      RECT  7.535000 1.015000  7.705000 2.380000 ;
      RECT  7.875000 0.945000  8.280000 1.115000 ;
      RECT  7.875000 1.115000  8.045000 2.125000 ;
      RECT  7.875000 2.125000  9.235000 2.295000 ;
      RECT  7.875000 2.295000  8.045000 2.730000 ;
      RECT  7.950000 0.605000  8.280000 0.945000 ;
      RECT  8.215000 1.285000  8.620000 1.955000 ;
      RECT  8.450000 0.435000  8.620000 0.605000 ;
      RECT  8.450000 0.605000  8.885000 0.935000 ;
      RECT  8.450000 1.110000  9.725000 1.280000 ;
      RECT  8.450000 1.280000  8.620000 1.285000 ;
      RECT  8.905000 1.950000  9.945000 2.120000 ;
      RECT  8.905000 2.120000  9.235000 2.125000 ;
      RECT  8.905000 2.295000  9.235000 2.980000 ;
      RECT  9.555000 0.260000 11.510000 0.430000 ;
      RECT  9.555000 0.430000  9.725000 1.110000 ;
      RECT  9.615000 1.580000  9.945000 1.950000 ;
      RECT  9.960000 0.600000 11.110000 0.850000 ;
      RECT 10.155000 1.180000 10.485000 1.280000 ;
      RECT 10.155000 1.280000 11.385000 1.580000 ;
      RECT 10.155000 1.580000 10.485000 1.755000 ;
      RECT 10.305000 2.100000 10.910000 2.270000 ;
      RECT 10.305000 2.270000 10.635000 2.980000 ;
      RECT 10.740000 1.750000 11.750000 1.920000 ;
      RECT 10.740000 1.920000 10.910000 2.100000 ;
      RECT 10.940000 0.850000 11.110000 0.940000 ;
      RECT 10.940000 0.940000 11.725000 1.110000 ;
      RECT 11.080000 2.090000 11.410000 2.260000 ;
      RECT 11.080000 2.260000 13.435000 2.430000 ;
      RECT 11.340000 0.430000 11.510000 0.600000 ;
      RECT 11.340000 0.600000 12.065000 0.770000 ;
      RECT 11.555000 1.110000 11.725000 1.750000 ;
      RECT 11.580000 1.920000 12.665000 2.090000 ;
      RECT 11.805000 2.430000 12.135000 2.980000 ;
      RECT 11.895000 0.770000 12.665000 0.940000 ;
      RECT 12.235000 0.255000 13.595000 0.425000 ;
      RECT 12.235000 0.425000 12.655000 0.600000 ;
      RECT 12.495000 0.940000 12.665000 1.130000 ;
      RECT 12.495000 1.130000 14.150000 1.300000 ;
      RECT 12.495000 1.300000 12.825000 1.550000 ;
      RECT 12.495000 1.720000 13.365000 1.890000 ;
      RECT 12.495000 1.890000 12.665000 1.920000 ;
      RECT 12.835000 0.595000 13.085000 0.665000 ;
      RECT 12.835000 0.665000 14.490000 0.835000 ;
      RECT 12.835000 0.835000 13.085000 0.960000 ;
      RECT 13.035000 1.470000 13.365000 1.720000 ;
      RECT 13.185000 2.060000 13.435000 2.260000 ;
      RECT 13.185000 2.430000 13.435000 2.505000 ;
      RECT 13.185000 2.505000 14.655000 2.675000 ;
      RECT 13.185000 2.675000 13.435000 2.980000 ;
      RECT 13.265000 0.425000 13.595000 0.495000 ;
      RECT 13.605000 1.005000 14.150000 1.130000 ;
      RECT 13.605000 1.300000 14.150000 1.335000 ;
      RECT 13.605000 1.335000 13.775000 2.005000 ;
      RECT 13.605000 2.005000 14.075000 2.335000 ;
      RECT 14.320000 0.835000 14.655000 1.005000 ;
      RECT 14.485000 1.005000 14.655000 1.430000 ;
      RECT 14.485000 1.430000 14.815000 1.760000 ;
      RECT 14.485000 1.760000 14.655000 2.505000 ;
      RECT 16.340000 0.540000 16.670000 1.220000 ;
      RECT 16.340000 1.220000 17.365000 1.550000 ;
      RECT 16.340000 1.550000 16.700000 2.940000 ;
    LAYER mcon ;
      RECT  5.915000 1.210000  6.085000 1.380000 ;
      RECT 10.235000 1.210000 10.405000 1.380000 ;
    LAYER met1 ;
      RECT  5.855000 1.180000  6.145000 1.225000 ;
      RECT  5.855000 1.225000 10.465000 1.365000 ;
      RECT  5.855000 1.365000  6.145000 1.410000 ;
      RECT 10.175000 1.180000 10.465000 1.225000 ;
      RECT 10.175000 1.365000 10.465000 1.410000 ;
  END
END sky130_fd_sc_ms__sdfbbn_2

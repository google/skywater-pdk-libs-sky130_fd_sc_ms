* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
X0 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X1 VPWR B_N a_354_252# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VPWR a_225_82# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 VPWR a_27_74# a_225_82# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_225_82# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 a_498_82# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND B_N a_354_252# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X7 a_390_82# C a_498_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 X a_225_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VPWR C a_225_82# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X10 VGND a_225_82# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_312_82# a_354_252# a_390_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_225_82# a_354_252# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 a_225_82# a_27_74# a_312_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X15 X a_225_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__dfxtp_2.pxi.spice
* Created: Fri Aug 28 17:25:17 2020
* 
x_PM_SKY130_FD_SC_MS__DFXTP_2%CLK N_CLK_M1010_g N_CLK_M1024_g CLK N_CLK_c_192_n
+ N_CLK_c_193_n PM_SKY130_FD_SC_MS__DFXTP_2%CLK
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_27_74# N_A_27_74#_M1024_s N_A_27_74#_M1010_s
+ N_A_27_74#_M1011_g N_A_27_74#_M1025_g N_A_27_74#_M1016_g N_A_27_74#_M1022_g
+ N_A_27_74#_M1018_g N_A_27_74#_c_255_n N_A_27_74#_c_256_n N_A_27_74#_M1017_g
+ N_A_27_74#_c_228_n N_A_27_74#_c_258_n N_A_27_74#_c_259_n N_A_27_74#_c_229_n
+ N_A_27_74#_c_230_n N_A_27_74#_c_274_n N_A_27_74#_c_231_n N_A_27_74#_c_232_n
+ N_A_27_74#_c_233_n N_A_27_74#_c_234_n N_A_27_74#_c_235_n N_A_27_74#_c_236_n
+ N_A_27_74#_c_237_n N_A_27_74#_c_238_n N_A_27_74#_c_239_n N_A_27_74#_c_240_n
+ N_A_27_74#_c_241_n N_A_27_74#_c_242_n N_A_27_74#_c_361_p N_A_27_74#_c_362_p
+ N_A_27_74#_c_243_n N_A_27_74#_c_244_n N_A_27_74#_c_321_p N_A_27_74#_c_245_n
+ N_A_27_74#_c_246_n N_A_27_74#_c_247_n N_A_27_74#_c_248_n N_A_27_74#_c_249_n
+ N_A_27_74#_c_250_n N_A_27_74#_c_262_n PM_SKY130_FD_SC_MS__DFXTP_2%A_27_74#
x_PM_SKY130_FD_SC_MS__DFXTP_2%D N_D_M1007_g N_D_c_488_n N_D_M1013_g N_D_c_494_n
+ N_D_c_490_n D N_D_c_496_n N_D_c_492_n PM_SKY130_FD_SC_MS__DFXTP_2%D
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_209_368# N_A_209_368#_M1025_d
+ N_A_209_368#_M1011_d N_A_209_368#_c_550_n N_A_209_368#_c_551_n
+ N_A_209_368#_c_561_n N_A_209_368#_M1012_g N_A_209_368#_M1015_g
+ N_A_209_368#_M1009_g N_A_209_368#_M1023_g N_A_209_368#_c_564_n
+ N_A_209_368#_c_565_n N_A_209_368#_c_554_n N_A_209_368#_c_566_n
+ N_A_209_368#_c_567_n N_A_209_368#_c_605_n N_A_209_368#_c_555_n
+ N_A_209_368#_c_556_n N_A_209_368#_c_569_n N_A_209_368#_c_570_n
+ N_A_209_368#_c_571_n N_A_209_368#_c_557_n N_A_209_368#_c_558_n
+ N_A_209_368#_c_655_n N_A_209_368#_c_623_n N_A_209_368#_c_559_n
+ N_A_209_368#_c_574_n N_A_209_368#_c_560_n
+ PM_SKY130_FD_SC_MS__DFXTP_2%A_209_368#
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_695_459# N_A_695_459#_M1003_d
+ N_A_695_459#_M1004_d N_A_695_459#_c_779_n N_A_695_459#_M1002_g
+ N_A_695_459#_c_773_n N_A_695_459#_M1000_g N_A_695_459#_c_781_n
+ N_A_695_459#_c_775_n N_A_695_459#_c_776_n N_A_695_459#_c_777_n
+ N_A_695_459#_c_803_n N_A_695_459#_c_778_n
+ PM_SKY130_FD_SC_MS__DFXTP_2%A_695_459#
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_541_429# N_A_541_429#_M1016_d
+ N_A_541_429#_M1012_d N_A_541_429#_M1004_g N_A_541_429#_c_858_n
+ N_A_541_429#_c_859_n N_A_541_429#_M1003_g N_A_541_429#_c_860_n
+ N_A_541_429#_c_868_n N_A_541_429#_c_861_n N_A_541_429#_c_869_n
+ N_A_541_429#_c_870_n N_A_541_429#_c_862_n N_A_541_429#_c_863_n
+ N_A_541_429#_c_864_n N_A_541_429#_c_865_n N_A_541_429#_c_866_n
+ PM_SKY130_FD_SC_MS__DFXTP_2%A_541_429#
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_1217_314# N_A_1217_314#_M1020_s
+ N_A_1217_314#_M1019_s N_A_1217_314#_M1006_g N_A_1217_314#_M1001_g
+ N_A_1217_314#_M1008_g N_A_1217_314#_M1005_g N_A_1217_314#_c_973_n
+ N_A_1217_314#_M1014_g N_A_1217_314#_M1021_g N_A_1217_314#_c_974_n
+ N_A_1217_314#_c_975_n N_A_1217_314#_c_976_n N_A_1217_314#_c_963_n
+ N_A_1217_314#_c_977_n N_A_1217_314#_c_978_n N_A_1217_314#_c_964_n
+ N_A_1217_314#_c_965_n N_A_1217_314#_c_966_n N_A_1217_314#_c_967_n
+ N_A_1217_314#_c_981_n N_A_1217_314#_c_968_n N_A_1217_314#_c_969_n
+ N_A_1217_314#_c_970_n PM_SKY130_FD_SC_MS__DFXTP_2%A_1217_314#
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_1022_424# N_A_1022_424#_M1009_d
+ N_A_1022_424#_M1018_d N_A_1022_424#_M1020_g N_A_1022_424#_M1019_g
+ N_A_1022_424#_c_1103_n N_A_1022_424#_c_1095_n N_A_1022_424#_c_1104_n
+ N_A_1022_424#_c_1105_n N_A_1022_424#_c_1096_n N_A_1022_424#_c_1097_n
+ N_A_1022_424#_c_1098_n N_A_1022_424#_c_1099_n N_A_1022_424#_c_1100_n
+ N_A_1022_424#_c_1101_n PM_SKY130_FD_SC_MS__DFXTP_2%A_1022_424#
x_PM_SKY130_FD_SC_MS__DFXTP_2%VPWR N_VPWR_M1010_d N_VPWR_M1007_s N_VPWR_M1002_d
+ N_VPWR_M1006_d N_VPWR_M1019_d N_VPWR_M1014_s N_VPWR_c_1196_n N_VPWR_c_1197_n
+ N_VPWR_c_1198_n N_VPWR_c_1199_n N_VPWR_c_1200_n VPWR N_VPWR_c_1201_n
+ N_VPWR_c_1202_n N_VPWR_c_1203_n N_VPWR_c_1204_n N_VPWR_c_1205_n
+ N_VPWR_c_1206_n N_VPWR_c_1207_n N_VPWR_c_1208_n N_VPWR_c_1209_n
+ N_VPWR_c_1210_n N_VPWR_c_1195_n PM_SKY130_FD_SC_MS__DFXTP_2%VPWR
x_PM_SKY130_FD_SC_MS__DFXTP_2%A_434_508# N_A_434_508#_M1013_d
+ N_A_434_508#_M1007_d N_A_434_508#_c_1302_n N_A_434_508#_c_1298_n
+ N_A_434_508#_c_1299_n N_A_434_508#_c_1300_n N_A_434_508#_c_1301_n
+ PM_SKY130_FD_SC_MS__DFXTP_2%A_434_508#
x_PM_SKY130_FD_SC_MS__DFXTP_2%Q N_Q_M1005_d N_Q_M1008_d N_Q_c_1346_n
+ N_Q_c_1354_n N_Q_c_1347_n N_Q_c_1348_n Q Q PM_SKY130_FD_SC_MS__DFXTP_2%Q
x_PM_SKY130_FD_SC_MS__DFXTP_2%VGND N_VGND_M1024_d N_VGND_M1013_s N_VGND_M1000_d
+ N_VGND_M1001_d N_VGND_M1020_d N_VGND_M1021_s N_VGND_c_1381_n N_VGND_c_1382_n
+ N_VGND_c_1383_n N_VGND_c_1384_n N_VGND_c_1385_n N_VGND_c_1386_n
+ N_VGND_c_1387_n N_VGND_c_1388_n N_VGND_c_1389_n VGND N_VGND_c_1390_n
+ N_VGND_c_1391_n N_VGND_c_1392_n N_VGND_c_1393_n N_VGND_c_1394_n
+ N_VGND_c_1395_n N_VGND_c_1396_n N_VGND_c_1397_n N_VGND_c_1398_n
+ N_VGND_c_1399_n PM_SKY130_FD_SC_MS__DFXTP_2%VGND
cc_1 VNB N_CLK_M1010_g 0.00192268f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_CLK_M1024_g 0.0303396f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_CLK_c_192_n 0.0163904f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_4 VNB N_CLK_c_193_n 0.0443414f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_5 VNB N_A_27_74#_M1011_g 0.00647031f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_74#_M1016_g 0.0498677f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_7 VNB N_A_27_74#_M1017_g 0.0382294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_228_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_229_n 0.0033521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_230_n 0.00891132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_231_n 0.00152612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_232_n 0.00775643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_233_n 0.0011177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_234_n 0.00348411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_235_n 0.00379259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_236_n 0.00224001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_237_n 0.00260191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_238_n 0.023115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_239_n 0.00163434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_240_n 0.00414722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_241_n 0.00129964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_242_n 0.00602315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_243_n 0.00251728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_244_n 0.00493702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_245_n 0.0334425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_246_n 0.0106563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_247_n 0.00404212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_248_n 0.0439085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_249_n 0.00605351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_250_n 0.0185348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_D_c_488_n 0.0160594f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_32 VNB N_D_M1013_g 0.0215042f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_D_c_490_n 0.00385947f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_34 VNB D 0.00368502f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_35 VNB N_D_c_492_n 0.0335085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_209_368#_c_550_n 0.126381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_A_209_368#_c_551_n 0.0124432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_209_368#_M1015_g 0.0281484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_209_368#_M1009_g 0.0246451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_209_368#_c_554_n 0.00373775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_209_368#_c_555_n 0.0131386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_209_368#_c_556_n 0.00259833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_209_368#_c_557_n 0.00731562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_209_368#_c_558_n 0.0270896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_209_368#_c_559_n 0.0344424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_209_368#_c_560_n 0.072622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_695_459#_c_773_n 0.0173655f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_48 VNB N_A_695_459#_M1000_g 0.0223643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_695_459#_c_775_n 0.00732475f $X=-0.19 $Y=-0.245 $X2=0.315
+ $Y2=1.665
cc_50 VNB N_A_695_459#_c_776_n 0.0134569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_695_459#_c_777_n 0.00513473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_695_459#_c_778_n 0.0557929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_541_429#_c_858_n 0.0253879f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_54 VNB N_A_541_429#_c_859_n 0.0170631f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_55 VNB N_A_541_429#_c_860_n 0.0163795f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_56 VNB N_A_541_429#_c_861_n 0.00432593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_541_429#_c_862_n 3.65459e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_541_429#_c_863_n 0.00705628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_541_429#_c_864_n 0.00228206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_541_429#_c_865_n 7.77907e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_541_429#_c_866_n 0.0133345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1217_314#_M1001_g 0.0468977f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_63 VNB N_A_1217_314#_M1005_g 0.0253468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1217_314#_M1021_g 0.0298331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1217_314#_c_963_n 0.0074104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1217_314#_c_964_n 0.00209332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1217_314#_c_965_n 0.00419184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1217_314#_c_966_n 0.00382769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1217_314#_c_967_n 0.0113781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1217_314#_c_968_n 0.00427438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1217_314#_c_969_n 0.00389508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1217_314#_c_970_n 0.0517972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1022_424#_M1020_g 0.0337753f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_74 VNB N_A_1022_424#_M1019_g 0.0100556f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.465
cc_75 VNB N_A_1022_424#_c_1095_n 0.00297687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1022_424#_c_1096_n 0.0017128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1022_424#_c_1097_n 0.0029215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1022_424#_c_1098_n 0.00104193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1022_424#_c_1099_n 0.00251939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1022_424#_c_1100_n 0.0361184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1022_424#_c_1101_n 0.0360683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VPWR_c_1195_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_434_508#_c_1298_n 0.00361891f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.465
cc_84 VNB N_A_434_508#_c_1299_n 0.00583226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_434_508#_c_1300_n 0.00232296f $X=-0.19 $Y=-0.245 $X2=0.315
+ $Y2=1.465
cc_86 VNB N_A_434_508#_c_1301_n 0.0085391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_Q_c_1346_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_88 VNB N_Q_c_1347_n 0.00127979f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_89 VNB N_Q_c_1348_n 0.00431429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1381_n 0.00529583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1382_n 0.00186565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1383_n 0.00684753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1384_n 0.0207706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1385_n 0.00937879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1386_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1387_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1388_n 0.0481606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1389_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1390_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1391_n 0.0284905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1392_n 0.0420639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1393_n 0.0210814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1394_n 0.0189349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1395_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1396_n 0.0025968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1397_n 0.00477982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1398_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1399_n 0.465903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VPB N_CLK_M1010_g 0.0298346f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_110 VPB N_CLK_c_192_n 0.00724255f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_111 VPB N_A_27_74#_M1011_g 0.0246707f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_112 VPB N_A_27_74#_M1016_g 0.00570065f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_113 VPB N_A_27_74#_M1022_g 0.0405724f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.665
cc_114 VPB N_A_27_74#_M1018_g 0.0301532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_74#_c_255_n 0.0466875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_74#_c_256_n 0.00908301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_74#_M1017_g 0.00178083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_74#_c_258_n 0.00758177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_74#_c_259_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_74#_c_231_n 0.00280413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_74#_c_240_n 0.0051246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_27_74#_c_262_n 0.0499872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_D_M1007_g 0.0288157f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_124 VPB N_D_c_494_n 0.00452018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_D_c_490_n 0.00477519f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_126 VPB N_D_c_496_n 0.045863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_209_368#_c_561_n 0.0553613f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_128 VPB N_A_209_368#_M1012_g 0.0320917f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_129 VPB N_A_209_368#_M1023_g 0.0226161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_209_368#_c_564_n 0.00803473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_209_368#_c_565_n 0.0106254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_209_368#_c_566_n 0.00608915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_209_368#_c_567_n 0.0109001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_209_368#_c_556_n 0.00341831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_209_368#_c_569_n 0.00537328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_209_368#_c_570_n 0.00428999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_209_368#_c_571_n 0.0390344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_209_368#_c_557_n 0.00877102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_209_368#_c_558_n 0.0260233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_209_368#_c_574_n 0.00224892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_695_459#_c_779_n 0.0175438f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_142 VPB N_A_695_459#_c_773_n 0.0344838f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_143 VPB N_A_695_459#_c_781_n 0.0202505f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.465
cc_144 VPB N_A_695_459#_c_777_n 0.00426196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_541_429#_M1004_g 0.0266437f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_146 VPB N_A_541_429#_c_868_n 0.0143735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_541_429#_c_869_n 0.00276587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_541_429#_c_870_n 0.00215598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_541_429#_c_862_n 0.0049133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_541_429#_c_865_n 0.00263638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_541_429#_c_866_n 0.038003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_1217_314#_M1006_g 0.0358383f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_153 VPB N_A_1217_314#_M1008_g 0.0216333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_1217_314#_c_973_n 0.0185413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_1217_314#_c_974_n 0.0326692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_1217_314#_c_975_n 0.0178663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_1217_314#_c_976_n 0.0155356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_1217_314#_c_977_n 0.0129456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_1217_314#_c_978_n 0.00293966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_1217_314#_c_966_n 0.00383426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_1217_314#_c_967_n 0.00520037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_1217_314#_c_981_n 0.0028231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_1217_314#_c_968_n 6.07799e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_1217_314#_c_970_n 0.0161311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_1022_424#_M1019_g 0.0237197f $X=-0.19 $Y=1.66 $X2=0.34 $Y2=1.465
cc_166 VPB N_A_1022_424#_c_1103_n 0.00821908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_1022_424#_c_1104_n 0.00685687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1022_424#_c_1105_n 2.35947e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_1022_424#_c_1097_n 4.74396e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1196_n 0.00797161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1197_n 0.014602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1198_n 0.0083809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1199_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1200_n 0.0644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1201_n 0.0203276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1202_n 0.0445709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1203_n 0.0535792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1204_n 0.0198858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1205_n 0.0195742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1206_n 0.0233502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1207_n 0.0151137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1208_n 0.0157363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1209_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1210_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1195_n 0.11158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_434_508#_c_1302_n 0.00543574f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_187 VPB N_A_434_508#_c_1300_n 4.75261e-19 $X=-0.19 $Y=1.66 $X2=0.315
+ $Y2=1.465
cc_188 VPB N_Q_c_1347_n 9.57035e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_189 VPB Q 0.00231613f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.465
cc_190 N_CLK_c_193_n N_A_27_74#_M1011_g 0.0336655f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_191 N_CLK_M1024_g N_A_27_74#_c_228_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_192 N_CLK_M1010_g N_A_27_74#_c_258_n 8.8334e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_193 N_CLK_c_192_n N_A_27_74#_c_258_n 0.0257548f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_194 N_CLK_c_193_n N_A_27_74#_c_258_n 0.0011953f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_195 N_CLK_M1010_g N_A_27_74#_c_259_n 0.0121004f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_196 N_CLK_M1024_g N_A_27_74#_c_229_n 0.0142287f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_197 N_CLK_c_192_n N_A_27_74#_c_229_n 0.010454f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_198 N_CLK_c_193_n N_A_27_74#_c_229_n 0.00142272f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_199 N_CLK_c_192_n N_A_27_74#_c_230_n 0.0209983f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_200 N_CLK_c_193_n N_A_27_74#_c_230_n 0.0015038f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_201 N_CLK_M1010_g N_A_27_74#_c_274_n 0.0152912f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_202 N_CLK_c_192_n N_A_27_74#_c_274_n 0.00433199f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_203 N_CLK_M1010_g N_A_27_74#_c_231_n 0.00365954f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_204 N_CLK_M1024_g N_A_27_74#_c_233_n 3.10948e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_205 N_CLK_M1024_g N_A_27_74#_c_244_n 0.00510574f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_206 N_CLK_c_192_n N_A_27_74#_c_244_n 0.0379192f $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_207 N_CLK_c_193_n N_A_27_74#_c_244_n 0.00365954f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_208 N_CLK_M1024_g N_A_27_74#_c_245_n 0.00404161f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_CLK_c_192_n N_A_27_74#_c_245_n 2.11025e-19 $X=0.34 $Y=1.465 $X2=0 $Y2=0
cc_210 N_CLK_c_193_n N_A_27_74#_c_245_n 0.0157402f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_211 N_CLK_M1024_g N_A_27_74#_c_250_n 0.0182143f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_212 N_CLK_M1010_g N_A_209_368#_c_565_n 6.54737e-19 $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_213 N_CLK_M1010_g N_VPWR_c_1196_n 0.0027763f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_214 N_CLK_M1010_g N_VPWR_c_1206_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_215 N_CLK_M1010_g N_VPWR_c_1195_n 0.00986118f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_216 N_CLK_M1024_g N_VGND_c_1381_n 0.0121339f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_217 N_CLK_M1024_g N_VGND_c_1390_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_218 N_CLK_M1024_g N_VGND_c_1399_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_27_74#_c_235_n N_D_c_488_n 0.00303023f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_220 N_A_27_74#_M1016_g N_D_M1013_g 0.0177252f $X=2.99 $Y=0.805 $X2=0 $Y2=0
cc_221 N_A_27_74#_c_234_n N_D_M1013_g 8.9778e-19 $X=1.73 $Y=0.81 $X2=0 $Y2=0
cc_222 N_A_27_74#_c_235_n N_D_M1013_g 0.0064381f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_237_n N_D_M1013_g 0.0108239f $X=2.435 $Y=0.81 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_238_n N_D_M1013_g 0.00283033f $X=3.585 $Y=0.34 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_235_n D 0.0293231f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_226 N_A_27_74#_M1011_g N_D_c_496_n 0.00196772f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_27_74#_M1016_g N_D_c_492_n 0.00227704f $X=2.99 $Y=0.805 $X2=0 $Y2=0
cc_228 N_A_27_74#_c_235_n N_D_c_492_n 0.00812532f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_232_n N_A_209_368#_M1025_d 0.00777821f $X=1.645 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_230 N_A_27_74#_M1016_g N_A_209_368#_c_550_n 0.00882199f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_231 N_A_27_74#_c_232_n N_A_209_368#_c_550_n 4.6256e-19 $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_232 N_A_27_74#_c_235_n N_A_209_368#_c_550_n 0.00764044f $X=2.35 $Y=0.895
+ $X2=0 $Y2=0
cc_233 N_A_27_74#_c_238_n N_A_209_368#_c_550_n 0.013889f $X=3.585 $Y=0.34 $X2=0
+ $Y2=0
cc_234 N_A_27_74#_c_239_n N_A_209_368#_c_550_n 0.0036181f $X=2.52 $Y=0.34 $X2=0
+ $Y2=0
cc_235 N_A_27_74#_c_232_n N_A_209_368#_c_551_n 9.85082e-19 $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_236 N_A_27_74#_c_250_n N_A_209_368#_c_551_n 0.010763f $X=0.982 $Y=1.22 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_M1016_g N_A_209_368#_c_561_n 0.00681571f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_238 N_A_27_74#_c_262_n N_A_209_368#_M1012_g 0.0248293f $X=3.145 $Y=1.92 $X2=0
+ $Y2=0
cc_239 N_A_27_74#_M1016_g N_A_209_368#_M1015_g 0.00842f $X=2.99 $Y=0.805 $X2=0
+ $Y2=0
cc_240 N_A_27_74#_c_238_n N_A_209_368#_M1015_g 0.0160142f $X=3.585 $Y=0.34 $X2=0
+ $Y2=0
cc_241 N_A_27_74#_c_241_n N_A_209_368#_M1015_g 0.00254317f $X=3.67 $Y=0.69 $X2=0
+ $Y2=0
cc_242 N_A_27_74#_c_242_n N_A_209_368#_M1015_g 0.00144191f $X=3.67 $Y=1.285
+ $X2=0 $Y2=0
cc_243 N_A_27_74#_c_246_n N_A_209_368#_M1015_g 0.00444424f $X=3.67 $Y=1.37 $X2=0
+ $Y2=0
cc_244 N_A_27_74#_c_262_n N_A_209_368#_M1015_g 8.37484e-19 $X=3.145 $Y=1.92
+ $X2=0 $Y2=0
cc_245 N_A_27_74#_M1017_g N_A_209_368#_M1009_g 0.012644f $X=5.785 $Y=0.83 $X2=0
+ $Y2=0
cc_246 N_A_27_74#_c_247_n N_A_209_368#_M1009_g 4.97101e-19 $X=5.725 $Y=0.345
+ $X2=0 $Y2=0
cc_247 N_A_27_74#_c_248_n N_A_209_368#_M1009_g 0.00853016f $X=5.725 $Y=0.345
+ $X2=0 $Y2=0
cc_248 N_A_27_74#_c_249_n N_A_209_368#_M1009_g 0.0133151f $X=5.56 $Y=0.382 $X2=0
+ $Y2=0
cc_249 N_A_27_74#_M1011_g N_A_209_368#_c_564_n 0.00483141f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_250 N_A_27_74#_M1011_g N_A_209_368#_c_565_n 0.0101098f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_251 N_A_27_74#_c_259_n N_A_209_368#_c_565_n 0.00481756f $X=0.28 $Y=2.815
+ $X2=0 $Y2=0
cc_252 N_A_27_74#_c_232_n N_A_209_368#_c_554_n 0.012787f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_253 N_A_27_74#_c_234_n N_A_209_368#_c_554_n 0.0150602f $X=1.73 $Y=0.81 $X2=0
+ $Y2=0
cc_254 N_A_27_74#_c_236_n N_A_209_368#_c_554_n 0.0133618f $X=1.815 $Y=0.895
+ $X2=0 $Y2=0
cc_255 N_A_27_74#_c_321_p N_A_209_368#_c_554_n 0.055389f $X=0.905 $Y=0.96 $X2=0
+ $Y2=0
cc_256 N_A_27_74#_c_250_n N_A_209_368#_c_554_n 0.00587111f $X=0.982 $Y=1.22
+ $X2=0 $Y2=0
cc_257 N_A_27_74#_M1022_g N_A_209_368#_c_567_n 0.0136395f $X=3.145 $Y=2.73 $X2=0
+ $Y2=0
cc_258 N_A_27_74#_M1018_g N_A_209_368#_c_605_n 4.19897e-19 $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_259 N_A_27_74#_c_256_n N_A_209_368#_c_555_n 0.00653142f $X=5.11 $Y=1.765
+ $X2=0 $Y2=0
cc_260 N_A_27_74#_M1017_g N_A_209_368#_c_555_n 6.96097e-19 $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_261 N_A_27_74#_M1018_g N_A_209_368#_c_556_n 0.0192626f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_262 N_A_27_74#_c_256_n N_A_209_368#_c_556_n 0.00529862f $X=5.11 $Y=1.765
+ $X2=0 $Y2=0
cc_263 N_A_27_74#_M1018_g N_A_209_368#_c_569_n 0.0106719f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_264 N_A_27_74#_M1018_g N_A_209_368#_c_570_n 7.9432e-19 $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_265 N_A_27_74#_c_255_n N_A_209_368#_c_570_n 7.71704e-19 $X=5.71 $Y=1.765
+ $X2=0 $Y2=0
cc_266 N_A_27_74#_M1018_g N_A_209_368#_c_571_n 0.0251524f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_267 N_A_27_74#_c_255_n N_A_209_368#_c_571_n 0.0262f $X=5.71 $Y=1.765 $X2=0
+ $Y2=0
cc_268 N_A_27_74#_M1011_g N_A_209_368#_c_557_n 0.00625126f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_269 N_A_27_74#_c_231_n N_A_209_368#_c_557_n 0.0204706f $X=0.76 $Y=1.95 $X2=0
+ $Y2=0
cc_270 N_A_27_74#_c_236_n N_A_209_368#_c_557_n 0.00301676f $X=1.815 $Y=0.895
+ $X2=0 $Y2=0
cc_271 N_A_27_74#_c_244_n N_A_209_368#_c_557_n 0.0270502f $X=0.905 $Y=1.045
+ $X2=0 $Y2=0
cc_272 N_A_27_74#_c_245_n N_A_209_368#_c_557_n 0.00326249f $X=0.97 $Y=1.385
+ $X2=0 $Y2=0
cc_273 N_A_27_74#_M1011_g N_A_209_368#_c_558_n 0.00914883f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_274 N_A_27_74#_c_244_n N_A_209_368#_c_558_n 2.01719e-19 $X=0.905 $Y=1.045
+ $X2=0 $Y2=0
cc_275 N_A_27_74#_c_245_n N_A_209_368#_c_558_n 0.0105541f $X=0.97 $Y=1.385 $X2=0
+ $Y2=0
cc_276 N_A_27_74#_M1022_g N_A_209_368#_c_623_n 0.0029552f $X=3.145 $Y=2.73 $X2=0
+ $Y2=0
cc_277 N_A_27_74#_c_256_n N_A_209_368#_c_559_n 0.0219614f $X=5.11 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_A_27_74#_M1017_g N_A_209_368#_c_559_n 0.0139565f $X=5.785 $Y=0.83 $X2=0
+ $Y2=0
cc_279 N_A_27_74#_M1018_g N_A_209_368#_c_574_n 0.012181f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_280 N_A_27_74#_c_232_n N_A_209_368#_c_560_n 0.00818799f $X=1.645 $Y=0.34
+ $X2=0 $Y2=0
cc_281 N_A_27_74#_c_234_n N_A_209_368#_c_560_n 0.0133241f $X=1.73 $Y=0.81 $X2=0
+ $Y2=0
cc_282 N_A_27_74#_c_236_n N_A_209_368#_c_560_n 0.0107758f $X=1.815 $Y=0.895
+ $X2=0 $Y2=0
cc_283 N_A_27_74#_c_237_n N_A_209_368#_c_560_n 0.00105808f $X=2.435 $Y=0.81
+ $X2=0 $Y2=0
cc_284 N_A_27_74#_c_321_p N_A_209_368#_c_560_n 7.84915e-19 $X=0.905 $Y=0.96
+ $X2=0 $Y2=0
cc_285 N_A_27_74#_c_245_n N_A_209_368#_c_560_n 0.010763f $X=0.97 $Y=1.385 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_249_n N_A_695_459#_M1003_d 0.00176461f $X=5.56 $Y=0.382
+ $X2=-0.19 $Y2=-0.245
cc_287 N_A_27_74#_M1022_g N_A_695_459#_c_773_n 0.00666974f $X=3.145 $Y=2.73
+ $X2=0 $Y2=0
cc_288 N_A_27_74#_c_240_n N_A_695_459#_c_773_n 0.0087111f $X=3.455 $Y=1.83 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_246_n N_A_695_459#_c_773_n 0.00576765f $X=3.67 $Y=1.37 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_c_262_n N_A_695_459#_c_773_n 0.0195013f $X=3.145 $Y=1.92 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_M1016_g N_A_695_459#_M1000_g 0.00190304f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_292 N_A_27_74#_c_238_n N_A_695_459#_M1000_g 4.66532e-19 $X=3.585 $Y=0.34
+ $X2=0 $Y2=0
cc_293 N_A_27_74#_c_241_n N_A_695_459#_M1000_g 0.00133931f $X=3.67 $Y=0.69 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_c_242_n N_A_695_459#_M1000_g 0.00608928f $X=3.67 $Y=1.285
+ $X2=0 $Y2=0
cc_295 N_A_27_74#_c_361_p N_A_695_459#_M1000_g 0.0165628f $X=4.405 $Y=0.775
+ $X2=0 $Y2=0
cc_296 N_A_27_74#_c_362_p N_A_695_459#_M1000_g 0.00152336f $X=4.49 $Y=0.69 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_M1022_g N_A_695_459#_c_781_n 0.0426774f $X=3.145 $Y=2.73 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_240_n N_A_695_459#_c_781_n 4.15763e-19 $X=3.455 $Y=1.83
+ $X2=0 $Y2=0
cc_299 N_A_27_74#_c_242_n N_A_695_459#_c_775_n 0.020179f $X=3.67 $Y=1.285 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_361_p N_A_695_459#_c_775_n 0.0422234f $X=4.405 $Y=0.775
+ $X2=0 $Y2=0
cc_301 N_A_27_74#_c_246_n N_A_695_459#_c_775_n 0.0103861f $X=3.67 $Y=1.37 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_M1017_g N_A_695_459#_c_776_n 5.90643e-19 $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_303 N_A_27_74#_c_361_p N_A_695_459#_c_776_n 0.00776603f $X=4.405 $Y=0.775
+ $X2=0 $Y2=0
cc_304 N_A_27_74#_c_249_n N_A_695_459#_c_776_n 0.0193861f $X=5.56 $Y=0.382 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_c_256_n N_A_695_459#_c_777_n 0.00115095f $X=5.11 $Y=1.765
+ $X2=0 $Y2=0
cc_306 N_A_27_74#_M1018_g N_A_695_459#_c_803_n 0.00109218f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_307 N_A_27_74#_M1016_g N_A_695_459#_c_778_n 0.00590602f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_308 N_A_27_74#_c_242_n N_A_695_459#_c_778_n 0.0027386f $X=3.67 $Y=1.285 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_361_p N_A_695_459#_c_778_n 0.00186236f $X=4.405 $Y=0.775
+ $X2=0 $Y2=0
cc_310 N_A_27_74#_c_246_n N_A_695_459#_c_778_n 0.00503498f $X=3.67 $Y=1.37 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_M1018_g N_A_541_429#_M1004_g 0.0132833f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_c_249_n N_A_541_429#_c_859_n 0.0117761f $X=5.56 $Y=0.382 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_c_361_p N_A_541_429#_c_860_n 0.00220972f $X=4.405 $Y=0.775
+ $X2=0 $Y2=0
cc_314 N_A_27_74#_M1022_g N_A_541_429#_c_868_n 0.0130279f $X=3.145 $Y=2.73 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_c_240_n N_A_541_429#_c_868_n 0.0293639f $X=3.455 $Y=1.83 $X2=0
+ $Y2=0
cc_316 N_A_27_74#_c_262_n N_A_541_429#_c_868_n 0.00773578f $X=3.145 $Y=1.92
+ $X2=0 $Y2=0
cc_317 N_A_27_74#_M1016_g N_A_541_429#_c_861_n 0.0138199f $X=2.99 $Y=0.805 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_240_n N_A_541_429#_c_861_n 0.00263532f $X=3.455 $Y=1.83
+ $X2=0 $Y2=0
cc_319 N_A_27_74#_c_242_n N_A_541_429#_c_861_n 0.0144307f $X=3.67 $Y=1.285 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_c_246_n N_A_541_429#_c_861_n 0.0135457f $X=3.67 $Y=1.37 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_240_n N_A_541_429#_c_869_n 0.00549631f $X=3.455 $Y=1.83
+ $X2=0 $Y2=0
cc_322 N_A_27_74#_M1022_g N_A_541_429#_c_870_n 0.00702984f $X=3.145 $Y=2.73
+ $X2=0 $Y2=0
cc_323 N_A_27_74#_M1016_g N_A_541_429#_c_862_n 0.00264997f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_324 N_A_27_74#_c_240_n N_A_541_429#_c_862_n 0.023857f $X=3.455 $Y=1.83 $X2=0
+ $Y2=0
cc_325 N_A_27_74#_c_262_n N_A_541_429#_c_862_n 0.00780837f $X=3.145 $Y=1.92
+ $X2=0 $Y2=0
cc_326 N_A_27_74#_M1016_g N_A_541_429#_c_863_n 0.015055f $X=2.99 $Y=0.805 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_240_n N_A_541_429#_c_863_n 0.0180492f $X=3.455 $Y=1.83 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_262_n N_A_541_429#_c_863_n 0.00425381f $X=3.145 $Y=1.92
+ $X2=0 $Y2=0
cc_329 N_A_27_74#_M1016_g N_A_541_429#_c_864_n 0.00395467f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_330 N_A_27_74#_c_238_n N_A_541_429#_c_864_n 0.0217287f $X=3.585 $Y=0.34 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_242_n N_A_541_429#_c_864_n 0.00392507f $X=3.67 $Y=1.285
+ $X2=0 $Y2=0
cc_332 N_A_27_74#_c_246_n N_A_541_429#_c_864_n 0.00210157f $X=3.67 $Y=1.37 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_c_240_n N_A_541_429#_c_865_n 0.0141197f $X=3.455 $Y=1.83 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_256_n N_A_541_429#_c_866_n 0.0116225f $X=5.11 $Y=1.765 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_M1017_g N_A_1217_314#_M1001_g 0.0548248f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_336 N_A_27_74#_c_248_n N_A_1217_314#_M1001_g 0.00120024f $X=5.725 $Y=0.345
+ $X2=0 $Y2=0
cc_337 N_A_27_74#_c_255_n N_A_1217_314#_c_974_n 0.00784778f $X=5.71 $Y=1.765
+ $X2=0 $Y2=0
cc_338 N_A_27_74#_M1017_g N_A_1217_314#_c_966_n 0.00106255f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_339 N_A_27_74#_M1017_g N_A_1217_314#_c_967_n 0.00784778f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_340 N_A_27_74#_c_249_n N_A_1022_424#_M1009_d 0.00253498f $X=5.56 $Y=0.382
+ $X2=-0.19 $Y2=-0.245
cc_341 N_A_27_74#_M1018_g N_A_1022_424#_c_1103_n 0.00566857f $X=5.02 $Y=2.54
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_M1017_g N_A_1022_424#_c_1095_n 0.00924351f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_c_247_n N_A_1022_424#_c_1095_n 0.0115372f $X=5.725 $Y=0.345
+ $X2=0 $Y2=0
cc_344 N_A_27_74#_c_248_n N_A_1022_424#_c_1095_n 0.00326587f $X=5.725 $Y=0.345
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_c_249_n N_A_1022_424#_c_1095_n 0.0145161f $X=5.56 $Y=0.382
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_c_255_n N_A_1022_424#_c_1104_n 0.0157792f $X=5.71 $Y=1.765
+ $X2=0 $Y2=0
cc_347 N_A_27_74#_M1018_g N_A_1022_424#_c_1105_n 9.33337e-19 $X=5.02 $Y=2.54
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_255_n N_A_1022_424#_c_1105_n 0.00878206f $X=5.71 $Y=1.765
+ $X2=0 $Y2=0
cc_349 N_A_27_74#_M1017_g N_A_1022_424#_c_1096_n 0.0079016f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_350 N_A_27_74#_c_255_n N_A_1022_424#_c_1097_n 0.00398323f $X=5.71 $Y=1.765
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_M1017_g N_A_1022_424#_c_1097_n 0.00891922f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_M1017_g N_A_1022_424#_c_1098_n 0.0019325f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_353 N_A_27_74#_M1017_g N_A_1022_424#_c_1101_n 0.0103633f $X=5.785 $Y=0.83
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_c_274_n N_VPWR_M1010_d 0.00284455f $X=0.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_27_74#_c_231_n N_VPWR_M1010_d 0.00140562f $X=0.76 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_356 N_A_27_74#_M1011_g N_VPWR_c_1196_n 0.00277602f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_259_n N_VPWR_c_1196_n 0.0233699f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_274_n N_VPWR_c_1196_n 0.0137812f $X=0.675 $Y=2.035 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_M1011_g N_VPWR_c_1201_n 0.00519767f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_M1022_g N_VPWR_c_1202_n 0.00486888f $X=3.145 $Y=2.73 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_M1018_g N_VPWR_c_1203_n 0.00335089f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_259_n N_VPWR_c_1206_n 0.014549f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_363 N_A_27_74#_M1011_g N_VPWR_c_1207_n 0.0028903f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_364 N_A_27_74#_M1011_g N_VPWR_c_1195_n 0.00983841f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_M1022_g N_VPWR_c_1195_n 0.00647345f $X=3.145 $Y=2.73 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_M1018_g N_VPWR_c_1195_n 0.00425046f $X=5.02 $Y=2.54 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_259_n N_VPWR_c_1195_n 0.0119743f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_M1016_g N_A_434_508#_c_1298_n 0.00106676f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_369 N_A_27_74#_c_238_n N_A_434_508#_c_1298_n 0.012736f $X=3.585 $Y=0.34 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_M1016_g N_A_434_508#_c_1299_n 0.0024813f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_371 N_A_27_74#_M1016_g N_A_434_508#_c_1300_n 2.75345e-19 $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_c_235_n N_A_434_508#_c_1300_n 0.0051689f $X=2.35 $Y=0.895
+ $X2=0 $Y2=0
cc_373 N_A_27_74#_M1016_g N_A_434_508#_c_1301_n 0.00134776f $X=2.99 $Y=0.805
+ $X2=0 $Y2=0
cc_374 N_A_27_74#_c_235_n N_A_434_508#_c_1301_n 0.003952f $X=2.35 $Y=0.895 $X2=0
+ $Y2=0
cc_375 N_A_27_74#_c_229_n N_VGND_M1024_d 8.91422e-19 $X=0.675 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_376 N_A_27_74#_c_244_n N_VGND_M1024_d 0.00910456f $X=0.905 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_377 N_A_27_74#_c_235_n N_VGND_M1013_s 0.0123591f $X=2.35 $Y=0.895 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_237_n N_VGND_M1013_s 0.00298707f $X=2.435 $Y=0.81 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_c_361_p N_VGND_M1000_d 0.015217f $X=4.405 $Y=0.775 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_362_p N_VGND_M1000_d 0.00466296f $X=4.49 $Y=0.69 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_243_n N_VGND_M1000_d 5.85761e-19 $X=4.575 $Y=0.34 $X2=0
+ $Y2=0
cc_382 N_A_27_74#_c_228_n N_VGND_c_1381_n 0.0158413f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_c_229_n N_VGND_c_1381_n 0.00573342f $X=0.675 $Y=1.045 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_233_n N_VGND_c_1381_n 0.0120522f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_244_n N_VGND_c_1381_n 0.0106391f $X=0.905 $Y=1.045 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_c_250_n N_VGND_c_1381_n 0.00213533f $X=0.982 $Y=1.22 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_232_n N_VGND_c_1382_n 0.0143635f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_c_234_n N_VGND_c_1382_n 0.0160274f $X=1.73 $Y=0.81 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_235_n N_VGND_c_1382_n 0.0153167f $X=2.35 $Y=0.895 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_c_237_n N_VGND_c_1382_n 0.0159675f $X=2.435 $Y=0.81 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_239_n N_VGND_c_1382_n 0.0143636f $X=2.52 $Y=0.34 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_238_n N_VGND_c_1383_n 0.01192f $X=3.585 $Y=0.34 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_241_n N_VGND_c_1383_n 0.00492412f $X=3.67 $Y=0.69 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_c_361_p N_VGND_c_1383_n 0.0191408f $X=4.405 $Y=0.775 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_362_p N_VGND_c_1383_n 0.00706899f $X=4.49 $Y=0.69 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_243_n N_VGND_c_1383_n 0.0144122f $X=4.575 $Y=0.34 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_M1017_g N_VGND_c_1384_n 0.00193748f $X=5.785 $Y=0.83 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_247_n N_VGND_c_1384_n 0.0124765f $X=5.725 $Y=0.345 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_248_n N_VGND_c_1384_n 0.00337434f $X=5.725 $Y=0.345 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_361_p N_VGND_c_1388_n 0.00262318f $X=4.405 $Y=0.775 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_243_n N_VGND_c_1388_n 0.0120795f $X=4.575 $Y=0.34 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_c_248_n N_VGND_c_1388_n 0.00653686f $X=5.725 $Y=0.345 $X2=0
+ $Y2=0
cc_403 N_A_27_74#_c_249_n N_VGND_c_1388_n 0.0833744f $X=5.56 $Y=0.382 $X2=0
+ $Y2=0
cc_404 N_A_27_74#_c_228_n N_VGND_c_1390_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_405 N_A_27_74#_c_232_n N_VGND_c_1391_n 0.0441828f $X=1.645 $Y=0.34 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_233_n N_VGND_c_1391_n 0.0117474f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_407 N_A_27_74#_c_250_n N_VGND_c_1391_n 0.00278149f $X=0.982 $Y=1.22 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_238_n N_VGND_c_1392_n 0.0802804f $X=3.585 $Y=0.34 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_239_n N_VGND_c_1392_n 0.0115893f $X=2.52 $Y=0.34 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_361_p N_VGND_c_1392_n 0.00283284f $X=4.405 $Y=0.775 $X2=0
+ $Y2=0
cc_411 N_A_27_74#_c_228_n N_VGND_c_1399_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_c_232_n N_VGND_c_1399_n 0.024692f $X=1.645 $Y=0.34 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_233_n N_VGND_c_1399_n 0.00603725f $X=1.135 $Y=0.34 $X2=0
+ $Y2=0
cc_414 N_A_27_74#_c_235_n N_VGND_c_1399_n 0.0114456f $X=2.35 $Y=0.895 $X2=0
+ $Y2=0
cc_415 N_A_27_74#_c_238_n N_VGND_c_1399_n 0.0424639f $X=3.585 $Y=0.34 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_239_n N_VGND_c_1399_n 0.00583135f $X=2.52 $Y=0.34 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_c_361_p N_VGND_c_1399_n 0.0118617f $X=4.405 $Y=0.775 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_243_n N_VGND_c_1399_n 0.00658903f $X=4.575 $Y=0.34 $X2=0
+ $Y2=0
cc_419 N_A_27_74#_c_248_n N_VGND_c_1399_n 0.0102677f $X=5.725 $Y=0.345 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_c_249_n N_VGND_c_1399_n 0.0466729f $X=5.56 $Y=0.382 $X2=0
+ $Y2=0
cc_421 N_A_27_74#_c_250_n N_VGND_c_1399_n 0.00356277f $X=0.982 $Y=1.22 $X2=0
+ $Y2=0
cc_422 N_D_M1013_g N_A_209_368#_c_550_n 0.00903828f $X=2.56 $Y=0.805 $X2=0 $Y2=0
cc_423 N_D_c_488_n N_A_209_368#_c_561_n 0.00857689f $X=2.485 $Y=1.225 $X2=0
+ $Y2=0
cc_424 N_D_c_490_n N_A_209_368#_c_561_n 0.0116011f $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_425 D N_A_209_368#_c_561_n 0.00173878f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_426 N_D_c_492_n N_A_209_368#_c_561_n 0.0210051f $X=2.165 $Y=1.225 $X2=0 $Y2=0
cc_427 N_D_c_490_n N_A_209_368#_M1012_g 7.72597e-19 $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_428 N_D_c_496_n N_A_209_368#_M1012_g 0.0153516f $X=2.08 $Y=2.215 $X2=0 $Y2=0
cc_429 N_D_M1007_g N_A_209_368#_c_564_n 0.00396362f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_430 N_D_M1007_g N_A_209_368#_c_565_n 0.00670104f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_431 N_D_c_494_n N_A_209_368#_c_565_n 0.0201346f $X=1.89 $Y=2.215 $X2=0 $Y2=0
cc_432 N_D_c_490_n N_A_209_368#_c_565_n 0.00438849f $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_433 N_D_c_496_n N_A_209_368#_c_565_n 0.003673f $X=2.08 $Y=2.215 $X2=0 $Y2=0
cc_434 D N_A_209_368#_c_554_n 0.00865774f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_435 N_D_M1007_g N_A_209_368#_c_566_n 0.0116906f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_436 N_D_c_494_n N_A_209_368#_c_566_n 0.0171661f $X=1.89 $Y=2.215 $X2=0 $Y2=0
cc_437 N_D_c_496_n N_A_209_368#_c_566_n 0.00157283f $X=2.08 $Y=2.215 $X2=0 $Y2=0
cc_438 N_D_M1007_g N_A_209_368#_c_567_n 0.00109206f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_439 N_D_c_490_n N_A_209_368#_c_557_n 0.0275441f $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_440 D N_A_209_368#_c_557_n 0.0106113f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_441 N_D_c_494_n N_A_209_368#_c_558_n 0.00109515f $X=1.89 $Y=2.215 $X2=0 $Y2=0
cc_442 N_D_c_490_n N_A_209_368#_c_558_n 0.0028864f $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_443 N_D_c_496_n N_A_209_368#_c_558_n 0.0289943f $X=2.08 $Y=2.215 $X2=0 $Y2=0
cc_444 N_D_M1007_g N_A_209_368#_c_655_n 0.0152836f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_445 D N_A_209_368#_c_560_n 0.00276667f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_446 N_D_c_492_n N_A_209_368#_c_560_n 0.0167825f $X=2.165 $Y=1.225 $X2=0 $Y2=0
cc_447 N_D_M1007_g N_VPWR_c_1202_n 0.0037204f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_448 N_D_M1007_g N_VPWR_c_1207_n 0.00537532f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_449 N_D_M1007_g N_VPWR_c_1195_n 0.00464944f $X=2.08 $Y=2.75 $X2=0 $Y2=0
cc_450 N_D_c_494_n N_A_434_508#_c_1302_n 0.0283695f $X=1.89 $Y=2.215 $X2=0 $Y2=0
cc_451 N_D_c_496_n N_A_434_508#_c_1302_n 0.00537053f $X=2.08 $Y=2.215 $X2=0
+ $Y2=0
cc_452 N_D_M1013_g N_A_434_508#_c_1298_n 0.00332421f $X=2.56 $Y=0.805 $X2=0
+ $Y2=0
cc_453 N_D_c_488_n N_A_434_508#_c_1299_n 7.12104e-19 $X=2.485 $Y=1.225 $X2=0
+ $Y2=0
cc_454 N_D_c_490_n N_A_434_508#_c_1299_n 0.00719172f $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_455 D N_A_434_508#_c_1299_n 0.0121624f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_456 N_D_c_492_n N_A_434_508#_c_1299_n 0.00172895f $X=2.165 $Y=1.225 $X2=0
+ $Y2=0
cc_457 N_D_c_488_n N_A_434_508#_c_1300_n 0.0011963f $X=2.485 $Y=1.225 $X2=0
+ $Y2=0
cc_458 N_D_c_490_n N_A_434_508#_c_1300_n 0.0283695f $X=1.89 $Y=2.05 $X2=0 $Y2=0
cc_459 D N_A_434_508#_c_1300_n 0.00413233f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_460 N_D_c_492_n N_A_434_508#_c_1300_n 0.00101622f $X=2.165 $Y=1.225 $X2=0
+ $Y2=0
cc_461 N_D_c_488_n N_A_434_508#_c_1301_n 0.0129042f $X=2.485 $Y=1.225 $X2=0
+ $Y2=0
cc_462 D N_A_434_508#_c_1301_n 0.0132098f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_463 N_D_c_492_n N_A_434_508#_c_1301_n 2.14136e-19 $X=2.165 $Y=1.225 $X2=0
+ $Y2=0
cc_464 N_D_M1013_g N_VGND_c_1382_n 9.04059e-19 $X=2.56 $Y=0.805 $X2=0 $Y2=0
cc_465 N_A_209_368#_c_605_n N_A_695_459#_M1004_d 0.0181399f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_466 N_A_209_368#_c_556_n N_A_695_459#_M1004_d 0.00571584f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_467 N_A_209_368#_c_574_n N_A_695_459#_M1004_d 0.00297458f $X=4.905 $Y=2.71
+ $X2=0 $Y2=0
cc_468 N_A_209_368#_c_567_n N_A_695_459#_c_779_n 2.02532e-19 $X=3.37 $Y=2.84
+ $X2=0 $Y2=0
cc_469 N_A_209_368#_c_605_n N_A_695_459#_c_779_n 0.00901849f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_470 N_A_209_368#_c_623_n N_A_695_459#_c_779_n 0.00796481f $X=3.455 $Y=2.71
+ $X2=0 $Y2=0
cc_471 N_A_209_368#_M1015_g N_A_695_459#_M1000_g 0.0306802f $X=3.465 $Y=0.715
+ $X2=0 $Y2=0
cc_472 N_A_209_368#_c_605_n N_A_695_459#_c_781_n 0.00429862f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_473 N_A_209_368#_M1009_g N_A_695_459#_c_776_n 0.00902589f $X=5.125 $Y=0.65
+ $X2=0 $Y2=0
cc_474 N_A_209_368#_c_555_n N_A_695_459#_c_776_n 0.0313132f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_475 N_A_209_368#_c_559_n N_A_695_459#_c_776_n 0.00153551f $X=5.25 $Y=1.315
+ $X2=0 $Y2=0
cc_476 N_A_209_368#_c_555_n N_A_695_459#_c_777_n 0.0104013f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_477 N_A_209_368#_c_556_n N_A_695_459#_c_777_n 0.0439905f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_478 N_A_209_368#_c_605_n N_A_695_459#_c_803_n 0.0217816f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_479 N_A_209_368#_c_556_n N_A_695_459#_c_803_n 0.025276f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_480 N_A_209_368#_c_567_n N_A_541_429#_M1012_d 0.00527995f $X=3.37 $Y=2.84
+ $X2=0 $Y2=0
cc_481 N_A_209_368#_c_605_n N_A_541_429#_M1004_g 0.0168155f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_482 N_A_209_368#_c_556_n N_A_541_429#_M1004_g 0.00266667f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_483 N_A_209_368#_c_623_n N_A_541_429#_M1004_g 6.76691e-19 $X=3.455 $Y=2.71
+ $X2=0 $Y2=0
cc_484 N_A_209_368#_c_574_n N_A_541_429#_M1004_g 0.00469102f $X=4.905 $Y=2.71
+ $X2=0 $Y2=0
cc_485 N_A_209_368#_c_555_n N_A_541_429#_c_858_n 0.00117602f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_486 N_A_209_368#_c_556_n N_A_541_429#_c_858_n 0.00186801f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_487 N_A_209_368#_c_559_n N_A_541_429#_c_858_n 0.00890637f $X=5.25 $Y=1.315
+ $X2=0 $Y2=0
cc_488 N_A_209_368#_M1009_g N_A_541_429#_c_859_n 0.0242638f $X=5.125 $Y=0.65
+ $X2=0 $Y2=0
cc_489 N_A_209_368#_c_567_n N_A_541_429#_c_868_n 0.0154247f $X=3.37 $Y=2.84
+ $X2=0 $Y2=0
cc_490 N_A_209_368#_c_605_n N_A_541_429#_c_868_n 0.0338822f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_491 N_A_209_368#_c_623_n N_A_541_429#_c_868_n 0.00916139f $X=3.455 $Y=2.71
+ $X2=0 $Y2=0
cc_492 N_A_209_368#_M1015_g N_A_541_429#_c_861_n 8.85132e-19 $X=3.465 $Y=0.715
+ $X2=0 $Y2=0
cc_493 N_A_209_368#_M1012_g N_A_541_429#_c_870_n 8.30632e-19 $X=2.615 $Y=2.355
+ $X2=0 $Y2=0
cc_494 N_A_209_368#_c_567_n N_A_541_429#_c_870_n 0.0155615f $X=3.37 $Y=2.84
+ $X2=0 $Y2=0
cc_495 N_A_209_368#_c_561_n N_A_541_429#_c_862_n 0.00337851f $X=2.525 $Y=1.765
+ $X2=0 $Y2=0
cc_496 N_A_209_368#_M1015_g N_A_541_429#_c_864_n 0.00419027f $X=3.465 $Y=0.715
+ $X2=0 $Y2=0
cc_497 N_A_209_368#_c_605_n N_A_541_429#_c_865_n 0.0036702f $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_498 N_A_209_368#_c_605_n N_A_541_429#_c_866_n 2.22941e-19 $X=4.82 $Y=2.71
+ $X2=0 $Y2=0
cc_499 N_A_209_368#_M1023_g N_A_1217_314#_M1006_g 0.0151946f $X=5.55 $Y=2.75
+ $X2=0 $Y2=0
cc_500 N_A_209_368#_c_569_n N_A_1217_314#_M1006_g 0.00176436f $X=5.545 $Y=2.99
+ $X2=0 $Y2=0
cc_501 N_A_209_368#_c_570_n N_A_1217_314#_M1006_g 0.0070221f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_502 N_A_209_368#_c_570_n N_A_1217_314#_c_974_n 0.00160392f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_503 N_A_209_368#_c_571_n N_A_1217_314#_c_974_n 0.0210017f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_504 N_A_209_368#_c_570_n N_A_1217_314#_c_966_n 0.0120093f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_505 N_A_209_368#_c_571_n N_A_1217_314#_c_966_n 6.90151e-19 $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_506 N_A_209_368#_c_569_n N_A_1022_424#_M1018_d 0.0045456f $X=5.545 $Y=2.99
+ $X2=0 $Y2=0
cc_507 N_A_209_368#_c_556_n N_A_1022_424#_c_1103_n 0.0378967f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_508 N_A_209_368#_c_569_n N_A_1022_424#_c_1103_n 0.0123303f $X=5.545 $Y=2.99
+ $X2=0 $Y2=0
cc_509 N_A_209_368#_c_570_n N_A_1022_424#_c_1103_n 0.042276f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_510 N_A_209_368#_c_571_n N_A_1022_424#_c_1103_n 0.00547001f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_511 N_A_209_368#_M1009_g N_A_1022_424#_c_1095_n 0.00183035f $X=5.125 $Y=0.65
+ $X2=0 $Y2=0
cc_512 N_A_209_368#_c_555_n N_A_1022_424#_c_1095_n 0.0116287f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_513 N_A_209_368#_c_559_n N_A_1022_424#_c_1095_n 0.00118967f $X=5.25 $Y=1.315
+ $X2=0 $Y2=0
cc_514 N_A_209_368#_c_555_n N_A_1022_424#_c_1104_n 0.00650602f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_515 N_A_209_368#_c_570_n N_A_1022_424#_c_1104_n 0.0181883f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_516 N_A_209_368#_c_571_n N_A_1022_424#_c_1104_n 0.00255675f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_517 N_A_209_368#_c_555_n N_A_1022_424#_c_1105_n 0.0145175f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_518 N_A_209_368#_c_556_n N_A_1022_424#_c_1105_n 0.0129484f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_519 N_A_209_368#_M1009_g N_A_1022_424#_c_1096_n 0.00176968f $X=5.125 $Y=0.65
+ $X2=0 $Y2=0
cc_520 N_A_209_368#_c_555_n N_A_1022_424#_c_1096_n 0.00600438f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_521 N_A_209_368#_c_559_n N_A_1022_424#_c_1096_n 2.52802e-19 $X=5.25 $Y=1.315
+ $X2=0 $Y2=0
cc_522 N_A_209_368#_c_555_n N_A_1022_424#_c_1097_n 0.0112992f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_523 N_A_209_368#_c_556_n N_A_1022_424#_c_1097_n 0.00518247f $X=4.905 $Y=2.625
+ $X2=0 $Y2=0
cc_524 N_A_209_368#_c_559_n N_A_1022_424#_c_1097_n 2.52802e-19 $X=5.25 $Y=1.315
+ $X2=0 $Y2=0
cc_525 N_A_209_368#_c_555_n N_A_1022_424#_c_1098_n 0.0145134f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_526 N_A_209_368#_c_559_n N_A_1022_424#_c_1098_n 6.86823e-19 $X=5.25 $Y=1.315
+ $X2=0 $Y2=0
cc_527 N_A_209_368#_c_570_n N_A_1022_424#_c_1101_n 0.0029887f $X=5.71 $Y=2.215
+ $X2=0 $Y2=0
cc_528 N_A_209_368#_c_566_n N_VPWR_M1007_s 0.0124309f $X=2.105 $Y=2.71 $X2=0
+ $Y2=0
cc_529 N_A_209_368#_c_605_n N_VPWR_M1002_d 0.00920965f $X=4.82 $Y=2.71 $X2=0
+ $Y2=0
cc_530 N_A_209_368#_c_564_n N_VPWR_c_1196_n 0.0130478f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_531 N_A_209_368#_M1023_g N_VPWR_c_1197_n 5.12146e-19 $X=5.55 $Y=2.75 $X2=0
+ $Y2=0
cc_532 N_A_209_368#_c_569_n N_VPWR_c_1197_n 0.00809712f $X=5.545 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_209_368#_c_570_n N_VPWR_c_1197_n 0.0168077f $X=5.71 $Y=2.215 $X2=0
+ $Y2=0
cc_534 N_A_209_368#_c_564_n N_VPWR_c_1201_n 0.0179277f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_535 N_A_209_368#_c_566_n N_VPWR_c_1201_n 0.00228036f $X=2.105 $Y=2.71 $X2=0
+ $Y2=0
cc_536 N_A_209_368#_c_566_n N_VPWR_c_1202_n 0.00310831f $X=2.105 $Y=2.71 $X2=0
+ $Y2=0
cc_537 N_A_209_368#_c_567_n N_VPWR_c_1202_n 0.0338287f $X=3.37 $Y=2.84 $X2=0
+ $Y2=0
cc_538 N_A_209_368#_c_605_n N_VPWR_c_1202_n 0.00310831f $X=4.82 $Y=2.71 $X2=0
+ $Y2=0
cc_539 N_A_209_368#_c_655_n N_VPWR_c_1202_n 0.00470377f $X=2.19 $Y=2.71 $X2=0
+ $Y2=0
cc_540 N_A_209_368#_c_623_n N_VPWR_c_1202_n 0.00470377f $X=3.455 $Y=2.71 $X2=0
+ $Y2=0
cc_541 N_A_209_368#_M1023_g N_VPWR_c_1203_n 0.00333833f $X=5.55 $Y=2.75 $X2=0
+ $Y2=0
cc_542 N_A_209_368#_c_605_n N_VPWR_c_1203_n 0.014661f $X=4.82 $Y=2.71 $X2=0
+ $Y2=0
cc_543 N_A_209_368#_c_569_n N_VPWR_c_1203_n 0.0584192f $X=5.545 $Y=2.99 $X2=0
+ $Y2=0
cc_544 N_A_209_368#_c_574_n N_VPWR_c_1203_n 0.011836f $X=4.905 $Y=2.71 $X2=0
+ $Y2=0
cc_545 N_A_209_368#_c_564_n N_VPWR_c_1207_n 0.00102152f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_546 N_A_209_368#_c_566_n N_VPWR_c_1207_n 0.026401f $X=2.105 $Y=2.71 $X2=0
+ $Y2=0
cc_547 N_A_209_368#_c_605_n N_VPWR_c_1208_n 0.0285558f $X=4.82 $Y=2.71 $X2=0
+ $Y2=0
cc_548 N_A_209_368#_M1023_g N_VPWR_c_1195_n 0.00425041f $X=5.55 $Y=2.75 $X2=0
+ $Y2=0
cc_549 N_A_209_368#_c_564_n N_VPWR_c_1195_n 0.0162859f $X=1.245 $Y=2.625 $X2=0
+ $Y2=0
cc_550 N_A_209_368#_c_566_n N_VPWR_c_1195_n 0.00980218f $X=2.105 $Y=2.71 $X2=0
+ $Y2=0
cc_551 N_A_209_368#_c_567_n N_VPWR_c_1195_n 0.0370929f $X=3.37 $Y=2.84 $X2=0
+ $Y2=0
cc_552 N_A_209_368#_c_605_n N_VPWR_c_1195_n 0.0286699f $X=4.82 $Y=2.71 $X2=0
+ $Y2=0
cc_553 N_A_209_368#_c_569_n N_VPWR_c_1195_n 0.0323207f $X=5.545 $Y=2.99 $X2=0
+ $Y2=0
cc_554 N_A_209_368#_c_655_n N_VPWR_c_1195_n 0.00551112f $X=2.19 $Y=2.71 $X2=0
+ $Y2=0
cc_555 N_A_209_368#_c_623_n N_VPWR_c_1195_n 0.0057678f $X=3.455 $Y=2.71 $X2=0
+ $Y2=0
cc_556 N_A_209_368#_c_574_n N_VPWR_c_1195_n 0.00626149f $X=4.905 $Y=2.71 $X2=0
+ $Y2=0
cc_557 N_A_209_368#_c_567_n N_A_434_508#_M1007_d 0.00487169f $X=3.37 $Y=2.84
+ $X2=0 $Y2=0
cc_558 N_A_209_368#_c_655_n N_A_434_508#_M1007_d 0.00479347f $X=2.19 $Y=2.71
+ $X2=0 $Y2=0
cc_559 N_A_209_368#_c_561_n N_A_434_508#_c_1302_n 0.00800027f $X=2.525 $Y=1.765
+ $X2=0 $Y2=0
cc_560 N_A_209_368#_M1012_g N_A_434_508#_c_1302_n 0.0133287f $X=2.615 $Y=2.355
+ $X2=0 $Y2=0
cc_561 N_A_209_368#_c_567_n N_A_434_508#_c_1302_n 0.013327f $X=3.37 $Y=2.84
+ $X2=0 $Y2=0
cc_562 N_A_209_368#_c_655_n N_A_434_508#_c_1302_n 0.00407411f $X=2.19 $Y=2.71
+ $X2=0 $Y2=0
cc_563 N_A_209_368#_c_558_n N_A_434_508#_c_1299_n 2.28565e-19 $X=1.565 $Y=1.515
+ $X2=0 $Y2=0
cc_564 N_A_209_368#_c_561_n N_A_434_508#_c_1300_n 0.0137402f $X=2.525 $Y=1.765
+ $X2=0 $Y2=0
cc_565 N_A_209_368#_c_561_n N_A_434_508#_c_1301_n 0.00286318f $X=2.525 $Y=1.765
+ $X2=0 $Y2=0
cc_566 N_A_209_368#_c_567_n A_647_504# 0.00241066f $X=3.37 $Y=2.84 $X2=-0.19
+ $Y2=-0.245
cc_567 N_A_209_368#_c_623_n A_647_504# 0.00297725f $X=3.455 $Y=2.71 $X2=-0.19
+ $Y2=-0.245
cc_568 N_A_209_368#_c_569_n A_1128_508# 8.3332e-19 $X=5.545 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_569 N_A_209_368#_c_570_n A_1128_508# 0.005339f $X=5.71 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_570 N_A_209_368#_c_550_n N_VGND_c_1382_n 0.0176819f $X=3.39 $Y=0.18 $X2=0
+ $Y2=0
cc_571 N_A_209_368#_c_560_n N_VGND_c_1382_n 0.001846f $X=1.58 $Y=1.35 $X2=0
+ $Y2=0
cc_572 N_A_209_368#_c_550_n N_VGND_c_1383_n 0.00296608f $X=3.39 $Y=0.18 $X2=0
+ $Y2=0
cc_573 N_A_209_368#_M1015_g N_VGND_c_1383_n 5.47932e-19 $X=3.465 $Y=0.715 $X2=0
+ $Y2=0
cc_574 N_A_209_368#_M1009_g N_VGND_c_1388_n 0.00275707f $X=5.125 $Y=0.65 $X2=0
+ $Y2=0
cc_575 N_A_209_368#_c_551_n N_VGND_c_1391_n 0.0109808f $X=1.76 $Y=0.18 $X2=0
+ $Y2=0
cc_576 N_A_209_368#_c_550_n N_VGND_c_1392_n 0.0308104f $X=3.39 $Y=0.18 $X2=0
+ $Y2=0
cc_577 N_A_209_368#_c_550_n N_VGND_c_1399_n 0.0411962f $X=3.39 $Y=0.18 $X2=0
+ $Y2=0
cc_578 N_A_209_368#_c_551_n N_VGND_c_1399_n 0.0060077f $X=1.76 $Y=0.18 $X2=0
+ $Y2=0
cc_579 N_A_209_368#_M1009_g N_VGND_c_1399_n 0.00544287f $X=5.125 $Y=0.65 $X2=0
+ $Y2=0
cc_580 N_A_695_459#_c_779_n N_A_541_429#_M1004_g 0.0149161f $X=3.565 $Y=2.445
+ $X2=0 $Y2=0
cc_581 N_A_695_459#_c_773_n N_A_541_429#_M1004_g 0.0150689f $X=3.755 $Y=2.295
+ $X2=0 $Y2=0
cc_582 N_A_695_459#_c_777_n N_A_541_429#_M1004_g 0.00186992f $X=4.565 $Y=2.125
+ $X2=0 $Y2=0
cc_583 N_A_695_459#_c_803_n N_A_541_429#_M1004_g 0.00552963f $X=4.565 $Y=2.29
+ $X2=0 $Y2=0
cc_584 N_A_695_459#_c_773_n N_A_541_429#_c_858_n 0.00253775f $X=3.755 $Y=2.295
+ $X2=0 $Y2=0
cc_585 N_A_695_459#_c_776_n N_A_541_429#_c_858_n 0.0082279f $X=4.565 $Y=1.415
+ $X2=0 $Y2=0
cc_586 N_A_695_459#_c_777_n N_A_541_429#_c_858_n 0.0072995f $X=4.565 $Y=2.125
+ $X2=0 $Y2=0
cc_587 N_A_695_459#_M1000_g N_A_541_429#_c_859_n 0.00751872f $X=3.855 $Y=0.715
+ $X2=0 $Y2=0
cc_588 N_A_695_459#_c_776_n N_A_541_429#_c_859_n 0.00965691f $X=4.565 $Y=1.415
+ $X2=0 $Y2=0
cc_589 N_A_695_459#_M1000_g N_A_541_429#_c_860_n 0.00168151f $X=3.855 $Y=0.715
+ $X2=0 $Y2=0
cc_590 N_A_695_459#_c_776_n N_A_541_429#_c_860_n 0.0137665f $X=4.565 $Y=1.415
+ $X2=0 $Y2=0
cc_591 N_A_695_459#_c_778_n N_A_541_429#_c_860_n 0.0181121f $X=3.855 $Y=1.25
+ $X2=0 $Y2=0
cc_592 N_A_695_459#_c_773_n N_A_541_429#_c_868_n 0.00823106f $X=3.755 $Y=2.295
+ $X2=0 $Y2=0
cc_593 N_A_695_459#_c_781_n N_A_541_429#_c_868_n 0.0138874f $X=3.755 $Y=2.37
+ $X2=0 $Y2=0
cc_594 N_A_695_459#_c_778_n N_A_541_429#_c_861_n 3.94393e-19 $X=3.855 $Y=1.25
+ $X2=0 $Y2=0
cc_595 N_A_695_459#_c_773_n N_A_541_429#_c_869_n 0.00496699f $X=3.755 $Y=2.295
+ $X2=0 $Y2=0
cc_596 N_A_695_459#_c_777_n N_A_541_429#_c_869_n 0.00767326f $X=4.565 $Y=2.125
+ $X2=0 $Y2=0
cc_597 N_A_695_459#_c_773_n N_A_541_429#_c_865_n 0.00296459f $X=3.755 $Y=2.295
+ $X2=0 $Y2=0
cc_598 N_A_695_459#_c_775_n N_A_541_429#_c_865_n 0.0226756f $X=4.48 $Y=1.222
+ $X2=0 $Y2=0
cc_599 N_A_695_459#_c_777_n N_A_541_429#_c_865_n 0.02363f $X=4.565 $Y=2.125
+ $X2=0 $Y2=0
cc_600 N_A_695_459#_c_803_n N_A_541_429#_c_865_n 3.75224e-19 $X=4.565 $Y=2.29
+ $X2=0 $Y2=0
cc_601 N_A_695_459#_c_778_n N_A_541_429#_c_865_n 0.00241698f $X=3.855 $Y=1.25
+ $X2=0 $Y2=0
cc_602 N_A_695_459#_c_773_n N_A_541_429#_c_866_n 0.0195148f $X=3.755 $Y=2.295
+ $X2=0 $Y2=0
cc_603 N_A_695_459#_c_775_n N_A_541_429#_c_866_n 0.00901557f $X=4.48 $Y=1.222
+ $X2=0 $Y2=0
cc_604 N_A_695_459#_c_777_n N_A_541_429#_c_866_n 0.0144265f $X=4.565 $Y=2.125
+ $X2=0 $Y2=0
cc_605 N_A_695_459#_c_803_n N_A_541_429#_c_866_n 0.00553753f $X=4.565 $Y=2.29
+ $X2=0 $Y2=0
cc_606 N_A_695_459#_c_778_n N_A_541_429#_c_866_n 0.0134837f $X=3.855 $Y=1.25
+ $X2=0 $Y2=0
cc_607 N_A_695_459#_c_776_n N_A_1022_424#_c_1095_n 0.0102101f $X=4.565 $Y=1.415
+ $X2=0 $Y2=0
cc_608 N_A_695_459#_c_776_n N_A_1022_424#_c_1096_n 0.00610459f $X=4.565 $Y=1.415
+ $X2=0 $Y2=0
cc_609 N_A_695_459#_c_779_n N_VPWR_c_1202_n 0.00499582f $X=3.565 $Y=2.445 $X2=0
+ $Y2=0
cc_610 N_A_695_459#_c_779_n N_VPWR_c_1208_n 0.00324862f $X=3.565 $Y=2.445 $X2=0
+ $Y2=0
cc_611 N_A_695_459#_c_779_n N_VPWR_c_1195_n 0.00647345f $X=3.565 $Y=2.445 $X2=0
+ $Y2=0
cc_612 N_A_695_459#_M1000_g N_VGND_c_1383_n 0.00178458f $X=3.855 $Y=0.715 $X2=0
+ $Y2=0
cc_613 N_A_695_459#_M1000_g N_VGND_c_1392_n 0.00376447f $X=3.855 $Y=0.715 $X2=0
+ $Y2=0
cc_614 N_A_695_459#_M1000_g N_VGND_c_1399_n 0.00503886f $X=3.855 $Y=0.715 $X2=0
+ $Y2=0
cc_615 N_A_541_429#_c_868_n N_VPWR_M1002_d 0.00530614f $X=3.965 $Y=2.34 $X2=0
+ $Y2=0
cc_616 N_A_541_429#_c_869_n N_VPWR_M1002_d 0.00210574f $X=4.05 $Y=2.255 $X2=0
+ $Y2=0
cc_617 N_A_541_429#_M1004_g N_VPWR_c_1203_n 0.00377953f $X=4.245 $Y=2.54 $X2=0
+ $Y2=0
cc_618 N_A_541_429#_M1004_g N_VPWR_c_1208_n 0.00408189f $X=4.245 $Y=2.54 $X2=0
+ $Y2=0
cc_619 N_A_541_429#_M1004_g N_VPWR_c_1195_n 0.00473901f $X=4.245 $Y=2.54 $X2=0
+ $Y2=0
cc_620 N_A_541_429#_c_870_n N_A_434_508#_c_1302_n 0.0115255f $X=2.855 $Y=2.34
+ $X2=0 $Y2=0
cc_621 N_A_541_429#_c_862_n N_A_434_508#_c_1302_n 0.0181841f $X=2.855 $Y=2.125
+ $X2=0 $Y2=0
cc_622 N_A_541_429#_c_861_n N_A_434_508#_c_1298_n 0.0119891f $X=3.115 $Y=1.49
+ $X2=0 $Y2=0
cc_623 N_A_541_429#_c_861_n N_A_434_508#_c_1299_n 0.00625146f $X=3.115 $Y=1.49
+ $X2=0 $Y2=0
cc_624 N_A_541_429#_c_863_n N_A_434_508#_c_1299_n 0.0136354f $X=3.115 $Y=1.575
+ $X2=0 $Y2=0
cc_625 N_A_541_429#_c_862_n N_A_434_508#_c_1300_n 0.0123059f $X=2.855 $Y=2.125
+ $X2=0 $Y2=0
cc_626 N_A_541_429#_c_861_n N_A_434_508#_c_1301_n 0.0129923f $X=3.115 $Y=1.49
+ $X2=0 $Y2=0
cc_627 N_A_541_429#_c_863_n N_A_434_508#_c_1301_n 0.00564757f $X=3.115 $Y=1.575
+ $X2=0 $Y2=0
cc_628 N_A_541_429#_c_859_n N_VGND_c_1383_n 0.00111902f $X=4.695 $Y=1 $X2=0
+ $Y2=0
cc_629 N_A_541_429#_c_859_n N_VGND_c_1388_n 0.00275707f $X=4.695 $Y=1 $X2=0
+ $Y2=0
cc_630 N_A_541_429#_c_859_n N_VGND_c_1399_n 0.00544287f $X=4.695 $Y=1 $X2=0
+ $Y2=0
cc_631 N_A_1217_314#_M1005_g N_A_1022_424#_M1020_g 0.0176639f $X=7.715 $Y=0.74
+ $X2=0 $Y2=0
cc_632 N_A_1217_314#_c_963_n N_A_1022_424#_M1020_g 0.00933371f $X=6.95 $Y=0.645
+ $X2=0 $Y2=0
cc_633 N_A_1217_314#_c_964_n N_A_1022_424#_M1020_g 0.00885592f $X=7.425 $Y=0.935
+ $X2=0 $Y2=0
cc_634 N_A_1217_314#_c_965_n N_A_1022_424#_M1020_g 0.00418246f $X=7.115 $Y=0.935
+ $X2=0 $Y2=0
cc_635 N_A_1217_314#_c_969_n N_A_1022_424#_M1020_g 0.00363238f $X=7.595 $Y=1.35
+ $X2=0 $Y2=0
cc_636 N_A_1217_314#_M1008_g N_A_1022_424#_M1019_g 0.0191529f $X=7.685 $Y=2.4
+ $X2=0 $Y2=0
cc_637 N_A_1217_314#_c_977_n N_A_1022_424#_M1019_g 4.69176e-19 $X=6.955 $Y=1.985
+ $X2=0 $Y2=0
cc_638 N_A_1217_314#_c_978_n N_A_1022_424#_M1019_g 0.0171642f $X=7.425 $Y=1.775
+ $X2=0 $Y2=0
cc_639 N_A_1217_314#_c_966_n N_A_1022_424#_M1019_g 5.82536e-19 $X=6.25 $Y=1.735
+ $X2=0 $Y2=0
cc_640 N_A_1217_314#_c_967_n N_A_1022_424#_M1019_g 0.00540101f $X=6.25 $Y=1.735
+ $X2=0 $Y2=0
cc_641 N_A_1217_314#_c_968_n N_A_1022_424#_M1019_g 0.00336854f $X=7.645 $Y=1.515
+ $X2=0 $Y2=0
cc_642 N_A_1217_314#_M1001_g N_A_1022_424#_c_1095_n 7.29352e-19 $X=6.175 $Y=0.83
+ $X2=0 $Y2=0
cc_643 N_A_1217_314#_c_974_n N_A_1022_424#_c_1104_n 5.62429e-19 $X=6.25 $Y=2.075
+ $X2=0 $Y2=0
cc_644 N_A_1217_314#_c_966_n N_A_1022_424#_c_1104_n 0.00841858f $X=6.25 $Y=1.735
+ $X2=0 $Y2=0
cc_645 N_A_1217_314#_M1001_g N_A_1022_424#_c_1096_n 0.00121928f $X=6.175 $Y=0.83
+ $X2=0 $Y2=0
cc_646 N_A_1217_314#_M1001_g N_A_1022_424#_c_1097_n 8.80397e-19 $X=6.175 $Y=0.83
+ $X2=0 $Y2=0
cc_647 N_A_1217_314#_c_966_n N_A_1022_424#_c_1097_n 0.0059056f $X=6.25 $Y=1.735
+ $X2=0 $Y2=0
cc_648 N_A_1217_314#_M1001_g N_A_1022_424#_c_1099_n 7.55095e-19 $X=6.175 $Y=0.83
+ $X2=0 $Y2=0
cc_649 N_A_1217_314#_c_978_n N_A_1022_424#_c_1099_n 0.0144321f $X=7.425 $Y=1.775
+ $X2=0 $Y2=0
cc_650 N_A_1217_314#_c_964_n N_A_1022_424#_c_1099_n 0.00889268f $X=7.425
+ $Y=0.935 $X2=0 $Y2=0
cc_651 N_A_1217_314#_c_965_n N_A_1022_424#_c_1099_n 0.0171547f $X=7.115 $Y=0.935
+ $X2=0 $Y2=0
cc_652 N_A_1217_314#_c_981_n N_A_1022_424#_c_1099_n 0.0109633f $X=6.915 $Y=1.775
+ $X2=0 $Y2=0
cc_653 N_A_1217_314#_c_969_n N_A_1022_424#_c_1099_n 0.0245629f $X=7.595 $Y=1.35
+ $X2=0 $Y2=0
cc_654 N_A_1217_314#_M1001_g N_A_1022_424#_c_1100_n 0.00390157f $X=6.175 $Y=0.83
+ $X2=0 $Y2=0
cc_655 N_A_1217_314#_M1005_g N_A_1022_424#_c_1100_n 0.00401851f $X=7.715 $Y=0.74
+ $X2=0 $Y2=0
cc_656 N_A_1217_314#_c_978_n N_A_1022_424#_c_1100_n 0.00111883f $X=7.425
+ $Y=1.775 $X2=0 $Y2=0
cc_657 N_A_1217_314#_c_964_n N_A_1022_424#_c_1100_n 9.38545e-19 $X=7.425
+ $Y=0.935 $X2=0 $Y2=0
cc_658 N_A_1217_314#_c_965_n N_A_1022_424#_c_1100_n 0.00418429f $X=7.115
+ $Y=0.935 $X2=0 $Y2=0
cc_659 N_A_1217_314#_c_981_n N_A_1022_424#_c_1100_n 0.00302844f $X=6.915
+ $Y=1.775 $X2=0 $Y2=0
cc_660 N_A_1217_314#_c_969_n N_A_1022_424#_c_1100_n 0.0031657f $X=7.595 $Y=1.35
+ $X2=0 $Y2=0
cc_661 N_A_1217_314#_c_970_n N_A_1022_424#_c_1100_n 0.0202913f $X=8.135 $Y=1.56
+ $X2=0 $Y2=0
cc_662 N_A_1217_314#_M1001_g N_A_1022_424#_c_1101_n 0.015418f $X=6.175 $Y=0.83
+ $X2=0 $Y2=0
cc_663 N_A_1217_314#_c_976_n N_A_1022_424#_c_1101_n 0.0194417f $X=6.79 $Y=1.775
+ $X2=0 $Y2=0
cc_664 N_A_1217_314#_c_965_n N_A_1022_424#_c_1101_n 0.00905319f $X=7.115
+ $Y=0.935 $X2=0 $Y2=0
cc_665 N_A_1217_314#_c_966_n N_A_1022_424#_c_1101_n 0.02578f $X=6.25 $Y=1.735
+ $X2=0 $Y2=0
cc_666 N_A_1217_314#_c_967_n N_A_1022_424#_c_1101_n 0.00125325f $X=6.25 $Y=1.735
+ $X2=0 $Y2=0
cc_667 N_A_1217_314#_c_981_n N_A_1022_424#_c_1101_n 0.00695811f $X=6.915
+ $Y=1.775 $X2=0 $Y2=0
cc_668 N_A_1217_314#_c_978_n N_VPWR_M1019_d 0.00108767f $X=7.425 $Y=1.775 $X2=0
+ $Y2=0
cc_669 N_A_1217_314#_c_968_n N_VPWR_M1019_d 0.00128514f $X=7.645 $Y=1.515 $X2=0
+ $Y2=0
cc_670 N_A_1217_314#_M1006_g N_VPWR_c_1197_n 0.0139303f $X=6.175 $Y=2.75 $X2=0
+ $Y2=0
cc_671 N_A_1217_314#_c_975_n N_VPWR_c_1197_n 0.00110038f $X=6.25 $Y=2.24 $X2=0
+ $Y2=0
cc_672 N_A_1217_314#_c_976_n N_VPWR_c_1197_n 0.004853f $X=6.79 $Y=1.775 $X2=0
+ $Y2=0
cc_673 N_A_1217_314#_c_977_n N_VPWR_c_1197_n 0.0227945f $X=6.955 $Y=1.985 $X2=0
+ $Y2=0
cc_674 N_A_1217_314#_c_966_n N_VPWR_c_1197_n 0.0107623f $X=6.25 $Y=1.735 $X2=0
+ $Y2=0
cc_675 N_A_1217_314#_M1008_g N_VPWR_c_1198_n 0.00612063f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_676 N_A_1217_314#_c_977_n N_VPWR_c_1198_n 0.0280207f $X=6.955 $Y=1.985 $X2=0
+ $Y2=0
cc_677 N_A_1217_314#_c_978_n N_VPWR_c_1198_n 0.0101401f $X=7.425 $Y=1.775 $X2=0
+ $Y2=0
cc_678 N_A_1217_314#_c_968_n N_VPWR_c_1198_n 0.0100981f $X=7.645 $Y=1.515 $X2=0
+ $Y2=0
cc_679 N_A_1217_314#_c_970_n N_VPWR_c_1198_n 3.95452e-19 $X=8.135 $Y=1.56 $X2=0
+ $Y2=0
cc_680 N_A_1217_314#_c_973_n N_VPWR_c_1200_n 0.00647357f $X=8.135 $Y=1.77 $X2=0
+ $Y2=0
cc_681 N_A_1217_314#_M1006_g N_VPWR_c_1203_n 0.00460063f $X=6.175 $Y=2.75 $X2=0
+ $Y2=0
cc_682 N_A_1217_314#_c_977_n N_VPWR_c_1204_n 0.00743562f $X=6.955 $Y=1.985 $X2=0
+ $Y2=0
cc_683 N_A_1217_314#_M1008_g N_VPWR_c_1205_n 0.005209f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_684 N_A_1217_314#_c_973_n N_VPWR_c_1205_n 0.0048691f $X=8.135 $Y=1.77 $X2=0
+ $Y2=0
cc_685 N_A_1217_314#_M1006_g N_VPWR_c_1195_n 0.00910094f $X=6.175 $Y=2.75 $X2=0
+ $Y2=0
cc_686 N_A_1217_314#_M1008_g N_VPWR_c_1195_n 0.00986839f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_687 N_A_1217_314#_c_973_n N_VPWR_c_1195_n 0.00875947f $X=8.135 $Y=1.77 $X2=0
+ $Y2=0
cc_688 N_A_1217_314#_c_977_n N_VPWR_c_1195_n 0.00847205f $X=6.955 $Y=1.985 $X2=0
+ $Y2=0
cc_689 N_A_1217_314#_M1005_g N_Q_c_1346_n 0.00908676f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_690 N_A_1217_314#_M1021_g N_Q_c_1346_n 0.0081896f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_691 N_A_1217_314#_c_963_n N_Q_c_1346_n 0.00416765f $X=6.95 $Y=0.645 $X2=0
+ $Y2=0
cc_692 N_A_1217_314#_M1008_g N_Q_c_1354_n 0.00283022f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_693 N_A_1217_314#_c_973_n N_Q_c_1354_n 0.00248758f $X=8.135 $Y=1.77 $X2=0
+ $Y2=0
cc_694 N_A_1217_314#_c_968_n N_Q_c_1354_n 0.00149108f $X=7.645 $Y=1.515 $X2=0
+ $Y2=0
cc_695 N_A_1217_314#_c_970_n N_Q_c_1354_n 0.00261762f $X=8.135 $Y=1.56 $X2=0
+ $Y2=0
cc_696 N_A_1217_314#_M1008_g N_Q_c_1347_n 0.00339637f $X=7.685 $Y=2.4 $X2=0
+ $Y2=0
cc_697 N_A_1217_314#_M1005_g N_Q_c_1347_n 0.00132265f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_698 N_A_1217_314#_c_973_n N_Q_c_1347_n 0.00606362f $X=8.135 $Y=1.77 $X2=0
+ $Y2=0
cc_699 N_A_1217_314#_M1021_g N_Q_c_1347_n 0.0110777f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_700 N_A_1217_314#_c_968_n N_Q_c_1347_n 0.0371177f $X=7.645 $Y=1.515 $X2=0
+ $Y2=0
cc_701 N_A_1217_314#_c_969_n N_Q_c_1347_n 0.00787517f $X=7.595 $Y=1.35 $X2=0
+ $Y2=0
cc_702 N_A_1217_314#_c_970_n N_Q_c_1347_n 0.0281936f $X=8.135 $Y=1.56 $X2=0
+ $Y2=0
cc_703 N_A_1217_314#_M1005_g N_Q_c_1348_n 0.00321427f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_704 N_A_1217_314#_M1021_g N_Q_c_1348_n 0.00215589f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_705 N_A_1217_314#_c_969_n N_Q_c_1348_n 0.00486121f $X=7.595 $Y=1.35 $X2=0
+ $Y2=0
cc_706 N_A_1217_314#_c_970_n N_Q_c_1348_n 0.00231623f $X=8.135 $Y=1.56 $X2=0
+ $Y2=0
cc_707 N_A_1217_314#_M1008_g Q 0.00927434f $X=7.685 $Y=2.4 $X2=0 $Y2=0
cc_708 N_A_1217_314#_c_973_n Q 0.0114306f $X=8.135 $Y=1.77 $X2=0 $Y2=0
cc_709 N_A_1217_314#_c_964_n N_VGND_M1020_d 0.00522191f $X=7.425 $Y=0.935 $X2=0
+ $Y2=0
cc_710 N_A_1217_314#_c_969_n N_VGND_M1020_d 0.00181629f $X=7.595 $Y=1.35 $X2=0
+ $Y2=0
cc_711 N_A_1217_314#_M1001_g N_VGND_c_1384_n 0.0140083f $X=6.175 $Y=0.83 $X2=0
+ $Y2=0
cc_712 N_A_1217_314#_c_963_n N_VGND_c_1384_n 0.0336757f $X=6.95 $Y=0.645 $X2=0
+ $Y2=0
cc_713 N_A_1217_314#_c_965_n N_VGND_c_1384_n 0.0121616f $X=7.115 $Y=0.935 $X2=0
+ $Y2=0
cc_714 N_A_1217_314#_M1005_g N_VGND_c_1385_n 0.00508404f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_715 N_A_1217_314#_c_963_n N_VGND_c_1385_n 0.0238225f $X=6.95 $Y=0.645 $X2=0
+ $Y2=0
cc_716 N_A_1217_314#_c_964_n N_VGND_c_1385_n 0.0237562f $X=7.425 $Y=0.935 $X2=0
+ $Y2=0
cc_717 N_A_1217_314#_c_970_n N_VGND_c_1385_n 3.25205e-19 $X=8.135 $Y=1.56 $X2=0
+ $Y2=0
cc_718 N_A_1217_314#_M1021_g N_VGND_c_1387_n 0.00646793f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_719 N_A_1217_314#_M1001_g N_VGND_c_1388_n 0.00347405f $X=6.175 $Y=0.83 $X2=0
+ $Y2=0
cc_720 N_A_1217_314#_c_963_n N_VGND_c_1393_n 0.0145482f $X=6.95 $Y=0.645 $X2=0
+ $Y2=0
cc_721 N_A_1217_314#_M1005_g N_VGND_c_1394_n 0.00434272f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_722 N_A_1217_314#_M1021_g N_VGND_c_1394_n 0.00422942f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_723 N_A_1217_314#_M1001_g N_VGND_c_1399_n 0.00395485f $X=6.175 $Y=0.83 $X2=0
+ $Y2=0
cc_724 N_A_1217_314#_M1005_g N_VGND_c_1399_n 0.00821165f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_725 N_A_1217_314#_M1021_g N_VGND_c_1399_n 0.00787255f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_726 N_A_1217_314#_c_963_n N_VGND_c_1399_n 0.0119922f $X=6.95 $Y=0.645 $X2=0
+ $Y2=0
cc_727 N_A_1217_314#_c_964_n N_VGND_c_1399_n 0.0064626f $X=7.425 $Y=0.935 $X2=0
+ $Y2=0
cc_728 N_A_1022_424#_M1019_g N_VPWR_c_1197_n 0.00242518f $X=7.18 $Y=2.34 $X2=0
+ $Y2=0
cc_729 N_A_1022_424#_M1019_g N_VPWR_c_1198_n 0.0167679f $X=7.18 $Y=2.34 $X2=0
+ $Y2=0
cc_730 N_A_1022_424#_M1019_g N_VPWR_c_1204_n 0.00492916f $X=7.18 $Y=2.34 $X2=0
+ $Y2=0
cc_731 N_A_1022_424#_M1019_g N_VPWR_c_1195_n 0.00511769f $X=7.18 $Y=2.34 $X2=0
+ $Y2=0
cc_732 N_A_1022_424#_M1020_g N_Q_c_1346_n 6.41234e-19 $X=7.165 $Y=0.645 $X2=0
+ $Y2=0
cc_733 N_A_1022_424#_M1019_g N_Q_c_1354_n 3.30752e-19 $X=7.18 $Y=2.34 $X2=0
+ $Y2=0
cc_734 N_A_1022_424#_M1020_g N_VGND_c_1384_n 0.00553153f $X=7.165 $Y=0.645 $X2=0
+ $Y2=0
cc_735 N_A_1022_424#_c_1095_n N_VGND_c_1384_n 0.00851381f $X=5.585 $Y=0.82 $X2=0
+ $Y2=0
cc_736 N_A_1022_424#_c_1096_n N_VGND_c_1384_n 0.00357959f $X=5.67 $Y=1.23 $X2=0
+ $Y2=0
cc_737 N_A_1022_424#_c_1101_n N_VGND_c_1384_n 0.0275041f $X=6.91 $Y=1.355 $X2=0
+ $Y2=0
cc_738 N_A_1022_424#_M1020_g N_VGND_c_1385_n 0.00426329f $X=7.165 $Y=0.645 $X2=0
+ $Y2=0
cc_739 N_A_1022_424#_M1020_g N_VGND_c_1393_n 0.00434272f $X=7.165 $Y=0.645 $X2=0
+ $Y2=0
cc_740 N_A_1022_424#_M1020_g N_VGND_c_1399_n 0.00453351f $X=7.165 $Y=0.645 $X2=0
+ $Y2=0
cc_741 N_VPWR_c_1198_n N_Q_c_1354_n 0.036031f $X=7.405 $Y=2.195 $X2=0 $Y2=0
cc_742 N_VPWR_c_1200_n N_Q_c_1347_n 0.0450788f $X=8.36 $Y=1.985 $X2=0 $Y2=0
cc_743 N_VPWR_c_1205_n Q 0.0157112f $X=8.275 $Y=3.33 $X2=0 $Y2=0
cc_744 N_VPWR_c_1195_n Q 0.0127977f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_745 N_Q_c_1346_n N_VGND_c_1385_n 0.0132163f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_746 N_Q_c_1346_n N_VGND_c_1387_n 0.0308798f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_747 N_Q_c_1346_n N_VGND_c_1394_n 0.0149085f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_748 N_Q_c_1346_n N_VGND_c_1399_n 0.0122037f $X=7.93 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__xor2_2.pxi.spice
* Created: Fri Aug 28 18:18:59 2020
* 
x_PM_SKY130_FD_SC_MS__XOR2_2%A N_A_M1001_g N_A_M1008_g N_A_M1007_g N_A_M1012_g
+ N_A_M1010_g N_A_M1013_g N_A_c_83_n N_A_c_92_n N_A_c_84_n A N_A_c_85_n
+ N_A_c_86_n N_A_c_87_n N_A_c_95_n PM_SKY130_FD_SC_MS__XOR2_2%A
x_PM_SKY130_FD_SC_MS__XOR2_2%B N_B_c_191_n N_B_M1005_g N_B_c_180_n N_B_M1004_g
+ N_B_c_181_n N_B_M1006_g N_B_M1002_g N_B_M1003_g N_B_c_184_n N_B_M1009_g
+ N_B_c_195_n N_B_c_185_n N_B_c_186_n B N_B_c_187_n N_B_c_188_n N_B_c_189_n
+ N_B_c_190_n PM_SKY130_FD_SC_MS__XOR2_2%B
x_PM_SKY130_FD_SC_MS__XOR2_2%A_183_74# N_A_183_74#_M1008_d N_A_183_74#_M1005_d
+ N_A_183_74#_M1000_g N_A_183_74#_M1011_g N_A_183_74#_M1014_g
+ N_A_183_74#_c_296_n N_A_183_74#_c_314_n N_A_183_74#_c_387_p
+ N_A_183_74#_c_317_n N_A_183_74#_c_321_n N_A_183_74#_c_303_n
+ N_A_183_74#_c_304_n N_A_183_74#_c_305_n N_A_183_74#_c_297_n
+ N_A_183_74#_c_306_n N_A_183_74#_c_298_n N_A_183_74#_c_299_n
+ PM_SKY130_FD_SC_MS__XOR2_2%A_183_74#
x_PM_SKY130_FD_SC_MS__XOR2_2%VPWR N_VPWR_M1001_s N_VPWR_M1012_d N_VPWR_M1002_d
+ N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n VPWR
+ N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_401_n N_VPWR_c_410_n
+ N_VPWR_c_411_n PM_SKY130_FD_SC_MS__XOR2_2%VPWR
x_PM_SKY130_FD_SC_MS__XOR2_2%A_313_368# N_A_313_368#_M1012_s
+ N_A_313_368#_M1013_s N_A_313_368#_M1014_d N_A_313_368#_M1003_s
+ N_A_313_368#_c_465_n N_A_313_368#_c_467_n N_A_313_368#_c_468_n
+ N_A_313_368#_c_461_n N_A_313_368#_c_462_n N_A_313_368#_c_488_n
+ N_A_313_368#_c_489_n N_A_313_368#_c_473_n N_A_313_368#_c_463_n
+ N_A_313_368#_c_464_n PM_SKY130_FD_SC_MS__XOR2_2%A_313_368#
x_PM_SKY130_FD_SC_MS__XOR2_2%X N_X_M1011_d N_X_M1009_d N_X_M1000_s N_X_c_518_n
+ N_X_c_527_n N_X_c_531_n N_X_c_532_n X X X X PM_SKY130_FD_SC_MS__XOR2_2%X
x_PM_SKY130_FD_SC_MS__XOR2_2%VGND N_VGND_M1008_s N_VGND_M1004_d N_VGND_M1010_s
+ N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n VGND
+ N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n
+ PM_SKY130_FD_SC_MS__XOR2_2%VGND
x_PM_SKY130_FD_SC_MS__XOR2_2%A_399_74# N_A_399_74#_M1007_d N_A_399_74#_M1006_s
+ N_A_399_74#_c_634_n N_A_399_74#_c_635_n N_A_399_74#_c_630_n
+ N_A_399_74#_c_631_n N_A_399_74#_c_632_n N_A_399_74#_c_633_n
+ PM_SKY130_FD_SC_MS__XOR2_2%A_399_74#
cc_1 VNB N_A_M1001_g 0.0101691f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_2 VNB N_A_M1008_g 0.0215071f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=0.69
cc_3 VNB N_A_M1007_g 0.0251369f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.74
cc_4 VNB N_A_M1010_g 0.029763f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=0.74
cc_5 VNB N_A_c_83_n 0.00355117f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.57
cc_6 VNB N_A_c_84_n 0.0143719f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.57
cc_7 VNB N_A_c_85_n 0.0035296f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.33
cc_8 VNB N_A_c_86_n 0.0492361f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.33
cc_9 VNB N_A_c_87_n 0.0394708f $X=-0.19 $Y=-0.245 $X2=2.435 $Y2=1.515
cc_10 VNB N_B_c_180_n 0.0137875f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.165
cc_11 VNB N_B_c_181_n 0.0166328f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.35
cc_12 VNB N_B_M1002_g 0.00621058f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=2.4
cc_13 VNB N_B_M1003_g 0.00728238f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=0.74
cc_14 VNB N_B_c_184_n 0.0230886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_185_n 0.00310902f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.515
cc_16 VNB N_B_c_186_n 0.0347201f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_B_c_187_n 0.0181516f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.33
cc_18 VNB N_B_c_188_n 0.00585017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_189_n 0.0522742f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.515
cc_20 VNB N_B_c_190_n 0.0209134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_183_74#_M1011_g 0.030475f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.68
cc_22 VNB N_A_183_74#_c_296_n 0.0307495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_183_74#_c_297_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_183_74#_c_298_n 0.00289376f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_25 VNB N_A_183_74#_c_299_n 0.0425942f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.33
cc_26 VNB N_VPWR_c_401_n 0.203486f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_27 VNB X 0.0551698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_563_n 0.00982167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_564_n 0.00770145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_565_n 0.0182584f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=0.74
cc_31 VNB N_VGND_c_566_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_567_n 0.0363605f $X=-0.19 $Y=-0.245 $X2=2.435 $Y2=2.4
cc_33 VNB N_VGND_c_568_n 0.0208042f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.57
cc_34 VNB N_VGND_c_569_n 0.0497191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.33
cc_35 VNB N_VGND_c_570_n 0.272347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_571_n 0.0065087f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.515
cc_37 VNB N_A_399_74#_c_630_n 0.00225138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_399_74#_c_631_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=2.4
cc_39 VNB N_A_399_74#_c_632_n 0.003709f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=0.74
cc_40 VNB N_A_399_74#_c_633_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_M1001_g 0.0317682f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_42 VPB N_A_M1012_g 0.0252785f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=2.4
cc_43 VPB N_A_M1013_g 0.0213198f $X=-0.19 $Y=1.66 $X2=2.435 $Y2=2.4
cc_44 VPB N_A_c_83_n 3.73539e-19 $X=-0.19 $Y=1.66 $X2=2.065 $Y2=1.57
cc_45 VPB N_A_c_92_n 0.00260543f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=1.515
cc_46 VPB N_A_c_84_n 0.0058102f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.57
cc_47 VPB N_A_c_87_n 0.00623051f $X=-0.19 $Y=1.66 $X2=2.435 $Y2=1.515
cc_48 VPB N_A_c_95_n 0.00225047f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.62
cc_49 VPB N_B_c_191_n 0.0226943f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.495
cc_50 VPB N_B_c_180_n 0.00433028f $X=-0.19 $Y=1.66 $X2=0.84 $Y2=1.165
cc_51 VPB N_B_M1002_g 0.0229594f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=2.4
cc_52 VPB N_B_M1003_g 0.0287554f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=0.74
cc_53 VPB N_B_c_195_n 0.0282403f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.705
cc_54 VPB N_A_183_74#_M1000_g 0.0198101f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.35
cc_55 VPB N_A_183_74#_M1014_g 0.020763f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=1.35
cc_56 VPB N_A_183_74#_c_296_n 0.0132546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_183_74#_c_303_n 0.0108843f $X=-0.19 $Y=1.66 $X2=2.065 $Y2=1.57
cc_58 VPB N_A_183_74#_c_304_n 0.0115014f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=1.515
cc_59 VPB N_A_183_74#_c_305_n 0.00144832f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.57
cc_60 VPB N_A_183_74#_c_306_n 0.00157687f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.33
cc_61 VPB N_A_183_74#_c_298_n 4.26294e-19 $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_62 VPB N_A_183_74#_c_299_n 0.00414736f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.33
cc_63 VPB N_VPWR_c_402_n 0.0119967f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=0.74
cc_64 VPB N_VPWR_c_403_n 0.0357725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_404_n 0.0059449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_405_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_406_n 0.0450697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_407_n 0.0366392f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.57
cc_69 VPB N_VPWR_c_408_n 0.0193916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_401_n 0.0813486f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_71 VPB N_VPWR_c_410_n 0.0061237f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.62
cc_72 VPB N_VPWR_c_411_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.6
cc_73 VPB N_A_313_368#_c_461_n 0.00467254f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=0.74
cc_74 VPB N_A_313_368#_c_462_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_313_368#_c_463_n 0.00858623f $X=-0.19 $Y=1.66 $X2=2.35 $Y2=1.515
cc_76 VPB N_A_313_368#_c_464_n 0.0335483f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.33
cc_77 VPB N_X_c_518_n 0.00722749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB X 0.00790891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_B_c_180_n 0.0035775f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_80 N_A_c_83_n N_B_c_180_n 8.76719e-19 $X=2.065 $Y=1.57 $X2=0 $Y2=0
cc_81 N_A_c_84_n N_B_c_180_n 0.00780989f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_82 N_A_c_85_n N_B_c_180_n 0.00298508f $X=0.75 $Y=1.33 $X2=0 $Y2=0
cc_83 N_A_c_86_n N_B_c_180_n 0.0101554f $X=0.84 $Y=1.33 $X2=0 $Y2=0
cc_84 N_A_c_87_n N_B_c_180_n 0.00434248f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_M1001_g N_B_c_195_n 0.0724811f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_86 N_A_M1012_g N_B_c_195_n 0.00434248f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_c_84_n N_B_c_195_n 0.0105252f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_88 N_A_c_86_n N_B_c_195_n 0.00444506f $X=0.84 $Y=1.33 $X2=0 $Y2=0
cc_89 N_A_c_95_n N_B_c_195_n 0.00295986f $X=0.75 $Y=1.62 $X2=0 $Y2=0
cc_90 N_A_M1008_g N_B_c_185_n 0.00380641f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_91 N_A_M1007_g N_B_c_185_n 0.00114688f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_c_83_n N_B_c_185_n 0.00431114f $X=2.065 $Y=1.57 $X2=0 $Y2=0
cc_93 N_A_c_84_n N_B_c_185_n 0.0247694f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_94 N_A_c_85_n N_B_c_185_n 0.0162366f $X=0.75 $Y=1.33 $X2=0 $Y2=0
cc_95 N_A_M1008_g N_B_c_186_n 0.0101554f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_96 N_A_M1007_g N_B_c_186_n 0.0114041f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_c_83_n N_B_c_186_n 4.0997e-19 $X=2.065 $Y=1.57 $X2=0 $Y2=0
cc_98 N_A_c_84_n N_B_c_186_n 0.00125809f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_99 N_A_c_85_n N_B_c_186_n 0.00133827f $X=0.75 $Y=1.33 $X2=0 $Y2=0
cc_100 N_A_M1008_g N_B_c_187_n 0.0222847f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_101 N_A_M1007_g N_B_c_187_n 0.0159573f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_M1007_g N_B_c_190_n 0.0148516f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_M1010_g N_B_c_190_n 0.0125184f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_c_83_n N_B_c_190_n 0.0503265f $X=2.065 $Y=1.57 $X2=0 $Y2=0
cc_105 N_A_c_84_n N_B_c_190_n 0.0140337f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_106 N_A_c_87_n N_B_c_190_n 0.00514776f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A_M1013_g N_A_183_74#_M1000_g 0.0244865f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_M1008_g N_A_183_74#_c_296_n 0.00915992f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_109 N_A_c_85_n N_A_183_74#_c_296_n 0.0341159f $X=0.75 $Y=1.33 $X2=0 $Y2=0
cc_110 N_A_c_86_n N_A_183_74#_c_296_n 0.0241688f $X=0.84 $Y=1.33 $X2=0 $Y2=0
cc_111 N_A_c_95_n N_A_183_74#_c_296_n 0.0135837f $X=0.75 $Y=1.62 $X2=0 $Y2=0
cc_112 N_A_M1008_g N_A_183_74#_c_314_n 0.01155f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_113 N_A_c_85_n N_A_183_74#_c_314_n 0.012793f $X=0.75 $Y=1.33 $X2=0 $Y2=0
cc_114 N_A_c_86_n N_A_183_74#_c_314_n 0.00693309f $X=0.84 $Y=1.33 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_A_183_74#_c_317_n 0.0192051f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_116 N_A_c_84_n N_A_183_74#_c_317_n 0.00840476f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_117 N_A_c_86_n N_A_183_74#_c_317_n 7.82553e-19 $X=0.84 $Y=1.33 $X2=0 $Y2=0
cc_118 N_A_c_95_n N_A_183_74#_c_317_n 0.022418f $X=0.75 $Y=1.62 $X2=0 $Y2=0
cc_119 N_A_M1001_g N_A_183_74#_c_321_n 0.00298755f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_120 N_A_M1012_g N_A_183_74#_c_303_n 0.0038924f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_M1012_g N_A_183_74#_c_304_n 0.0140828f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_M1013_g N_A_183_74#_c_304_n 0.0122082f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_c_84_n N_A_183_74#_c_304_n 0.0843289f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_124 N_A_c_87_n N_A_183_74#_c_304_n 7.41451e-19 $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_M1013_g N_A_183_74#_c_305_n 0.00418128f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_c_92_n N_A_183_74#_c_305_n 0.00866859f $X=2.35 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A_M1008_g N_A_183_74#_c_297_n 0.0118202f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_128 N_A_c_85_n N_A_183_74#_c_297_n 0.00111819f $X=0.75 $Y=1.33 $X2=0 $Y2=0
cc_129 N_A_c_84_n N_A_183_74#_c_306_n 0.019491f $X=1.845 $Y=1.57 $X2=0 $Y2=0
cc_130 N_A_c_92_n N_A_183_74#_c_298_n 0.0282435f $X=2.35 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_c_87_n N_A_183_74#_c_298_n 0.00243584f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_c_92_n N_A_183_74#_c_299_n 3.31787e-19 $X=2.35 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_87_n N_A_183_74#_c_299_n 0.0244865f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_M1001_g N_VPWR_c_403_n 0.0190872f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_135 N_A_M1012_g N_VPWR_c_404_n 0.0114727f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_M1013_g N_VPWR_c_404_n 0.00141551f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_M1001_g N_VPWR_c_406_n 0.00460063f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_138 N_A_M1012_g N_VPWR_c_406_n 0.00460063f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_M1013_g N_VPWR_c_407_n 0.00517089f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_M1001_g N_VPWR_c_401_n 0.00908371f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_141 N_A_M1012_g N_VPWR_c_401_n 0.00471f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1013_g N_VPWR_c_401_n 0.00537649f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_M1012_g N_A_313_368#_c_465_n 0.0114498f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_M1013_g N_A_313_368#_c_465_n 0.0101462f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_M1013_g N_A_313_368#_c_467_n 8.84614e-19 $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_M1012_g N_A_313_368#_c_468_n 7.35764e-19 $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_M1013_g N_A_313_368#_c_468_n 0.00632616f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_M1013_g N_A_313_368#_c_462_n 0.00337536f $X=2.435 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_M1012_g N_A_313_368#_c_463_n 4.69176e-19 $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_VGND_c_563_n 0.00783745f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_M1010_g N_VGND_c_564_n 0.00754401f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_M1008_g N_VGND_c_565_n 0.00324657f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_153 N_A_M1008_g N_VGND_c_567_n 0.00790139f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_154 N_A_M1007_g N_VGND_c_568_n 0.00434272f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_M1010_g N_VGND_c_568_n 0.00324657f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_M1008_g N_VGND_c_570_n 0.00414829f $X=0.84 $Y=0.69 $X2=0 $Y2=0
cc_157 N_A_M1007_g N_VGND_c_570_n 0.00823061f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_M1010_g N_VGND_c_570_n 0.00414754f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_M1010_g N_A_399_74#_c_634_n 0.0115434f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_M1010_g N_A_399_74#_c_635_n 0.00392441f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_M1007_g N_A_399_74#_c_631_n 0.00782447f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_M1010_g N_A_399_74#_c_631_n 0.0117268f $X=2.35 $Y=0.74 $X2=0 $Y2=0
cc_163 N_B_c_185_n N_A_183_74#_M1008_d 4.25891e-19 $X=1.32 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_164 N_B_c_181_n N_A_183_74#_M1011_g 0.0320922f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_165 N_B_c_188_n N_A_183_74#_M1011_g 0.00482264f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_166 N_B_c_190_n N_A_183_74#_M1011_g 0.0164208f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_167 N_B_c_191_n N_A_183_74#_c_317_n 0.0148401f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_168 N_B_c_191_n N_A_183_74#_c_303_n 5.76194e-19 $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_169 N_B_c_185_n N_A_183_74#_c_297_n 0.00356533f $X=1.32 $Y=1.095 $X2=0 $Y2=0
cc_170 N_B_c_187_n N_A_183_74#_c_297_n 0.00683951f $X=1.32 $Y=1.12 $X2=0 $Y2=0
cc_171 N_B_c_195_n N_A_183_74#_c_306_n 0.00657502f $X=1.23 $Y=1.81 $X2=0 $Y2=0
cc_172 N_B_M1002_g N_A_183_74#_c_298_n 4.705e-19 $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B_c_188_n N_A_183_74#_c_298_n 0.00972241f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_174 N_B_c_190_n N_A_183_74#_c_298_n 0.0335231f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_175 N_B_M1002_g N_A_183_74#_c_299_n 0.0394208f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_176 N_B_c_188_n N_A_183_74#_c_299_n 0.00235767f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_177 N_B_c_189_n N_A_183_74#_c_299_n 0.013022f $X=4.285 $Y=1.385 $X2=0 $Y2=0
cc_178 N_B_c_190_n N_A_183_74#_c_299_n 0.0130365f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_179 N_B_c_191_n N_VPWR_c_403_n 0.00253889f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_180 N_B_M1002_g N_VPWR_c_405_n 0.0102406f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_181 N_B_M1003_g N_VPWR_c_405_n 0.00398325f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_182 N_B_c_191_n N_VPWR_c_406_n 0.00553757f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_183 N_B_M1002_g N_VPWR_c_407_n 0.00460063f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_184 N_B_M1003_g N_VPWR_c_408_n 0.005209f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_185 N_B_c_191_n N_VPWR_c_401_n 0.0109471f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_186 N_B_M1002_g N_VPWR_c_401_n 0.00908665f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_187 N_B_M1003_g N_VPWR_c_401_n 0.00985858f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_188 N_B_M1002_g N_A_313_368#_c_461_n 0.00100119f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_189 N_B_M1002_g N_A_313_368#_c_473_n 0.0145524f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_190 N_B_M1003_g N_A_313_368#_c_473_n 0.0132272f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_191 N_B_M1002_g N_A_313_368#_c_464_n 5.08493e-19 $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_192 N_B_M1003_g N_A_313_368#_c_464_n 0.0132016f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_193 N_B_c_188_n N_X_M1011_d 0.00102686f $X=3.98 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_194 N_B_c_190_n N_X_M1011_d 7.6724e-19 $X=3.485 $Y=1.28 $X2=-0.19 $Y2=-0.245
cc_195 N_B_M1002_g N_X_c_518_n 0.0128082f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_196 N_B_M1003_g N_X_c_518_n 0.0180064f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_197 N_B_c_188_n N_X_c_518_n 0.0300986f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_198 N_B_c_189_n N_X_c_518_n 0.00413654f $X=4.285 $Y=1.385 $X2=0 $Y2=0
cc_199 N_B_c_190_n N_X_c_518_n 0.00557038f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_200 N_B_c_181_n N_X_c_527_n 0.00852146f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_201 N_B_c_184_n N_X_c_527_n 0.0130838f $X=4.305 $Y=1.22 $X2=0 $Y2=0
cc_202 N_B_c_188_n N_X_c_527_n 0.0249583f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_203 N_B_c_189_n N_X_c_527_n 0.00113975f $X=4.285 $Y=1.385 $X2=0 $Y2=0
cc_204 N_B_c_190_n N_X_c_531_n 0.00199421f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_205 N_B_c_181_n N_X_c_532_n 0.00258525f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_206 N_B_c_184_n N_X_c_532_n 3.33737e-19 $X=4.305 $Y=1.22 $X2=0 $Y2=0
cc_207 N_B_c_190_n N_X_c_532_n 0.0249583f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_208 N_B_c_181_n X 0.00174786f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_209 N_B_M1002_g X 0.0013716f $X=3.785 $Y=2.4 $X2=0 $Y2=0
cc_210 N_B_M1003_g X 0.0117559f $X=4.285 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B_c_184_n X 0.0154377f $X=4.305 $Y=1.22 $X2=0 $Y2=0
cc_212 N_B_c_188_n X 0.0369267f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_213 N_B_c_189_n X 0.0126211f $X=4.285 $Y=1.385 $X2=0 $Y2=0
cc_214 N_B_c_185_n N_VGND_M1004_d 0.00298526f $X=1.32 $Y=1.095 $X2=0 $Y2=0
cc_215 N_B_c_190_n N_VGND_M1004_d 0.00395088f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_216 N_B_c_190_n N_VGND_M1010_s 0.00939434f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_217 N_B_c_185_n N_VGND_c_563_n 0.00762697f $X=1.32 $Y=1.095 $X2=0 $Y2=0
cc_218 N_B_c_186_n N_VGND_c_563_n 5.32428e-19 $X=1.32 $Y=1.285 $X2=0 $Y2=0
cc_219 N_B_c_187_n N_VGND_c_563_n 0.00677708f $X=1.32 $Y=1.12 $X2=0 $Y2=0
cc_220 N_B_c_190_n N_VGND_c_563_n 0.0191843f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_221 N_B_c_187_n N_VGND_c_565_n 0.00434272f $X=1.32 $Y=1.12 $X2=0 $Y2=0
cc_222 N_B_c_181_n N_VGND_c_569_n 0.00278271f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_223 N_B_c_184_n N_VGND_c_569_n 0.00323524f $X=4.305 $Y=1.22 $X2=0 $Y2=0
cc_224 N_B_c_181_n N_VGND_c_570_n 0.00354947f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_225 N_B_c_184_n N_VGND_c_570_n 0.00416766f $X=4.305 $Y=1.22 $X2=0 $Y2=0
cc_226 N_B_c_187_n N_VGND_c_570_n 0.00821949f $X=1.32 $Y=1.12 $X2=0 $Y2=0
cc_227 N_B_c_190_n N_A_399_74#_M1007_d 0.00176461f $X=3.485 $Y=1.28 $X2=-0.19
+ $Y2=-0.245
cc_228 N_B_c_188_n N_A_399_74#_M1006_s 0.00450749f $X=3.98 $Y=1.385 $X2=0 $Y2=0
cc_229 N_B_c_190_n N_A_399_74#_c_634_n 0.0580321f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_230 N_B_c_190_n N_A_399_74#_c_631_n 0.0167101f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_231 N_B_c_184_n N_A_399_74#_c_632_n 0.00417469f $X=4.305 $Y=1.22 $X2=0 $Y2=0
cc_232 N_B_c_181_n N_A_399_74#_c_633_n 0.0100142f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_233 N_B_c_190_n N_A_399_74#_c_633_n 0.00305575f $X=3.485 $Y=1.28 $X2=0 $Y2=0
cc_234 N_A_183_74#_c_321_n N_VPWR_M1001_s 0.00891927f $X=0.415 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_235 N_A_183_74#_c_304_n N_VPWR_M1012_d 0.00412003f $X=2.685 $Y=2.045 $X2=0
+ $Y2=0
cc_236 N_A_183_74#_c_317_n N_VPWR_c_403_n 0.00213291f $X=1.065 $Y=2.045 $X2=0
+ $Y2=0
cc_237 N_A_183_74#_c_321_n N_VPWR_c_403_n 0.0101883f $X=0.415 $Y=2.045 $X2=0
+ $Y2=0
cc_238 N_A_183_74#_c_303_n N_VPWR_c_403_n 0.00901567f $X=1.15 $Y=2.815 $X2=0
+ $Y2=0
cc_239 N_A_183_74#_M1014_g N_VPWR_c_405_n 3.18965e-19 $X=3.335 $Y=2.4 $X2=0
+ $Y2=0
cc_240 N_A_183_74#_c_303_n N_VPWR_c_406_n 0.011066f $X=1.15 $Y=2.815 $X2=0 $Y2=0
cc_241 N_A_183_74#_M1000_g N_VPWR_c_407_n 0.00333896f $X=2.885 $Y=2.4 $X2=0
+ $Y2=0
cc_242 N_A_183_74#_M1014_g N_VPWR_c_407_n 0.00333896f $X=3.335 $Y=2.4 $X2=0
+ $Y2=0
cc_243 N_A_183_74#_M1000_g N_VPWR_c_401_n 0.00422796f $X=2.885 $Y=2.4 $X2=0
+ $Y2=0
cc_244 N_A_183_74#_M1014_g N_VPWR_c_401_n 0.00422796f $X=3.335 $Y=2.4 $X2=0
+ $Y2=0
cc_245 N_A_183_74#_c_303_n N_VPWR_c_401_n 0.00915947f $X=1.15 $Y=2.815 $X2=0
+ $Y2=0
cc_246 N_A_183_74#_c_317_n A_119_392# 0.00598462f $X=1.065 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_183_74#_c_304_n N_A_313_368#_M1012_s 0.00567673f $X=2.685 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_248 N_A_183_74#_c_304_n N_A_313_368#_M1013_s 0.00554439f $X=2.685 $Y=2.045
+ $X2=0 $Y2=0
cc_249 N_A_183_74#_c_305_n N_A_313_368#_M1013_s 0.00137127f $X=2.77 $Y=1.96
+ $X2=0 $Y2=0
cc_250 N_A_183_74#_c_304_n N_A_313_368#_c_465_n 0.0372622f $X=2.685 $Y=2.045
+ $X2=0 $Y2=0
cc_251 N_A_183_74#_M1000_g N_A_313_368#_c_467_n 0.00244571f $X=2.885 $Y=2.4
+ $X2=0 $Y2=0
cc_252 N_A_183_74#_c_304_n N_A_313_368#_c_467_n 0.0176007f $X=2.685 $Y=2.045
+ $X2=0 $Y2=0
cc_253 N_A_183_74#_M1000_g N_A_313_368#_c_468_n 0.0063721f $X=2.885 $Y=2.4 $X2=0
+ $Y2=0
cc_254 N_A_183_74#_M1014_g N_A_313_368#_c_468_n 5.15815e-19 $X=3.335 $Y=2.4
+ $X2=0 $Y2=0
cc_255 N_A_183_74#_M1000_g N_A_313_368#_c_461_n 0.0115958f $X=2.885 $Y=2.4 $X2=0
+ $Y2=0
cc_256 N_A_183_74#_M1014_g N_A_313_368#_c_461_n 0.0133188f $X=3.335 $Y=2.4 $X2=0
+ $Y2=0
cc_257 N_A_183_74#_M1000_g N_A_313_368#_c_462_n 0.001916f $X=2.885 $Y=2.4 $X2=0
+ $Y2=0
cc_258 N_A_183_74#_M1014_g N_A_313_368#_c_488_n 0.00244698f $X=3.335 $Y=2.4
+ $X2=0 $Y2=0
cc_259 N_A_183_74#_M1000_g N_A_313_368#_c_489_n 5.51649e-19 $X=2.885 $Y=2.4
+ $X2=0 $Y2=0
cc_260 N_A_183_74#_M1014_g N_A_313_368#_c_489_n 0.00908606f $X=3.335 $Y=2.4
+ $X2=0 $Y2=0
cc_261 N_A_183_74#_c_303_n N_A_313_368#_c_463_n 0.0448606f $X=1.15 $Y=2.815
+ $X2=0 $Y2=0
cc_262 N_A_183_74#_c_304_n N_A_313_368#_c_463_n 0.0198322f $X=2.685 $Y=2.045
+ $X2=0 $Y2=0
cc_263 N_A_183_74#_M1014_g N_X_c_518_n 0.0166981f $X=3.335 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_183_74#_c_298_n N_X_c_531_n 0.00794396f $X=2.96 $Y=1.515 $X2=0 $Y2=0
cc_265 N_A_183_74#_c_299_n N_X_c_531_n 0.00230303f $X=3.335 $Y=1.515 $X2=0 $Y2=0
cc_266 N_A_183_74#_M1011_g N_X_c_532_n 0.00325715f $X=3.28 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_183_74#_c_296_n N_VGND_M1008_s 0.010282f $X=0.33 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_183_74#_c_314_n N_VGND_M1008_s 0.0082279f $X=0.89 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_183_74#_c_387_p N_VGND_M1008_s 0.0109498f $X=0.415 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_270 N_A_183_74#_c_297_n N_VGND_c_563_n 0.0191765f $X=1.055 $Y=0.595 $X2=0
+ $Y2=0
cc_271 N_A_183_74#_M1011_g N_VGND_c_564_n 0.00132236f $X=3.28 $Y=0.74 $X2=0
+ $Y2=0
cc_272 N_A_183_74#_c_314_n N_VGND_c_565_n 0.0023667f $X=0.89 $Y=0.755 $X2=0
+ $Y2=0
cc_273 N_A_183_74#_c_297_n N_VGND_c_565_n 0.0141563f $X=1.055 $Y=0.595 $X2=0
+ $Y2=0
cc_274 N_A_183_74#_c_314_n N_VGND_c_567_n 0.022543f $X=0.89 $Y=0.755 $X2=0 $Y2=0
cc_275 N_A_183_74#_c_387_p N_VGND_c_567_n 0.014469f $X=0.415 $Y=0.755 $X2=0
+ $Y2=0
cc_276 N_A_183_74#_c_297_n N_VGND_c_567_n 0.00623386f $X=1.055 $Y=0.595 $X2=0
+ $Y2=0
cc_277 N_A_183_74#_M1011_g N_VGND_c_569_n 0.00278271f $X=3.28 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_183_74#_M1011_g N_VGND_c_570_n 0.00358525f $X=3.28 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_183_74#_c_314_n N_VGND_c_570_n 0.00561864f $X=0.89 $Y=0.755 $X2=0
+ $Y2=0
cc_280 N_A_183_74#_c_387_p N_VGND_c_570_n 8.1202e-19 $X=0.415 $Y=0.755 $X2=0
+ $Y2=0
cc_281 N_A_183_74#_c_297_n N_VGND_c_570_n 0.0117515f $X=1.055 $Y=0.595 $X2=0
+ $Y2=0
cc_282 N_A_183_74#_M1011_g N_A_399_74#_c_633_n 0.0119265f $X=3.28 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_VPWR_M1012_d N_A_313_368#_c_465_n 0.0042374f $X=2.025 $Y=1.84 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_404_n N_A_313_368#_c_465_n 0.018542f $X=2.16 $Y=2.81 $X2=0 $Y2=0
cc_285 N_VPWR_c_401_n N_A_313_368#_c_465_n 0.0114452f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_405_n N_A_313_368#_c_461_n 0.0117236f $X=4.01 $Y=2.645 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_407_n N_A_313_368#_c_461_n 0.0557595f $X=3.845 $Y=3.33 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_401_n N_A_313_368#_c_461_n 0.0308071f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_404_n N_A_313_368#_c_462_n 0.0119238f $X=2.16 $Y=2.81 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_407_n N_A_313_368#_c_462_n 0.0234458f $X=3.845 $Y=3.33 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_401_n N_A_313_368#_c_462_n 0.0125551f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_M1002_d N_A_313_368#_c_473_n 0.00427048f $X=3.875 $Y=1.84 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_405_n N_A_313_368#_c_473_n 0.0189268f $X=4.01 $Y=2.645 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_404_n N_A_313_368#_c_463_n 0.0118774f $X=2.16 $Y=2.81 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_406_n N_A_313_368#_c_463_n 0.011066f $X=1.995 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_401_n N_A_313_368#_c_463_n 0.00915947f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_405_n N_A_313_368#_c_464_n 0.0177529f $X=4.01 $Y=2.645 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_408_n N_A_313_368#_c_464_n 0.0149952f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_401_n N_A_313_368#_c_464_n 0.0123436f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_M1002_d N_X_c_518_n 0.00466501f $X=3.875 $Y=1.84 $X2=0 $Y2=0
cc_301 N_A_313_368#_c_461_n N_X_M1000_s 0.00165831f $X=3.395 $Y=2.99 $X2=0 $Y2=0
cc_302 N_A_313_368#_M1014_d N_X_c_518_n 0.00373373f $X=3.425 $Y=1.84 $X2=0 $Y2=0
cc_303 N_A_313_368#_M1003_s N_X_c_518_n 0.00361349f $X=4.375 $Y=1.84 $X2=0 $Y2=0
cc_304 N_A_313_368#_c_488_n N_X_c_518_n 0.0149351f $X=3.535 $Y=2.36 $X2=0 $Y2=0
cc_305 N_A_313_368#_c_473_n N_X_c_518_n 0.0372622f $X=4.345 $Y=2.275 $X2=0 $Y2=0
cc_306 N_A_313_368#_c_464_n N_X_c_518_n 0.025124f $X=4.515 $Y=2.275 $X2=0 $Y2=0
cc_307 N_A_313_368#_c_461_n N_X_c_531_n 0.0118736f $X=3.395 $Y=2.99 $X2=0 $Y2=0
cc_308 N_X_c_527_n N_VGND_c_569_n 0.00236949f $X=4.355 $Y=0.755 $X2=0 $Y2=0
cc_309 X N_VGND_c_569_n 0.0146502f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_310 N_X_c_527_n N_VGND_c_570_n 0.0053981f $X=4.355 $Y=0.755 $X2=0 $Y2=0
cc_311 X N_VGND_c_570_n 0.0120674f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_312 N_X_c_527_n N_A_399_74#_M1006_s 0.00808075f $X=4.355 $Y=0.755 $X2=0 $Y2=0
cc_313 N_X_c_527_n N_A_399_74#_c_632_n 0.0236098f $X=4.355 $Y=0.755 $X2=0 $Y2=0
cc_314 X N_A_399_74#_c_632_n 0.00624725f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_315 N_X_M1011_d N_A_399_74#_c_633_n 0.00176891f $X=3.355 $Y=0.37 $X2=0 $Y2=0
cc_316 N_X_c_527_n N_A_399_74#_c_633_n 0.00570513f $X=4.355 $Y=0.755 $X2=0 $Y2=0
cc_317 N_X_c_532_n N_A_399_74#_c_633_n 0.0148574f $X=3.66 $Y=0.717 $X2=0 $Y2=0
cc_318 N_VGND_M1010_s N_A_399_74#_c_634_n 0.0182056f $X=2.425 $Y=0.37 $X2=0
+ $Y2=0
cc_319 N_VGND_c_564_n N_A_399_74#_c_634_n 0.0259664f $X=2.65 $Y=0.335 $X2=0
+ $Y2=0
cc_320 N_VGND_c_568_n N_A_399_74#_c_634_n 0.0023667f $X=2.48 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_569_n N_A_399_74#_c_634_n 0.00273597f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_570_n N_A_399_74#_c_634_n 0.0106036f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_M1010_s N_A_399_74#_c_635_n 0.00436696f $X=2.425 $Y=0.37 $X2=0
+ $Y2=0
cc_324 N_VGND_c_564_n N_A_399_74#_c_635_n 0.00570874f $X=2.65 $Y=0.335 $X2=0
+ $Y2=0
cc_325 N_VGND_M1010_s N_A_399_74#_c_630_n 6.5924e-19 $X=2.425 $Y=0.37 $X2=0
+ $Y2=0
cc_326 N_VGND_c_564_n N_A_399_74#_c_630_n 0.0148884f $X=2.65 $Y=0.335 $X2=0
+ $Y2=0
cc_327 N_VGND_c_569_n N_A_399_74#_c_630_n 0.0120491f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_570_n N_A_399_74#_c_630_n 0.00658331f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_563_n N_A_399_74#_c_631_n 0.0283283f $X=1.555 $Y=0.595 $X2=0
+ $Y2=0
cc_330 N_VGND_c_564_n N_A_399_74#_c_631_n 0.00613886f $X=2.65 $Y=0.335 $X2=0
+ $Y2=0
cc_331 N_VGND_c_568_n N_A_399_74#_c_631_n 0.0141563f $X=2.48 $Y=0 $X2=0 $Y2=0
cc_332 N_VGND_c_570_n N_A_399_74#_c_631_n 0.0117515f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_569_n N_A_399_74#_c_633_n 0.0650102f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_c_570_n N_A_399_74#_c_633_n 0.0368892f $X=4.56 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__sdfbbp_1.spice
* Created: Fri Aug 28 18:11:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfbbp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfbbp_1  VNB VPB SCD D SCE CLK SET_B RESET_B VPWR Q_N
+ Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1006 A_119_119# N_SCD_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_197_119#_M1033_d N_SCE_M1033_g A_119_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1011 A_299_119# N_D_M1011_g N_A_197_119#_M1033_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_341_93#_M1016_g A_299_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1155 AS=0.0441 PD=0.97 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1043 N_A_341_93#_M1043_d N_SCE_M1043_g N_VGND_M1016_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1155 PD=1.41 PS=0.97 NRD=0 NRS=77.136 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1044 N_VGND_M1044_d N_CLK_M1044_g N_A_622_98#_M1044_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.30025 AS=0.2109 PD=1.74 PS=2.05 NRD=56.868 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_877_98#_M1002_d N_A_622_98#_M1002_g N_VGND_M1044_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2516 AS=0.30025 PD=2.16 PS=1.74 NRD=4.044 NRS=56.868 M=1 R=4.93333
+ SA=75001.1 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1038 N_A_1092_96#_M1038_d N_A_622_98#_M1038_g N_A_197_119#_M1038_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1034 A_1192_96# N_A_877_98#_M1034_g N_A_1092_96#_M1038_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0809375 AS=0.0735 PD=0.89 PS=0.77 NRD=39.336 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_1250_231#_M1000_g A_1192_96# VNB NLOWVT L=0.15 W=0.42
+ AD=0.151254 AS=0.0809375 PD=1.16907 PS=0.89 NRD=87.168 NRS=39.336 M=1 R=2.8
+ SA=75000.8 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_1418_125#_M1025_d N_SET_B_M1025_g N_VGND_M1000_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.229287 AS=0.198071 PD=1.45 PS=1.53093 NRD=78.948 NRS=66.564 M=1
+ R=3.66667 SA=75001.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1021 N_A_1250_231#_M1021_d N_A_1092_96#_M1021_g N_A_1418_125#_M1025_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.229287 PD=0.83 PS=1.45 NRD=0 NRS=78.948 M=1
+ R=3.66667 SA=75001.9 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1022 N_A_1418_125#_M1022_d N_A_1625_93#_M1022_g N_A_1250_231#_M1021_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.322425 AS=0.077 PD=2.47 PS=0.83 NRD=115.896 NRS=0
+ M=1 R=3.66667 SA=75002.3 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1017 A_1880_119# N_A_1250_231#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.15675 PD=0.76 PS=1.67 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1003 N_A_1881_420#_M1003_d N_A_877_98#_M1003_g A_1880_119# VNB NLOWVT L=0.15
+ W=0.55 AD=0.132936 AS=0.05775 PD=1.3268 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1026 A_2061_74# N_A_622_98#_M1026_g N_A_1881_420#_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0819 AS=0.101514 PD=0.81 PS=1.0132 NRD=39.996 NRS=53.34 M=1 R=2.8
+ SA=75000.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_2037_442#_M1001_g A_2061_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0819 PD=0.796552 PS=0.81 NRD=23.568 NRS=39.996 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_2271_74#_M1004_d N_SET_B_M1004_g N_VGND_M1001_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.154634 PD=1.02 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_2037_442#_M1035_d N_A_1881_420#_M1035_g N_A_2271_74#_M1004_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1443 AS=0.1036 PD=1.13 PS=1.02 NRD=17.832 NRS=0 M=1
+ R=4.93333 SA=75001.5 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1045 N_A_2271_74#_M1045_d N_A_1625_93#_M1045_g N_A_2037_442#_M1035_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.2146 AS=0.1443 PD=2.06 PS=1.13 NRD=0.804 NRS=0 M=1
+ R=4.93333 SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g N_A_1625_93#_M1007_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0783879 AS=0.1197 PD=0.771207 PS=1.41 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_Q_N_M1036_d N_A_2037_442#_M1036_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.138112 PD=2.05 PS=1.35879 NRD=0 NRS=4.044 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_2037_442#_M1027_g N_A_2881_74#_M1027_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1005 N_Q_M1005_d N_A_2881_74#_M1005_g N_VGND_M1027_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_SCD_M1010_g N_A_27_464#_M1010_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1056 AS=0.1792 PD=0.97 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.6 A=0.1152 P=1.64 MULT=1
MM1028 A_221_464# N_SCE_M1028_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1056 PD=0.88 PS=0.97 NRD=19.9955 NRS=1.5366 M=1 R=3.55556
+ SA=90000.7 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1039 N_A_197_119#_M1039_d N_D_M1039_g A_221_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.1
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1042 N_A_27_464#_M1042_d N_A_341_93#_M1042_g N_A_197_119#_M1039_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.1792 AS=0.0864 PD=1.84 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90001.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1032 N_A_341_93#_M1032_d N_SCE_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.1792 PD=1.84 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1014 N_VPWR_M1014_d N_CLK_M1014_g N_A_622_98#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1019 N_A_877_98#_M1019_d N_A_622_98#_M1019_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1029 N_A_1092_96#_M1029_d N_A_877_98#_M1029_g N_A_197_119#_M1029_s VPB PSHORT
+ L=0.18 W=0.64 AD=0.130838 AS=0.1792 PD=1.23774 PS=1.84 NRD=23.0687 NRS=0 M=1
+ R=3.55556 SA=90000.2 SB=90002.7 A=0.1152 P=1.64 MULT=1
MM1037 A_1224_419# N_A_622_98#_M1037_g N_A_1092_96#_M1029_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0858623 PD=0.66 PS=0.812264 NRD=30.4759 NRS=14.0658 M=1
+ R=2.33333 SA=90000.8 SB=90003.5 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1250_231#_M1020_g A_1224_419# VPB PSHORT L=0.18 W=0.42
+ AD=0.1509 AS=0.0504 PD=0.996667 PS=0.66 NRD=38.6908 NRS=30.4759 M=1 R=2.33333
+ SA=90001.2 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1015 N_A_1250_231#_M1015_d N_SET_B_M1015_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1512 AS=0.3018 PD=1.2 PS=1.99333 NRD=19.9167 NRS=69.1667 M=1
+ R=4.66667 SA=90001.2 SB=90002.8 A=0.1512 P=2.04 MULT=1
MM1030 A_1583_379# N_A_1092_96#_M1030_g N_A_1250_231#_M1015_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1008 AS=0.1512 PD=1.08 PS=1.2 NRD=15.2281 NRS=0 M=1 R=4.66667
+ SA=90001.7 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1008_d N_A_1625_93#_M1008_g A_1583_379# VPB PSHORT L=0.18 W=0.84
+ AD=0.1386 AS=0.1008 PD=1.17 PS=1.08 NRD=5.8509 NRS=15.2281 M=1 R=4.66667
+ SA=90002.1 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1031 A_1769_379# N_A_1250_231#_M1031_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1719 AS=0.1386 PD=1.425 PS=1.17 NRD=35.0857 NRS=5.8509 M=1 R=4.66667
+ SA=90002.6 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1012 N_A_1881_420#_M1012_d N_A_622_98#_M1012_g A_1769_379# VPB PSHORT L=0.18
+ W=0.84 AD=0.1806 AS=0.1719 PD=1.6 PS=1.425 NRD=0 NRS=35.0857 M=1 R=4.66667
+ SA=90002.7 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1040 A_1989_504# N_A_877_98#_M1040_g N_A_1881_420#_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0903 PD=0.66 PS=0.8 NRD=30.4759 NRS=39.8531 M=1
+ R=2.33333 SA=90001.9 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_2037_442#_M1024_g A_1989_504# VPB PSHORT L=0.18 W=0.42
+ AD=0.152191 AS=0.0504 PD=1.09437 PS=0.66 NRD=44.5417 NRS=30.4759 M=1 R=2.33333
+ SA=90002.3 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1046 N_A_2037_442#_M1046_d N_SET_B_M1046_g N_VPWR_M1024_d VPB PSHORT L=0.18
+ W=1 AD=0.185 AS=0.362359 PD=1.37 PS=2.60563 NRD=18.715 NRS=15.7403 M=1
+ R=5.55556 SA=90001.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1041 A_2387_392# N_A_1881_420#_M1041_g N_A_2037_442#_M1046_d VPB PSHORT L=0.18
+ W=1 AD=0.105 AS=0.185 PD=1.21 PS=1.37 NRD=9.8303 NRS=0 M=1 R=5.55556
+ SA=90002.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_1625_93#_M1009_g A_2387_392# VPB PSHORT L=0.18 W=1
+ AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1047 N_VPWR_M1047_d N_RESET_B_M1047_g N_A_1625_93#_M1047_s VPB PSHORT L=0.18
+ W=0.64 AD=0.123345 AS=0.1696 PD=1.05818 PS=1.81 NRD=42.3747 NRS=0 M=1
+ R=3.55556 SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1013 N_Q_N_M1013_d N_A_2037_442#_M1013_g N_VPWR_M1047_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.215855 PD=2.76 PS=1.85182 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1018 N_VPWR_M1018_d N_A_2037_442#_M1018_g N_A_2881_74#_M1018_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1488 AS=0.2352 PD=1.24286 PS=2.24 NRD=11.7215 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1023 N_Q_M1023_d N_A_2881_74#_M1023_g N_VPWR_M1018_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.1984 PD=2.78 PS=1.65714 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX48_noxref VNB VPB NWDIODE A=30.3272 P=36.36
c_180 VNB 0 3.53193e-20 $X=0 $Y=0
c_2350 A_1769_379# 0 9.6863e-20 $X=8.845 $Y=1.895
*
.include "sky130_fd_sc_ms__sdfbbp_1.pxi.spice"
*
.ends
*
*

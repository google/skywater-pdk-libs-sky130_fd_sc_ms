* File: sky130_fd_sc_ms__a211o_4.pex.spice
* Created: Fri Aug 28 16:56:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A211O_4%A_105_280# 1 2 3 4 15 17 18 21 25 29 31 33
+ 36 38 40 41 43 44 47 50 51 53 55 59 61 63 65 67 71 77
c175 77 0 1.0197e-19 $X=5.89 $Y=1.105
c176 63 0 1.45535e-19 $X=5.725 $Y=1.195
c177 59 0 1.44395e-19 $X=3.195 $Y=0.615
c178 47 0 6.27654e-20 $X=2.13 $Y=1.385
r179 85 86 19.6524 $w=2.33e-07 $l=9.5e-08 $layer=POLY_cond $X=1.965 $Y=1.385
+ $X2=2.06 $Y2=1.385
r180 84 85 69.3004 $w=2.33e-07 $l=3.35e-07 $layer=POLY_cond $X=1.63 $Y=1.385
+ $X2=1.965 $Y2=1.385
r181 77 79 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.89 $Y=1.105
+ $X2=5.89 $Y2=1.195
r182 67 68 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.16 $Y=0.955
+ $X2=3.16 $Y2=1.215
r183 64 74 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.245 $Y=1.195
+ $X2=4.102 $Y2=1.195
r184 63 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=1.195
+ $X2=5.89 $Y2=1.195
r185 63 64 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=5.725 $Y=1.195
+ $X2=4.245 $Y2=1.195
r186 62 67 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.28 $Y=0.955
+ $X2=3.16 $Y2=0.955
r187 61 74 9.70478 $w=2.83e-07 $l=2.4e-07 $layer=LI1_cond $X=4.102 $Y=0.955
+ $X2=4.102 $Y2=1.195
r188 61 71 2.4262 $w=2.83e-07 $l=6e-08 $layer=LI1_cond $X=4.102 $Y=0.955
+ $X2=4.102 $Y2=0.895
r189 61 62 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.96 $Y=0.955
+ $X2=3.28 $Y2=0.955
r190 57 67 4.08157 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=0.87
+ $X2=3.16 $Y2=0.955
r191 57 59 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=3.16 $Y=0.87
+ $X2=3.16 $Y2=0.615
r192 53 55 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=2.615 $Y=2.145
+ $X2=3.66 $Y2=2.145
r193 52 65 3.19717 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.615 $Y=1.215
+ $X2=2.53 $Y2=1.34
r194 51 68 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.04 $Y=1.215
+ $X2=3.16 $Y2=1.215
r195 51 52 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.04 $Y=1.215
+ $X2=2.615 $Y2=1.215
r196 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.53 $Y=2.06
+ $X2=2.615 $Y2=2.145
r197 49 65 3.3845 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.53 $Y=1.55 $X2=2.53
+ $Y2=1.34
r198 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.53 $Y=1.55
+ $X2=2.53 $Y2=2.06
r199 47 86 14.4807 $w=2.33e-07 $l=7e-08 $layer=POLY_cond $X=2.13 $Y=1.385
+ $X2=2.06 $Y2=1.385
r200 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.385 $X2=2.13 $Y2=1.385
r201 44 65 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.34
+ $X2=2.53 $Y2=1.34
r202 44 46 8.64332 $w=4.18e-07 $l=3.15e-07 $layer=LI1_cond $X=2.445 $Y=1.34
+ $X2=2.13 $Y2=1.34
r203 41 47 74.4721 $w=2.33e-07 $l=4.34741e-07 $layer=POLY_cond $X=2.49 $Y=1.22
+ $X2=2.13 $Y2=1.385
r204 41 43 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.49 $Y=1.22
+ $X2=2.49 $Y2=0.74
r205 38 86 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.22
+ $X2=2.06 $Y2=1.385
r206 38 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.06 $Y=1.22
+ $X2=2.06 $Y2=0.74
r207 34 85 8.89359 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.55
+ $X2=1.965 $Y2=1.385
r208 34 36 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.965 $Y=1.55
+ $X2=1.965 $Y2=2.4
r209 31 84 13.0941 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.22
+ $X2=1.63 $Y2=1.385
r210 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.63 $Y=1.22
+ $X2=1.63 $Y2=0.74
r211 27 84 23.7897 $w=2.33e-07 $l=2.14942e-07 $layer=POLY_cond $X=1.515 $Y=1.55
+ $X2=1.63 $Y2=1.385
r212 27 29 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.515 $Y=1.55
+ $X2=1.515 $Y2=2.4
r213 23 27 65.1631 $w=2.33e-07 $l=3.82721e-07 $layer=POLY_cond $X=1.2 $Y=1.4
+ $X2=1.515 $Y2=1.55
r214 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.2 $Y=1.4 $X2=1.2
+ $Y2=0.74
r215 19 23 27.927 $w=2.33e-07 $l=2.06761e-07 $layer=POLY_cond $X=1.065 $Y=1.55
+ $X2=1.2 $Y2=1.4
r216 19 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.065 $Y=1.55
+ $X2=1.065 $Y2=2.4
r217 17 19 24.7186 $w=2.33e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.975 $Y=1.475
+ $X2=1.065 $Y2=1.55
r218 17 18 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.975 $Y=1.475
+ $X2=0.705 $Y2=1.475
r219 13 18 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.615 $Y=1.55
+ $X2=0.705 $Y2=1.475
r220 13 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.615 $Y=1.55
+ $X2=0.615 $Y2=2.4
r221 4 55 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.96 $X2=3.66 $Y2=2.145
r222 3 77 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.615 $X2=5.89 $Y2=1.105
r223 2 71 182 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_NDIFF $count=1 $X=3.975
+ $Y=0.54 $X2=4.14 $Y2=0.895
r224 1 67 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.47 $X2=3.195 $Y2=0.965
r225 1 59 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.47 $X2=3.195 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%B1 3 7 11 15 17 20 21 25 26 33
c100 33 0 6.11229e-20 $X=4.35 $Y=1.635
c101 20 0 6.27654e-20 $X=2.94 $Y=1.635
c102 15 0 7.83994e-20 $X=4.375 $Y=0.935
r103 33 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.635
+ $X2=4.35 $Y2=1.8
r104 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.635
+ $X2=4.35 $Y2=1.47
r105 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.35
+ $Y=1.635 $X2=4.35 $Y2=1.635
r106 26 40 6.74519 $w=4.16e-07 $l=2.995e-07 $layer=LI1_cond $X=4.08 $Y=2.035
+ $X2=4.24 $Y2=1.805
r107 25 40 4.10577 $w=4.16e-07 $l=1.4e-07 $layer=LI1_cond $X=4.24 $Y=1.665
+ $X2=4.24 $Y2=1.805
r108 25 34 0.879808 $w=4.16e-07 $l=3e-08 $layer=LI1_cond $X=4.24 $Y=1.665
+ $X2=4.24 $Y2=1.635
r109 21 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.94 $Y=1.635
+ $X2=2.94 $Y2=1.8
r110 21 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.94 $Y=1.635
+ $X2=2.94 $Y2=1.47
r111 20 23 6.12235 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.945 $Y=1.635
+ $X2=2.945 $Y2=1.805
r112 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.635 $X2=2.94 $Y2=1.635
r113 18 23 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.105 $Y=1.805
+ $X2=2.945 $Y2=1.805
r114 17 40 6.01746 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=4.24 $Y2=1.805
r115 17 18 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=3.105 $Y2=1.805
r116 15 35 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.375 $Y=0.935
+ $X2=4.375 $Y2=1.47
r117 11 36 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.36 $Y=2.46
+ $X2=4.36 $Y2=1.8
r118 7 30 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.98 $Y=0.79
+ $X2=2.98 $Y2=1.47
r119 3 31 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.935 $Y=2.46
+ $X2=2.935 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%C1 3 7 11 13 15 16 25
c58 16 0 5.16691e-20 $X=3.6 $Y=1.295
c59 13 0 1.3059e-19 $X=3.9 $Y=1.29
c60 3 0 1.44395e-19 $X=3.41 $Y=0.79
r61 24 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.885 $Y=1.455
+ $X2=3.9 $Y2=1.455
r62 22 24 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.615 $Y=1.455
+ $X2=3.885 $Y2=1.455
r63 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.455 $X2=3.615 $Y2=1.455
r64 20 22 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.435 $Y=1.455
+ $X2=3.615 $Y2=1.455
r65 18 20 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.41 $Y=1.455
+ $X2=3.435 $Y2=1.455
r66 16 23 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.615 $Y=1.295
+ $X2=3.615 $Y2=1.455
r67 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.29 $X2=3.9
+ $Y2=1.455
r68 13 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.9 $Y=1.29 $X2=3.9
+ $Y2=0.86
r69 9 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.885 $Y=1.62
+ $X2=3.885 $Y2=1.455
r70 9 11 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=3.885 $Y=1.62
+ $X2=3.885 $Y2=2.46
r71 5 20 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=1.62
+ $X2=3.435 $Y2=1.455
r72 5 7 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=3.435 $Y=1.62
+ $X2=3.435 $Y2=2.46
r73 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.29
+ $X2=3.41 $Y2=1.455
r74 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.41 $Y=1.29 $X2=3.41
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%A1 3 7 11 15 17 18 19 30
c51 19 0 8.78532e-20 $X=6 $Y=1.665
c52 15 0 1.54739e-19 $X=6.105 $Y=0.935
c53 11 0 2.28503e-19 $X=6.07 $Y=2.46
c54 7 0 1.25287e-19 $X=5.675 $Y=0.935
c55 3 0 1.60809e-19 $X=5.62 $Y=2.46
r56 29 30 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.07 $Y=1.615
+ $X2=6.105 $Y2=1.615
r57 27 29 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.695 $Y=1.615
+ $X2=6.07 $Y2=1.615
r58 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.695
+ $Y=1.615 $X2=5.695 $Y2=1.615
r59 25 27 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.675 $Y=1.615
+ $X2=5.695 $Y2=1.615
r60 23 25 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=5.62 $Y=1.615
+ $X2=5.675 $Y2=1.615
r61 19 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6 $Y=1.615
+ $X2=5.695 $Y2=1.615
r62 18 28 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.695 $Y2=1.615
r63 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r64 13 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.105 $Y2=1.615
r65 13 15 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.105 $Y2=0.935
r66 9 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.07 $Y=1.78
+ $X2=6.07 $Y2=1.615
r67 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.07 $Y=1.78 $X2=6.07
+ $Y2=2.46
r68 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.45
+ $X2=5.675 $Y2=1.615
r69 5 7 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.675 $Y=1.45
+ $X2=5.675 $Y2=0.935
r70 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.62 $Y=1.78
+ $X2=5.62 $Y2=1.615
r71 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.62 $Y=1.78 $X2=5.62
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%A2 3 5 6 10 11 13 15 20 22 24
c64 22 0 1.25287e-19 $X=5.04 $Y=0.555
c65 20 0 3.8172e-19 $X=6.535 $Y=0.935
r66 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=0.34
+ $X2=5.155 $Y2=0.505
r67 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=0.34 $X2=5.155 $Y2=0.34
r68 24 27 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.155 $Y=0.2
+ $X2=5.155 $Y2=0.34
r69 22 28 8.27445 $w=3.17e-07 $l=2.15e-07 $layer=LI1_cond $X=5.122 $Y=0.555
+ $X2=5.122 $Y2=0.34
r70 20 21 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.535 $Y=0.935
+ $X2=6.535 $Y2=1.385
r71 17 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.535 $Y=0.275
+ $X2=6.535 $Y2=0.935
r72 13 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.52 $Y=1.475 $X2=6.52
+ $Y2=1.385
r73 13 15 382.879 $w=1.8e-07 $l=9.85e-07 $layer=POLY_cond $X=6.52 $Y=1.475
+ $X2=6.52 $Y2=2.46
r74 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=0.2
+ $X2=5.155 $Y2=0.2
r75 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.46 $Y=0.2
+ $X2=6.535 $Y2=0.275
r76 11 12 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=6.46 $Y=0.2
+ $X2=5.32 $Y2=0.2
r77 10 29 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.245 $Y=0.935
+ $X2=5.245 $Y2=0.505
r78 8 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.245 $Y=1.33
+ $X2=5.245 $Y2=0.935
r79 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.17 $Y=1.405
+ $X2=5.245 $Y2=1.33
r80 5 6 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=5.17 $Y=1.405
+ $X2=4.905 $Y2=1.405
r81 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.815 $Y=1.48
+ $X2=4.905 $Y2=1.405
r82 1 3 380.935 $w=1.8e-07 $l=9.8e-07 $layer=POLY_cond $X=4.815 $Y=1.48
+ $X2=4.815 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%VPWR 1 2 3 4 5 16 18 22 26 28 32 38 42 45 46
+ 47 49 62 63 69 72 75
r93 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r97 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r98 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r100 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r101 60 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r102 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 57 75 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=5.555 $Y=3.33
+ $X2=5.217 $Y2=3.33
r104 57 59 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.555 $Y=3.33
+ $X2=6 $Y2=3.33
r105 56 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r107 53 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 50 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.19 $Y2=3.33
r111 50 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 49 75 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=5.217 $Y2=3.33
r113 49 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 47 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 47 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 45 59 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=3.33 $X2=6
+ $Y2=3.33
r117 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.13 $Y=3.33
+ $X2=6.295 $Y2=3.33
r118 44 62 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.46 $Y=3.33 $X2=6.96
+ $Y2=3.33
r119 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=3.33
+ $X2=6.295 $Y2=3.33
r120 40 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=3.245
+ $X2=6.295 $Y2=3.33
r121 40 42 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.295 $Y=3.245
+ $X2=6.295 $Y2=2.375
r122 36 75 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.217 $Y=3.245
+ $X2=5.217 $Y2=3.33
r123 36 38 13.467 $w=6.73e-07 $l=7.6e-07 $layer=LI1_cond $X=5.217 $Y=3.245
+ $X2=5.217 $Y2=2.485
r124 32 35 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.19 $Y=1.985
+ $X2=2.19 $Y2=2.815
r125 30 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r126 30 35 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.815
r127 29 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.25 $Y2=3.33
r128 28 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=3.33
+ $X2=2.19 $Y2=3.33
r129 28 29 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.105 $Y=3.33
+ $X2=1.375 $Y2=3.33
r130 24 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=3.245
+ $X2=1.25 $Y2=3.33
r131 24 26 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=1.25 $Y=3.245
+ $X2=1.25 $Y2=2.225
r132 23 66 3.89925 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.237 $Y2=3.33
r133 22 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=1.25 $Y2=3.33
r134 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=0.475 $Y2=3.33
r135 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.35 $Y=1.985
+ $X2=0.35 $Y2=2.815
r136 16 66 3.24391 $w=2.5e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.237 $Y2=3.33
r137 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.35 $Y2=2.815
r138 5 42 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=6.16
+ $Y=1.96 $X2=6.295 $Y2=2.375
r139 4 38 150 $w=1.7e-07 $l=7.28183e-07 $layer=licon1_PDIFF $count=4 $X=4.905
+ $Y=1.96 $X2=5.39 $Y2=2.485
r140 3 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.84 $X2=2.19 $Y2=2.815
r141 3 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.84 $X2=2.19 $Y2=1.985
r142 2 26 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.155
+ $Y=1.84 $X2=1.29 $Y2=2.225
r143 1 21 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.39 $Y2=2.815
r144 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.39 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%X 1 2 3 4 14 17 21 22 23 27 31 35 37 39 43
+ 44 50 52
r71 49 52 0.128611 $w=4.63e-07 $l=5e-09 $layer=LI1_cond $X=1.562 $Y=0.96
+ $X2=1.562 $Y2=0.965
r72 44 50 2.39545 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.562 $Y=1.325
+ $X2=1.562 $Y2=1.24
r73 44 50 0.385832 $w=4.63e-07 $l=1.5e-08 $layer=LI1_cond $X=1.562 $Y=1.225
+ $X2=1.562 $Y2=1.24
r74 43 49 2.99104 $w=3.17e-07 $l=8.5e-08 $layer=LI1_cond $X=1.562 $Y=0.875
+ $X2=1.562 $Y2=0.96
r75 43 44 6.17331 $w=4.63e-07 $l=2.4e-07 $layer=LI1_cond $X=1.562 $Y=0.985
+ $X2=1.562 $Y2=1.225
r76 43 52 0.514442 $w=4.63e-07 $l=2e-08 $layer=LI1_cond $X=1.562 $Y=0.985
+ $X2=1.562 $Y2=0.965
r77 39 41 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.275 $Y=0.745
+ $X2=2.275 $Y2=0.875
r78 36 43 3.66292 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=1.795 $Y=0.875
+ $X2=1.562 $Y2=0.875
r79 35 41 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.18 $Y=0.875 $X2=2.275
+ $Y2=0.875
r80 35 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.18 $Y=0.875
+ $X2=1.795 $Y2=0.875
r81 31 33 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.74 $Y=1.985
+ $X2=1.74 $Y2=2.815
r82 29 31 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.74 $Y=1.89
+ $X2=1.74 $Y2=1.985
r83 25 43 2.99104 $w=3.17e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.415 $Y=0.79
+ $X2=1.562 $Y2=0.875
r84 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.415 $Y=0.79
+ $X2=1.415 $Y2=0.515
r85 24 37 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.925 $Y=1.805
+ $X2=0.8 $Y2=1.805
r86 23 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.575 $Y=1.805
+ $X2=1.74 $Y2=1.89
r87 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.575 $Y=1.805
+ $X2=0.925 $Y2=1.805
r88 21 44 6.53816 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=1.33 $Y=1.325
+ $X2=1.562 $Y2=1.325
r89 21 22 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.33 $Y=1.325
+ $X2=0.925 $Y2=1.325
r90 17 19 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.8 $Y=1.985 $X2=0.8
+ $Y2=2.815
r91 15 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.89 $X2=0.8
+ $Y2=1.805
r92 15 17 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=1.89 $X2=0.8
+ $Y2=1.985
r93 14 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.72 $X2=0.8
+ $Y2=1.805
r94 13 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.8 $Y=1.41
+ $X2=0.925 $Y2=1.325
r95 13 14 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.8 $Y=1.41 $X2=0.8
+ $Y2=1.72
r96 4 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.84 $X2=1.74 $Y2=2.815
r97 4 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.84 $X2=1.74 $Y2=1.985
r98 3 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.84 $X2=0.84 $Y2=2.815
r99 3 17 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.84 $X2=0.84 $Y2=1.985
r100 2 39 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.37 $X2=2.275 $Y2=0.745
r101 1 52 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=0.37 $X2=1.415 $Y2=0.965
r102 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=0.37 $X2=1.415 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%A_517_392# 1 2 3 4 13 15 16 19 21 25 27 29
+ 31 33 41 42
c73 42 0 2.8071e-20 $X=5.82 $Y=2.035
c74 29 0 4.76839e-20 $X=6.77 $Y=2.12
c75 27 0 6.42024e-21 $X=6.58 $Y=2.035
c76 25 0 3.07137e-19 $X=5.845 $Y=2.465
r77 46 47 3.8299 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.145
+ $X2=5.82 $Y2=2.23
r78 45 46 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=5.82 $Y=2.115 $X2=5.82
+ $Y2=2.145
r79 42 45 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=5.82 $Y=2.035 $X2=5.82
+ $Y2=2.115
r80 33 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.71 $Y=2.485 $X2=2.71
+ $Y2=2.565
r81 29 49 2.96985 $w=2.8e-07 $l=1.01735e-07 $layer=LI1_cond $X=6.77 $Y=2.12
+ $X2=6.745 $Y2=2.03
r82 29 31 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=6.77 $Y=2.12
+ $X2=6.77 $Y2=2.815
r83 28 42 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.96 $Y=2.035
+ $X2=5.82 $Y2=2.035
r84 27 49 4.39021 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.58 $Y=2.035
+ $X2=6.745 $Y2=2.03
r85 27 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.58 $Y=2.035
+ $X2=5.96 $Y2=2.035
r86 25 47 11.5244 $w=2.33e-07 $l=2.35e-07 $layer=LI1_cond $X=5.842 $Y=2.465
+ $X2=5.842 $Y2=2.23
r87 22 39 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.71 $Y=2.145
+ $X2=4.565 $Y2=2.145
r88 21 46 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.68 $Y=2.145
+ $X2=5.82 $Y2=2.145
r89 21 22 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=5.68 $Y=2.145
+ $X2=4.71 $Y2=2.145
r90 17 41 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.605 $Y=2.57
+ $X2=4.565 $Y2=2.485
r91 17 19 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=4.605 $Y=2.57
+ $X2=4.605 $Y2=2.825
r92 16 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=2.4
+ $X2=4.565 $Y2=2.485
r93 15 39 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=2.23
+ $X2=4.565 $Y2=2.145
r94 15 16 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=4.565 $Y=2.23
+ $X2=4.565 $Y2=2.4
r95 14 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=2.485
+ $X2=2.71 $Y2=2.485
r96 13 41 2.76166 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.42 $Y=2.485
+ $X2=4.565 $Y2=2.485
r97 13 14 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=4.42 $Y=2.485
+ $X2=2.875 $Y2=2.485
r98 4 49 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=1.96 $X2=6.745 $Y2=2.105
r99 4 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.61
+ $Y=1.96 $X2=6.745 $Y2=2.815
r100 3 45 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.71
+ $Y=1.96 $X2=5.845 $Y2=2.115
r101 3 25 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=5.71
+ $Y=1.96 $X2=5.845 $Y2=2.465
r102 2 41 600 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=1.96 $X2=4.585 $Y2=2.485
r103 2 39 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=1.96 $X2=4.585 $Y2=2.145
r104 2 19 600 $w=1.7e-07 $l=9.30054e-07 $layer=licon1_PDIFF $count=1 $X=4.45
+ $Y=1.96 $X2=4.585 $Y2=2.825
r105 1 36 600 $w=1.7e-07 $l=6.64568e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.96 $X2=2.71 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%A_605_392# 1 2 11
r14 8 11 41.9489 $w=2.48e-07 $l=9.1e-07 $layer=LI1_cond $X=3.21 $Y=2.865
+ $X2=4.12 $Y2=2.865
r15 2 11 600 $w=1.7e-07 $l=9.34692e-07 $layer=licon1_PDIFF $count=1 $X=3.975
+ $Y=1.96 $X2=4.12 $Y2=2.825
r16 1 8 600 $w=1.7e-07 $l=9.53021e-07 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.96 $X2=3.21 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%VGND 1 2 3 4 5 6 21 23 27 31 37 41 45 47 48
+ 49 50 51 52 58 63 68 82 84 87 90 93
r101 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r102 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r103 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r104 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r105 79 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r106 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r107 76 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r108 76 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r109 75 78 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r110 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 73 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.59
+ $Y2=0
r112 73 75 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=5.04 $Y2=0
r113 72 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r114 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r115 69 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=0 $X2=3.625
+ $Y2=0
r116 69 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.79 $Y=0 $X2=4.08
+ $Y2=0
r117 68 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.59
+ $Y2=0
r118 68 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.08
+ $Y2=0
r119 67 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r120 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r121 64 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.705
+ $Y2=0
r122 64 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.12
+ $Y2=0
r123 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.625
+ $Y2=0
r124 63 66 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.12
+ $Y2=0
r125 62 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r126 62 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r127 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 59 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.845
+ $Y2=0
r129 59 61 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.16
+ $Y2=0
r130 58 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.705
+ $Y2=0
r131 58 61 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.16
+ $Y2=0
r132 56 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r133 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r134 52 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r135 52 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r136 52 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r137 50 78 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=6.48 $Y2=0
r138 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.75
+ $Y2=0
r139 49 81 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.96
+ $Y2=0
r140 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.75
+ $Y2=0
r141 47 55 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.72
+ $Y2=0
r142 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.985
+ $Y2=0
r143 43 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0
r144 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0.76
r145 39 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0
r146 39 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0.765
r147 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0
r148 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0.615
r149 31 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.705 $Y=0.515
+ $X2=2.705 $Y2=0.855
r150 29 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0
r151 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0.515
r152 25 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0
r153 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0.525
r154 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.985
+ $Y2=0
r155 23 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.845
+ $Y2=0
r156 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.15
+ $Y2=0
r157 19 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0
r158 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0.515
r159 6 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.61
+ $Y=0.615 $X2=6.75 $Y2=0.76
r160 5 41 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.615 $X2=4.59 $Y2=0.765
r161 4 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.47 $X2=3.625 $Y2=0.615
r162 3 33 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.37 $X2=2.705 $Y2=0.855
r163 3 31 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.37 $X2=2.705 $Y2=0.515
r164 2 27 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.37 $X2=1.845 $Y2=0.525
r165 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.86
+ $Y=0.37 $X2=0.985 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A211O_4%A_1064_123# 1 2 7 11 13
c23 13 0 2.7959e-19 $X=6.32 $Y=1.11
c24 11 0 1.39955e-19 $X=6.32 $Y=0.845
r25 11 16 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.32 $Y=0.845
+ $X2=6.32 $Y2=0.72
r26 11 13 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.32 $Y=0.845
+ $X2=6.32 $Y2=1.11
r27 7 16 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.235 $Y=0.76
+ $X2=6.32 $Y2=0.72
r28 7 9 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.235 $Y=0.76
+ $X2=5.46 $Y2=0.76
r29 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.615 $X2=6.32 $Y2=0.76
r30 2 13 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.615 $X2=6.32 $Y2=1.11
r31 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.615 $X2=5.46 $Y2=0.76
.ends


* NGSPICE file created from sky130_fd_sc_ms__nand2_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand2_2 A B VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.408e+11p ps=8.4e+06u
M1001 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=6.438e+11p ps=6.18e+06u
M1003 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.442e+11p ps=2.14e+06u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


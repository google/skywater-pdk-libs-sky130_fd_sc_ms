* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 VPWR GATE a_261_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 a_261_392# a_309_338# a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 VPWR CLK a_990_393# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 VPWR a_315_54# a_309_338# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X4 a_267_80# a_315_54# a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 VGND CLK a_984_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_477_124# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VGND GATE a_267_80# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VPWR a_990_393# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND a_315_54# a_309_338# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_27_74# a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 a_984_125# a_27_74# a_990_393# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_83_260# a_309_338# a_477_124# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_83_260# a_315_54# a_487_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X14 a_990_393# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X15 a_315_54# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X16 a_487_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X17 a_27_74# a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND a_990_393# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_315_54# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

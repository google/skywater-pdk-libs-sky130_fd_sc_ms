* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 VPWR a_418_74# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=2.97415e+12p pd=2.322e+07u as=6.048e+11p ps=5.56e+06u
M1001 a_418_74# CIN a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=4.181e+11p ps=4.09e+06u
M1002 VGND A a_1238_74# VNB nlowvt w=740000u l=150000u
+  ad=2.9966e+12p pd=2.115e+07u as=2.664e+11p ps=2.2e+06u
M1003 VPWR A a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.23132e+12p ps=6.6e+06u
M1004 a_740_347# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1005 VPWR A a_538_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1006 a_740_347# CIN VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 SUM a_1024_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1008 SUM a_1024_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1144_347# CIN a_1024_74# VPB pshort w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=3.2e+11p ps=2.64e+06u
M1010 VPWR a_1024_74# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 COUT a_418_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1012 VPWR B a_740_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1024_74# a_418_74# a_740_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_418_74# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_734_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1016 a_1024_74# a_418_74# a_734_74# VNB nlowvt w=740000u l=150000u
+  ad=3.922e+11p pd=2.54e+06u as=0p ps=0u
M1017 a_27_392# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_1238_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.747e+11p ps=2.93e+06u
M1019 COUT a_418_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1024_74# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 COUT a_418_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1024_74# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1023 VPWR a_418_74# COUT VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 SUM a_1024_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 COUT a_418_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_532_74# B a_418_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1027 a_418_74# CIN a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1028 a_1160_74# CIN a_1024_74# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1029 a_538_347# B a_418_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1238_347# B a_1144_347# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_734_74# CIN VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND B a_734_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND A a_532_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_1024_74# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_418_74# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 SUM a_1024_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1238_74# B a_1160_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

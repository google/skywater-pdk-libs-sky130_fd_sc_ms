* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_229_398# B_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5055e+11p pd=1.69e+06u as=5.10375e+11p ps=4.39e+06u
M1001 a_513_74# a_229_398# a_435_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=1.776e+11p ps=1.96e+06u
M1002 VGND A_N a_27_398# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.50975e+11p ps=1.67e+06u
M1003 VGND D a_627_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=3.108e+11p ps=2.32e+06u
M1004 VPWR a_27_398# Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.1844e+12p pd=8.46e+06u as=9.856e+11p ps=8.48e+06u
M1005 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_229_398# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1007 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_229_398# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_435_74# a_27_398# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.9585e+11p ps=2.05e+06u
M1010 VPWR A_N a_27_398# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1011 a_627_74# C a_513_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4_2 A B C D VGND VNB VPB VPWR Y
X0 a_493_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_493_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VGND D Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_119_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 VPWR A a_493_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_27_368# C a_119_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_119_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_27_368# B a_493_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 Y D a_119_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

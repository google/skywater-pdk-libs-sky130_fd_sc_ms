* File: sky130_fd_sc_ms__o32ai_1.pxi.spice
* Created: Fri Aug 28 18:04:07 2020
* 
x_PM_SKY130_FD_SC_MS__O32AI_1%B1 N_B1_c_53_n N_B1_M1009_g N_B1_M1006_g B1
+ N_B1_c_56_n PM_SKY130_FD_SC_MS__O32AI_1%B1
x_PM_SKY130_FD_SC_MS__O32AI_1%B2 N_B2_M1008_g N_B2_M1003_g B2 N_B2_c_81_n
+ N_B2_c_82_n PM_SKY130_FD_SC_MS__O32AI_1%B2
x_PM_SKY130_FD_SC_MS__O32AI_1%A3 N_A3_M1002_g N_A3_M1000_g A3 A3 A3 N_A3_c_113_n
+ N_A3_c_114_n PM_SKY130_FD_SC_MS__O32AI_1%A3
x_PM_SKY130_FD_SC_MS__O32AI_1%A2 N_A2_M1005_g N_A2_M1007_g A2 A2 A2 A2
+ N_A2_c_152_n N_A2_c_153_n PM_SKY130_FD_SC_MS__O32AI_1%A2
x_PM_SKY130_FD_SC_MS__O32AI_1%A1 N_A1_c_190_n N_A1_M1001_g N_A1_M1004_g A1
+ N_A1_c_193_n PM_SKY130_FD_SC_MS__O32AI_1%A1
x_PM_SKY130_FD_SC_MS__O32AI_1%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_c_216_n
+ N_VPWR_c_217_n N_VPWR_c_218_n N_VPWR_c_219_n VPWR N_VPWR_c_220_n
+ N_VPWR_c_215_n PM_SKY130_FD_SC_MS__O32AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O32AI_1%Y N_Y_M1009_d N_Y_M1008_d N_Y_c_248_n Y
+ N_Y_c_250_n N_Y_c_249_n PM_SKY130_FD_SC_MS__O32AI_1%Y
x_PM_SKY130_FD_SC_MS__O32AI_1%A_27_74# N_A_27_74#_M1009_s N_A_27_74#_M1003_d
+ N_A_27_74#_M1007_d N_A_27_74#_c_283_n N_A_27_74#_c_284_n N_A_27_74#_c_296_n
+ N_A_27_74#_c_285_n N_A_27_74#_c_286_n N_A_27_74#_c_287_n N_A_27_74#_c_288_n
+ PM_SKY130_FD_SC_MS__O32AI_1%A_27_74#
x_PM_SKY130_FD_SC_MS__O32AI_1%VGND N_VGND_M1000_d N_VGND_M1001_d N_VGND_c_328_n
+ N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n VGND
+ N_VGND_c_333_n N_VGND_c_334_n PM_SKY130_FD_SC_MS__O32AI_1%VGND
cc_1 VNB N_B1_c_53_n 0.0254704f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_B1_M1006_g 0.00857766f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_3 VNB B1 0.0084694f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_c_56_n 0.0641433f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_5 VNB N_B2_M1003_g 0.0290226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B2_c_81_n 0.00473922f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_7 VNB N_B2_c_82_n 0.0300742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A3_M1000_g 0.0270536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_c_113_n 0.0269877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A3_c_114_n 0.00166948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_M1007_g 0.0260977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_152_n 0.0251326f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_13 VNB N_A2_c_153_n 0.00421825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_190_n 0.0198499f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_15 VNB N_A1_M1004_g 0.00922335f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_16 VNB A1 0.0260696f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A1_c_193_n 0.0557102f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_18 VNB N_VPWR_c_215_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_248_n 0.00685991f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_20 VNB N_Y_c_249_n 0.00701282f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_21 VNB N_A_27_74#_c_283_n 0.005426f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_22 VNB N_A_27_74#_c_284_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_23 VNB N_A_27_74#_c_285_n 0.018049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_286_n 0.00949292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_287_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_288_n 0.0284201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_328_n 0.00977355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_329_n 0.0142197f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_29 VNB N_VGND_c_330_n 0.0361072f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_30 VNB N_VGND_c_331_n 0.0488022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_332_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_333_n 0.0196495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_334_n 0.211748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_B1_M1006_g 0.0272286f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_35 VPB N_B2_M1008_g 0.0231699f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_36 VPB N_B2_c_81_n 0.00305026f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_37 VPB N_B2_c_82_n 0.00802714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A3_M1002_g 0.0246532f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_39 VPB N_A3_c_113_n 0.00566893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A3_c_114_n 0.00100674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A2_M1005_g 0.0230562f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_42 VPB N_A2_c_152_n 0.00554661f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_43 VPB N_A2_c_153_n 0.00292113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A1_M1004_g 0.0307479f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_45 VPB N_VPWR_c_216_n 0.0128289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_217_n 0.0594609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_218_n 0.0145486f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_48 VPB N_VPWR_c_219_n 0.0556281f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_49 VPB N_VPWR_c_220_n 0.0668259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_215_n 0.0808933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_Y_c_250_n 0.00493928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_Y_c_249_n 0.00125128f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_53 N_B1_M1006_g N_B2_M1008_g 0.0453251f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_54 N_B1_c_53_n N_B2_M1003_g 0.0177514f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_55 N_B1_c_56_n N_B2_c_81_n 3.23937e-19 $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_56 N_B1_c_56_n N_B2_c_82_n 0.0469832f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_57 N_B1_M1006_g N_VPWR_c_217_n 0.00694389f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_58 B1 N_VPWR_c_217_n 0.0186019f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_59 N_B1_c_56_n N_VPWR_c_217_n 0.00317208f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_60 N_B1_M1006_g N_VPWR_c_220_n 0.0053223f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_61 N_B1_M1006_g N_VPWR_c_215_n 0.0102181f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_62 N_B1_c_53_n N_Y_c_248_n 0.00369403f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_63 N_B1_c_56_n N_Y_c_248_n 9.24686e-19 $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_64 N_B1_M1006_g N_Y_c_250_n 0.0221689f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_65 N_B1_c_53_n N_Y_c_249_n 0.0038858f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_66 N_B1_M1006_g N_Y_c_249_n 0.0148368f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_67 B1 N_Y_c_249_n 0.0249687f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_B1_c_56_n N_Y_c_249_n 0.00377991f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_69 N_B1_c_53_n N_A_27_74#_c_283_n 0.0118798f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_70 N_B1_c_53_n N_A_27_74#_c_288_n 0.0130776f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_71 B1 N_A_27_74#_c_288_n 0.0260103f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B1_c_56_n N_A_27_74#_c_288_n 0.00198538f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_73 N_B1_c_53_n N_VGND_c_331_n 0.00291626f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_74 N_B1_c_53_n N_VGND_c_334_n 0.00365046f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_75 N_B2_M1008_g N_A3_M1002_g 0.0187284f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_76 N_B2_M1003_g N_A3_M1000_g 0.0247403f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_77 N_B2_c_81_n N_A3_c_113_n 0.00280188f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B2_c_82_n N_A3_c_113_n 0.0176022f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B2_M1008_g N_A3_c_114_n 9.47293e-19 $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_80 N_B2_c_81_n N_A3_c_114_n 0.0271942f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B2_c_82_n N_A3_c_114_n 4.13661e-19 $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B2_M1008_g N_VPWR_c_220_n 0.00349816f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_83 N_B2_M1008_g N_VPWR_c_215_n 0.00430919f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_84 N_B2_M1003_g N_Y_c_248_n 0.00351046f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_85 N_B2_c_81_n N_Y_c_248_n 0.0111437f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B2_c_82_n N_Y_c_248_n 0.00466348f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_87 N_B2_M1008_g N_Y_c_250_n 0.0353476f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_88 N_B2_c_81_n N_Y_c_250_n 0.0267117f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B2_c_82_n N_Y_c_250_n 0.0012618f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B2_M1003_g N_Y_c_249_n 0.00364258f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B2_c_81_n N_Y_c_249_n 0.0323503f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B2_c_82_n N_Y_c_249_n 0.00674683f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B2_M1003_g N_A_27_74#_c_283_n 0.0160377f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B2_M1003_g N_A_27_74#_c_286_n 0.0015383f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_95 N_B2_M1003_g N_VGND_c_331_n 0.00291649f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_96 N_B2_M1003_g N_VGND_c_334_n 0.00362117f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A3_M1002_g N_A2_M1005_g 0.0418006f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A3_c_114_n N_A2_M1005_g 0.00270938f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A3_M1000_g N_A2_M1007_g 0.0239043f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A3_c_113_n N_A2_c_152_n 0.0173872f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A3_c_114_n N_A2_c_152_n 3.65288e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A3_M1002_g N_A2_c_153_n 0.0060915f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A3_c_113_n N_A2_c_153_n 0.00202953f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A3_c_114_n N_A2_c_153_n 0.0953745f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A3_M1002_g N_VPWR_c_220_n 0.00553757f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A3_M1002_g N_VPWR_c_215_n 0.00548045f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A3_c_114_n N_VPWR_c_215_n 0.0118917f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A3_M1002_g N_Y_c_250_n 0.0131951f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A3_c_114_n N_Y_c_250_n 0.0468572f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A3_c_114_n A_345_368# 0.0080887f $X=1.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_111 N_A3_M1000_g N_A_27_74#_c_284_n 0.00227966f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A3_M1000_g N_A_27_74#_c_296_n 0.00785824f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A3_M1000_g N_A_27_74#_c_285_n 0.0119119f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A3_c_113_n N_A_27_74#_c_285_n 4.86414e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A3_c_114_n N_A_27_74#_c_285_n 0.0150021f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A3_M1000_g N_A_27_74#_c_286_n 0.00158144f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A3_c_113_n N_A_27_74#_c_286_n 8.52409e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A3_c_114_n N_A_27_74#_c_286_n 0.0118341f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A3_M1000_g N_A_27_74#_c_287_n 9.95504e-19 $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A3_M1000_g N_VGND_c_328_n 0.00624419f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A3_M1000_g N_VGND_c_331_n 0.00433139f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A3_M1000_g N_VGND_c_334_n 0.00818567f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A2_M1007_g N_A1_c_190_n 0.0199226f $X=2.33 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_124 N_A2_M1005_g N_A1_M1004_g 0.03848f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A2_c_153_n N_A1_M1004_g 0.0129267f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A2_M1007_g A1 5.55987e-19 $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A2_c_152_n A1 5.4813e-19 $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A2_c_153_n A1 0.00716206f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A2_c_152_n N_A1_c_193_n 0.0184923f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A2_c_153_n N_A1_c_193_n 0.00174259f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A2_M1005_g N_VPWR_c_219_n 0.00184516f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A2_c_153_n N_VPWR_c_219_n 0.0445659f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A2_M1005_g N_VPWR_c_220_n 0.00363952f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A2_c_153_n N_VPWR_c_220_n 0.010629f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A2_M1005_g N_VPWR_c_215_n 0.00446867f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A2_c_153_n N_VPWR_c_215_n 0.01298f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A2_c_153_n N_Y_c_250_n 0.0112401f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A2_c_153_n A_345_368# 0.0124161f $X=2.28 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_139 N_A2_c_153_n A_459_368# 0.0144081f $X=2.28 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_140 N_A2_M1007_g N_A_27_74#_c_296_n 9.49738e-19 $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A2_M1007_g N_A_27_74#_c_285_n 0.013469f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A2_c_152_n N_A_27_74#_c_285_n 0.00128242f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A2_c_153_n N_A_27_74#_c_285_n 0.0320971f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A2_M1007_g N_A_27_74#_c_287_n 0.0104013f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_M1007_g N_VGND_c_328_n 0.00754067f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1007_g N_VGND_c_333_n 0.00434272f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_M1007_g N_VGND_c_334_n 0.00822293f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_VPWR_c_219_n 0.0277571f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_149 A1 N_VPWR_c_219_n 0.017092f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A1_c_193_n N_VPWR_c_219_n 0.00275616f $X=3.045 $Y=1.385 $X2=0 $Y2=0
cc_151 N_A1_M1004_g N_VPWR_c_220_n 0.00460063f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A1_M1004_g N_VPWR_c_215_n 0.00909693f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A1_c_190_n N_A_27_74#_c_285_n 0.0101123f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A1_c_190_n N_A_27_74#_c_287_n 0.0081858f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A1_c_190_n N_VGND_c_330_n 0.00495522f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_156 A1 N_VGND_c_330_n 0.0221981f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A1_c_193_n N_VGND_c_330_n 0.00180116f $X=3.045 $Y=1.385 $X2=0 $Y2=0
cc_158 N_A1_c_190_n N_VGND_c_333_n 0.00434272f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A1_c_190_n N_VGND_c_334_n 0.00824124f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_160 N_VPWR_c_220_n N_Y_c_250_n 0.0323354f $X=2.835 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_215_n N_Y_c_250_n 0.026297f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_c_217_n N_Y_c_249_n 0.0491356f $X=0.3 $Y=1.985 $X2=0 $Y2=0
cc_163 A_131_368# N_Y_c_250_n 0.00148865f $X=0.655 $Y=1.84 $X2=1.21 $Y2=2.115
cc_164 A_131_368# N_Y_c_249_n 0.00121106f $X=0.655 $Y=1.84 $X2=1.005 $Y2=1.95
cc_165 N_Y_M1009_d N_A_27_74#_c_283_n 0.00723582f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_166 N_Y_c_248_n N_A_27_74#_c_283_n 0.0305034f $X=0.895 $Y=0.91 $X2=0 $Y2=0
cc_167 N_Y_c_248_n N_A_27_74#_c_286_n 0.00142263f $X=0.895 $Y=0.91 $X2=0 $Y2=0
cc_168 N_Y_c_249_n N_A_27_74#_c_286_n 0.00186133f $X=1.005 $Y=1.95 $X2=0 $Y2=0
cc_169 N_A_27_74#_c_285_n N_VGND_M1000_d 0.0048312f $X=2.38 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_27_74#_c_284_n N_VGND_c_328_n 0.00795492f $X=1.515 $Y=0.52 $X2=0
+ $Y2=0
cc_171 N_A_27_74#_c_285_n N_VGND_c_328_n 0.0228485f $X=2.38 $Y=1.095 $X2=0 $Y2=0
cc_172 N_A_27_74#_c_287_n N_VGND_c_328_n 0.031539f $X=2.545 $Y=0.515 $X2=0 $Y2=0
cc_173 N_A_27_74#_c_287_n N_VGND_c_330_n 0.0254897f $X=2.545 $Y=0.515 $X2=0
+ $Y2=0
cc_174 N_A_27_74#_c_283_n N_VGND_c_331_n 0.0358046f $X=1.35 $Y=0.435 $X2=0 $Y2=0
cc_175 N_A_27_74#_c_284_n N_VGND_c_331_n 0.0146502f $X=1.515 $Y=0.52 $X2=0 $Y2=0
cc_176 N_A_27_74#_c_288_n N_VGND_c_331_n 0.0146186f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_177 N_A_27_74#_c_287_n N_VGND_c_333_n 0.0144922f $X=2.545 $Y=0.515 $X2=0
+ $Y2=0
cc_178 N_A_27_74#_c_283_n N_VGND_c_334_n 0.0306817f $X=1.35 $Y=0.435 $X2=0 $Y2=0
cc_179 N_A_27_74#_c_284_n N_VGND_c_334_n 0.0120674f $X=1.515 $Y=0.52 $X2=0 $Y2=0
cc_180 N_A_27_74#_c_287_n N_VGND_c_334_n 0.0118826f $X=2.545 $Y=0.515 $X2=0
+ $Y2=0
cc_181 N_A_27_74#_c_288_n N_VGND_c_334_n 0.0120551f $X=0.28 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__and4_2.spice
* Created: Wed Sep  2 11:58:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4_2.pex.spice"
.subckt sky130_fd_sc_ms__and4_2  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_143_74# N_A_M1005_g N_A_56_74#_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1000 A_221_74# N_B_M1000_g A_143_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1011 A_335_74# N_C_M1011_g A_221_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75001.2
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_D_M1004_g A_335_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=7.296 NRS=25.128 M=1 R=4.93333 SA=75001.7
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1004_d N_A_56_74#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=15.396 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_56_74#_M1008_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2738 AS=0.1036 PD=2.22 PS=1.02 NRD=8.508 NRS=0 M=1 R=4.93333 SA=75002.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_A_56_74#_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.37 PD=1.27 PS=2.74 NRD=0 NRS=16.7253 M=1 R=5.55556 SA=90000.3
+ SB=90002.9 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_56_74#_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.24 AS=0.135 PD=1.48 PS=1.27 NRD=20.685 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1006 N_A_56_74#_M1006_d N_C_M1006_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.24 PD=1.27 PS=1.48 NRD=0 NRS=18.715 M=1 R=5.55556 SA=90001.4
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_D_M1007_g N_A_56_74#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.221698 AS=0.135 PD=1.4717 PS=1.27 NRD=15.7403 NRS=0 M=1 R=5.55556
+ SA=90001.8 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1009 N_X_M1009_d N_A_56_74#_M1009_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.248302 PD=1.39 PS=1.6483 NRD=0 NRS=14.0658 M=1 R=6.22222
+ SA=90002.2 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1010 N_X_M1009_d N_A_56_74#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.4368 PD=1.39 PS=3.02 NRD=0 NRS=15.8191 M=1 R=6.22222 SA=90002.7
+ SB=90000.3 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__and4_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfstp_4.spice
* Created: Wed Sep  2 12:03:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfstp_4.pex.spice"
.subckt sky130_fd_sc_ms__dfstp_4  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1032 N_VGND_M1032_d N_D_M1032_g N_A_27_74#_M1032_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_CLK_M1035_g N_A_225_74#_M1035_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_398_74#_M1018_d N_A_225_74#_M1018_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_612_74#_M1023_d N_A_225_74#_M1023_g N_A_27_74#_M1023_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0945 AS=0.18665 PD=0.87 PS=1.8 NRD=48.564 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1013 A_732_74# N_A_398_74#_M1013_g N_A_612_74#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0945 PD=0.66 PS=0.87 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_767_402#_M1003_g A_732_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.147 AS=0.0504 PD=1.54 PS=0.66 NRD=8.568 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1026 A_1035_118# N_A_612_74#_M1026_g N_A_767_402#_M1026_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1491 PD=0.66 PS=1.55 NRD=18.564 NRS=9.996 M=1 R=2.8
+ SA=75000.3 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_SET_B_M1016_g A_1035_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0930736 AS=0.0504 PD=0.832075 PS=0.66 NRD=37.848 NRS=18.564 M=1 R=2.8
+ SA=75000.7 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1028 A_1225_74# N_A_612_74#_M1028_g N_VGND_M1016_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1264 AS=0.141826 PD=1.035 PS=1.26792 NRD=26.712 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_1324_392#_M1006_d N_A_398_74#_M1006_g A_1225_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.127668 AS=0.1264 PD=1.20755 PS=1.035 NRD=0 NRS=26.712 M=1
+ R=4.26667 SA=75001.4 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1015 A_1436_88# N_A_225_74#_M1015_g N_A_1324_392#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0837821 PD=0.66 PS=0.792453 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75001.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1007 A_1514_88# N_A_1484_62#_M1007_g A_1436_88# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SET_B_M1004_g A_1514_88# VNB NLOWVT L=0.15 W=0.42
+ AD=0.21735 AS=0.0504 PD=1.455 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_A_1484_62#_M1005_d N_A_1324_392#_M1005_g N_VGND_M1004_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.21735 PD=1.41 PS=1.455 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75003.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_1324_392#_M1000_g N_A_1940_74#_M1000_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1295 AS=0.2627 PD=1.09 PS=2.19 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.3 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1008 N_Q_M1008_d N_A_1940_74#_M1008_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1009 N_Q_M1008_d N_A_1940_74#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=1.45 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_Q_M1017_d N_A_1940_74#_M1017_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.2627 PD=1.065 PS=1.45 NRD=7.296 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1034 N_Q_M1017_d N_A_1940_74#_M1034_g N_VGND_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.2627 PD=1.065 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1031 N_VPWR_M1031_d N_D_M1031_g N_A_27_74#_M1031_s VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_CLK_M1024_g N_A_225_74#_M1024_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1027 N_A_398_74#_M1027_d N_A_225_74#_M1027_g N_VPWR_M1024_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_612_74#_M1001_d N_A_398_74#_M1001_g N_A_27_74#_M1001_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90004.5 A=0.0756 P=1.2 MULT=1
MM1002 A_719_463# N_A_225_74#_M1002_g N_A_612_74#_M1001_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0672 PD=0.66 PS=0.74 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90004 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_767_402#_M1010_g A_719_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.15855 AS=0.0504 PD=1.175 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90003.6 A=0.0756 P=1.2 MULT=1
MM1038 N_A_767_402#_M1038_d N_A_612_74#_M1038_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.15855 PD=0.69 PS=1.175 NRD=0 NRS=218.099 M=1 R=2.33333
+ SA=90002 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_SET_B_M1011_g N_A_767_402#_M1038_d VPB PSHORT L=0.18
+ W=0.42 AD=0.109348 AS=0.0567 PD=0.908028 PS=0.69 NRD=107.877 NRS=0 M=1
+ R=2.33333 SA=90002.5 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1033 A_1223_347# N_A_612_74#_M1033_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.182187 AS=0.260352 PD=1.55 PS=2.16197 NRD=25.0387 NRS=4.9053 M=1
+ R=5.55556 SA=90001.4 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1025 N_A_1324_392#_M1025_d N_A_225_74#_M1025_g A_1223_347# VPB PSHORT L=0.18
+ W=1 AD=0.290141 AS=0.182187 PD=2.27465 PS=1.55 NRD=0 NRS=25.0387 M=1 R=5.55556
+ SA=90001.8 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1036 A_1483_508# N_A_398_74#_M1036_g N_A_1324_392#_M1025_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.121859 PD=0.66 PS=0.955352 NRD=30.4759 NRS=79.7259 M=1
+ R=2.33333 SA=90002.6 SB=90001 A=0.0756 P=1.2 MULT=1
MM1014 N_VPWR_M1014_d N_A_1484_62#_M1014_g A_1483_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.0504 PD=0.69 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90003
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1019 N_A_1324_392#_M1019_d N_SET_B_M1019_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90003.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1012 N_A_1484_62#_M1012_d N_A_1324_392#_M1012_g N_VPWR_M1012_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.1092 AS=0.1113 PD=1.36 PS=1.37 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1020 N_A_1940_74#_M1020_d N_A_1324_392#_M1020_g N_VPWR_M1020_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.2226 PD=1.11 PS=2.21 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1021 N_A_1940_74#_M1020_d N_A_1324_392#_M1021_g N_VPWR_M1021_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.1542 PD=1.11 PS=1.25143 NRD=0 NRS=15.2281 M=1
+ R=4.66667 SA=90000.6 SB=90002 A=0.1512 P=2.04 MULT=1
MM1022 N_Q_M1022_d N_A_1940_74#_M1022_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2056 PD=1.39 PS=1.66857 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.9
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1029 N_Q_M1022_d N_A_1940_74#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.4
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1030 N_Q_M1030_d N_A_1940_74#_M1030_g N_VPWR_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.8
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1037 N_Q_M1030_d N_A_1940_74#_M1037_g N_VPWR_M1037_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX39_noxref VNB VPB NWDIODE A=24.9216 P=30.61
c_142 VNB 0 7.64129e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dfstp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlxtn_2.pex.spice
* Created: Fri Aug 28 17:29:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLXTN_2%D 3 7 9 13 16
c29 3 0 1.87332e-19 $X=0.495 $Y=0.875
r30 15 16 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.655 $Y2=1.465
r31 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.495 $Y2=1.465
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r33 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r34 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.63
+ $X2=0.655 $Y2=1.465
r35 5 7 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.655 $Y=1.63
+ $X2=0.655 $Y2=2.54
r36 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r37 1 3 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%GATE_N 3 7 9 12
c44 12 0 1.38982e-19 $X=1.15 $Y=1.615
r45 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.615
+ $X2=1.15 $Y2=1.78
r46 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.615
+ $X2=1.15 $Y2=1.45
r47 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.615 $X2=1.15 $Y2=1.615
r48 7 15 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=1.205 $Y=2.54
+ $X2=1.205 $Y2=1.78
r49 3 14 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.085 $Y=0.78
+ $X2=1.085 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%A_232_82# 1 2 7 11 13 15 16 18 20 23 27 29
+ 33 35 39 40 43 46 47 48 50 52 53 58 60 61 64 65
c158 65 0 4.79549e-20 $X=4.185 $Y=1.65
c159 64 0 1.38828e-19 $X=4.185 $Y=1.65
c160 52 0 1.38982e-19 $X=1.43 $Y=2.265
c161 35 0 1.87332e-19 $X=1.485 $Y=1.045
c162 23 0 1.93416e-19 $X=3.88 $Y=2.725
r163 72 74 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.825 $Y=1.65
+ $X2=3.88 $Y2=1.65
r164 65 74 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=4.185 $Y=1.65
+ $X2=3.88 $Y2=1.65
r165 64 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=1.65
+ $X2=4.185 $Y2=1.815
r166 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.65 $X2=4.185 $Y2=1.65
r167 60 62 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.605
+ $X2=1.685 $Y2=1.77
r168 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.605 $X2=1.72 $Y2=1.605
r169 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=0.925 $X2=1.72 $Y2=0.925
r170 53 62 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.57 $Y=2.1
+ $X2=1.57 $Y2=1.77
r171 52 54 7.68295 $w=3.88e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=2.265
+ $X2=1.46 $Y2=2.525
r172 52 53 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=2.265
+ $X2=1.46 $Y2=2.1
r173 50 67 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.105 $Y=2.905
+ $X2=4.105 $Y2=1.815
r174 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=2.99
+ $X2=4.105 $Y2=2.905
r175 47 48 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=4.02 $Y=2.99
+ $X2=3.045 $Y2=2.99
r176 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.96 $Y=2.905
+ $X2=3.045 $Y2=2.99
r177 45 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=2.61
+ $X2=2.96 $Y2=2.905
r178 44 54 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.655 $Y=2.525
+ $X2=1.46 $Y2=2.525
r179 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.875 $Y=2.525
+ $X2=2.96 $Y2=2.61
r180 43 44 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=2.875 $Y=2.525
+ $X2=1.655 $Y2=2.525
r181 40 60 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.685 $Y=1.57
+ $X2=1.685 $Y2=1.605
r182 39 57 3.08538 $w=4e-07 $l=2.05e-07 $layer=LI1_cond $X=1.685 $Y=1.17
+ $X2=1.685 $Y2=0.965
r183 39 40 11.5244 $w=3.98e-07 $l=4e-07 $layer=LI1_cond $X=1.685 $Y=1.17
+ $X2=1.685 $Y2=1.57
r184 35 57 4.21417 $w=2.5e-07 $l=2.36643e-07 $layer=LI1_cond $X=1.485 $Y=1.045
+ $X2=1.685 $Y2=0.965
r185 35 37 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.485 $Y=1.045
+ $X2=1.3 $Y2=1.045
r186 31 33 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.605 $Y=1.185
+ $X2=3.825 $Y2=1.185
r187 26 61 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.72 $Y=1.335
+ $X2=1.72 $Y2=1.605
r188 26 27 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.72 $Y=1.335
+ $X2=1.72 $Y2=1.26
r189 25 58 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.72 $Y=1.185
+ $X2=1.72 $Y2=0.925
r190 25 27 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.72 $Y=1.185
+ $X2=1.72 $Y2=1.26
r191 21 74 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.88 $Y=1.815
+ $X2=3.88 $Y2=1.65
r192 21 23 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=3.88 $Y=1.815
+ $X2=3.88 $Y2=2.725
r193 20 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.485
+ $X2=3.825 $Y2=1.65
r194 19 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.825 $Y=1.26
+ $X2=3.825 $Y2=1.185
r195 19 20 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.825 $Y=1.26
+ $X2=3.825 $Y2=1.485
r196 16 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.605 $Y=1.11
+ $X2=3.605 $Y2=1.185
r197 16 18 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=1.11
+ $X2=3.605 $Y2=0.715
r198 13 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=1.26
r199 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.74
r200 9 29 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.215 $Y=1.26
+ $X2=2.355 $Y2=1.26
r201 9 11 406.202 $w=1.8e-07 $l=1.045e-06 $layer=POLY_cond $X=2.215 $Y=1.335
+ $X2=2.215 $Y2=2.38
r202 8 27 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.26
+ $X2=1.72 $Y2=1.26
r203 7 9 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.125 $Y=1.26 $X2=2.215
+ $Y2=1.26
r204 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.125 $Y=1.26
+ $X2=1.885 $Y2=1.26
r205 2 52 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.295
+ $Y=2.12 $X2=1.43 $Y2=2.265
r206 1 37 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.41 $X2=1.3 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%A_27_120# 1 2 7 9 11 13 15 18 21 22 25 26 27
+ 29 34 37 42
r114 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.465 $X2=2.805 $Y2=1.465
r115 39 42 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.56 $Y=1.465
+ $X2=2.805 $Y2=1.465
r116 33 34 8.09223 $w=5.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.855
+ $X2=0.795 $Y2=0.855
r117 31 33 9.35116 $w=5.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.855
+ $X2=0.71 $Y2=0.855
r118 29 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=1.3
+ $X2=2.56 $Y2=1.465
r119 28 29 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=1.3
r120 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=2.56 $Y2=0.425
r121 26 27 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=1.315 $Y2=0.34
r122 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.315 $Y2=0.34
r123 24 25 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.58
r124 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=0.665
+ $X2=1.23 $Y2=0.58
r125 22 34 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.145 $Y=0.665
+ $X2=0.795 $Y2=0.665
r126 21 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.71 $Y2=2.035
r127 20 33 7.75927 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=0.855
r128 20 21 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r129 16 37 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.43 $Y=2.035
+ $X2=0.71 $Y2=2.035
r130 16 18 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.43 $Y=2.12
+ $X2=0.43 $Y2=2.265
r131 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.215 $Y=1.11
+ $X2=3.215 $Y2=0.715
r132 12 43 48.5468 $w=2.78e-07 $l=3.52987e-07 $layer=POLY_cond $X=2.97 $Y=1.185
+ $X2=2.805 $Y2=1.465
r133 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.14 $Y=1.185
+ $X2=3.215 $Y2=1.11
r134 11 12 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.14 $Y=1.185
+ $X2=2.97 $Y2=1.185
r135 7 43 34.5863 $w=2.78e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.85 $Y=1.63
+ $X2=2.805 $Y2=1.465
r136 7 9 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=2.85 $Y=1.63 $X2=2.85
+ $Y2=2.46
r137 2 18 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=2.12 $X2=0.43 $Y2=2.265
r138 1 31 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.6 $X2=0.28 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%A_369_392# 1 2 9 13 16 18 19 22 24 25 31 32
+ 33 41
c105 41 0 1.38828e-19 $X=4.21 $Y=0.585
c106 31 0 4.79549e-20 $X=3.345 $Y=1.635
c107 24 0 6.89381e-20 $X=4.21 $Y=0.42
c108 22 0 3.15497e-20 $X=3.485 $Y=0.42
r109 32 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.635
+ $X2=3.345 $Y2=1.8
r110 31 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.345 $Y=1.635
+ $X2=3.345 $Y2=1.885
r111 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=1.635
+ $X2=3.345 $Y2=1.47
r112 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.635 $X2=3.345 $Y2=1.635
r113 28 29 6.58523 $w=3.52e-07 $l=1.9e-07 $layer=LI1_cond $X=1.99 $Y=2.035
+ $X2=2.18 $Y2=2.035
r114 25 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=0.42
+ $X2=4.21 $Y2=0.585
r115 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=0.42 $X2=4.21 $Y2=0.42
r116 22 24 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=3.485 $Y=0.42
+ $X2=4.21 $Y2=0.42
r117 20 22 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.4 $Y=0.585
+ $X2=3.485 $Y2=0.42
r118 20 33 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.4 $Y=0.585
+ $X2=3.4 $Y2=1.47
r119 19 29 7.60401 $w=3.52e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.305 $Y=1.885
+ $X2=2.18 $Y2=2.035
r120 18 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.885
+ $X2=3.345 $Y2=1.885
r121 18 19 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.18 $Y=1.885
+ $X2=2.305 $Y2=1.885
r122 14 29 2.74175 $w=2.5e-07 $l=2.35e-07 $layer=LI1_cond $X=2.18 $Y=1.8
+ $X2=2.18 $Y2=2.035
r123 14 16 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.18 $Y=1.8
+ $X2=2.18 $Y2=0.86
r124 13 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.3 $Y=0.905
+ $X2=4.3 $Y2=0.585
r125 9 38 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.27 $Y=2.46
+ $X2=3.27 $Y2=1.8
r126 2 28 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.105
r127 1 16 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.37 $X2=2.14 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%A_842_405# 1 2 9 13 17 21 25 29 31 34 36 41
+ 43 47 50 52 55 62 63 69
c101 52 0 1.98766e-19 $X=5.59 $Y=1.795
c102 13 0 6.89381e-20 $X=4.69 $Y=0.905
r103 61 62 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.502 $Y=0.955
+ $X2=5.502 $Y2=1.125
r104 59 60 7.83799 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.462 $Y=1.96
+ $X2=5.462 $Y2=2.19
r105 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.08
+ $Y=1.46 $X2=6.08 $Y2=1.46
r106 53 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.46
+ $X2=5.59 $Y2=1.46
r107 53 55 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.675 $Y=1.46
+ $X2=6.08 $Y2=1.46
r108 52 59 9.00471 $w=3.58e-07 $l=2.19875e-07 $layer=LI1_cond $X=5.59 $Y=1.795
+ $X2=5.462 $Y2=1.96
r109 51 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=1.625
+ $X2=5.59 $Y2=1.46
r110 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.59 $Y=1.625
+ $X2=5.59 $Y2=1.795
r111 50 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=5.59 $Y2=1.46
r112 50 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=5.59 $Y2=1.125
r113 47 61 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=5.455 $Y=0.52
+ $X2=5.455 $Y2=0.955
r114 41 60 5.71829 $w=3.58e-07 $l=1.87029e-07 $layer=LI1_cond $X=5.415 $Y=2.355
+ $X2=5.462 $Y2=2.19
r115 41 43 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.415 $Y=2.355
+ $X2=5.415 $Y2=2.79
r116 39 69 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.525 $Y=2.19
+ $X2=4.69 $Y2=2.19
r117 39 66 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.525 $Y=2.19
+ $X2=4.3 $Y2=2.19
r118 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.525
+ $Y=2.19 $X2=4.525 $Y2=2.19
r119 36 60 1.20828 $w=3.3e-07 $l=2.12e-07 $layer=LI1_cond $X=5.25 $Y=2.19
+ $X2=5.462 $Y2=2.19
r120 36 38 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=5.25 $Y=2.19
+ $X2=4.525 $Y2=2.19
r121 34 35 2.23839 $w=3.23e-07 $l=1.5e-08 $layer=POLY_cond $X=6.68 $Y=1.46
+ $X2=6.695 $Y2=1.46
r122 33 34 71.6285 $w=3.23e-07 $l=4.8e-07 $layer=POLY_cond $X=6.2 $Y=1.46
+ $X2=6.68 $Y2=1.46
r123 32 33 1.49226 $w=3.23e-07 $l=1e-08 $layer=POLY_cond $X=6.19 $Y=1.46 $X2=6.2
+ $Y2=1.46
r124 31 56 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.11 $Y=1.46 $X2=6.08
+ $Y2=1.46
r125 31 32 11.6848 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.11 $Y=1.46 $X2=6.19
+ $Y2=1.46
r126 27 35 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.625
+ $X2=6.695 $Y2=1.46
r127 27 29 301.25 $w=1.8e-07 $l=7.75e-07 $layer=POLY_cond $X=6.695 $Y=1.625
+ $X2=6.695 $Y2=2.4
r128 23 34 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.68 $Y=1.295
+ $X2=6.68 $Y2=1.46
r129 23 25 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.68 $Y=1.295
+ $X2=6.68 $Y2=0.74
r130 19 32 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.19 $Y=1.295
+ $X2=6.19 $Y2=1.46
r131 19 21 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.19 $Y=1.295
+ $X2=6.19 $Y2=0.74
r132 15 33 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.2 $Y=1.625
+ $X2=6.2 $Y2=1.46
r133 15 17 301.25 $w=1.8e-07 $l=7.75e-07 $layer=POLY_cond $X=6.2 $Y=1.625
+ $X2=6.2 $Y2=2.4
r134 11 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=2.025
+ $X2=4.69 $Y2=2.19
r135 11 13 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=4.69 $Y=2.025
+ $X2=4.69 $Y2=0.905
r136 7 66 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=2.355
+ $X2=4.3 $Y2=2.19
r137 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.3 $Y=2.355 $X2=4.3
+ $Y2=2.725
r138 2 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.815 $X2=5.415 $Y2=1.96
r139 2 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.815 $X2=5.415 $Y2=2.79
r140 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.275
+ $Y=0.375 $X2=5.415 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%A_672_392# 1 2 9 13 17 18 20 21 29
r74 29 32 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.17 $Y=1.46
+ $X2=5.17 $Y2=1.625
r75 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.17 $Y=1.46
+ $X2=5.17 $Y2=1.295
r76 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.17
+ $Y=1.46 $X2=5.17 $Y2=1.46
r77 20 21 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=2.225
+ $X2=3.59 $Y2=2.14
r78 18 25 14.0393 $w=3.24e-07 $l=3.77492e-07 $layer=LI1_cond $X=4.25 $Y=1.23
+ $X2=3.95 $Y2=1.055
r79 17 28 9.67586 $w=2.9e-07 $l=3.04072e-07 $layer=LI1_cond $X=4.99 $Y=1.23
+ $X2=5.162 $Y2=1.46
r80 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.99 $Y=1.23
+ $X2=4.25 $Y2=1.23
r81 15 25 6.96605 $w=3.24e-07 $l=1.85e-07 $layer=LI1_cond $X=3.765 $Y=1.055
+ $X2=3.95 $Y2=1.055
r82 15 21 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.765 $Y=1.055
+ $X2=3.765 $Y2=2.14
r83 13 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.2 $Y=0.745 $X2=5.2
+ $Y2=1.295
r84 9 32 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.19 $Y=2.375
+ $X2=5.19 $Y2=1.625
r85 2 20 300 $w=1.7e-07 $l=3.39522e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.96 $X2=3.53 $Y2=2.225
r86 1 25 182 $w=1.7e-07 $l=6.15366e-07 $layer=licon1_NDIFF $count=1 $X=3.68
+ $Y=0.395 $X2=3.95 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%VPWR 1 2 3 4 5 18 22 26 30 32 37 38 40 41 42
+ 48 64 69 74 77 80
c78 77 0 1.93416e-19 $X=5.08 $Y=3.02
r79 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r80 76 77 10.6911 $w=7.88e-07 $l=1.2e-07 $layer=LI1_cond $X=4.96 $Y=3.02
+ $X2=5.08 $Y2=3.02
r81 72 76 6.05609 $w=7.88e-07 $l=4e-07 $layer=LI1_cond $X=4.56 $Y=3.02 $X2=4.96
+ $Y2=3.02
r82 72 74 11.9023 $w=7.88e-07 $l=2e-07 $layer=LI1_cond $X=4.56 $Y=3.02 $X2=4.36
+ $Y2=3.02
r83 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 67 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r87 64 79 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=7.017 $Y2=3.33
r88 64 66 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 63 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r90 63 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 62 77 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=5.08 $Y2=3.33
r92 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 58 74 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=4.36 $Y2=3.33
r95 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 56 69 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.532 $Y2=3.33
r97 56 58 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r98 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r102 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 48 69 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.532 $Y2=3.33
r104 48 53 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r105 46 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 42 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 42 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 40 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 40 41 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.952 $Y2=3.33
r111 39 66 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 39 41 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=5.952 $Y2=3.33
r113 37 45 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.93 $Y2=3.33
r115 36 50 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r116 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.93 $Y2=3.33
r117 32 35 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=6.96 $Y=1.985
+ $X2=6.96 $Y2=2.815
r118 30 79 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=7.017 $Y2=3.33
r119 30 35 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=6.96 $Y2=2.815
r120 26 29 44.4897 $w=2.13e-07 $l=8.3e-07 $layer=LI1_cond $X=5.952 $Y=1.985
+ $X2=5.952 $Y2=2.815
r121 24 41 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.952 $Y=3.245
+ $X2=5.952 $Y2=3.33
r122 24 29 23.0489 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=5.952 $Y=3.245
+ $X2=5.952 $Y2=2.815
r123 20 69 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.532 $Y=3.245
+ $X2=2.532 $Y2=3.33
r124 20 22 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=2.532 $Y=3.245
+ $X2=2.532 $Y2=2.945
r125 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=3.33
r126 16 18 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=2.395
r127 5 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.84 $X2=6.92 $Y2=2.815
r128 5 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.84 $X2=6.92 $Y2=1.985
r129 4 29 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.975 $Y2=2.815
r130 4 26 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.975 $Y2=1.985
r131 3 76 300 $w=1.7e-07 $l=6.9401e-07 $layer=licon1_PDIFF $count=2 $X=4.39
+ $Y=2.515 $X2=4.96 $Y2=2.79
r132 2 22 600 $w=1.7e-07 $l=1.09172e-06 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.96 $X2=2.53 $Y2=2.945
r133 1 18 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=0.745
+ $Y=2.12 $X2=0.93 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%Q 1 2 9 13 14 15 16 29 31
r23 21 31 2.21269 $w=3.73e-07 $l=7.2e-08 $layer=LI1_cond $X=6.447 $Y=2.107
+ $X2=6.447 $Y2=2.035
r24 15 16 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=6.447 $Y=2.405
+ $X2=6.447 $Y2=2.775
r25 14 31 0.215123 $w=3.73e-07 $l=7e-09 $layer=LI1_cond $X=6.447 $Y=2.028
+ $X2=6.447 $Y2=2.035
r26 14 29 6.80275 $w=3.73e-07 $l=1.08e-07 $layer=LI1_cond $X=6.447 $Y=2.028
+ $X2=6.447 $Y2=1.92
r27 14 15 8.97369 $w=3.73e-07 $l=2.92e-07 $layer=LI1_cond $X=6.447 $Y=2.113
+ $X2=6.447 $Y2=2.405
r28 14 21 0.184391 $w=3.73e-07 $l=6e-09 $layer=LI1_cond $X=6.447 $Y=2.113
+ $X2=6.447 $Y2=2.107
r29 13 29 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.5 $Y=1.125
+ $X2=6.5 $Y2=1.92
r30 7 13 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=6.452 $Y=0.993
+ $X2=6.452 $Y2=1.125
r31 7 9 20.7875 $w=2.63e-07 $l=4.78e-07 $layer=LI1_cond $X=6.452 $Y=0.993
+ $X2=6.452 $Y2=0.515
r32 2 31 600 $w=1.7e-07 $l=3.1305e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.445 $Y2=2.085
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.265
+ $Y=0.37 $X2=6.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTN_2%VGND 1 2 3 4 5 18 22 28 30 32 34 36 41 49 54
+ 59 66 72 75 78 82
r85 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r86 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r87 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r88 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r89 66 69 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r90 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r92 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r93 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 60 78 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=5.992
+ $Y2=0
r95 60 62 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.48
+ $Y2=0
r96 59 81 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r97 59 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r98 58 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r99 58 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r100 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r101 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.985
+ $Y2=0
r102 55 57 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.52
+ $Y2=0
r103 54 78 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=5.845 $Y=0
+ $X2=5.992 $Y2=0
r104 54 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=0
+ $X2=5.52 $Y2=0
r105 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r106 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r107 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=2.98
+ $Y2=0
r108 50 52 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.145 $Y=0
+ $X2=4.56 $Y2=0
r109 49 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.985
+ $Y2=0
r110 49 52 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.56
+ $Y2=0
r111 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r112 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r113 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r114 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r115 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r116 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 42 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r118 42 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r119 41 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.98
+ $Y2=0
r120 41 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=0
+ $X2=2.64 $Y2=0
r121 39 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 36 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r124 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r125 34 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r126 34 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r127 30 81 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r128 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r129 26 78 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.992 $Y=0.085
+ $X2=5.992 $Y2=0
r130 26 28 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=5.992 $Y=0.085
+ $X2=5.992 $Y2=0.515
r131 22 24 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.985 $Y=0.515
+ $X2=4.985 $Y2=0.89
r132 20 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0
r133 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0.515
r134 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0
r135 16 18 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0.54
r136 5 32 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.37 $X2=6.92 $Y2=0.515
r137 4 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.83
+ $Y=0.37 $X2=5.975 $Y2=0.515
r138 3 24 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.695 $X2=4.985 $Y2=0.89
r139 3 22 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.695 $X2=4.985 $Y2=0.515
r140 2 18 91 $w=1.7e-07 $l=6.29285e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.37 $X2=2.98 $Y2=0.54
r141 1 69 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.6 $X2=0.79 $Y2=0.325
.ends


* File: sky130_fd_sc_ms__a21oi_1.pxi.spice
* Created: Fri Aug 28 16:59:52 2020
* 
x_PM_SKY130_FD_SC_MS__A21OI_1%A2 N_A2_M1003_g N_A2_c_40_n N_A2_M1005_g A2
+ N_A2_c_42_n PM_SKY130_FD_SC_MS__A21OI_1%A2
x_PM_SKY130_FD_SC_MS__A21OI_1%A1 N_A1_M1002_g N_A1_M1000_g A1 N_A1_c_65_n
+ N_A1_c_66_n PM_SKY130_FD_SC_MS__A21OI_1%A1
x_PM_SKY130_FD_SC_MS__A21OI_1%B1 N_B1_c_101_n N_B1_M1004_g N_B1_M1001_g B1
+ N_B1_c_104_n PM_SKY130_FD_SC_MS__A21OI_1%B1
x_PM_SKY130_FD_SC_MS__A21OI_1%A_29_368# N_A_29_368#_M1003_s N_A_29_368#_M1000_d
+ N_A_29_368#_c_130_n N_A_29_368#_c_131_n N_A_29_368#_c_137_n
+ N_A_29_368#_c_132_n PM_SKY130_FD_SC_MS__A21OI_1%A_29_368#
x_PM_SKY130_FD_SC_MS__A21OI_1%VPWR N_VPWR_M1003_d N_VPWR_c_156_n VPWR
+ N_VPWR_c_157_n N_VPWR_c_158_n N_VPWR_c_155_n N_VPWR_c_160_n
+ PM_SKY130_FD_SC_MS__A21OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A21OI_1%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_180_n N_Y_c_181_n
+ N_Y_c_184_n N_Y_c_185_n N_Y_c_182_n Y Y Y PM_SKY130_FD_SC_MS__A21OI_1%Y
x_PM_SKY130_FD_SC_MS__A21OI_1%VGND N_VGND_M1005_s N_VGND_M1004_d N_VGND_c_219_n
+ N_VGND_c_220_n N_VGND_c_221_n N_VGND_c_222_n VGND N_VGND_c_223_n
+ N_VGND_c_224_n PM_SKY130_FD_SC_MS__A21OI_1%VGND
cc_1 VNB N_A2_M1003_g 0.00908106f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A2_c_40_n 0.0204319f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_3 VNB A2 0.00894107f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A2_c_42_n 0.05777f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.385
cc_5 VNB N_A1_M1002_g 0.0248365f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_A1_c_65_n 0.0237158f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_7 VNB N_A1_c_66_n 0.00959608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_101_n 0.0209416f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.55
cc_9 VNB N_B1_M1001_g 0.00842224f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_10 VNB B1 0.00662327f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_B1_c_104_n 0.0580426f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_12 VNB N_VPWR_c_155_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_180_n 0.00320135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_181_n 0.0035645f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_15 VNB N_Y_c_182_n 0.00543429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_219_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_17 VNB N_VGND_c_220_n 0.0350088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_221_n 0.0107718f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_19 VNB N_VGND_c_222_n 0.0358154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_223_n 0.0319078f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_21 VNB N_VGND_c_224_n 0.146074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A2_M1003_g 0.0310996f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_23 VPB N_A1_M1000_g 0.0213465f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_24 VPB N_A1_c_65_n 0.00548342f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_25 VPB N_A1_c_66_n 0.00399982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_26 VPB N_B1_M1001_g 0.0285034f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_27 VPB N_A_29_368#_c_130_n 0.0190505f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_28 VPB N_A_29_368#_c_131_n 0.0314181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_A_29_368#_c_132_n 0.00242978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_156_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_31 VPB N_VPWR_c_157_n 0.0178349f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_32 VPB N_VPWR_c_158_n 0.0302175f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_33 VPB N_VPWR_c_155_n 0.0531649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_160_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_Y_c_181_n 3.49014e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_36 VPB N_Y_c_184_n 0.00934184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_Y_c_185_n 0.00103426f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_38 VPB Y 0.0431963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 N_A2_c_40_n N_A1_M1002_g 0.0428551f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_40 A2 N_A1_M1002_g 6.23327e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 N_A2_M1003_g N_A1_M1000_g 0.030344f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_42 N_A2_c_42_n N_A1_c_65_n 0.0428551f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_43 A2 N_A1_c_66_n 0.0162065f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A2_c_42_n N_A1_c_66_n 0.00847156f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_45 N_A2_M1003_g N_A_29_368#_c_130_n 0.00674321f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_46 A2 N_A_29_368#_c_130_n 0.0195989f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A2_c_42_n N_A_29_368#_c_130_n 0.00223475f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_48 N_A2_M1003_g N_A_29_368#_c_131_n 0.00101635f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_49 N_A2_M1003_g N_A_29_368#_c_137_n 0.0197181f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_50 N_A2_M1003_g N_VPWR_c_156_n 0.0128939f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_51 N_A2_M1003_g N_VPWR_c_157_n 0.0050621f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_52 N_A2_M1003_g N_VPWR_c_155_n 0.0100258f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_53 N_A2_c_40_n N_Y_c_180_n 0.0026419f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_54 N_A2_c_40_n N_VGND_c_220_n 0.0167319f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_55 A2 N_VGND_c_220_n 0.024157f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A2_c_42_n N_VGND_c_220_n 0.00199226f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_57 N_A2_c_40_n N_VGND_c_223_n 0.00383152f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A2_c_40_n N_VGND_c_224_n 0.0075694f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_59 N_A1_M1002_g N_B1_c_101_n 0.0197297f $X=0.87 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_60 N_A1_M1000_g N_B1_M1001_g 0.0304799f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A1_c_65_n N_B1_c_104_n 0.0204028f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_62 N_A1_c_66_n N_B1_c_104_n 3.9345e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_63 N_A1_M1000_g N_A_29_368#_c_130_n 7.78664e-19 $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_64 N_A1_c_66_n N_A_29_368#_c_137_n 0.014876f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_65 N_A1_M1000_g N_A_29_368#_c_132_n 0.0197005f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A1_c_65_n N_A_29_368#_c_132_n 0.00103037f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_67 N_A1_c_66_n N_A_29_368#_c_132_n 0.0111874f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_68 N_A1_M1000_g N_VPWR_c_156_n 0.00995356f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A1_M1000_g N_VPWR_c_158_n 0.0050621f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A1_M1000_g N_VPWR_c_155_n 0.00998985f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_71 N_A1_M1002_g N_Y_c_180_n 0.0117918f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A1_M1002_g N_Y_c_181_n 0.00323848f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A1_M1000_g N_Y_c_181_n 2.2305e-19 $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_74 N_A1_c_65_n N_Y_c_181_n 0.0020371f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_75 N_A1_c_66_n N_Y_c_181_n 0.0284379f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A1_M1000_g N_Y_c_185_n 0.00338076f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A1_c_66_n N_Y_c_185_n 0.00504905f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A1_M1002_g N_Y_c_182_n 0.00444011f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_79 N_A1_c_65_n N_Y_c_182_n 0.00625244f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A1_c_66_n N_Y_c_182_n 0.0109718f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A1_M1002_g N_VGND_c_220_n 0.00236525f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_82 N_A1_M1002_g N_VGND_c_223_n 0.00434272f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A1_M1002_g N_VGND_c_224_n 0.00821699f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B1_M1001_g N_A_29_368#_c_132_n 0.0145067f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_85 N_B1_M1001_g N_VPWR_c_156_n 7.62978e-19 $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_86 N_B1_M1001_g N_VPWR_c_158_n 0.005209f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_87 N_B1_M1001_g N_VPWR_c_155_n 0.00987181f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_88 N_B1_c_101_n N_Y_c_180_n 0.0038671f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_89 N_B1_c_101_n N_Y_c_181_n 0.00108982f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_90 N_B1_M1001_g N_Y_c_181_n 0.00810997f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_91 B1 N_Y_c_181_n 0.0252697f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_92 N_B1_c_104_n N_Y_c_181_n 0.00827951f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_93 N_B1_M1001_g N_Y_c_184_n 0.0151829f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_94 B1 N_Y_c_184_n 0.0212273f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B1_c_104_n N_Y_c_184_n 0.00369882f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_96 N_B1_M1001_g N_Y_c_185_n 0.00362788f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_97 N_B1_c_101_n N_Y_c_182_n 0.0131024f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_98 N_B1_M1001_g Y 0.00147311f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_99 N_B1_c_101_n N_VGND_c_222_n 0.0075574f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_100 B1 N_VGND_c_222_n 0.0200189f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B1_c_104_n N_VGND_c_222_n 0.00166151f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_102 N_B1_c_101_n N_VGND_c_223_n 0.00461464f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_103 N_B1_c_101_n N_VGND_c_224_n 0.00913518f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_104 N_A_29_368#_c_137_n N_VPWR_M1003_d 0.00410339f $X=0.833 $Y=2.107
+ $X2=-0.19 $Y2=1.66
cc_105 N_A_29_368#_c_131_n N_VPWR_c_156_n 0.0225402f $X=0.27 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_29_368#_c_137_n N_VPWR_c_156_n 0.0165663f $X=0.833 $Y=2.107 $X2=0
+ $Y2=0
cc_107 N_A_29_368#_c_132_n N_VPWR_c_156_n 0.0235977f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_108 N_A_29_368#_c_131_n N_VPWR_c_157_n 0.0130739f $X=0.27 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_29_368#_c_132_n N_VPWR_c_158_n 0.0129872f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_110 N_A_29_368#_c_131_n N_VPWR_c_155_n 0.0108215f $X=0.27 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_29_368#_c_132_n N_VPWR_c_155_n 0.0106816f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_112 N_A_29_368#_M1000_d N_Y_c_185_n 0.00130971f $X=1.065 $Y=1.84 $X2=0 $Y2=0
cc_113 N_A_29_368#_c_132_n N_Y_c_185_n 0.00772658f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_114 N_A_29_368#_c_132_n Y 0.024932f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_115 N_VPWR_c_158_n Y 0.011066f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_c_155_n Y 0.00915947f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_117 N_Y_c_180_n N_VGND_c_220_n 0.0222599f $X=1.105 $Y=0.515 $X2=0 $Y2=0
cc_118 N_Y_c_180_n N_VGND_c_222_n 0.0184459f $X=1.105 $Y=0.515 $X2=0 $Y2=0
cc_119 N_Y_c_182_n N_VGND_c_222_n 7.76044e-19 $X=1.155 $Y=1.18 $X2=0 $Y2=0
cc_120 N_Y_c_180_n N_VGND_c_223_n 0.0163488f $X=1.105 $Y=0.515 $X2=0 $Y2=0
cc_121 N_Y_c_180_n N_VGND_c_224_n 0.0134757f $X=1.105 $Y=0.515 $X2=0 $Y2=0

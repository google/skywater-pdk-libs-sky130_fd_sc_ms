* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A1 a_280_107# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_280_107# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_131_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y B1 a_131_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_280_107# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR A2 a_131_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VPWR A1 a_131_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_131_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND A2 a_280_107# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_131_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o221ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o221ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.210000 1.260000 6.575000 1.590000 ;
        RECT 6.405000 1.090000 8.455000 1.260000 ;
        RECT 8.285000 1.260000 9.955000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.430000 8.035000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.350000 3.555000 1.710000 ;
        RECT 2.545000 1.710000 6.000000 1.880000 ;
        RECT 5.405000 1.350000 6.000000 1.710000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.185000 1.180000 5.195000 1.540000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.405000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.312800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 1.010000 ;
        RECT 0.545000 1.010000 1.745000 1.180000 ;
        RECT 0.565000 1.950000 1.825000 2.050000 ;
        RECT 0.565000 2.050000 8.160000 2.120000 ;
        RECT 0.565000 2.120000 0.895000 2.980000 ;
        RECT 1.405000 0.595000 1.745000 1.010000 ;
        RECT 1.575000 1.180000 1.745000 1.820000 ;
        RECT 1.575000 1.820000 1.825000 1.950000 ;
        RECT 1.575000 2.120000 7.260000 2.220000 ;
        RECT 1.575000 2.220000 1.825000 2.980000 ;
        RECT 4.055000 2.220000 4.225000 2.735000 ;
        RECT 4.925000 2.220000 5.255000 2.735000 ;
        RECT 6.845000 1.950000 8.160000 2.050000 ;
        RECT 6.845000 2.220000 7.260000 2.520000 ;
        RECT 6.930000 2.520000 7.260000 2.735000 ;
        RECT 7.830000 2.120000 8.160000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.255000  2.165000 0.425000 ;
      RECT 0.115000  0.425000  0.375000 1.180000 ;
      RECT 0.115000  1.950000  0.365000 3.245000 ;
      RECT 1.045000  0.425000  1.235000 0.840000 ;
      RECT 1.065000  2.290000  1.395000 3.245000 ;
      RECT 1.915000  0.425000  2.165000 0.770000 ;
      RECT 1.915000  0.770000  3.155000 1.010000 ;
      RECT 1.915000  1.010000  4.015000 1.180000 ;
      RECT 2.025000  2.390000  2.355000 3.245000 ;
      RECT 2.395000  0.350000  6.235000 0.600000 ;
      RECT 2.525000  2.390000  3.855000 2.560000 ;
      RECT 2.525000  2.560000  2.855000 2.980000 ;
      RECT 3.025000  2.730000  3.355000 3.245000 ;
      RECT 3.335000  0.600000  3.505000 0.840000 ;
      RECT 3.525000  2.560000  3.855000 2.905000 ;
      RECT 3.525000  2.905000  5.755000 3.075000 ;
      RECT 3.685000  0.770000  5.735000 1.010000 ;
      RECT 4.425000  2.390000  4.755000 2.905000 ;
      RECT 5.405000  1.010000  5.735000 1.050000 ;
      RECT 5.425000  2.390000  5.755000 2.905000 ;
      RECT 5.905000  0.600000  6.235000 0.750000 ;
      RECT 5.905000  0.750000  9.025000 0.920000 ;
      RECT 5.905000  0.920000  6.235000 1.090000 ;
      RECT 5.925000  2.390000  6.255000 3.245000 ;
      RECT 6.405000  0.085000  6.735000 0.580000 ;
      RECT 6.425000  2.650000  6.675000 2.730000 ;
      RECT 6.425000  2.730000  6.760000 2.905000 ;
      RECT 6.425000  2.905000  8.530000 3.075000 ;
      RECT 6.905000  0.350000  7.155000 0.750000 ;
      RECT 7.335000  0.085000  7.665000 0.580000 ;
      RECT 7.460000  2.290000  7.630000 2.905000 ;
      RECT 7.835000  0.350000  8.085000 0.750000 ;
      RECT 8.265000  0.085000  8.605000 0.580000 ;
      RECT 8.360000  1.950000  9.510000 2.120000 ;
      RECT 8.360000  2.120000  8.530000 2.905000 ;
      RECT 8.730000  2.290000  8.980000 3.245000 ;
      RECT 8.775000  0.350000  9.025000 0.750000 ;
      RECT 8.775000  0.920000  9.965000 1.090000 ;
      RECT 9.180000  2.120000  9.510000 2.980000 ;
      RECT 9.205000  0.085000  9.535000 0.750000 ;
      RECT 9.710000  1.950000  9.960000 3.245000 ;
      RECT 9.715000  0.350000  9.965000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_ms__o221ai_4
END LIBRARY

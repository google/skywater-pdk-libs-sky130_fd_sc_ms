* File: sky130_fd_sc_ms__a311oi_2.pxi.spice
* Created: Wed Sep  2 11:54:49 2020
* 
x_PM_SKY130_FD_SC_MS__A311OI_2%A3 N_A3_M1016_g N_A3_c_92_n N_A3_M1009_g
+ N_A3_c_93_n N_A3_M1010_g N_A3_M1017_g A3 N_A3_c_96_n
+ PM_SKY130_FD_SC_MS__A311OI_2%A3
x_PM_SKY130_FD_SC_MS__A311OI_2%A2 N_A2_c_132_n N_A2_M1008_g N_A2_M1001_g
+ N_A2_c_134_n N_A2_M1013_g N_A2_M1003_g N_A2_c_136_n A2 N_A2_c_137_n
+ N_A2_c_138_n PM_SKY130_FD_SC_MS__A311OI_2%A2
x_PM_SKY130_FD_SC_MS__A311OI_2%A1 N_A1_M1002_g N_A1_M1004_g N_A1_M1011_g
+ N_A1_M1015_g N_A1_c_190_n A1 N_A1_c_191_n PM_SKY130_FD_SC_MS__A311OI_2%A1
x_PM_SKY130_FD_SC_MS__A311OI_2%B1 N_B1_M1014_g N_B1_M1005_g N_B1_M1006_g B1 B1
+ B1 N_B1_c_244_n PM_SKY130_FD_SC_MS__A311OI_2%B1
x_PM_SKY130_FD_SC_MS__A311OI_2%C1 N_C1_M1000_g N_C1_M1007_g N_C1_M1012_g C1
+ N_C1_c_292_n N_C1_c_293_n PM_SKY130_FD_SC_MS__A311OI_2%C1
x_PM_SKY130_FD_SC_MS__A311OI_2%VPWR N_VPWR_M1016_s N_VPWR_M1017_s N_VPWR_M1003_s
+ N_VPWR_M1004_s N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n
+ N_VPWR_c_335_n N_VPWR_c_336_n VPWR N_VPWR_c_337_n N_VPWR_c_338_n
+ N_VPWR_c_339_n N_VPWR_c_330_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n
+ PM_SKY130_FD_SC_MS__A311OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A311OI_2%A_130_368# N_A_130_368#_M1016_d
+ N_A_130_368#_M1001_d N_A_130_368#_M1002_d N_A_130_368#_M1005_d
+ N_A_130_368#_c_402_n N_A_130_368#_c_403_n N_A_130_368#_c_404_n
+ N_A_130_368#_c_405_n N_A_130_368#_c_406_n N_A_130_368#_c_407_n
+ N_A_130_368#_c_408_n N_A_130_368#_c_409_n N_A_130_368#_c_410_n
+ N_A_130_368#_c_445_n PM_SKY130_FD_SC_MS__A311OI_2%A_130_368#
x_PM_SKY130_FD_SC_MS__A311OI_2%A_692_368# N_A_692_368#_M1005_s
+ N_A_692_368#_M1006_s N_A_692_368#_M1012_s N_A_692_368#_c_471_n
+ N_A_692_368#_c_472_n N_A_692_368#_c_473_n N_A_692_368#_c_484_n
+ N_A_692_368#_c_474_n N_A_692_368#_c_475_n N_A_692_368#_c_476_n
+ PM_SKY130_FD_SC_MS__A311OI_2%A_692_368#
x_PM_SKY130_FD_SC_MS__A311OI_2%Y N_Y_M1011_d N_Y_M1015_d N_Y_M1000_d N_Y_M1007_d
+ N_Y_c_515_n N_Y_c_516_n N_Y_c_521_n N_Y_c_517_n N_Y_c_539_n Y Y Y N_Y_c_520_n
+ PM_SKY130_FD_SC_MS__A311OI_2%Y
x_PM_SKY130_FD_SC_MS__A311OI_2%A_45_74# N_A_45_74#_M1009_d N_A_45_74#_M1010_d
+ N_A_45_74#_M1013_d N_A_45_74#_c_568_n N_A_45_74#_c_573_n N_A_45_74#_c_569_n
+ N_A_45_74#_c_570_n N_A_45_74#_c_579_n N_A_45_74#_c_571_n N_A_45_74#_c_583_n
+ PM_SKY130_FD_SC_MS__A311OI_2%A_45_74#
x_PM_SKY130_FD_SC_MS__A311OI_2%VGND N_VGND_M1009_s N_VGND_M1014_d N_VGND_c_603_n
+ N_VGND_c_604_n VGND N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n
+ N_VGND_c_608_n N_VGND_c_609_n N_VGND_c_610_n PM_SKY130_FD_SC_MS__A311OI_2%VGND
x_PM_SKY130_FD_SC_MS__A311OI_2%A_300_74# N_A_300_74#_M1008_s N_A_300_74#_M1011_s
+ N_A_300_74#_c_653_n N_A_300_74#_c_654_n PM_SKY130_FD_SC_MS__A311OI_2%A_300_74#
cc_1 VNB N_A3_M1016_g 0.00916985f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.4
cc_2 VNB N_A3_c_92_n 0.022852f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_3 VNB N_A3_c_93_n 0.0168728f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_4 VNB N_A3_M1017_g 0.00104571f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_5 VNB A3 0.0155644f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A3_c_96_n 0.0488463f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.43
cc_7 VNB N_A2_c_132_n 0.0174681f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.55
cc_8 VNB N_A2_M1001_g 0.00599907f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_9 VNB N_A2_c_134_n 0.022624f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.22
cc_10 VNB N_A2_M1003_g 0.0061241f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_11 VNB N_A2_c_136_n 0.00595132f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_12 VNB N_A2_c_137_n 0.0464088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_138_n 0.00814841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_M1011_g 0.0285804f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.64
cc_15 VNB N_A1_M1015_g 0.0236097f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A1_c_190_n 0.003533f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.43
cc_17 VNB N_A1_c_191_n 0.0812203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_M1014_g 0.0281458f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.4
cc_19 VNB B1 0.00612637f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_B1_c_244_n 0.0434029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C1_M1000_g 0.0346834f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.4
cc_22 VNB N_C1_c_292_n 0.00305603f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_23 VNB N_C1_c_293_n 0.0487634f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_24 VNB N_VPWR_c_330_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_515_n 0.0126151f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_26 VNB N_Y_c_516_n 0.00206055f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.43
cc_27 VNB N_Y_c_517_n 0.00198283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.0734368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB Y 0.0265258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_520_n 0.00555748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_45_74#_c_568_n 0.0207156f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_32 VNB N_A_45_74#_c_569_n 0.0102706f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_33 VNB N_A_45_74#_c_570_n 0.00216743f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.43
cc_34 VNB N_A_45_74#_c_571_n 0.00469816f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.295
cc_35 VNB N_VGND_c_603_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_36 VNB N_VGND_c_604_n 0.0127126f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_37 VNB N_VGND_c_605_n 0.0196185f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.43
cc_38 VNB N_VGND_c_606_n 0.0766417f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.43
cc_39 VNB N_VGND_c_607_n 0.0343549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_608_n 0.323383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_609_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_610_n 0.0115409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_300_74#_c_653_n 0.002374f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_44 VNB N_A_300_74#_c_654_n 0.0263182f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_45 VPB N_A3_M1016_g 0.0276728f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=2.4
cc_46 VPB N_A3_M1017_g 0.0217377f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_47 VPB N_A2_M1001_g 0.0217377f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_48 VPB N_A2_M1003_g 0.0220915f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_49 VPB N_A1_M1002_g 0.0201072f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=2.4
cc_50 VPB N_A1_M1004_g 0.025668f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_51 VPB N_A1_c_190_n 0.00380343f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.43
cc_52 VPB N_A1_c_191_n 0.0125306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_B1_M1005_g 0.0250818f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_54 VPB N_B1_M1006_g 0.0197821f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.64
cc_55 VPB B1 0.00974621f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_56 VPB N_B1_c_244_n 0.00573543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_C1_M1007_g 0.0201623f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_58 VPB N_C1_M1012_g 0.023109f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.64
cc_59 VPB N_C1_c_292_n 0.00262436f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_60 VPB N_C1_c_293_n 0.00646983f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_61 VPB N_VPWR_c_331_n 0.0124065f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_62 VPB N_VPWR_c_332_n 0.0653866f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_63 VPB N_VPWR_c_333_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.43
cc_64 VPB N_VPWR_c_334_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.43
cc_65 VPB N_VPWR_c_335_n 0.00520669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_336_n 0.0119204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_337_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_338_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_339_n 0.0619448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_330_n 0.0872843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_341_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_342_n 0.00516566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_343_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_130_368#_c_402_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_75 VPB N_A_130_368#_c_403_n 0.00242893f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.43
cc_76 VPB N_A_130_368#_c_404_n 0.00490377f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.385
cc_77 VPB N_A_130_368#_c_405_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.43
cc_78 VPB N_A_130_368#_c_406_n 0.0059024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_130_368#_c_407_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_130_368#_c_408_n 0.0125008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_130_368#_c_409_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_130_368#_c_410_n 0.00241466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_692_368#_c_471_n 0.00583913f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_84 VPB N_A_692_368#_c_472_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_692_368#_c_473_n 0.00405878f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_86 VPB N_A_692_368#_c_474_n 0.0116218f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.43
cc_87 VPB N_A_692_368#_c_475_n 0.0241341f $X=-0.19 $Y=1.66 $X2=0.652 $Y2=1.385
cc_88 VPB N_A_692_368#_c_476_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_Y_c_521_n 0.011537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB Y 0.0136452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 N_A3_c_93_n N_A2_c_132_n 0.0103348f $X=0.995 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_92 N_A3_c_96_n N_A2_M1001_g 0.0358562f $X=0.995 $Y=1.43 $X2=0 $Y2=0
cc_93 A3 N_A2_c_137_n 2.0669e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A3_c_96_n N_A2_c_137_n 0.0176201f $X=0.995 $Y=1.43 $X2=0 $Y2=0
cc_95 N_A3_c_93_n N_A2_c_138_n 0.00444493f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_96 A3 N_A2_c_138_n 0.0233695f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A3_c_96_n N_A2_c_138_n 4.92803e-19 $X=0.995 $Y=1.43 $X2=0 $Y2=0
cc_98 N_A3_M1016_g N_VPWR_c_332_n 0.00649184f $X=0.56 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A3_M1016_g N_VPWR_c_333_n 0.005209f $X=0.56 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A3_M1017_g N_VPWR_c_333_n 0.005209f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A3_M1017_g N_VPWR_c_334_n 0.00363491f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A3_M1016_g N_VPWR_c_330_n 0.00986184f $X=0.56 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A3_M1017_g N_VPWR_c_330_n 0.00982376f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A3_M1016_g N_A_130_368#_c_402_n 0.014728f $X=0.56 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A3_M1017_g N_A_130_368#_c_402_n 0.0152527f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A3_M1017_g N_A_130_368#_c_403_n 0.0168394f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A3_M1016_g N_A_130_368#_c_404_n 0.00749011f $X=0.56 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A3_M1017_g N_A_130_368#_c_404_n 0.00341009f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_109 A3 N_A_130_368#_c_404_n 0.0182301f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A3_c_96_n N_A_130_368#_c_404_n 7.12326e-19 $X=0.995 $Y=1.43 $X2=0 $Y2=0
cc_111 N_A3_M1017_g N_A_130_368#_c_405_n 7.23242e-19 $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A3_c_92_n N_A_45_74#_c_568_n 4.43891e-19 $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A3_c_92_n N_A_45_74#_c_573_n 0.00979433f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A3_c_93_n N_A_45_74#_c_573_n 0.014168f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_115 A3 N_A_45_74#_c_573_n 0.0234443f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A3_c_96_n N_A_45_74#_c_573_n 6.29572e-19 $X=0.995 $Y=1.43 $X2=0 $Y2=0
cc_117 N_A3_c_93_n N_A_45_74#_c_570_n 2.82517e-19 $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_118 N_A3_c_92_n N_VGND_c_603_n 0.010528f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_119 N_A3_c_93_n N_VGND_c_603_n 0.00755236f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A3_c_92_n N_VGND_c_605_n 0.00383152f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_121 N_A3_c_93_n N_VGND_c_606_n 0.00383152f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A3_c_92_n N_VGND_c_608_n 0.00387841f $X=0.565 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A3_c_93_n N_VGND_c_608_n 0.00384065f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_124 N_A2_c_136_n N_A1_c_190_n 0.0139406f $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A2_c_137_n N_A1_c_190_n 2.46355e-19 $X=1.91 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A2_M1003_g N_A1_c_191_n 0.0338081f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A2_c_136_n N_A1_c_191_n 6.33995e-19 $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A2_c_137_n N_A1_c_191_n 0.0164469f $X=1.91 $Y=1.385 $X2=0 $Y2=0
cc_129 N_A2_M1001_g N_VPWR_c_334_n 0.00363491f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A2_M1003_g N_VPWR_c_335_n 0.00403758f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A2_M1001_g N_VPWR_c_337_n 0.005209f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A2_M1003_g N_VPWR_c_337_n 0.005209f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A2_M1001_g N_VPWR_c_330_n 0.00982376f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_VPWR_c_330_n 0.00982655f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A2_M1001_g N_A_130_368#_c_402_n 7.23242e-19 $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A2_M1001_g N_A_130_368#_c_403_n 0.0128923f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A2_c_138_n N_A_130_368#_c_403_n 0.0333429f $X=1.315 $Y=1.365 $X2=0
+ $Y2=0
cc_138 N_A2_M1001_g N_A_130_368#_c_405_n 0.0152527f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A2_M1003_g N_A_130_368#_c_405_n 0.0153709f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A2_M1003_g N_A_130_368#_c_406_n 0.0130683f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A2_c_136_n N_A_130_368#_c_406_n 0.0174421f $X=1.925 $Y=1.385 $X2=0
+ $Y2=0
cc_142 N_A2_c_137_n N_A_130_368#_c_406_n 0.00201785f $X=1.91 $Y=1.385 $X2=0
+ $Y2=0
cc_143 N_A2_M1001_g N_A_130_368#_c_409_n 0.00228751f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A2_M1003_g N_A_130_368#_c_409_n 0.00228751f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A2_c_136_n N_A_130_368#_c_409_n 0.0275631f $X=1.925 $Y=1.385 $X2=0
+ $Y2=0
cc_146 N_A2_c_137_n N_A_130_368#_c_409_n 0.00225438f $X=1.91 $Y=1.385 $X2=0
+ $Y2=0
cc_147 N_A2_c_134_n N_Y_c_515_n 0.00316716f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A2_c_132_n N_A_45_74#_c_570_n 6.33564e-19 $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A2_c_138_n N_A_45_74#_c_579_n 0.014682f $X=1.315 $Y=1.365 $X2=0 $Y2=0
cc_150 N_A2_c_134_n N_A_45_74#_c_571_n 0.00192588f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A2_c_136_n N_A_45_74#_c_571_n 0.0118504f $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A2_c_137_n N_A_45_74#_c_571_n 0.00376554f $X=1.91 $Y=1.385 $X2=0 $Y2=0
cc_153 N_A2_c_132_n N_A_45_74#_c_583_n 0.0116093f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A2_c_134_n N_A_45_74#_c_583_n 0.00924272f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A2_c_136_n N_A_45_74#_c_583_n 0.0324746f $X=1.925 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A2_c_137_n N_A_45_74#_c_583_n 0.00239267f $X=1.91 $Y=1.385 $X2=0 $Y2=0
cc_157 N_A2_c_132_n N_VGND_c_603_n 5.54504e-19 $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A2_c_132_n N_VGND_c_606_n 0.00433162f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A2_c_134_n N_VGND_c_606_n 0.00291649f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_160 N_A2_c_132_n N_VGND_c_608_n 0.00432528f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A2_c_134_n N_VGND_c_608_n 0.0036412f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_162 N_A2_c_132_n N_A_300_74#_c_654_n 0.00337267f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A2_c_134_n N_A_300_74#_c_654_n 0.0132302f $X=1.855 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A1_M1015_g N_B1_M1014_g 0.0200484f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_c_190_n N_B1_M1005_g 4.38787e-19 $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_166 N_A1_M1004_g B1 4.21136e-19 $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A1_c_190_n B1 0.0284542f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_168 N_A1_c_191_n B1 0.00243885f $X=3.035 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A1_c_190_n N_B1_c_244_n 6.20541e-19 $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_170 N_A1_c_191_n N_B1_c_244_n 0.0120684f $X=3.035 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A1_M1002_g N_VPWR_c_335_n 0.0173282f $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A1_M1004_g N_VPWR_c_335_n 5.96618e-19 $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_M1002_g N_VPWR_c_336_n 5.41206e-19 $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A1_M1004_g N_VPWR_c_336_n 0.014289f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A1_M1002_g N_VPWR_c_338_n 0.00460063f $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A1_M1004_g N_VPWR_c_338_n 0.00460063f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A1_M1002_g N_VPWR_c_330_n 0.00908554f $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A1_M1004_g N_VPWR_c_330_n 0.00908554f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A1_M1002_g N_A_130_368#_c_405_n 0.00109504f $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A1_M1002_g N_A_130_368#_c_406_n 0.0149303f $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A1_c_190_n N_A_130_368#_c_406_n 0.0159748f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_182 N_A1_M1002_g N_A_130_368#_c_407_n 3.62369e-19 $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A1_M1004_g N_A_130_368#_c_407_n 3.62369e-19 $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A1_M1004_g N_A_130_368#_c_408_n 0.0173389f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_c_190_n N_A_130_368#_c_408_n 0.0316217f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_186 N_A1_c_191_n N_A_130_368#_c_408_n 0.00784816f $X=3.035 $Y=1.515 $X2=0
+ $Y2=0
cc_187 N_A1_M1002_g N_A_130_368#_c_410_n 2.3892e-19 $X=2.39 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_M1004_g N_A_130_368#_c_410_n 0.00184981f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A1_c_190_n N_A_130_368#_c_410_n 0.0182439f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_190 N_A1_c_191_n N_A_130_368#_c_410_n 0.00252774f $X=3.035 $Y=1.515 $X2=0
+ $Y2=0
cc_191 N_A1_M1004_g N_A_692_368#_c_471_n 0.0010136f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A1_M1004_g N_A_692_368#_c_473_n 5.89323e-19 $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A1_M1011_g N_Y_c_515_n 0.0144828f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1015_g N_Y_c_515_n 0.0192938f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_c_190_n N_Y_c_515_n 0.0528772f $X=2.87 $Y=1.45 $X2=0 $Y2=0
cc_196 N_A1_c_191_n N_Y_c_515_n 0.0090734f $X=3.035 $Y=1.515 $X2=0 $Y2=0
cc_197 N_A1_M1015_g N_Y_c_516_n 4.15473e-19 $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A1_M1011_g N_VGND_c_606_n 0.00291649f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_M1015_g N_VGND_c_606_n 0.00433162f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A1_M1011_g N_VGND_c_608_n 0.0036412f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A1_M1015_g N_VGND_c_608_n 0.00449183f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A1_M1011_g N_A_300_74#_c_653_n 0.00479781f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A1_M1015_g N_A_300_74#_c_653_n 0.00420713f $X=3.365 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_M1011_g N_A_300_74#_c_654_n 0.0122192f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B1_M1014_g N_C1_M1000_g 0.0105379f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B1_M1006_g N_C1_M1007_g 0.0160413f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_207 B1 N_C1_M1007_g 0.00408271f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_208 B1 N_C1_c_292_n 0.0345267f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_209 B1 N_C1_c_293_n 0.0139618f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_210 N_B1_c_244_n N_C1_c_293_n 0.0215898f $X=4.26 $Y=1.515 $X2=0 $Y2=0
cc_211 N_B1_M1005_g N_VPWR_c_336_n 0.00186424f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_212 N_B1_M1005_g N_VPWR_c_339_n 0.00333891f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_213 N_B1_M1006_g N_VPWR_c_339_n 0.00333896f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B1_M1005_g N_VPWR_c_330_n 0.00427818f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_215 N_B1_M1006_g N_VPWR_c_330_n 0.00422796f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_216 N_B1_M1005_g N_A_130_368#_c_408_n 0.0162264f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_217 B1 N_A_130_368#_c_408_n 0.0308308f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_218 B1 N_A_130_368#_c_445_n 0.0154871f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B1_c_244_n N_A_130_368#_c_445_n 5.54777e-19 $X=4.26 $Y=1.515 $X2=0
+ $Y2=0
cc_220 N_B1_M1005_g N_A_692_368#_c_471_n 0.00899279f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B1_M1006_g N_A_692_368#_c_471_n 5.58167e-19 $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B1_M1005_g N_A_692_368#_c_472_n 0.0113093f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_223 N_B1_M1006_g N_A_692_368#_c_472_n 0.0116345f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_224 N_B1_M1005_g N_A_692_368#_c_473_n 0.00302214f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_225 N_B1_M1005_g N_A_692_368#_c_484_n 6.26133e-19 $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_226 N_B1_M1006_g N_A_692_368#_c_484_n 0.0129291f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_227 B1 N_A_692_368#_c_484_n 0.0233867f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_M1006_g N_A_692_368#_c_476_n 0.001916f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_229 B1 N_Y_c_515_n 8.08061e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B1_M1014_g N_Y_c_516_n 0.00654828f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B1_M1014_g N_Y_c_517_n 0.00909025f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_232 B1 N_Y_c_517_n 0.0221514f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B1_c_244_n N_Y_c_517_n 9.31826e-19 $X=4.26 $Y=1.515 $X2=0 $Y2=0
cc_234 N_B1_M1014_g N_Y_c_520_n 0.0104686f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_235 B1 N_Y_c_520_n 0.0720188f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B1_c_244_n N_Y_c_520_n 0.0122984f $X=4.26 $Y=1.515 $X2=0 $Y2=0
cc_237 N_B1_M1014_g N_VGND_c_604_n 0.00509642f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_M1014_g N_VGND_c_606_n 0.00434272f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_M1014_g N_VGND_c_608_n 0.00822954f $X=3.795 $Y=0.74 $X2=0 $Y2=0
cc_240 N_C1_M1007_g N_VPWR_c_339_n 0.00333896f $X=4.71 $Y=2.4 $X2=0 $Y2=0
cc_241 N_C1_M1012_g N_VPWR_c_339_n 0.00333896f $X=5.16 $Y=2.4 $X2=0 $Y2=0
cc_242 N_C1_M1007_g N_VPWR_c_330_n 0.00422796f $X=4.71 $Y=2.4 $X2=0 $Y2=0
cc_243 N_C1_M1012_g N_VPWR_c_330_n 0.00426715f $X=5.16 $Y=2.4 $X2=0 $Y2=0
cc_244 N_C1_M1007_g N_A_692_368#_c_484_n 0.0129423f $X=4.71 $Y=2.4 $X2=0 $Y2=0
cc_245 N_C1_M1012_g N_A_692_368#_c_484_n 6.27116e-19 $X=5.16 $Y=2.4 $X2=0 $Y2=0
cc_246 N_C1_c_293_n N_A_692_368#_c_484_n 2.22637e-19 $X=5.16 $Y=1.515 $X2=0
+ $Y2=0
cc_247 N_C1_M1007_g N_A_692_368#_c_474_n 0.0116345f $X=4.71 $Y=2.4 $X2=0 $Y2=0
cc_248 N_C1_M1012_g N_A_692_368#_c_474_n 0.014552f $X=5.16 $Y=2.4 $X2=0 $Y2=0
cc_249 N_C1_M1007_g N_A_692_368#_c_475_n 5.73047e-19 $X=4.71 $Y=2.4 $X2=0 $Y2=0
cc_250 N_C1_M1012_g N_A_692_368#_c_475_n 0.00892729f $X=5.16 $Y=2.4 $X2=0 $Y2=0
cc_251 N_C1_M1007_g N_A_692_368#_c_476_n 0.001916f $X=4.71 $Y=2.4 $X2=0 $Y2=0
cc_252 N_C1_M1012_g N_Y_c_521_n 0.0180748f $X=5.16 $Y=2.4 $X2=0 $Y2=0
cc_253 N_C1_c_292_n N_Y_c_521_n 0.00977036f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_254 N_C1_c_292_n N_Y_c_539_n 0.0144665f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_255 N_C1_c_293_n N_Y_c_539_n 5.53536e-19 $X=5.16 $Y=1.515 $X2=0 $Y2=0
cc_256 N_C1_M1000_g Y 0.0186914f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_257 N_C1_c_292_n Y 0.0281815f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_258 N_C1_c_293_n Y 0.0128182f $X=5.16 $Y=1.515 $X2=0 $Y2=0
cc_259 N_C1_M1000_g Y 0.00350742f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_260 N_C1_c_292_n Y 0.0263529f $X=5.01 $Y=1.515 $X2=0 $Y2=0
cc_261 N_C1_c_293_n Y 0.0174096f $X=5.16 $Y=1.515 $X2=0 $Y2=0
cc_262 N_C1_M1000_g N_Y_c_520_n 0.010805f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_263 N_C1_M1000_g N_VGND_c_604_n 0.00511882f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_264 N_C1_M1000_g N_VGND_c_607_n 0.00433162f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_265 N_C1_M1000_g N_VGND_c_608_n 0.00824204f $X=4.635 $Y=0.74 $X2=0 $Y2=0
cc_266 N_VPWR_c_332_n N_A_130_368#_c_402_n 0.0365535f $X=0.335 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_333_n N_A_130_368#_c_402_n 0.0144623f $X=1.15 $Y=3.33 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_334_n N_A_130_368#_c_402_n 0.0309473f $X=1.235 $Y=2.225 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_330_n N_A_130_368#_c_402_n 0.0118344f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_270 N_VPWR_M1017_s N_A_130_368#_c_403_n 0.00165831f $X=1.1 $Y=1.84 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_334_n N_A_130_368#_c_403_n 0.0126919f $X=1.235 $Y=2.225 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_332_n N_A_130_368#_c_404_n 0.00326551f $X=0.335 $Y=1.985 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_334_n N_A_130_368#_c_405_n 0.0309473f $X=1.235 $Y=2.225 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_335_n N_A_130_368#_c_405_n 0.0309974f $X=2.15 $Y=2.225 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_337_n N_A_130_368#_c_405_n 0.0144623f $X=2.05 $Y=3.33 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_330_n N_A_130_368#_c_405_n 0.0118344f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_277 N_VPWR_M1003_s N_A_130_368#_c_406_n 0.00197722f $X=2 $Y=1.84 $X2=0 $Y2=0
cc_278 N_VPWR_c_335_n N_A_130_368#_c_406_n 0.0172996f $X=2.15 $Y=2.225 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_335_n N_A_130_368#_c_407_n 0.030194f $X=2.15 $Y=2.225 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_336_n N_A_130_368#_c_407_n 0.0233699f $X=3.065 $Y=2.405 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_338_n N_A_130_368#_c_407_n 0.00749631f $X=2.9 $Y=3.33 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_330_n N_A_130_368#_c_407_n 0.0062048f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_283 N_VPWR_M1004_s N_A_130_368#_c_408_n 0.00466209f $X=2.93 $Y=1.84 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_336_n N_A_130_368#_c_408_n 0.0219767f $X=3.065 $Y=2.405 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_336_n N_A_692_368#_c_471_n 0.0473717f $X=3.065 $Y=2.405 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_339_n N_A_692_368#_c_472_n 0.0354851f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_330_n N_A_692_368#_c_472_n 0.0198934f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_336_n N_A_692_368#_c_473_n 0.0139f $X=3.065 $Y=2.405 $X2=0 $Y2=0
cc_289 N_VPWR_c_339_n N_A_692_368#_c_473_n 0.0238921f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_330_n N_A_692_368#_c_473_n 0.0128639f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_339_n N_A_692_368#_c_474_n 0.0593439f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_330_n N_A_692_368#_c_474_n 0.032751f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_293 N_VPWR_c_339_n N_A_692_368#_c_476_n 0.0234458f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_330_n N_A_692_368#_c_476_n 0.0125551f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_A_130_368#_c_408_n N_A_692_368#_M1005_s 0.00575251f $X=3.925 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_296 N_A_130_368#_c_408_n N_A_692_368#_c_471_n 0.0223576f $X=3.925 $Y=2.035
+ $X2=0 $Y2=0
cc_297 N_A_130_368#_M1005_d N_A_692_368#_c_472_n 0.00165831f $X=3.9 $Y=1.84
+ $X2=0 $Y2=0
cc_298 N_A_130_368#_c_445_n N_A_692_368#_c_472_n 0.0118736f $X=4.035 $Y=2.115
+ $X2=0 $Y2=0
cc_299 N_A_130_368#_c_406_n N_A_45_74#_c_571_n 0.00418019f $X=2.53 $Y=1.805
+ $X2=0 $Y2=0
cc_300 N_A_692_368#_c_474_n N_Y_M1007_d 0.00165831f $X=5.22 $Y=2.99 $X2=0 $Y2=0
cc_301 N_A_692_368#_M1012_s N_Y_c_521_n 0.00663587f $X=5.25 $Y=1.84 $X2=0 $Y2=0
cc_302 N_A_692_368#_c_475_n N_Y_c_521_n 0.0231797f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_303 N_A_692_368#_c_474_n N_Y_c_539_n 0.0118736f $X=5.22 $Y=2.99 $X2=0 $Y2=0
cc_304 N_A_692_368#_M1012_s Y 0.0017814f $X=5.25 $Y=1.84 $X2=0 $Y2=0
cc_305 N_Y_c_515_n N_A_45_74#_c_571_n 0.0118023f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_306 N_Y_c_520_n N_VGND_M1014_d 0.00793129f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_307 N_Y_c_516_n N_VGND_c_604_n 0.0184853f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_308 Y N_VGND_c_604_n 0.0214218f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_309 N_Y_c_520_n N_VGND_c_604_n 0.0468625f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_310 N_Y_c_516_n N_VGND_c_606_n 0.0109942f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_311 Y N_VGND_c_607_n 0.0421459f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_312 N_Y_c_515_n N_VGND_c_608_n 0.00699508f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_313 N_Y_c_516_n N_VGND_c_608_n 0.00904371f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_314 Y N_VGND_c_608_n 0.0349449f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_315 N_Y_c_515_n N_A_300_74#_M1011_s 0.00178215f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_316 N_Y_c_515_n N_A_300_74#_c_653_n 0.0165836f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_317 N_Y_c_516_n N_A_300_74#_c_653_n 0.0135554f $X=3.58 $Y=0.515 $X2=0 $Y2=0
cc_318 N_Y_M1011_d N_A_300_74#_c_654_n 0.00374227f $X=2.595 $Y=0.37 $X2=0 $Y2=0
cc_319 N_Y_c_515_n N_A_300_74#_c_654_n 0.0201119f $X=3.495 $Y=1.015 $X2=0 $Y2=0
cc_320 N_A_45_74#_c_573_n N_VGND_M1009_s 0.00406005f $X=1.125 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_321 N_A_45_74#_c_568_n N_VGND_c_603_n 0.0121972f $X=0.35 $Y=0.515 $X2=0 $Y2=0
cc_322 N_A_45_74#_c_573_n N_VGND_c_603_n 0.0167019f $X=1.125 $Y=0.925 $X2=0
+ $Y2=0
cc_323 N_A_45_74#_c_570_n N_VGND_c_603_n 0.0135953f $X=1.21 $Y=0.495 $X2=0 $Y2=0
cc_324 N_A_45_74#_c_568_n N_VGND_c_605_n 0.0110895f $X=0.35 $Y=0.515 $X2=0 $Y2=0
cc_325 N_A_45_74#_c_570_n N_VGND_c_606_n 0.00814895f $X=1.21 $Y=0.495 $X2=0
+ $Y2=0
cc_326 N_A_45_74#_c_568_n N_VGND_c_608_n 0.00916858f $X=0.35 $Y=0.515 $X2=0
+ $Y2=0
cc_327 N_A_45_74#_c_573_n N_VGND_c_608_n 0.0116543f $X=1.125 $Y=0.925 $X2=0
+ $Y2=0
cc_328 N_A_45_74#_c_570_n N_VGND_c_608_n 0.00627841f $X=1.21 $Y=0.495 $X2=0
+ $Y2=0
cc_329 N_A_45_74#_c_583_n N_VGND_c_608_n 0.0070825f $X=1.905 $Y=0.91 $X2=0 $Y2=0
cc_330 N_A_45_74#_c_583_n N_A_300_74#_M1008_s 0.0034629f $X=1.905 $Y=0.91
+ $X2=-0.19 $Y2=-0.245
cc_331 N_A_45_74#_M1013_d N_A_300_74#_c_654_n 0.0032303f $X=1.93 $Y=0.37 $X2=0
+ $Y2=0
cc_332 N_A_45_74#_c_570_n N_A_300_74#_c_654_n 0.010629f $X=1.21 $Y=0.495 $X2=0
+ $Y2=0
cc_333 N_A_45_74#_c_583_n N_A_300_74#_c_654_n 0.0430812f $X=1.905 $Y=0.91 $X2=0
+ $Y2=0
cc_334 N_VGND_c_606_n N_A_300_74#_c_654_n 0.0755134f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_608_n N_A_300_74#_c_654_n 0.064201f $X=5.52 $Y=0 $X2=0 $Y2=0

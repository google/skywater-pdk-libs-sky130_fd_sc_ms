* File: sky130_fd_sc_ms__fah_4.pxi.spice
* Created: Fri Aug 28 17:35:50 2020
* 
x_PM_SKY130_FD_SC_MS__FAH_4%A N_A_M1005_g N_A_M1037_g N_A_M1038_g N_A_M1006_g A
+ N_A_c_298_n N_A_c_299_n PM_SKY130_FD_SC_MS__FAH_4%A
x_PM_SKY130_FD_SC_MS__FAH_4%A_27_74# N_A_27_74#_M1037_s N_A_27_74#_M1005_s
+ N_A_27_74#_c_340_n N_A_27_74#_M1003_g N_A_27_74#_c_342_n N_A_27_74#_M1007_g
+ N_A_27_74#_c_343_n N_A_27_74#_c_344_n N_A_27_74#_c_351_n N_A_27_74#_c_352_n
+ N_A_27_74#_c_345_n N_A_27_74#_c_346_n N_A_27_74#_c_347_n N_A_27_74#_c_348_n
+ N_A_27_74#_c_349_n PM_SKY130_FD_SC_MS__FAH_4%A_27_74#
x_PM_SKY130_FD_SC_MS__FAH_4%A_586_257# N_A_586_257#_M1025_d N_A_586_257#_M1026_d
+ N_A_586_257#_M1010_d N_A_586_257#_c_411_n N_A_586_257#_M1019_g
+ N_A_586_257#_M1030_g N_A_586_257#_c_414_n N_A_586_257#_c_415_n
+ N_A_586_257#_M1035_g N_A_586_257#_M1029_g N_A_586_257#_c_418_n
+ N_A_586_257#_c_419_n N_A_586_257#_c_420_n N_A_586_257#_c_421_n
+ N_A_586_257#_c_422_n N_A_586_257#_c_423_n N_A_586_257#_c_430_n
+ N_A_586_257#_c_431_n N_A_586_257#_c_424_n N_A_586_257#_c_425_n
+ N_A_586_257#_c_470_p N_A_586_257#_c_432_n N_A_586_257#_c_426_n
+ PM_SKY130_FD_SC_MS__FAH_4%A_586_257#
x_PM_SKY130_FD_SC_MS__FAH_4%B N_B_M1033_g N_B_M1018_g N_B_c_588_n N_B_c_589_n
+ N_B_M1027_g N_B_M1023_g N_B_c_591_n N_B_M1025_g N_B_c_581_n N_B_c_593_n
+ N_B_M1010_g N_B_c_582_n N_B_c_583_n N_B_c_595_n N_B_c_596_n N_B_c_584_n
+ N_B_c_585_n N_B_c_598_n B B N_B_c_586_n PM_SKY130_FD_SC_MS__FAH_4%B
x_PM_SKY130_FD_SC_MS__FAH_4%A_531_362# N_A_531_362#_M1027_d N_A_531_362#_M1033_d
+ N_A_531_362#_c_726_n N_A_531_362#_M1000_g N_A_531_362#_c_728_n
+ N_A_531_362#_M1021_g N_A_531_362#_c_744_n N_A_531_362#_c_745_n
+ N_A_531_362#_c_729_n N_A_531_362#_M1041_g N_A_531_362#_M1043_g
+ N_A_531_362#_c_731_n N_A_531_362#_c_748_n N_A_531_362#_c_732_n
+ N_A_531_362#_c_749_n N_A_531_362#_c_733_n N_A_531_362#_c_734_n
+ N_A_531_362#_c_735_n N_A_531_362#_c_736_n N_A_531_362#_c_737_n
+ N_A_531_362#_c_738_n N_A_531_362#_c_739_n N_A_531_362#_c_740_n
+ N_A_531_362#_c_741_n N_A_531_362#_c_742_n PM_SKY130_FD_SC_MS__FAH_4%A_531_362#
x_PM_SKY130_FD_SC_MS__FAH_4%A_536_114# N_A_536_114#_M1018_d N_A_536_114#_M1023_d
+ N_A_536_114#_M1040_g N_A_536_114#_M1004_g N_A_536_114#_c_932_n
+ N_A_536_114#_c_933_n N_A_536_114#_M1026_g N_A_536_114#_c_935_n
+ N_A_536_114#_c_944_n N_A_536_114#_c_945_n N_A_536_114#_c_946_n
+ N_A_536_114#_M1001_g N_A_536_114#_c_936_n N_A_536_114#_c_954_n
+ N_A_536_114#_c_937_n N_A_536_114#_c_938_n N_A_536_114#_c_939_n
+ N_A_536_114#_c_962_n N_A_536_114#_c_948_n N_A_536_114#_c_968_n
+ N_A_536_114#_c_1019_n N_A_536_114#_c_940_n N_A_536_114#_c_941_n
+ N_A_536_114#_c_969_n PM_SKY130_FD_SC_MS__FAH_4%A_536_114#
x_PM_SKY130_FD_SC_MS__FAH_4%A_1378_125# N_A_1378_125#_M1040_d
+ N_A_1378_125#_M1017_s N_A_1378_125#_M1004_d N_A_1378_125#_M1034_s
+ N_A_1378_125#_M1016_g N_A_1378_125#_c_1128_n N_A_1378_125#_c_1129_n
+ N_A_1378_125#_M1020_g N_A_1378_125#_c_1130_n N_A_1378_125#_c_1131_n
+ N_A_1378_125#_c_1140_n N_A_1378_125#_c_1132_n N_A_1378_125#_c_1155_n
+ N_A_1378_125#_c_1156_n N_A_1378_125#_c_1142_n N_A_1378_125#_c_1143_n
+ N_A_1378_125#_c_1133_n N_A_1378_125#_c_1192_n N_A_1378_125#_c_1145_n
+ N_A_1378_125#_c_1134_n N_A_1378_125#_c_1230_p N_A_1378_125#_c_1146_n
+ N_A_1378_125#_c_1147_n N_A_1378_125#_c_1135_n N_A_1378_125#_c_1136_n
+ N_A_1378_125#_c_1157_n N_A_1378_125#_c_1172_n N_A_1378_125#_c_1203_n
+ N_A_1378_125#_c_1148_n N_A_1378_125#_c_1149_n N_A_1378_125#_c_1137_n
+ N_A_1378_125#_c_1150_n N_A_1378_125#_c_1151_n N_A_1378_125#_c_1138_n
+ PM_SKY130_FD_SC_MS__FAH_4%A_1378_125#
x_PM_SKY130_FD_SC_MS__FAH_4%A_1268_379# N_A_1268_379#_M1041_d
+ N_A_1268_379#_M1000_d N_A_1268_379#_M1008_g N_A_1268_379#_M1024_g
+ N_A_1268_379#_c_1348_n N_A_1268_379#_M1009_g N_A_1268_379#_c_1349_n
+ N_A_1268_379#_M1011_g N_A_1268_379#_M1036_g N_A_1268_379#_M1039_g
+ N_A_1268_379#_c_1350_n N_A_1268_379#_M1014_g N_A_1268_379#_c_1351_n
+ N_A_1268_379#_M1022_g N_A_1268_379#_c_1368_n N_A_1268_379#_c_1352_n
+ N_A_1268_379#_c_1353_n N_A_1268_379#_c_1354_n N_A_1268_379#_c_1355_n
+ N_A_1268_379#_c_1356_n N_A_1268_379#_c_1418_n N_A_1268_379#_c_1438_p
+ N_A_1268_379#_c_1419_n N_A_1268_379#_c_1357_n N_A_1268_379#_c_1446_p
+ N_A_1268_379#_c_1365_n N_A_1268_379#_c_1358_n N_A_1268_379#_c_1359_n
+ PM_SKY130_FD_SC_MS__FAH_4%A_1268_379#
x_PM_SKY130_FD_SC_MS__FAH_4%CI N_CI_M1034_g N_CI_M1017_g CI N_CI_c_1522_n
+ N_CI_c_1523_n N_CI_c_1524_n PM_SKY130_FD_SC_MS__FAH_4%CI
x_PM_SKY130_FD_SC_MS__FAH_4%A_1278_102# N_A_1278_102#_M1021_d
+ N_A_1278_102#_M1043_d N_A_1278_102#_M1012_g N_A_1278_102#_c_1560_n
+ N_A_1278_102#_M1002_g N_A_1278_102#_M1013_g N_A_1278_102#_c_1561_n
+ N_A_1278_102#_M1028_g N_A_1278_102#_M1015_g N_A_1278_102#_c_1562_n
+ N_A_1278_102#_M1031_g N_A_1278_102#_c_1563_n N_A_1278_102#_M1042_g
+ N_A_1278_102#_M1032_g N_A_1278_102#_c_1564_n N_A_1278_102#_c_1565_n
+ N_A_1278_102#_c_1579_n N_A_1278_102#_c_1566_n N_A_1278_102#_c_1567_n
+ N_A_1278_102#_c_1568_n N_A_1278_102#_c_1645_n N_A_1278_102#_c_1615_n
+ N_A_1278_102#_c_1569_n N_A_1278_102#_c_1570_n N_A_1278_102#_c_1571_n
+ N_A_1278_102#_c_1572_n N_A_1278_102#_c_1702_p N_A_1278_102#_c_1573_n
+ N_A_1278_102#_c_1582_n N_A_1278_102#_c_1739_p N_A_1278_102#_c_1574_n
+ PM_SKY130_FD_SC_MS__FAH_4%A_1278_102#
x_PM_SKY130_FD_SC_MS__FAH_4%VPWR N_VPWR_M1005_d N_VPWR_M1003_s N_VPWR_M1010_s
+ N_VPWR_M1016_d N_VPWR_M1024_s N_VPWR_M1039_s N_VPWR_M1034_d N_VPWR_M1013_s
+ N_VPWR_M1032_s N_VPWR_c_1777_n N_VPWR_c_1778_n N_VPWR_c_1779_n N_VPWR_c_1780_n
+ N_VPWR_c_1781_n N_VPWR_c_1782_n N_VPWR_c_1783_n N_VPWR_c_1784_n
+ N_VPWR_c_1785_n N_VPWR_c_1786_n VPWR N_VPWR_c_1787_n N_VPWR_c_1788_n
+ N_VPWR_c_1789_n N_VPWR_c_1790_n N_VPWR_c_1791_n N_VPWR_c_1792_n
+ N_VPWR_c_1793_n N_VPWR_c_1794_n N_VPWR_c_1795_n N_VPWR_c_1796_n
+ N_VPWR_c_1797_n N_VPWR_c_1798_n N_VPWR_c_1799_n N_VPWR_c_1776_n
+ PM_SKY130_FD_SC_MS__FAH_4%VPWR
x_PM_SKY130_FD_SC_MS__FAH_4%A_200_74# N_A_200_74#_M1038_d N_A_200_74#_M1030_d
+ N_A_200_74#_M1006_d N_A_200_74#_M1019_d N_A_200_74#_c_1943_n
+ N_A_200_74#_c_1951_n N_A_200_74#_c_1952_n N_A_200_74#_c_1944_n
+ N_A_200_74#_c_1945_n N_A_200_74#_c_1953_n N_A_200_74#_c_1946_n
+ N_A_200_74#_c_1947_n N_A_200_74#_c_1955_n N_A_200_74#_c_1948_n
+ N_A_200_74#_c_1949_n N_A_200_74#_c_1950_n N_A_200_74#_c_1980_n
+ N_A_200_74#_c_1981_n N_A_200_74#_c_1956_n PM_SKY130_FD_SC_MS__FAH_4%A_200_74#
x_PM_SKY130_FD_SC_MS__FAH_4%A_430_362# N_A_430_362#_M1007_d N_A_430_362#_M1035_d
+ N_A_430_362#_M1003_d N_A_430_362#_M1029_d N_A_430_362#_c_2067_n
+ N_A_430_362#_c_2056_n N_A_430_362#_c_2053_n N_A_430_362#_c_2058_n
+ N_A_430_362#_c_2086_n N_A_430_362#_c_2059_n N_A_430_362#_c_2060_n
+ N_A_430_362#_c_2054_n N_A_430_362#_c_2055_n
+ PM_SKY130_FD_SC_MS__FAH_4%A_430_362#
x_PM_SKY130_FD_SC_MS__FAH_4%A_1183_102# N_A_1183_102#_M1021_s
+ N_A_1183_102#_M1020_s N_A_1183_102#_M1001_d N_A_1183_102#_c_2137_n
+ N_A_1183_102#_c_2145_n N_A_1183_102#_c_2138_n N_A_1183_102#_c_2139_n
+ N_A_1183_102#_c_2140_n N_A_1183_102#_c_2141_n N_A_1183_102#_c_2142_n
+ N_A_1183_102#_c_2143_n N_A_1183_102#_c_2144_n
+ PM_SKY130_FD_SC_MS__FAH_4%A_1183_102#
x_PM_SKY130_FD_SC_MS__FAH_4%COUT N_COUT_M1009_d N_COUT_M1014_d N_COUT_M1008_d
+ N_COUT_M1036_d N_COUT_c_2249_n N_COUT_c_2255_n N_COUT_c_2244_n N_COUT_c_2245_n
+ N_COUT_c_2265_n COUT PM_SKY130_FD_SC_MS__FAH_4%COUT
x_PM_SKY130_FD_SC_MS__FAH_4%SUM N_SUM_M1002_s N_SUM_M1031_s N_SUM_M1012_d
+ N_SUM_M1015_d N_SUM_c_2296_n N_SUM_c_2293_n N_SUM_c_2290_n N_SUM_c_2306_n
+ N_SUM_c_2310_n N_SUM_c_2314_n N_SUM_c_2291_n N_SUM_c_2292_n N_SUM_c_2325_n SUM
+ SUM SUM SUM PM_SKY130_FD_SC_MS__FAH_4%SUM
x_PM_SKY130_FD_SC_MS__FAH_4%VGND N_VGND_M1037_d N_VGND_M1007_s N_VGND_M1025_s
+ N_VGND_M1020_d N_VGND_M1011_s N_VGND_M1022_s N_VGND_M1017_d N_VGND_M1028_d
+ N_VGND_M1042_d N_VGND_c_2353_n N_VGND_c_2354_n N_VGND_c_2355_n N_VGND_c_2356_n
+ N_VGND_c_2357_n N_VGND_c_2358_n N_VGND_c_2359_n N_VGND_c_2360_n
+ N_VGND_c_2361_n N_VGND_c_2362_n N_VGND_c_2363_n N_VGND_c_2364_n
+ N_VGND_c_2365_n N_VGND_c_2366_n N_VGND_c_2367_n N_VGND_c_2368_n
+ N_VGND_c_2369_n N_VGND_c_2370_n N_VGND_c_2371_n N_VGND_c_2372_n VGND
+ N_VGND_c_2373_n N_VGND_c_2374_n N_VGND_c_2375_n N_VGND_c_2376_n
+ N_VGND_c_2377_n N_VGND_c_2378_n N_VGND_c_2379_n N_VGND_c_2380_n
+ PM_SKY130_FD_SC_MS__FAH_4%VGND
cc_1 VNB N_A_M1037_g 0.0412524f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_A_M1038_g 0.0426015f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.69
cc_3 VNB N_A_c_298_n 0.026091f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.635
cc_4 VNB N_A_c_299_n 0.00139506f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.635
cc_5 VNB N_A_27_74#_c_340_n 0.0245076f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_6 VNB N_A_27_74#_M1003_g 0.00858251f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.69
cc_7 VNB N_A_27_74#_c_342_n 0.0200397f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.8
cc_8 VNB N_A_27_74#_c_343_n 0.0116462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_344_n 0.036209f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.635
cc_10 VNB N_A_27_74#_c_345_n 0.0177754f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.655
cc_11 VNB N_A_27_74#_c_346_n 0.00948845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_347_n 0.0151628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_348_n 0.00597812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_349_n 0.0319921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_586_257#_c_411_n 0.00513041f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.69
cc_16 VNB N_A_586_257#_M1019_g 0.0139335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_586_257#_M1030_g 0.0224714f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_A_586_257#_c_414_n 0.123671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_586_257#_c_415_n 0.0126957f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.635
cc_20 VNB N_A_586_257#_M1035_g 0.0115669f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.635
cc_21 VNB N_A_586_257#_M1029_g 0.00650845f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.655
cc_22 VNB N_A_586_257#_c_418_n 0.0143455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_586_257#_c_419_n 0.00241727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_586_257#_c_420_n 0.00970608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_586_257#_c_421_n 4.43882e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_586_257#_c_422_n 0.00799781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_586_257#_c_423_n 0.00360986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_586_257#_c_424_n 0.00279228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_586_257#_c_425_n 0.0455158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_586_257#_c_426_n 0.0041569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_M1033_g 0.00169103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_M1018_g 0.0230225f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_33 VNB N_B_M1027_g 0.0257908f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.8
cc_34 VNB N_B_c_581_n 0.0177375f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.635
cc_35 VNB N_B_c_582_n 0.0129725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_c_583_n 0.00823579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_584_n 0.00309161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_c_585_n 0.0491482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_c_586_n 0.0210497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_531_362#_c_726_n 0.0262425f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_41 VNB N_A_531_362#_M1000_g 0.0140818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_531_362#_c_728_n 0.0182193f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.8
cc_43 VNB N_A_531_362#_c_729_n 0.00524739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_531_362#_M1041_g 0.0310732f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.635
cc_45 VNB N_A_531_362#_c_731_n 0.0107711f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.655
cc_46 VNB N_A_531_362#_c_732_n 0.00616063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_531_362#_c_733_n 0.00355979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_531_362#_c_734_n 0.0367291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_531_362#_c_735_n 7.86527e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_531_362#_c_736_n 0.00142874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_531_362#_c_737_n 0.00941364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_531_362#_c_738_n 0.00171766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_531_362#_c_739_n 0.00329535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_531_362#_c_740_n 0.0025665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_531_362#_c_741_n 0.00305769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_531_362#_c_742_n 0.00341732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_536_114#_M1040_g 0.0326569f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.69
cc_58 VNB N_A_536_114#_c_932_n 0.0629254f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_59 VNB N_A_536_114#_c_933_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_536_114#_M1026_g 0.038262f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.635
cc_61 VNB N_A_536_114#_c_935_n 0.0067347f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.635
cc_62 VNB N_A_536_114#_c_936_n 0.0190896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_536_114#_c_937_n 0.00479265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_536_114#_c_938_n 0.00312166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_536_114#_c_939_n 0.00208534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_536_114#_c_940_n 0.0194231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_536_114#_c_941_n 0.00461116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1378_125#_M1016_g 6.87871e-19 $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_69 VNB N_A_1378_125#_c_1128_n 0.029712f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_70 VNB N_A_1378_125#_c_1129_n 0.0194911f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.635
cc_71 VNB N_A_1378_125#_c_1130_n 0.0606606f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=1.635
cc_72 VNB N_A_1378_125#_c_1131_n 0.0166148f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=1.635
cc_73 VNB N_A_1378_125#_c_1132_n 0.00318612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1378_125#_c_1133_n 2.18548e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1378_125#_c_1134_n 0.00182852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1378_125#_c_1135_n 0.00381942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1378_125#_c_1136_n 0.00390559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1378_125#_c_1137_n 0.00521068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1378_125#_c_1138_n 0.0099962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1268_379#_c_1348_n 0.0178234f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_81 VNB N_A_1268_379#_c_1349_n 0.0173227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1268_379#_c_1350_n 0.0167614f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=1.655
cc_83 VNB N_A_1268_379#_c_1351_n 0.0171709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1268_379#_c_1352_n 0.00547584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1268_379#_c_1353_n 0.0158008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1268_379#_c_1354_n 0.00837569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1268_379#_c_1355_n 0.00647118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1268_379#_c_1356_n 0.00406402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1268_379#_c_1357_n 0.0023506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1268_379#_c_1358_n 2.00779e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1268_379#_c_1359_n 0.117337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_CI_c_1522_n 0.0309874f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.69
cc_93 VNB N_CI_c_1523_n 0.00469037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_CI_c_1524_n 0.0226132f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.8
cc_95 VNB N_A_1278_102#_c_1560_n 0.0175886f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.69
cc_96 VNB N_A_1278_102#_c_1561_n 0.0157917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1278_102#_c_1562_n 0.0157666f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.635
cc_98 VNB N_A_1278_102#_c_1563_n 0.0190146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1278_102#_c_1564_n 0.0138786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1278_102#_c_1565_n 0.00907818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1278_102#_c_1566_n 0.0318645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1278_102#_c_1567_n 0.00356064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1278_102#_c_1568_n 0.00562295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1278_102#_c_1569_n 0.00945148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1278_102#_c_1570_n 0.00816918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1278_102#_c_1571_n 0.00207724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1278_102#_c_1572_n 0.00218313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1278_102#_c_1573_n 3.26534e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1278_102#_c_1574_n 0.0902967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VPWR_c_1776_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_200_74#_c_1943_n 0.0083354f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_112 VNB N_A_200_74#_c_1944_n 0.00766276f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.635
cc_113 VNB N_A_200_74#_c_1945_n 3.33625e-19 $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=1.635
cc_114 VNB N_A_200_74#_c_1946_n 0.00273312f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.655
cc_115 VNB N_A_200_74#_c_1947_n 4.04208e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_200_74#_c_1948_n 0.022654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_200_74#_c_1949_n 0.00283451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_200_74#_c_1950_n 0.00423936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_430_362#_c_2053_n 0.00847888f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.635
cc_120 VNB N_A_430_362#_c_2054_n 0.00796915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_430_362#_c_2055_n 0.00646182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1183_102#_c_2137_n 0.00400184f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.8
cc_123 VNB N_A_1183_102#_c_2138_n 0.00416306f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.635
cc_124 VNB N_A_1183_102#_c_2139_n 0.00511891f $X=-0.19 $Y=-0.245 $X2=0.93
+ $Y2=1.635
cc_125 VNB N_A_1183_102#_c_2140_n 0.00498462f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.655
cc_126 VNB N_A_1183_102#_c_2141_n 0.00241138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1183_102#_c_2142_n 0.0045185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1183_102#_c_2143_n 0.00376343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_1183_102#_c_2144_n 0.00218094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_COUT_c_2244_n 0.00744718f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.635
cc_131 VNB N_COUT_c_2245_n 2.03526e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.655
cc_132 VNB COUT 9.02517e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_SUM_c_2290_n 0.00252589f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.635
cc_134 VNB N_SUM_c_2291_n 0.00252451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_SUM_c_2292_n 0.00103798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2353_n 0.00559476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2354_n 0.0111162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2355_n 0.00949613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2356_n 0.00714062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2357_n 0.0110399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2358_n 0.0172286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2359_n 0.0168841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2360_n 0.0076199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2361_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2362_n 0.0570466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2363_n 0.0171566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2364_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2365_n 0.0699813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2366_n 0.00631846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2367_n 0.117702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2368_n 0.00477896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2369_n 0.0179354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2370_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2371_n 0.0184888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2372_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2373_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2374_n 0.0204264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2375_n 0.0178099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2376_n 0.0175291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2377_n 0.0049761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2378_n 0.0065087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2379_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2380_n 0.788711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VPB N_A_M1005_g 0.0260646f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_165 VPB N_A_M1006_g 0.0279343f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_166 VPB N_A_c_298_n 0.0211049f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_167 VPB N_A_c_299_n 0.00565092f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_168 VPB N_A_27_74#_M1003_g 0.0251123f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.69
cc_169 VPB N_A_27_74#_c_351_n 0.00536733f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_170 VPB N_A_27_74#_c_352_n 0.0359862f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.635
cc_171 VPB N_A_27_74#_c_347_n 0.0146823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_27_74#_c_348_n 0.00972014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_27_74#_c_349_n 0.00801318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_586_257#_M1019_g 0.017725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_586_257#_M1029_g 0.0211386f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.655
cc_176 VPB N_A_586_257#_c_423_n 0.00197822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_586_257#_c_430_n 0.00289646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_586_257#_c_431_n 0.00502683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_586_257#_c_432_n 0.00179224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_B_M1033_g 0.0339571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_B_c_588_n 0.0593489f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.47
cc_182 VPB N_B_c_589_n 0.0136144f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.69
cc_183 VPB N_B_M1023_g 0.035202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_B_c_591_n 0.0636826f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.635
cc_185 VPB N_B_c_581_n 0.0225824f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_186 VPB N_B_c_593_n 0.0197521f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.655
cc_187 VPB N_B_c_583_n 0.00824806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_B_c_595_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_B_c_596_n 0.0575079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_B_c_585_n 0.00947325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_B_c_598_n 0.0869696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB B 0.00842404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_531_362#_M1000_g 0.03667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_531_362#_c_744_n 0.0842742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_531_362#_c_745_n 0.0138928f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_196 VPB N_A_531_362#_c_729_n 0.0298219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_531_362#_M1043_g 0.0162556f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.635
cc_198 VPB N_A_531_362#_c_748_n 8.68553e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_531_362#_c_749_n 0.00119535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_531_362#_c_735_n 0.00122028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_531_362#_c_736_n 0.00200282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_531_362#_c_737_n 0.00156811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_531_362#_c_738_n 9.34773e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_531_362#_c_739_n 0.00312165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_531_362#_c_740_n 5.94209e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_531_362#_c_741_n 0.00103142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_531_362#_c_742_n 6.95589e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_536_114#_M1004_g 0.0196975f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.8
cc_209 VPB N_A_536_114#_c_935_n 0.0134841f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_210 VPB N_A_536_114#_c_944_n 0.0336047f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_211 VPB N_A_536_114#_c_945_n 0.0107368f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_212 VPB N_A_536_114#_c_946_n 0.0211047f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.635
cc_213 VPB N_A_536_114#_c_939_n 0.0013019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_536_114#_c_948_n 0.00579394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_536_114#_c_940_n 0.0106635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_536_114#_c_941_n 0.00229624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1378_125#_M1016_g 0.0295826f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_218 VPB N_A_1378_125#_c_1140_n 0.0018385f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=1.635
cc_219 VPB N_A_1378_125#_c_1132_n 0.00137024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1378_125#_c_1142_n 0.00242283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1378_125#_c_1143_n 0.00324866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1378_125#_c_1133_n 0.00313877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1378_125#_c_1145_n 0.00508016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1378_125#_c_1146_n 0.00924466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1378_125#_c_1147_n 0.0191248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1378_125#_c_1148_n 0.0156487f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1378_125#_c_1149_n 0.00176287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1378_125#_c_1150_n 0.00295895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1378_125#_c_1151_n 0.00280614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1378_125#_c_1138_n 0.00548583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1268_379#_M1008_g 0.0243183f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.47
cc_232 VPB N_A_1268_379#_M1024_g 0.0231837f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.8
cc_233 VPB N_A_1268_379#_M1036_g 0.0224204f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_234 VPB N_A_1268_379#_M1039_g 0.0230488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1268_379#_c_1352_n 0.00158722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1268_379#_c_1365_n 9.52746e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1268_379#_c_1359_n 0.0338462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_CI_M1034_g 0.0264516f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_239 VPB N_CI_c_1522_n 0.0059217f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.69
cc_240 VPB N_CI_c_1523_n 0.00542064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1278_102#_M1012_g 0.0230595f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.47
cc_242 VPB N_A_1278_102#_M1013_g 0.022308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1278_102#_M1015_g 0.0223861f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_244 VPB N_A_1278_102#_M1032_g 0.0258625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1278_102#_c_1579_n 0.00158464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1278_102#_c_1569_n 0.00788264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1278_102#_c_1572_n 0.00137598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1278_102#_c_1582_n 0.00233749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1278_102#_c_1574_n 0.014623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1777_n 0.0055443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1778_n 0.0122591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1779_n 0.0134912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1780_n 0.0089971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1781_n 0.0120875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1782_n 0.0583744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1783_n 0.0138213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1784_n 0.0196302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1785_n 0.0217477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1786_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1787_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1788_n 0.0203166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1789_n 0.0947465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1790_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1791_n 0.0196104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1792_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1793_n 0.0147666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1794_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1795_n 0.0823222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1796_n 0.0196476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1797_n 0.0196302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1798_n 0.024486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1799_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1776_n 0.12093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_200_74#_c_1951_n 0.00562616f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_275 VPB N_A_200_74#_c_1952_n 0.00715555f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.635
cc_276 VPB N_A_200_74#_c_1953_n 0.012804f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_277 VPB N_A_200_74#_c_1946_n 0.00561673f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.655
cc_278 VPB N_A_200_74#_c_1955_n 0.00511378f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.655
cc_279 VPB N_A_200_74#_c_1956_n 0.00782515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_430_362#_c_2056_n 0.00462982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_430_362#_c_2053_n 0.00207464f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.635
cc_282 VPB N_A_430_362#_c_2058_n 0.00561071f $X=-0.19 $Y=1.66 $X2=0.925
+ $Y2=1.635
cc_283 VPB N_A_430_362#_c_2059_n 7.2733e-19 $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.635
cc_284 VPB N_A_430_362#_c_2060_n 0.00149358f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.655
cc_285 VPB N_A_430_362#_c_2055_n 0.00352699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_1183_102#_c_2145_n 0.00255151f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=2.46
cc_287 VPB N_A_1183_102#_c_2140_n 0.0155832f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.655
cc_288 VPB N_A_1183_102#_c_2141_n 0.00252098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_A_1183_102#_c_2142_n 0.00483988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_1183_102#_c_2143_n 0.00522976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_A_1183_102#_c_2144_n 0.00458784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_SUM_c_2293_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_293 VPB N_SUM_c_2292_n 0.00151412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB SUM 0.00240191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 N_A_M1037_g N_A_27_74#_c_344_n 0.0069942f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_296 N_A_M1005_g N_A_27_74#_c_352_n 4.7096e-19 $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_297 N_A_M1037_g N_A_27_74#_c_345_n 0.0158996f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_298 N_A_M1038_g N_A_27_74#_c_345_n 0.0156348f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_299 N_A_c_298_n N_A_27_74#_c_345_n 0.00505519f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_300 N_A_c_299_n N_A_27_74#_c_345_n 0.0487599f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_301 N_A_M1037_g N_A_27_74#_c_347_n 0.00728315f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_302 N_A_c_298_n N_A_27_74#_c_347_n 0.00897861f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_303 N_A_c_299_n N_A_27_74#_c_347_n 0.0229882f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_304 N_A_M1038_g N_A_27_74#_c_348_n 0.00127558f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_305 N_A_c_298_n N_A_27_74#_c_348_n 4.84451e-19 $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_306 N_A_c_299_n N_A_27_74#_c_348_n 0.00840148f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_307 N_A_M1038_g N_A_27_74#_c_349_n 0.00625278f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_308 N_A_c_298_n N_A_27_74#_c_349_n 0.00997888f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_309 N_A_c_299_n N_A_27_74#_c_349_n 5.10923e-19 $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_310 N_A_M1005_g N_VPWR_c_1777_n 0.0193916f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_311 N_A_M1006_g N_VPWR_c_1777_n 0.00297869f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_312 N_A_c_298_n N_VPWR_c_1777_n 0.00215577f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_313 N_A_c_299_n N_VPWR_c_1777_n 0.0173474f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_314 N_A_M1005_g N_VPWR_c_1787_n 0.00460063f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_315 N_A_M1006_g N_VPWR_c_1788_n 0.00519767f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_316 N_A_M1006_g N_VPWR_c_1793_n 0.00285056f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_317 N_A_M1005_g N_VPWR_c_1776_n 0.00912296f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_318 N_A_M1006_g N_VPWR_c_1776_n 0.0098373f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_319 N_A_M1038_g N_A_200_74#_c_1943_n 0.00515882f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_320 N_A_M1006_g N_A_200_74#_c_1951_n 0.00485231f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_321 N_A_M1006_g N_A_200_74#_c_1952_n 0.00823125f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_322 N_A_c_299_n N_A_200_74#_c_1952_n 0.00409946f $X=0.93 $Y=1.635 $X2=0 $Y2=0
cc_323 N_A_M1038_g N_A_200_74#_c_1945_n 0.00251256f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_324 N_A_M1037_g N_VGND_c_2353_n 0.0136178f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_325 N_A_M1038_g N_VGND_c_2353_n 0.00294833f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_326 N_A_M1038_g N_VGND_c_2354_n 0.00314342f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_327 N_A_M1037_g N_VGND_c_2363_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_328 N_A_M1038_g N_VGND_c_2373_n 0.00434272f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_329 N_A_M1037_g N_VGND_c_2380_n 0.00761198f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_330 N_A_M1038_g N_VGND_c_2380_n 0.00825283f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_342_n N_B_M1018_g 0.0199186f $X=2.13 $Y=1.32 $X2=0 $Y2=0
cc_332 N_A_27_74#_M1003_g N_B_c_582_n 0.0315596f $X=2.06 $Y=2.37 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_343_n N_B_c_582_n 8.55344e-19 $X=2.087 $Y=1.395 $X2=0 $Y2=0
cc_334 N_A_27_74#_c_352_n N_VPWR_c_1777_n 0.0325765f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_352_n N_VPWR_c_1787_n 0.0124046f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_M1003_g N_VPWR_c_1789_n 0.00498031f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_M1003_g N_VPWR_c_1793_n 0.00387214f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_M1003_g N_VPWR_c_1776_n 0.00643509f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_352_n N_VPWR_c_1776_n 0.0102675f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_M1003_g N_A_200_74#_c_1951_n 0.00403522f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_M1003_g N_A_200_74#_c_1952_n 0.00320339f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_345_n N_A_200_74#_c_1952_n 0.00755559f $X=1.335 $Y=1.255
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_c_348_n N_A_200_74#_c_1952_n 4.33375e-19 $X=1.5 $Y=1.255 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_345_n N_A_200_74#_c_1944_n 0.00225701f $X=1.335 $Y=1.255
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_c_348_n N_A_200_74#_c_1944_n 0.0269944f $X=1.5 $Y=1.255 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_349_n N_A_200_74#_c_1944_n 0.00671447f $X=1.5 $Y=1.395 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_345_n N_A_200_74#_c_1945_n 0.0244789f $X=1.335 $Y=1.255
+ $X2=0 $Y2=0
cc_348 N_A_27_74#_c_340_n N_A_200_74#_c_1946_n 0.0100734f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_M1003_g N_A_200_74#_c_1946_n 0.033785f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_342_n N_A_200_74#_c_1946_n 0.00665243f $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_343_n N_A_200_74#_c_1946_n 0.00325556f $X=2.087 $Y=1.395
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_348_n N_A_200_74#_c_1946_n 0.0360181f $X=1.5 $Y=1.255 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_349_n N_A_200_74#_c_1946_n 0.00117139f $X=1.5 $Y=1.395 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_342_n N_A_200_74#_c_1947_n 0.0127769f $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_M1003_g N_A_200_74#_c_1955_n 0.0133514f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_356 N_A_27_74#_c_342_n N_A_200_74#_c_1948_n 0.00671582f $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_342_n N_A_200_74#_c_1949_n 0.00327201f $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_342_n N_A_200_74#_c_1980_n 0.0106459f $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_M1003_g N_A_200_74#_c_1981_n 0.00526159f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_M1003_g N_A_430_362#_c_2056_n 2.25052e-19 $X=2.06 $Y=2.37
+ $X2=0 $Y2=0
cc_361 N_A_27_74#_c_343_n N_A_430_362#_c_2056_n 0.00118597f $X=2.087 $Y=1.395
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_M1003_g N_A_430_362#_c_2053_n 0.0025091f $X=2.06 $Y=2.37 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_342_n N_A_430_362#_c_2053_n 0.00524153f $X=2.13 $Y=1.32
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_c_348_n N_VGND_M1007_s 0.00156848f $X=1.5 $Y=1.255 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_344_n N_VGND_c_2353_n 0.023067f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_345_n N_VGND_c_2353_n 0.0177054f $X=1.335 $Y=1.255 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_342_n N_VGND_c_2354_n 0.00164705f $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_344_n N_VGND_c_2363_n 0.0124046f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_342_n N_VGND_c_2365_n 7.81861e-19 $X=2.13 $Y=1.32 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_344_n N_VGND_c_2380_n 0.0102675f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_371 N_A_586_257#_M1019_g N_B_M1033_g 0.0392344f $X=3.02 $Y=2.23 $X2=0 $Y2=0
cc_372 N_A_586_257#_c_411_n N_B_M1018_g 0.00796434f $X=3.02 $Y=1.375 $X2=0 $Y2=0
cc_373 N_A_586_257#_M1030_g N_B_M1018_g 0.00936875f $X=3.035 $Y=0.89 $X2=0 $Y2=0
cc_374 N_A_586_257#_M1019_g N_B_c_588_n 0.00909182f $X=3.02 $Y=2.23 $X2=0 $Y2=0
cc_375 N_A_586_257#_M1030_g N_B_M1027_g 0.0147851f $X=3.035 $Y=0.89 $X2=0 $Y2=0
cc_376 N_A_586_257#_c_414_n N_B_M1027_g 0.0202577f $X=3.94 $Y=0.205 $X2=0 $Y2=0
cc_377 N_A_586_257#_M1029_g N_B_M1027_g 0.00169039f $X=4.09 $Y=2.23 $X2=0 $Y2=0
cc_378 N_A_586_257#_c_419_n N_B_M1027_g 3.66293e-19 $X=4.22 $Y=0.375 $X2=0 $Y2=0
cc_379 N_A_586_257#_M1019_g N_B_M1023_g 0.0268898f $X=3.02 $Y=2.23 $X2=0 $Y2=0
cc_380 N_A_586_257#_M1029_g N_B_c_591_n 0.0104341f $X=4.09 $Y=2.23 $X2=0 $Y2=0
cc_381 N_A_586_257#_c_423_n N_B_c_581_n 0.00916868f $X=5.18 $Y=1.95 $X2=0 $Y2=0
cc_382 N_A_586_257#_c_430_n N_B_c_581_n 0.00619499f $X=5.855 $Y=2.035 $X2=0
+ $Y2=0
cc_383 N_A_586_257#_c_426_n N_B_c_581_n 0.00269178f $X=5.25 $Y=0.812 $X2=0 $Y2=0
cc_384 N_A_586_257#_c_423_n N_B_c_593_n 0.0031496f $X=5.18 $Y=1.95 $X2=0 $Y2=0
cc_385 N_A_586_257#_c_430_n N_B_c_593_n 0.0165f $X=5.855 $Y=2.035 $X2=0 $Y2=0
cc_386 N_A_586_257#_M1019_g N_B_c_582_n 0.00796434f $X=3.02 $Y=2.23 $X2=0 $Y2=0
cc_387 N_A_586_257#_c_411_n N_B_c_583_n 0.0147851f $X=3.02 $Y=1.375 $X2=0 $Y2=0
cc_388 N_A_586_257#_M1029_g N_B_c_583_n 0.0387754f $X=4.09 $Y=2.23 $X2=0 $Y2=0
cc_389 N_A_586_257#_c_420_n N_B_c_584_n 0.0106025f $X=5.095 $Y=0.79 $X2=0 $Y2=0
cc_390 N_A_586_257#_c_423_n N_B_c_584_n 0.0499366f $X=5.18 $Y=1.95 $X2=0 $Y2=0
cc_391 N_A_586_257#_c_431_n N_B_c_584_n 0.0115604f $X=5.265 $Y=2.035 $X2=0 $Y2=0
cc_392 N_A_586_257#_M1035_g N_B_c_585_n 0.00164105f $X=4.015 $Y=0.97 $X2=0 $Y2=0
cc_393 N_A_586_257#_c_418_n N_B_c_585_n 0.012188f $X=4.06 $Y=1.515 $X2=0 $Y2=0
cc_394 N_A_586_257#_c_420_n N_B_c_585_n 0.00280668f $X=5.095 $Y=0.79 $X2=0 $Y2=0
cc_395 N_A_586_257#_c_423_n N_B_c_585_n 0.0125365f $X=5.18 $Y=1.95 $X2=0 $Y2=0
cc_396 N_A_586_257#_M1029_g N_B_c_598_n 0.012188f $X=4.09 $Y=2.23 $X2=0 $Y2=0
cc_397 N_A_586_257#_c_423_n N_B_c_598_n 0.00481635f $X=5.18 $Y=1.95 $X2=0 $Y2=0
cc_398 N_A_586_257#_c_431_n N_B_c_598_n 0.00471f $X=5.265 $Y=2.035 $X2=0 $Y2=0
cc_399 N_A_586_257#_M1029_g B 6.22863e-19 $X=4.09 $Y=2.23 $X2=0 $Y2=0
cc_400 N_A_586_257#_c_431_n B 0.00491516f $X=5.265 $Y=2.035 $X2=0 $Y2=0
cc_401 N_A_586_257#_c_414_n N_B_c_586_n 0.00407633f $X=3.94 $Y=0.205 $X2=0 $Y2=0
cc_402 N_A_586_257#_c_419_n N_B_c_586_n 0.00413008f $X=4.22 $Y=0.375 $X2=0 $Y2=0
cc_403 N_A_586_257#_c_420_n N_B_c_586_n 0.016111f $X=5.095 $Y=0.79 $X2=0 $Y2=0
cc_404 N_A_586_257#_c_422_n N_B_c_586_n 0.00803714f $X=5.24 $Y=0.495 $X2=0 $Y2=0
cc_405 N_A_586_257#_c_423_n N_B_c_586_n 0.0101534f $X=5.18 $Y=1.95 $X2=0 $Y2=0
cc_406 N_A_586_257#_c_424_n N_B_c_586_n 0.00440876f $X=5.405 $Y=0.34 $X2=0 $Y2=0
cc_407 N_A_586_257#_c_426_n N_B_c_586_n 0.00193266f $X=5.25 $Y=0.812 $X2=0 $Y2=0
cc_408 N_A_586_257#_c_470_p N_A_531_362#_c_726_n 8.30687e-19 $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_409 N_A_586_257#_c_470_p N_A_531_362#_M1000_g 0.00112325f $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_410 N_A_586_257#_c_432_n N_A_531_362#_M1000_g 0.00597566f $X=5.94 $Y=2.815
+ $X2=0 $Y2=0
cc_411 N_A_586_257#_c_425_n N_A_531_362#_c_728_n 0.00999979f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_412 N_A_586_257#_c_425_n N_A_531_362#_M1041_g 0.00116683f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_413 N_A_586_257#_M1019_g N_A_531_362#_c_748_n 0.00646307f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_414 N_A_586_257#_c_414_n N_A_531_362#_c_732_n 0.00269116f $X=3.94 $Y=0.205
+ $X2=0 $Y2=0
cc_415 N_A_586_257#_M1035_g N_A_531_362#_c_732_n 0.00268889f $X=4.015 $Y=0.97
+ $X2=0 $Y2=0
cc_416 N_A_586_257#_M1029_g N_A_531_362#_c_732_n 3.68163e-19 $X=4.09 $Y=2.23
+ $X2=0 $Y2=0
cc_417 N_A_586_257#_c_419_n N_A_531_362#_c_732_n 0.00349151f $X=4.22 $Y=0.375
+ $X2=0 $Y2=0
cc_418 N_A_586_257#_c_423_n N_A_531_362#_c_733_n 0.022718f $X=5.18 $Y=1.95 $X2=0
+ $Y2=0
cc_419 N_A_586_257#_c_430_n N_A_531_362#_c_733_n 0.00316141f $X=5.855 $Y=2.035
+ $X2=0 $Y2=0
cc_420 N_A_586_257#_c_425_n N_A_531_362#_c_733_n 0.00987192f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_421 N_A_586_257#_c_423_n N_A_531_362#_c_734_n 0.00185163f $X=5.18 $Y=1.95
+ $X2=0 $Y2=0
cc_422 N_A_586_257#_c_430_n N_A_531_362#_c_734_n 4.59916e-19 $X=5.855 $Y=2.035
+ $X2=0 $Y2=0
cc_423 N_A_586_257#_c_425_n N_A_531_362#_c_734_n 0.00528412f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_424 N_A_586_257#_M1019_g N_A_531_362#_c_736_n 0.00316228f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_425 N_A_586_257#_c_423_n N_A_531_362#_c_737_n 0.0170417f $X=5.18 $Y=1.95
+ $X2=0 $Y2=0
cc_426 N_A_586_257#_c_430_n N_A_531_362#_c_737_n 0.00271436f $X=5.855 $Y=2.035
+ $X2=0 $Y2=0
cc_427 N_A_586_257#_M1029_g N_A_531_362#_c_738_n 0.00667835f $X=4.09 $Y=2.23
+ $X2=0 $Y2=0
cc_428 N_A_586_257#_c_418_n N_A_531_362#_c_738_n 0.00192343f $X=4.06 $Y=1.515
+ $X2=0 $Y2=0
cc_429 N_A_586_257#_M1019_g N_A_531_362#_c_739_n 0.0122378f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_430 N_A_586_257#_M1029_g N_A_531_362#_c_740_n 0.0109826f $X=4.09 $Y=2.23
+ $X2=0 $Y2=0
cc_431 N_A_586_257#_c_418_n N_A_531_362#_c_740_n 0.00274966f $X=4.06 $Y=1.515
+ $X2=0 $Y2=0
cc_432 N_A_586_257#_c_423_n N_A_531_362#_c_741_n 0.00262178f $X=5.18 $Y=1.95
+ $X2=0 $Y2=0
cc_433 N_A_586_257#_c_430_n N_A_531_362#_c_741_n 0.00260289f $X=5.855 $Y=2.035
+ $X2=0 $Y2=0
cc_434 N_A_586_257#_c_423_n N_A_531_362#_c_742_n 0.0282409f $X=5.18 $Y=1.95
+ $X2=0 $Y2=0
cc_435 N_A_586_257#_c_430_n N_A_531_362#_c_742_n 0.0113501f $X=5.855 $Y=2.035
+ $X2=0 $Y2=0
cc_436 N_A_586_257#_c_425_n N_A_536_114#_M1040_g 0.0133649f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_437 N_A_586_257#_c_425_n N_A_536_114#_c_932_n 0.0114204f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_438 N_A_586_257#_c_425_n N_A_536_114#_M1026_g 0.0133313f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_439 N_A_586_257#_M1030_g N_A_536_114#_c_954_n 0.00789174f $X=3.035 $Y=0.89
+ $X2=0 $Y2=0
cc_440 N_A_586_257#_c_411_n N_A_536_114#_c_937_n 0.00233382f $X=3.02 $Y=1.375
+ $X2=0 $Y2=0
cc_441 N_A_586_257#_M1019_g N_A_536_114#_c_937_n 0.0016671f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_442 N_A_586_257#_M1030_g N_A_536_114#_c_937_n 0.00737443f $X=3.035 $Y=0.89
+ $X2=0 $Y2=0
cc_443 N_A_586_257#_c_411_n N_A_536_114#_c_938_n 0.00212801f $X=3.02 $Y=1.375
+ $X2=0 $Y2=0
cc_444 N_A_586_257#_M1019_g N_A_536_114#_c_938_n 7.91705e-19 $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_445 N_A_586_257#_M1030_g N_A_536_114#_c_938_n 0.00102588f $X=3.035 $Y=0.89
+ $X2=0 $Y2=0
cc_446 N_A_586_257#_M1019_g N_A_536_114#_c_939_n 0.00514678f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_447 N_A_586_257#_M1019_g N_A_536_114#_c_962_n 0.00182484f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_448 N_A_586_257#_M1010_d N_A_536_114#_c_948_n 0.00582967f $X=5.805 $Y=1.84
+ $X2=0 $Y2=0
cc_449 N_A_586_257#_M1029_g N_A_536_114#_c_948_n 0.00230085f $X=4.09 $Y=2.23
+ $X2=0 $Y2=0
cc_450 N_A_586_257#_c_430_n N_A_536_114#_c_948_n 0.0297432f $X=5.855 $Y=2.035
+ $X2=0 $Y2=0
cc_451 N_A_586_257#_c_431_n N_A_536_114#_c_948_n 0.0121663f $X=5.265 $Y=2.035
+ $X2=0 $Y2=0
cc_452 N_A_586_257#_c_470_p N_A_536_114#_c_948_n 0.0141241f $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_453 N_A_586_257#_M1019_g N_A_536_114#_c_968_n 4.3363e-19 $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_454 N_A_586_257#_M1029_g N_A_536_114#_c_969_n 0.00252029f $X=4.09 $Y=2.23
+ $X2=0 $Y2=0
cc_455 N_A_586_257#_c_432_n N_A_1378_125#_c_1140_n 0.0529708f $X=5.94 $Y=2.815
+ $X2=0 $Y2=0
cc_456 N_A_586_257#_c_470_p N_A_1378_125#_c_1132_n 0.00135599f $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_457 N_A_586_257#_c_432_n N_A_1378_125#_c_1155_n 0.00592118f $X=5.94 $Y=2.815
+ $X2=0 $Y2=0
cc_458 N_A_586_257#_c_425_n N_A_1378_125#_c_1156_n 0.00155742f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_459 N_A_586_257#_c_470_p N_A_1378_125#_c_1157_n 0.00976375f $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_460 N_A_586_257#_c_432_n N_A_1378_125#_c_1157_n 0.00209431f $X=5.94 $Y=2.815
+ $X2=0 $Y2=0
cc_461 N_A_586_257#_M1026_d N_A_1268_379#_c_1353_n 0.00930497f $X=7.81 $Y=0.735
+ $X2=0 $Y2=0
cc_462 N_A_586_257#_M1026_d N_A_1278_102#_c_1564_n 0.00762323f $X=7.81 $Y=0.735
+ $X2=0 $Y2=0
cc_463 N_A_586_257#_c_425_n N_A_1278_102#_c_1567_n 0.0157411f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_464 N_A_586_257#_c_425_n N_A_1278_102#_c_1573_n 0.123842f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_465 N_A_586_257#_c_430_n N_VPWR_M1010_s 0.00470819f $X=5.855 $Y=2.035 $X2=0
+ $Y2=0
cc_466 N_A_586_257#_c_430_n N_VPWR_c_1778_n 0.0197151f $X=5.855 $Y=2.035 $X2=0
+ $Y2=0
cc_467 N_A_586_257#_c_432_n N_VPWR_c_1778_n 0.0233699f $X=5.94 $Y=2.815 $X2=0
+ $Y2=0
cc_468 N_A_586_257#_c_432_n N_VPWR_c_1795_n 0.00749631f $X=5.94 $Y=2.815 $X2=0
+ $Y2=0
cc_469 N_A_586_257#_M1029_g N_VPWR_c_1776_n 0.00106495f $X=4.09 $Y=2.23 $X2=0
+ $Y2=0
cc_470 N_A_586_257#_c_432_n N_VPWR_c_1776_n 0.0062048f $X=5.94 $Y=2.815 $X2=0
+ $Y2=0
cc_471 N_A_586_257#_M1019_g N_A_200_74#_c_1955_n 0.00834507f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_472 N_A_586_257#_M1030_g N_A_200_74#_c_1948_n 0.0142833f $X=3.035 $Y=0.89
+ $X2=0 $Y2=0
cc_473 N_A_586_257#_c_414_n N_A_200_74#_c_1948_n 0.0119842f $X=3.94 $Y=0.205
+ $X2=0 $Y2=0
cc_474 N_A_586_257#_c_415_n N_A_200_74#_c_1948_n 0.00214615f $X=3.11 $Y=0.205
+ $X2=0 $Y2=0
cc_475 N_A_586_257#_c_419_n N_A_200_74#_c_1948_n 0.0051397f $X=4.22 $Y=0.375
+ $X2=0 $Y2=0
cc_476 N_A_586_257#_M1030_g N_A_200_74#_c_1950_n 0.00566822f $X=3.035 $Y=0.89
+ $X2=0 $Y2=0
cc_477 N_A_586_257#_c_414_n N_A_200_74#_c_1950_n 0.00203445f $X=3.94 $Y=0.205
+ $X2=0 $Y2=0
cc_478 N_A_586_257#_c_419_n N_A_200_74#_c_1950_n 0.00575387f $X=4.22 $Y=0.375
+ $X2=0 $Y2=0
cc_479 N_A_586_257#_M1019_g N_A_200_74#_c_1956_n 4.30617e-19 $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_480 N_A_586_257#_c_421_n N_A_430_362#_M1035_d 0.00298848f $X=4.385 $Y=0.79
+ $X2=0 $Y2=0
cc_481 N_A_586_257#_M1019_g N_A_430_362#_c_2067_n 7.41077e-19 $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_482 N_A_586_257#_M1019_g N_A_430_362#_c_2058_n 0.013998f $X=3.02 $Y=2.23
+ $X2=0 $Y2=0
cc_483 N_A_586_257#_M1029_g N_A_430_362#_c_2058_n 0.0123666f $X=4.09 $Y=2.23
+ $X2=0 $Y2=0
cc_484 N_A_586_257#_c_414_n N_A_430_362#_c_2054_n 9.69313e-19 $X=3.94 $Y=0.205
+ $X2=0 $Y2=0
cc_485 N_A_586_257#_M1035_g N_A_430_362#_c_2054_n 0.00378878f $X=4.015 $Y=0.97
+ $X2=0 $Y2=0
cc_486 N_A_586_257#_c_418_n N_A_430_362#_c_2054_n 0.00310738f $X=4.06 $Y=1.515
+ $X2=0 $Y2=0
cc_487 N_A_586_257#_c_420_n N_A_430_362#_c_2054_n 0.00931342f $X=5.095 $Y=0.79
+ $X2=0 $Y2=0
cc_488 N_A_586_257#_c_421_n N_A_430_362#_c_2054_n 0.0218245f $X=4.385 $Y=0.79
+ $X2=0 $Y2=0
cc_489 N_A_586_257#_c_423_n N_A_430_362#_c_2054_n 0.00528634f $X=5.18 $Y=1.95
+ $X2=0 $Y2=0
cc_490 N_A_586_257#_M1035_g N_A_430_362#_c_2055_n 5.25265e-19 $X=4.015 $Y=0.97
+ $X2=0 $Y2=0
cc_491 N_A_586_257#_c_418_n N_A_430_362#_c_2055_n 0.00714519f $X=4.06 $Y=1.515
+ $X2=0 $Y2=0
cc_492 N_A_586_257#_c_426_n N_A_1183_102#_c_2137_n 0.00145282f $X=5.25 $Y=0.812
+ $X2=0 $Y2=0
cc_493 N_A_586_257#_c_422_n N_A_1183_102#_c_2139_n 0.00449343f $X=5.24 $Y=0.495
+ $X2=0 $Y2=0
cc_494 N_A_586_257#_c_425_n N_A_1183_102#_c_2139_n 0.0239506f $X=8.03 $Y=0.34
+ $X2=0 $Y2=0
cc_495 N_A_586_257#_c_426_n N_A_1183_102#_c_2139_n 0.007426f $X=5.25 $Y=0.812
+ $X2=0 $Y2=0
cc_496 N_A_586_257#_c_470_p N_A_1183_102#_c_2141_n 0.00201273f $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_497 N_A_586_257#_c_470_p N_A_1183_102#_c_2144_n 0.0101183f $X=5.94 $Y=2.12
+ $X2=0 $Y2=0
cc_498 N_A_586_257#_c_420_n N_VGND_M1025_s 0.00766383f $X=5.095 $Y=0.79 $X2=0
+ $Y2=0
cc_499 N_A_586_257#_c_414_n N_VGND_c_2355_n 0.0064857f $X=3.94 $Y=0.205 $X2=0
+ $Y2=0
cc_500 N_A_586_257#_c_419_n N_VGND_c_2355_n 0.0196201f $X=4.22 $Y=0.375 $X2=0
+ $Y2=0
cc_501 N_A_586_257#_c_420_n N_VGND_c_2355_n 0.0240041f $X=5.095 $Y=0.79 $X2=0
+ $Y2=0
cc_502 N_A_586_257#_c_424_n N_VGND_c_2355_n 0.0114116f $X=5.405 $Y=0.34 $X2=0
+ $Y2=0
cc_503 N_A_586_257#_c_415_n N_VGND_c_2365_n 0.0372813f $X=3.11 $Y=0.205 $X2=0
+ $Y2=0
cc_504 N_A_586_257#_c_419_n N_VGND_c_2365_n 0.0222109f $X=4.22 $Y=0.375 $X2=0
+ $Y2=0
cc_505 N_A_586_257#_c_420_n N_VGND_c_2365_n 0.0031456f $X=5.095 $Y=0.79 $X2=0
+ $Y2=0
cc_506 N_A_586_257#_c_420_n N_VGND_c_2367_n 0.00229474f $X=5.095 $Y=0.79 $X2=0
+ $Y2=0
cc_507 N_A_586_257#_c_424_n N_VGND_c_2367_n 0.0221883f $X=5.405 $Y=0.34 $X2=0
+ $Y2=0
cc_508 N_A_586_257#_c_425_n N_VGND_c_2367_n 0.178512f $X=8.03 $Y=0.34 $X2=0
+ $Y2=0
cc_509 N_A_586_257#_M1026_d N_VGND_c_2380_n 0.00264327f $X=7.81 $Y=0.735 $X2=0
+ $Y2=0
cc_510 N_A_586_257#_c_414_n N_VGND_c_2380_n 0.0454724f $X=3.94 $Y=0.205 $X2=0
+ $Y2=0
cc_511 N_A_586_257#_c_415_n N_VGND_c_2380_n 0.00565852f $X=3.11 $Y=0.205 $X2=0
+ $Y2=0
cc_512 N_A_586_257#_c_419_n N_VGND_c_2380_n 0.0112205f $X=4.22 $Y=0.375 $X2=0
+ $Y2=0
cc_513 N_A_586_257#_c_420_n N_VGND_c_2380_n 0.010926f $X=5.095 $Y=0.79 $X2=0
+ $Y2=0
cc_514 N_A_586_257#_c_424_n N_VGND_c_2380_n 0.012026f $X=5.405 $Y=0.34 $X2=0
+ $Y2=0
cc_515 N_A_586_257#_c_425_n N_VGND_c_2380_n 0.100401f $X=8.03 $Y=0.34 $X2=0
+ $Y2=0
cc_516 N_B_c_581_n N_A_531_362#_M1000_g 0.0146357f $X=5.625 $Y=1.69 $X2=0 $Y2=0
cc_517 N_B_c_593_n N_A_531_362#_c_745_n 0.0146357f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_518 N_B_M1033_g N_A_531_362#_c_748_n 2.39329e-19 $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_519 N_B_M1023_g N_A_531_362#_c_748_n 2.19181e-19 $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_520 N_B_M1027_g N_A_531_362#_c_732_n 0.00705094f $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_521 N_B_M1027_g N_A_531_362#_c_749_n 2.84119e-19 $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_522 N_B_M1023_g N_A_531_362#_c_749_n 8.31533e-19 $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_523 N_B_c_583_n N_A_531_362#_c_749_n 0.00348379f $X=3.6 $Y=1.735 $X2=0 $Y2=0
cc_524 N_B_c_581_n N_A_531_362#_c_733_n 0.00107287f $X=5.625 $Y=1.69 $X2=0 $Y2=0
cc_525 N_B_c_586_n N_A_531_362#_c_733_n 7.39786e-19 $X=4.867 $Y=1.22 $X2=0 $Y2=0
cc_526 N_B_c_581_n N_A_531_362#_c_734_n 0.0188089f $X=5.625 $Y=1.69 $X2=0 $Y2=0
cc_527 N_B_c_586_n N_A_531_362#_c_734_n 0.0100376f $X=4.867 $Y=1.22 $X2=0 $Y2=0
cc_528 N_B_c_583_n N_A_531_362#_c_735_n 0.00746851f $X=3.6 $Y=1.735 $X2=0 $Y2=0
cc_529 N_B_c_581_n N_A_531_362#_c_737_n 0.00123133f $X=5.625 $Y=1.69 $X2=0 $Y2=0
cc_530 N_B_c_584_n N_A_531_362#_c_737_n 0.0225642f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_531 N_B_c_585_n N_A_531_362#_c_737_n 0.0116427f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_532 N_B_M1023_g N_A_531_362#_c_738_n 2.36581e-19 $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_533 N_B_M1033_g N_A_531_362#_c_739_n 0.00162406f $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_534 N_B_M1027_g N_A_531_362#_c_739_n 4.37976e-19 $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_535 N_B_c_582_n N_A_531_362#_c_739_n 4.57847e-19 $X=2.577 $Y=1.6 $X2=0 $Y2=0
cc_536 N_B_c_581_n N_A_531_362#_c_741_n 0.00184864f $X=5.625 $Y=1.69 $X2=0 $Y2=0
cc_537 N_B_c_593_n N_A_531_362#_c_741_n 2.8248e-19 $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_538 N_B_c_581_n N_A_531_362#_c_742_n 0.00880327f $X=5.625 $Y=1.69 $X2=0 $Y2=0
cc_539 N_B_c_593_n N_A_531_362#_c_742_n 3.43025e-19 $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_540 N_B_c_585_n N_A_531_362#_c_742_n 0.00111121f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_541 N_B_M1018_g N_A_536_114#_c_954_n 0.00632239f $X=2.605 $Y=0.89 $X2=0 $Y2=0
cc_542 N_B_M1027_g N_A_536_114#_c_954_n 8.92633e-19 $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_543 N_B_M1027_g N_A_536_114#_c_937_n 0.00863311f $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_544 N_B_M1018_g N_A_536_114#_c_938_n 0.00481202f $X=2.605 $Y=0.89 $X2=0 $Y2=0
cc_545 N_B_M1027_g N_A_536_114#_c_939_n 0.00430669f $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_546 N_B_M1023_g N_A_536_114#_c_939_n 0.00254002f $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_547 N_B_c_583_n N_A_536_114#_c_939_n 0.00494864f $X=3.6 $Y=1.735 $X2=0 $Y2=0
cc_548 N_B_c_584_n N_A_536_114#_c_948_n 0.0239682f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_549 N_B_c_598_n N_A_536_114#_c_948_n 0.00678069f $X=4.8 $Y=2.065 $X2=0 $Y2=0
cc_550 B N_A_536_114#_c_948_n 0.00790442f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_551 N_B_M1023_g N_A_536_114#_c_968_n 0.00345155f $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_552 N_B_M1023_g N_A_536_114#_c_969_n 0.0103625f $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_553 N_B_c_593_n N_A_1378_125#_c_1132_n 7.84657e-19 $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_554 N_B_c_593_n N_A_1378_125#_c_1155_n 3.70581e-19 $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_555 N_B_c_593_n N_VPWR_c_1778_n 0.0146218f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_556 N_B_c_596_n N_VPWR_c_1778_n 0.00611087f $X=4.867 $Y=2.678 $X2=0 $Y2=0
cc_557 N_B_c_598_n N_VPWR_c_1778_n 0.00223913f $X=4.8 $Y=2.065 $X2=0 $Y2=0
cc_558 B N_VPWR_c_1778_n 0.053123f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_559 N_B_c_589_n N_VPWR_c_1789_n 0.0612047f $X=2.655 $Y=3.095 $X2=0 $Y2=0
cc_560 N_B_c_596_n N_VPWR_c_1789_n 0.00162283f $X=4.867 $Y=2.678 $X2=0 $Y2=0
cc_561 B N_VPWR_c_1789_n 0.0154309f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_562 N_B_M1033_g N_VPWR_c_1793_n 0.00228023f $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_563 N_B_c_593_n N_VPWR_c_1795_n 0.00460063f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_564 N_B_c_588_n N_VPWR_c_1776_n 0.0247373f $X=3.55 $Y=3.095 $X2=0 $Y2=0
cc_565 N_B_c_589_n N_VPWR_c_1776_n 0.00637935f $X=2.655 $Y=3.095 $X2=0 $Y2=0
cc_566 N_B_c_591_n N_VPWR_c_1776_n 0.0396807f $X=4.635 $Y=3.095 $X2=0 $Y2=0
cc_567 N_B_c_593_n N_VPWR_c_1776_n 0.00909416f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_568 N_B_c_595_n N_VPWR_c_1776_n 0.0111982f $X=3.64 $Y=3.095 $X2=0 $Y2=0
cc_569 N_B_c_596_n N_VPWR_c_1776_n 0.00681954f $X=4.867 $Y=2.678 $X2=0 $Y2=0
cc_570 B N_VPWR_c_1776_n 0.0160249f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_571 N_B_M1033_g N_A_200_74#_c_1946_n 7.73078e-19 $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_572 N_B_M1018_g N_A_200_74#_c_1947_n 0.00103514f $X=2.605 $Y=0.89 $X2=0 $Y2=0
cc_573 N_B_M1033_g N_A_200_74#_c_1955_n 0.0130742f $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_574 N_B_c_588_n N_A_200_74#_c_1955_n 0.00628297f $X=3.55 $Y=3.095 $X2=0 $Y2=0
cc_575 N_B_M1018_g N_A_200_74#_c_1948_n 0.00696728f $X=2.605 $Y=0.89 $X2=0 $Y2=0
cc_576 N_B_M1027_g N_A_200_74#_c_1950_n 0.0038515f $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_577 N_B_M1033_g N_A_200_74#_c_1956_n 0.00435791f $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_578 N_B_c_588_n N_A_200_74#_c_1956_n 0.00710348f $X=3.55 $Y=3.095 $X2=0 $Y2=0
cc_579 N_B_M1023_g N_A_200_74#_c_1956_n 0.0116368f $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_580 N_B_M1033_g N_A_430_362#_c_2067_n 0.00530181f $X=2.565 $Y=2.23 $X2=0
+ $Y2=0
cc_581 N_B_M1033_g N_A_430_362#_c_2056_n 0.00355096f $X=2.565 $Y=2.23 $X2=0
+ $Y2=0
cc_582 N_B_M1018_g N_A_430_362#_c_2053_n 0.00394831f $X=2.605 $Y=0.89 $X2=0
+ $Y2=0
cc_583 N_B_c_582_n N_A_430_362#_c_2053_n 0.00500723f $X=2.577 $Y=1.6 $X2=0 $Y2=0
cc_584 N_B_M1033_g N_A_430_362#_c_2058_n 0.0129226f $X=2.565 $Y=2.23 $X2=0 $Y2=0
cc_585 N_B_c_588_n N_A_430_362#_c_2058_n 3.25194e-19 $X=3.55 $Y=3.095 $X2=0
+ $Y2=0
cc_586 N_B_M1023_g N_A_430_362#_c_2058_n 0.0178158f $X=3.64 $Y=2.23 $X2=0 $Y2=0
cc_587 N_B_c_591_n N_A_430_362#_c_2058_n 0.00963729f $X=4.635 $Y=3.095 $X2=0
+ $Y2=0
cc_588 N_B_M1033_g N_A_430_362#_c_2086_n 8.69859e-19 $X=2.565 $Y=2.23 $X2=0
+ $Y2=0
cc_589 N_B_c_598_n N_A_430_362#_c_2060_n 0.00625368f $X=4.8 $Y=2.065 $X2=0 $Y2=0
cc_590 B N_A_430_362#_c_2060_n 0.0506083f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_591 N_B_c_584_n N_A_430_362#_c_2054_n 0.00710254f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_592 N_B_c_585_n N_A_430_362#_c_2054_n 9.95678e-19 $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_593 N_B_c_586_n N_A_430_362#_c_2054_n 0.00305391f $X=4.867 $Y=1.22 $X2=0
+ $Y2=0
cc_594 N_B_c_584_n N_A_430_362#_c_2055_n 0.0506083f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_595 N_B_c_585_n N_A_430_362#_c_2055_n 0.00625368f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_596 N_B_c_581_n N_A_1183_102#_c_2141_n 0.0012536f $X=5.625 $Y=1.69 $X2=0
+ $Y2=0
cc_597 N_B_c_581_n N_A_1183_102#_c_2144_n 0.00166313f $X=5.625 $Y=1.69 $X2=0
+ $Y2=0
cc_598 N_B_c_586_n N_VGND_c_2355_n 0.00304098f $X=4.867 $Y=1.22 $X2=0 $Y2=0
cc_599 N_B_c_586_n N_VGND_c_2367_n 0.00331702f $X=4.867 $Y=1.22 $X2=0 $Y2=0
cc_600 N_B_M1027_g N_VGND_c_2380_n 9.20682e-19 $X=3.545 $Y=0.97 $X2=0 $Y2=0
cc_601 N_B_c_586_n N_VGND_c_2380_n 0.00434026f $X=4.867 $Y=1.22 $X2=0 $Y2=0
cc_602 N_A_531_362#_M1000_g N_A_536_114#_M1040_g 7.26991e-19 $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_603 N_A_531_362#_c_728_n N_A_536_114#_M1040_g 0.0279332f $X=6.315 $Y=1.225
+ $X2=0 $Y2=0
cc_604 N_A_531_362#_M1041_g N_A_536_114#_M1040_g 0.0260519f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_605 N_A_531_362#_M1000_g N_A_536_114#_M1004_g 0.0241315f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_606 N_A_531_362#_c_744_n N_A_536_114#_M1004_g 0.0105864f $X=7.395 $Y=3.15
+ $X2=0 $Y2=0
cc_607 N_A_531_362#_c_729_n N_A_536_114#_M1004_g 0.0103287f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_608 N_A_531_362#_M1043_g N_A_536_114#_M1004_g 0.0175733f $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_609 N_A_531_362#_M1041_g N_A_536_114#_c_932_n 0.00737859f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_610 N_A_531_362#_M1041_g N_A_536_114#_M1026_g 0.0299929f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_611 N_A_531_362#_c_729_n N_A_536_114#_c_935_n 0.00977874f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_612 N_A_531_362#_M1041_g N_A_536_114#_c_935_n 0.00155237f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_613 N_A_531_362#_M1043_g N_A_536_114#_c_945_n 0.00515444f $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_614 N_A_531_362#_c_732_n N_A_536_114#_c_937_n 0.0134796f $X=3.8 $Y=0.795
+ $X2=0 $Y2=0
cc_615 N_A_531_362#_c_735_n N_A_536_114#_c_937_n 0.00473204f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_616 N_A_531_362#_c_736_n N_A_536_114#_c_937_n 0.00836826f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_617 N_A_531_362#_c_739_n N_A_536_114#_c_937_n 0.0137557f $X=3.12 $Y=1.665
+ $X2=0 $Y2=0
cc_618 N_A_531_362#_c_736_n N_A_536_114#_c_938_n 2.40749e-19 $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_619 N_A_531_362#_c_739_n N_A_536_114#_c_938_n 0.0235736f $X=3.12 $Y=1.665
+ $X2=0 $Y2=0
cc_620 N_A_531_362#_c_748_n N_A_536_114#_c_939_n 0.00557146f $X=2.79 $Y=1.955
+ $X2=0 $Y2=0
cc_621 N_A_531_362#_c_732_n N_A_536_114#_c_939_n 0.0120864f $X=3.8 $Y=0.795
+ $X2=0 $Y2=0
cc_622 N_A_531_362#_c_749_n N_A_536_114#_c_939_n 0.0143722f $X=3.885 $Y=1.657
+ $X2=0 $Y2=0
cc_623 N_A_531_362#_c_735_n N_A_536_114#_c_939_n 0.0150315f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_624 N_A_531_362#_c_736_n N_A_536_114#_c_939_n 0.00279507f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_625 N_A_531_362#_c_738_n N_A_536_114#_c_939_n 9.29394e-19 $X=4.225 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_531_362#_c_739_n N_A_536_114#_c_939_n 0.0159739f $X=3.12 $Y=1.665
+ $X2=0 $Y2=0
cc_627 N_A_531_362#_c_748_n N_A_536_114#_c_962_n 0.00642163f $X=2.79 $Y=1.955
+ $X2=0 $Y2=0
cc_628 N_A_531_362#_M1000_g N_A_536_114#_c_948_n 0.00417072f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_629 N_A_531_362#_c_749_n N_A_536_114#_c_948_n 6.05036e-19 $X=3.885 $Y=1.657
+ $X2=0 $Y2=0
cc_630 N_A_531_362#_c_733_n N_A_536_114#_c_948_n 8.13645e-19 $X=5.64 $Y=1.21
+ $X2=0 $Y2=0
cc_631 N_A_531_362#_c_735_n N_A_536_114#_c_948_n 0.0129499f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_632 N_A_531_362#_c_737_n N_A_536_114#_c_948_n 0.0825934f $X=5.375 $Y=1.665
+ $X2=0 $Y2=0
cc_633 N_A_531_362#_c_738_n N_A_536_114#_c_948_n 0.0248843f $X=4.225 $Y=1.665
+ $X2=0 $Y2=0
cc_634 N_A_531_362#_c_740_n N_A_536_114#_c_948_n 0.00116792f $X=4.08 $Y=1.665
+ $X2=0 $Y2=0
cc_635 N_A_531_362#_c_741_n N_A_536_114#_c_948_n 0.0233591f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_636 N_A_531_362#_c_742_n N_A_536_114#_c_948_n 2.40735e-19 $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_637 N_A_531_362#_c_748_n N_A_536_114#_c_968_n 0.00106211f $X=2.79 $Y=1.955
+ $X2=0 $Y2=0
cc_638 N_A_531_362#_c_735_n N_A_536_114#_c_968_n 0.0241992f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_639 N_A_531_362#_c_729_n N_A_536_114#_c_1019_n 0.00125149f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_640 N_A_531_362#_M1000_g N_A_536_114#_c_940_n 0.0142342f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_641 N_A_531_362#_M1041_g N_A_536_114#_c_940_n 0.0205221f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_642 N_A_531_362#_M1000_g N_A_536_114#_c_941_n 0.0014699f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_643 N_A_531_362#_c_729_n N_A_536_114#_c_941_n 0.00136801f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_644 N_A_531_362#_M1041_g N_A_536_114#_c_941_n 0.00317368f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_645 N_A_531_362#_M1043_g N_A_536_114#_c_941_n 4.81894e-19 $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_646 N_A_531_362#_c_749_n N_A_536_114#_c_969_n 0.0102151f $X=3.885 $Y=1.657
+ $X2=0 $Y2=0
cc_647 N_A_531_362#_c_735_n N_A_536_114#_c_969_n 0.00306143f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_648 N_A_531_362#_c_738_n N_A_536_114#_c_969_n 5.80029e-19 $X=4.225 $Y=1.665
+ $X2=0 $Y2=0
cc_649 N_A_531_362#_c_740_n N_A_536_114#_c_969_n 0.00740799f $X=4.08 $Y=1.665
+ $X2=0 $Y2=0
cc_650 N_A_531_362#_M1000_g N_A_1378_125#_c_1140_n 0.0199884f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_651 N_A_531_362#_M1000_g N_A_1378_125#_c_1132_n 0.0128376f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_652 N_A_531_362#_c_731_n N_A_1378_125#_c_1132_n 0.00536743f $X=6.275 $Y=1.3
+ $X2=0 $Y2=0
cc_653 N_A_531_362#_M1000_g N_A_1378_125#_c_1155_n 0.00804942f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_654 N_A_531_362#_c_744_n N_A_1378_125#_c_1155_n 2.05582e-19 $X=7.395 $Y=3.15
+ $X2=0 $Y2=0
cc_655 N_A_531_362#_c_745_n N_A_1378_125#_c_1155_n 0.00124206f $X=6.34 $Y=3.15
+ $X2=0 $Y2=0
cc_656 N_A_531_362#_c_728_n N_A_1378_125#_c_1156_n 0.00672781f $X=6.315 $Y=1.225
+ $X2=0 $Y2=0
cc_657 N_A_531_362#_M1043_g N_A_1378_125#_c_1142_n 0.0222111f $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_658 N_A_531_362#_M1000_g N_A_1378_125#_c_1143_n 2.96297e-19 $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_659 N_A_531_362#_c_729_n N_A_1378_125#_c_1133_n 0.0195087f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_660 N_A_531_362#_M1000_g N_A_1378_125#_c_1157_n 0.00777904f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_661 N_A_531_362#_M1041_g N_A_1378_125#_c_1172_n 0.00289517f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_662 N_A_531_362#_c_744_n N_A_1378_125#_c_1148_n 0.0177136f $X=7.395 $Y=3.15
+ $X2=0 $Y2=0
cc_663 N_A_531_362#_c_729_n N_A_1268_379#_c_1368_n 0.00576827f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_664 N_A_531_362#_M1043_g N_A_1268_379#_c_1368_n 0.00850357f $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_665 N_A_531_362#_c_729_n N_A_1268_379#_c_1352_n 0.0136784f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_666 N_A_531_362#_M1043_g N_A_1268_379#_c_1352_n 0.00868701f $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_667 N_A_531_362#_M1000_g N_A_1268_379#_c_1365_n 0.00146275f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_668 N_A_531_362#_M1043_g N_A_1268_379#_c_1365_n 8.40045e-19 $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_669 N_A_531_362#_c_729_n N_A_1268_379#_c_1358_n 0.00119706f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_670 N_A_531_362#_M1041_g N_A_1268_379#_c_1358_n 0.00775771f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_671 N_A_531_362#_M1041_g N_A_1278_102#_c_1564_n 0.0136367f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_672 N_A_531_362#_c_728_n N_A_1278_102#_c_1573_n 0.00288518f $X=6.315 $Y=1.225
+ $X2=0 $Y2=0
cc_673 N_A_531_362#_M1043_g N_A_1278_102#_c_1582_n 9.7128e-19 $X=7.485 $Y=2.535
+ $X2=0 $Y2=0
cc_674 N_A_531_362#_M1000_g N_VPWR_c_1778_n 5.45431e-19 $X=6.25 $Y=2.315 $X2=0
+ $Y2=0
cc_675 N_A_531_362#_c_745_n N_VPWR_c_1778_n 0.00232909f $X=6.34 $Y=3.15 $X2=0
+ $Y2=0
cc_676 N_A_531_362#_c_745_n N_VPWR_c_1795_n 0.0309847f $X=6.34 $Y=3.15 $X2=0
+ $Y2=0
cc_677 N_A_531_362#_c_744_n N_VPWR_c_1776_n 0.0315693f $X=7.395 $Y=3.15 $X2=0
+ $Y2=0
cc_678 N_A_531_362#_c_745_n N_VPWR_c_1776_n 0.00803917f $X=6.34 $Y=3.15 $X2=0
+ $Y2=0
cc_679 N_A_531_362#_M1033_d N_A_200_74#_c_1955_n 0.00171563f $X=2.655 $Y=1.81
+ $X2=0 $Y2=0
cc_680 N_A_531_362#_c_732_n N_A_200_74#_c_1950_n 0.0103425f $X=3.8 $Y=0.795
+ $X2=0 $Y2=0
cc_681 N_A_531_362#_c_735_n N_A_200_74#_c_1950_n 3.85053e-19 $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_682 N_A_531_362#_c_748_n N_A_430_362#_c_2056_n 0.0115171f $X=2.79 $Y=1.955
+ $X2=0 $Y2=0
cc_683 N_A_531_362#_c_748_n N_A_430_362#_c_2053_n 5.97682e-19 $X=2.79 $Y=1.955
+ $X2=0 $Y2=0
cc_684 N_A_531_362#_c_736_n N_A_430_362#_c_2053_n 9.67639e-19 $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_685 N_A_531_362#_c_739_n N_A_430_362#_c_2053_n 0.014194f $X=3.12 $Y=1.665
+ $X2=0 $Y2=0
cc_686 N_A_531_362#_M1033_d N_A_430_362#_c_2058_n 0.00329713f $X=2.655 $Y=1.81
+ $X2=0 $Y2=0
cc_687 N_A_531_362#_c_748_n N_A_430_362#_c_2058_n 0.0144417f $X=2.79 $Y=1.955
+ $X2=0 $Y2=0
cc_688 N_A_531_362#_c_735_n N_A_430_362#_c_2058_n 0.00377063f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_689 N_A_531_362#_c_736_n N_A_430_362#_c_2058_n 0.00654775f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_690 N_A_531_362#_c_739_n N_A_430_362#_c_2058_n 0.0039944f $X=3.12 $Y=1.665
+ $X2=0 $Y2=0
cc_691 N_A_531_362#_c_740_n N_A_430_362#_c_2058_n 0.00172575f $X=4.08 $Y=1.665
+ $X2=0 $Y2=0
cc_692 N_A_531_362#_c_737_n N_A_430_362#_c_2059_n 0.0015291f $X=5.375 $Y=1.665
+ $X2=0 $Y2=0
cc_693 N_A_531_362#_c_732_n N_A_430_362#_c_2054_n 0.0105543f $X=3.8 $Y=0.795
+ $X2=0 $Y2=0
cc_694 N_A_531_362#_c_737_n N_A_430_362#_c_2054_n 0.00376865f $X=5.375 $Y=1.665
+ $X2=0 $Y2=0
cc_695 N_A_531_362#_c_738_n N_A_430_362#_c_2054_n 0.00500911f $X=4.225 $Y=1.665
+ $X2=0 $Y2=0
cc_696 N_A_531_362#_c_740_n N_A_430_362#_c_2054_n 0.00443325f $X=4.08 $Y=1.665
+ $X2=0 $Y2=0
cc_697 N_A_531_362#_c_732_n N_A_430_362#_c_2055_n 0.00914317f $X=3.8 $Y=0.795
+ $X2=0 $Y2=0
cc_698 N_A_531_362#_c_737_n N_A_430_362#_c_2055_n 0.0105541f $X=5.375 $Y=1.665
+ $X2=0 $Y2=0
cc_699 N_A_531_362#_c_738_n N_A_430_362#_c_2055_n 0.00311445f $X=4.225 $Y=1.665
+ $X2=0 $Y2=0
cc_700 N_A_531_362#_c_740_n N_A_430_362#_c_2055_n 0.0141676f $X=4.08 $Y=1.665
+ $X2=0 $Y2=0
cc_701 N_A_531_362#_c_726_n N_A_1183_102#_c_2137_n 0.0133355f $X=6.16 $Y=1.3
+ $X2=0 $Y2=0
cc_702 N_A_531_362#_M1000_g N_A_1183_102#_c_2137_n 0.00416118f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_703 N_A_531_362#_c_728_n N_A_1183_102#_c_2137_n 0.0040557f $X=6.315 $Y=1.225
+ $X2=0 $Y2=0
cc_704 N_A_531_362#_c_733_n N_A_1183_102#_c_2137_n 0.0209267f $X=5.64 $Y=1.21
+ $X2=0 $Y2=0
cc_705 N_A_531_362#_c_734_n N_A_1183_102#_c_2137_n 0.00154856f $X=5.64 $Y=1.21
+ $X2=0 $Y2=0
cc_706 N_A_531_362#_c_742_n N_A_1183_102#_c_2137_n 0.00825969f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_707 N_A_531_362#_c_726_n N_A_1183_102#_c_2139_n 0.00374179f $X=6.16 $Y=1.3
+ $X2=0 $Y2=0
cc_708 N_A_531_362#_c_726_n N_A_1183_102#_c_2140_n 2.87966e-19 $X=6.16 $Y=1.3
+ $X2=0 $Y2=0
cc_709 N_A_531_362#_M1000_g N_A_1183_102#_c_2140_n 0.00803195f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_710 N_A_531_362#_c_729_n N_A_1183_102#_c_2140_n 0.00468925f $X=7.245 $Y=1.67
+ $X2=0 $Y2=0
cc_711 N_A_531_362#_M1041_g N_A_1183_102#_c_2140_n 0.00679529f $X=7.245 $Y=0.945
+ $X2=0 $Y2=0
cc_712 N_A_531_362#_c_726_n N_A_1183_102#_c_2141_n 0.00277597f $X=6.16 $Y=1.3
+ $X2=0 $Y2=0
cc_713 N_A_531_362#_c_741_n N_A_1183_102#_c_2141_n 0.0222478f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_714 N_A_531_362#_c_742_n N_A_1183_102#_c_2141_n 0.00121051f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_715 N_A_531_362#_c_726_n N_A_1183_102#_c_2144_n 0.00288449f $X=6.16 $Y=1.3
+ $X2=0 $Y2=0
cc_716 N_A_531_362#_M1000_g N_A_1183_102#_c_2144_n 0.00278366f $X=6.25 $Y=2.315
+ $X2=0 $Y2=0
cc_717 N_A_531_362#_c_741_n N_A_1183_102#_c_2144_n 8.8892e-19 $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_718 N_A_531_362#_c_742_n N_A_1183_102#_c_2144_n 0.0106479f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_719 N_A_531_362#_c_732_n N_VGND_c_2365_n 0.00343252f $X=3.8 $Y=0.795 $X2=0
+ $Y2=0
cc_720 N_A_531_362#_c_728_n N_VGND_c_2367_n 6.91459e-19 $X=6.315 $Y=1.225 $X2=0
+ $Y2=0
cc_721 N_A_531_362#_c_732_n N_VGND_c_2380_n 0.00445579f $X=3.8 $Y=0.795 $X2=0
+ $Y2=0
cc_722 N_A_536_114#_c_1019_n N_A_1378_125#_M1004_d 0.00345455f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_723 N_A_536_114#_c_941_n N_A_1378_125#_M1004_d 0.00243306f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_724 N_A_536_114#_c_944_n N_A_1378_125#_M1016_g 0.0298911f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_725 N_A_536_114#_M1026_g N_A_1378_125#_c_1130_n 0.00348748f $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_726 N_A_536_114#_c_944_n N_A_1378_125#_c_1130_n 0.01821f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_727 N_A_536_114#_c_936_n N_A_1378_125#_c_1130_n 0.0109628f $X=7.89 $Y=1.525
+ $X2=0 $Y2=0
cc_728 N_A_536_114#_M1004_g N_A_1378_125#_c_1140_n 0.00101754f $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_729 N_A_536_114#_c_948_n N_A_1378_125#_c_1140_n 0.00190547f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_730 N_A_536_114#_M1040_g N_A_1378_125#_c_1132_n 0.00365823f $X=6.815 $Y=0.945
+ $X2=0 $Y2=0
cc_731 N_A_536_114#_M1004_g N_A_1378_125#_c_1132_n 6.67674e-19 $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_732 N_A_536_114#_c_948_n N_A_1378_125#_c_1132_n 0.00350009f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_733 N_A_536_114#_c_1019_n N_A_1378_125#_c_1132_n 2.31446e-19 $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_734 N_A_536_114#_c_940_n N_A_1378_125#_c_1132_n 0.00197208f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_735 N_A_536_114#_c_941_n N_A_1378_125#_c_1132_n 0.0430354f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_736 N_A_536_114#_M1004_g N_A_1378_125#_c_1143_n 0.00243847f $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_737 N_A_536_114#_c_935_n N_A_1378_125#_c_1133_n 0.0106656f $X=7.89 $Y=1.89
+ $X2=0 $Y2=0
cc_738 N_A_536_114#_c_945_n N_A_1378_125#_c_1133_n 0.00953145f $X=7.965 $Y=1.965
+ $X2=0 $Y2=0
cc_739 N_A_536_114#_c_946_n N_A_1378_125#_c_1133_n 0.00222845f $X=8.435 $Y=2.04
+ $X2=0 $Y2=0
cc_740 N_A_536_114#_c_935_n N_A_1378_125#_c_1192_n 7.88981e-19 $X=7.89 $Y=1.89
+ $X2=0 $Y2=0
cc_741 N_A_536_114#_c_936_n N_A_1378_125#_c_1192_n 0.00842362f $X=7.89 $Y=1.525
+ $X2=0 $Y2=0
cc_742 N_A_536_114#_c_946_n N_A_1378_125#_c_1145_n 0.0135627f $X=8.435 $Y=2.04
+ $X2=0 $Y2=0
cc_743 N_A_536_114#_M1026_g N_A_1378_125#_c_1134_n 5.07384e-19 $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_744 N_A_536_114#_c_944_n N_A_1378_125#_c_1134_n 0.00188466f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_745 N_A_536_114#_M1004_g N_A_1378_125#_c_1157_n 4.25583e-19 $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_746 N_A_536_114#_c_948_n N_A_1378_125#_c_1157_n 0.0148436f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_A_536_114#_c_1019_n N_A_1378_125#_c_1157_n 2.36937e-19 $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_A_536_114#_c_941_n N_A_1378_125#_c_1157_n 0.0120703f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_749 N_A_536_114#_M1040_g N_A_1378_125#_c_1172_n 0.00169538f $X=6.815 $Y=0.945
+ $X2=0 $Y2=0
cc_750 N_A_536_114#_c_940_n N_A_1378_125#_c_1172_n 3.46431e-19 $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_751 N_A_536_114#_M1040_g N_A_1378_125#_c_1203_n 0.0082901f $X=6.815 $Y=0.945
+ $X2=0 $Y2=0
cc_752 N_A_536_114#_c_940_n N_A_1378_125#_c_1203_n 0.00140147f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_753 N_A_536_114#_c_941_n N_A_1378_125#_c_1203_n 0.0252002f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_754 N_A_536_114#_M1004_g N_A_1378_125#_c_1148_n 0.00190574f $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_755 N_A_536_114#_c_946_n N_A_1378_125#_c_1149_n 0.0017775f $X=8.435 $Y=2.04
+ $X2=0 $Y2=0
cc_756 N_A_536_114#_c_935_n N_A_1378_125#_c_1137_n 0.00287462f $X=7.89 $Y=1.89
+ $X2=0 $Y2=0
cc_757 N_A_536_114#_c_944_n N_A_1378_125#_c_1137_n 0.00525621f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_758 N_A_536_114#_c_936_n N_A_1378_125#_c_1137_n 0.00320778f $X=7.89 $Y=1.525
+ $X2=0 $Y2=0
cc_759 N_A_536_114#_c_946_n N_A_1378_125#_c_1150_n 0.00171724f $X=8.435 $Y=2.04
+ $X2=0 $Y2=0
cc_760 N_A_536_114#_c_948_n N_A_1268_379#_M1000_d 0.00453557f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_A_536_114#_c_941_n N_A_1268_379#_M1000_d 0.00215817f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_762 N_A_536_114#_M1004_g N_A_1268_379#_c_1368_n 0.0103795f $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_763 N_A_536_114#_c_1019_n N_A_1268_379#_c_1368_n 0.00340501f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_A_536_114#_c_941_n N_A_1268_379#_c_1368_n 0.0157976f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_765 N_A_536_114#_M1004_g N_A_1268_379#_c_1352_n 6.03697e-19 $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_766 N_A_536_114#_M1026_g N_A_1268_379#_c_1352_n 0.00353047f $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_767 N_A_536_114#_c_935_n N_A_1268_379#_c_1352_n 7.84728e-19 $X=7.89 $Y=1.89
+ $X2=0 $Y2=0
cc_768 N_A_536_114#_c_1019_n N_A_1268_379#_c_1352_n 0.00687373f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_A_536_114#_c_941_n N_A_1268_379#_c_1352_n 0.0336475f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_770 N_A_536_114#_M1026_g N_A_1268_379#_c_1353_n 0.0108313f $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_771 N_A_536_114#_c_936_n N_A_1268_379#_c_1353_n 0.00326105f $X=7.89 $Y=1.525
+ $X2=0 $Y2=0
cc_772 N_A_536_114#_M1004_g N_A_1268_379#_c_1365_n 0.00703373f $X=6.845 $Y=2.315
+ $X2=0 $Y2=0
cc_773 N_A_536_114#_c_948_n N_A_1268_379#_c_1365_n 0.0066578f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_774 N_A_536_114#_c_940_n N_A_1268_379#_c_1365_n 7.94282e-19 $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_775 N_A_536_114#_c_941_n N_A_1268_379#_c_1365_n 0.0055304f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_776 N_A_536_114#_M1026_g N_A_1268_379#_c_1358_n 0.00944858f $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_777 N_A_536_114#_M1040_g N_A_1278_102#_c_1564_n 0.0113534f $X=6.815 $Y=0.945
+ $X2=0 $Y2=0
cc_778 N_A_536_114#_M1026_g N_A_1278_102#_c_1564_n 0.0127697f $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_779 N_A_536_114#_M1026_g N_A_1278_102#_c_1565_n 0.00387243f $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_780 N_A_536_114#_c_946_n N_A_1278_102#_c_1579_n 0.012045f $X=8.435 $Y=2.04
+ $X2=0 $Y2=0
cc_781 N_A_536_114#_M1026_g N_A_1278_102#_c_1567_n 6.08134e-19 $X=7.735 $Y=1.055
+ $X2=0 $Y2=0
cc_782 N_A_536_114#_c_944_n N_A_1278_102#_c_1582_n 0.00832282f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_783 N_A_536_114#_c_946_n N_A_1278_102#_c_1582_n 0.0105739f $X=8.435 $Y=2.04
+ $X2=0 $Y2=0
cc_784 N_A_536_114#_c_948_n N_VPWR_c_1778_n 0.00272918f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_785 N_A_536_114#_c_946_n N_VPWR_c_1795_n 0.00330849f $X=8.435 $Y=2.04 $X2=0
+ $Y2=0
cc_786 N_A_536_114#_c_946_n N_VPWR_c_1796_n 2.76574e-19 $X=8.435 $Y=2.04 $X2=0
+ $Y2=0
cc_787 N_A_536_114#_c_946_n N_VPWR_c_1776_n 0.00653145f $X=8.435 $Y=2.04 $X2=0
+ $Y2=0
cc_788 N_A_536_114#_c_937_n N_A_200_74#_M1030_d 0.00205757f $X=3.375 $Y=1.295
+ $X2=0 $Y2=0
cc_789 N_A_536_114#_c_939_n N_A_200_74#_M1019_d 0.00156646f $X=3.46 $Y=1.935
+ $X2=0 $Y2=0
cc_790 N_A_536_114#_c_962_n N_A_200_74#_M1019_d 0.00347062f $X=3.545 $Y=2.027
+ $X2=0 $Y2=0
cc_791 N_A_536_114#_c_968_n N_A_200_74#_M1019_d 0.00129587f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_792 N_A_536_114#_c_954_n N_A_200_74#_c_1948_n 0.0180331f $X=2.82 $Y=0.745
+ $X2=0 $Y2=0
cc_793 N_A_536_114#_c_937_n N_A_200_74#_c_1950_n 0.0201241f $X=3.375 $Y=1.295
+ $X2=0 $Y2=0
cc_794 N_A_536_114#_c_948_n N_A_430_362#_M1029_d 7.72498e-19 $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_795 N_A_536_114#_c_938_n N_A_430_362#_c_2053_n 0.0129693f $X=2.985 $Y=1.295
+ $X2=0 $Y2=0
cc_796 N_A_536_114#_M1023_d N_A_430_362#_c_2058_n 0.00476982f $X=3.73 $Y=1.81
+ $X2=0 $Y2=0
cc_797 N_A_536_114#_c_962_n N_A_430_362#_c_2058_n 0.00970512f $X=3.545 $Y=2.027
+ $X2=0 $Y2=0
cc_798 N_A_536_114#_c_948_n N_A_430_362#_c_2058_n 0.00811886f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_799 N_A_536_114#_c_968_n N_A_430_362#_c_2058_n 0.00741469f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_800 N_A_536_114#_c_969_n N_A_430_362#_c_2058_n 0.0232705f $X=3.865 $Y=2.025
+ $X2=0 $Y2=0
cc_801 N_A_536_114#_c_948_n N_A_430_362#_c_2059_n 0.00934256f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_802 N_A_536_114#_c_969_n N_A_430_362#_c_2059_n 0.00756748f $X=3.865 $Y=2.025
+ $X2=0 $Y2=0
cc_803 N_A_536_114#_c_948_n N_A_430_362#_c_2060_n 0.0162661f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_804 N_A_536_114#_c_968_n N_A_430_362#_c_2060_n 0.00119381f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_805 N_A_536_114#_c_968_n N_A_430_362#_c_2055_n 4.59904e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_806 N_A_536_114#_c_944_n N_A_1183_102#_c_2145_n 0.00661671f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_807 N_A_536_114#_c_935_n N_A_1183_102#_c_2140_n 0.00469594f $X=7.89 $Y=1.89
+ $X2=0 $Y2=0
cc_808 N_A_536_114#_c_944_n N_A_1183_102#_c_2140_n 0.0093148f $X=8.345 $Y=1.965
+ $X2=0 $Y2=0
cc_809 N_A_536_114#_c_936_n N_A_1183_102#_c_2140_n 0.00101843f $X=7.89 $Y=1.525
+ $X2=0 $Y2=0
cc_810 N_A_536_114#_c_948_n N_A_1183_102#_c_2140_n 0.0488037f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_811 N_A_536_114#_c_1019_n N_A_1183_102#_c_2140_n 0.0232331f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_812 N_A_536_114#_c_940_n N_A_1183_102#_c_2140_n 0.00118099f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_813 N_A_536_114#_c_941_n N_A_1183_102#_c_2140_n 0.0225784f $X=6.795 $Y=1.57
+ $X2=0 $Y2=0
cc_814 N_A_536_114#_c_948_n N_A_1183_102#_c_2141_n 0.0249507f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_815 N_A_536_114#_c_948_n N_A_1183_102#_c_2144_n 0.00105696f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_816 N_A_536_114#_c_933_n N_VGND_c_2367_n 0.0232872f $X=6.89 $Y=0.18 $X2=0
+ $Y2=0
cc_817 N_A_536_114#_c_932_n N_VGND_c_2380_n 0.0241942f $X=7.66 $Y=0.18 $X2=0
+ $Y2=0
cc_818 N_A_536_114#_c_933_n N_VGND_c_2380_n 0.00604517f $X=6.89 $Y=0.18 $X2=0
+ $Y2=0
cc_819 N_A_1378_125#_c_1132_n N_A_1268_379#_M1000_d 6.59425e-19 $X=6.4 $Y=1.98
+ $X2=0 $Y2=0
cc_820 N_A_1378_125#_c_1157_n N_A_1268_379#_M1000_d 0.0042726f $X=6.4 $Y=2.065
+ $X2=0 $Y2=0
cc_821 N_A_1378_125#_M1016_g N_A_1268_379#_M1008_g 0.011271f $X=8.97 $Y=2.34
+ $X2=0 $Y2=0
cc_822 N_A_1378_125#_c_1146_n N_A_1268_379#_M1008_g 0.0140294f $X=12.295
+ $Y=2.695 $X2=0 $Y2=0
cc_823 N_A_1378_125#_c_1146_n N_A_1268_379#_M1024_g 0.0133968f $X=12.295
+ $Y=2.695 $X2=0 $Y2=0
cc_824 N_A_1378_125#_c_1146_n N_A_1268_379#_M1036_g 0.0133831f $X=12.295
+ $Y=2.695 $X2=0 $Y2=0
cc_825 N_A_1378_125#_c_1146_n N_A_1268_379#_M1039_g 0.0146423f $X=12.295
+ $Y=2.695 $X2=0 $Y2=0
cc_826 N_A_1378_125#_M1004_d N_A_1268_379#_c_1368_n 0.00849579f $X=6.935
+ $Y=1.895 $X2=0 $Y2=0
cc_827 N_A_1378_125#_c_1142_n N_A_1268_379#_c_1368_n 0.00808319f $X=7.705 $Y=2.9
+ $X2=0 $Y2=0
cc_828 N_A_1378_125#_c_1143_n N_A_1268_379#_c_1368_n 0.0193349f $X=7.165 $Y=2.9
+ $X2=0 $Y2=0
cc_829 N_A_1378_125#_c_1133_n N_A_1268_379#_c_1368_n 0.0133618f $X=7.79 $Y=2.725
+ $X2=0 $Y2=0
cc_830 N_A_1378_125#_c_1148_n N_A_1268_379#_c_1368_n 0.00588296f $X=6.99 $Y=2.9
+ $X2=0 $Y2=0
cc_831 N_A_1378_125#_c_1133_n N_A_1268_379#_c_1352_n 0.0474384f $X=7.79 $Y=2.725
+ $X2=0 $Y2=0
cc_832 N_A_1378_125#_c_1192_n N_A_1268_379#_c_1352_n 0.0131597f $X=7.875
+ $Y=1.565 $X2=0 $Y2=0
cc_833 N_A_1378_125#_c_1134_n N_A_1268_379#_c_1352_n 0.00429305f $X=8.37
+ $Y=1.485 $X2=0 $Y2=0
cc_834 N_A_1378_125#_c_1130_n N_A_1268_379#_c_1353_n 0.0147022f $X=8.88 $Y=1.485
+ $X2=0 $Y2=0
cc_835 N_A_1378_125#_c_1192_n N_A_1268_379#_c_1353_n 0.005212f $X=7.875 $Y=1.565
+ $X2=0 $Y2=0
cc_836 N_A_1378_125#_c_1134_n N_A_1268_379#_c_1353_n 0.0294386f $X=8.37 $Y=1.485
+ $X2=0 $Y2=0
cc_837 N_A_1378_125#_c_1230_p N_A_1268_379#_c_1353_n 0.0109343f $X=8.71 $Y=1.485
+ $X2=0 $Y2=0
cc_838 N_A_1378_125#_c_1137_n N_A_1268_379#_c_1353_n 0.0115008f $X=8.205
+ $Y=1.485 $X2=0 $Y2=0
cc_839 N_A_1378_125#_c_1129_n N_A_1268_379#_c_1354_n 0.00264848f $X=9.425
+ $Y=1.32 $X2=0 $Y2=0
cc_840 N_A_1378_125#_c_1128_n N_A_1268_379#_c_1355_n 0.00244367f $X=9.35
+ $Y=1.395 $X2=0 $Y2=0
cc_841 N_A_1378_125#_c_1129_n N_A_1268_379#_c_1355_n 0.0115199f $X=9.425 $Y=1.32
+ $X2=0 $Y2=0
cc_842 N_A_1378_125#_c_1130_n N_A_1268_379#_c_1355_n 0.00471226f $X=8.88
+ $Y=1.485 $X2=0 $Y2=0
cc_843 N_A_1378_125#_c_1131_n N_A_1268_379#_c_1355_n 5.33801e-19 $X=8.97
+ $Y=1.485 $X2=0 $Y2=0
cc_844 N_A_1378_125#_c_1129_n N_A_1268_379#_c_1418_n 0.00916304f $X=9.425
+ $Y=1.32 $X2=0 $Y2=0
cc_845 N_A_1378_125#_c_1129_n N_A_1268_379#_c_1419_n 0.00857086f $X=9.425
+ $Y=1.32 $X2=0 $Y2=0
cc_846 N_A_1378_125#_c_1128_n N_A_1268_379#_c_1357_n 5.43742e-19 $X=9.35
+ $Y=1.395 $X2=0 $Y2=0
cc_847 N_A_1378_125#_c_1129_n N_A_1268_379#_c_1357_n 0.0035906f $X=9.425 $Y=1.32
+ $X2=0 $Y2=0
cc_848 N_A_1378_125#_c_1148_n N_A_1268_379#_c_1365_n 0.0163439f $X=6.99 $Y=2.9
+ $X2=0 $Y2=0
cc_849 N_A_1378_125#_c_1128_n N_A_1268_379#_c_1359_n 0.0074675f $X=9.35 $Y=1.395
+ $X2=0 $Y2=0
cc_850 N_A_1378_125#_c_1131_n N_A_1268_379#_c_1359_n 0.011271f $X=8.97 $Y=1.485
+ $X2=0 $Y2=0
cc_851 N_A_1378_125#_c_1147_n N_CI_M1034_g 0.00934009f $X=12.505 $Y=2.61 $X2=0
+ $Y2=0
cc_852 N_A_1378_125#_c_1151_n N_CI_M1034_g 0.00297355f $X=12.55 $Y=2.035 $X2=0
+ $Y2=0
cc_853 N_A_1378_125#_c_1138_n N_CI_M1034_g 0.00439592f $X=12.505 $Y=1.95 $X2=0
+ $Y2=0
cc_854 N_A_1378_125#_c_1136_n N_CI_c_1522_n 0.00113088f $X=12.69 $Y=1.095 $X2=0
+ $Y2=0
cc_855 N_A_1378_125#_c_1138_n N_CI_c_1522_n 0.00223089f $X=12.505 $Y=1.95 $X2=0
+ $Y2=0
cc_856 N_A_1378_125#_c_1136_n N_CI_c_1523_n 0.0144777f $X=12.69 $Y=1.095 $X2=0
+ $Y2=0
cc_857 N_A_1378_125#_c_1151_n N_CI_c_1523_n 0.00447259f $X=12.55 $Y=2.035 $X2=0
+ $Y2=0
cc_858 N_A_1378_125#_c_1138_n N_CI_c_1523_n 0.0342075f $X=12.505 $Y=1.95 $X2=0
+ $Y2=0
cc_859 N_A_1378_125#_c_1136_n N_CI_c_1524_n 0.00315064f $X=12.69 $Y=1.095 $X2=0
+ $Y2=0
cc_860 N_A_1378_125#_c_1138_n N_CI_c_1524_n 0.00387942f $X=12.505 $Y=1.95 $X2=0
+ $Y2=0
cc_861 N_A_1378_125#_c_1156_n N_A_1278_102#_M1021_d 4.52186e-19 $X=6.485 $Y=1.13
+ $X2=-0.19 $Y2=-0.245
cc_862 N_A_1378_125#_c_1203_n N_A_1278_102#_M1021_d 0.0048891f $X=6.865 $Y=1.115
+ $X2=-0.19 $Y2=-0.245
cc_863 N_A_1378_125#_c_1142_n N_A_1278_102#_M1043_d 0.00299756f $X=7.705 $Y=2.9
+ $X2=0 $Y2=0
cc_864 N_A_1378_125#_c_1133_n N_A_1278_102#_M1043_d 0.015495f $X=7.79 $Y=2.725
+ $X2=0 $Y2=0
cc_865 N_A_1378_125#_c_1145_n N_A_1278_102#_M1043_d 0.00984277f $X=8.545 $Y=2.99
+ $X2=0 $Y2=0
cc_866 N_A_1378_125#_c_1149_n N_A_1278_102#_M1043_d 0.00438009f $X=7.79 $Y=2.9
+ $X2=0 $Y2=0
cc_867 N_A_1378_125#_M1040_d N_A_1278_102#_c_1564_n 0.00208687f $X=6.89 $Y=0.625
+ $X2=0 $Y2=0
cc_868 N_A_1378_125#_c_1172_n N_A_1278_102#_c_1564_n 0.0116568f $X=7.03 $Y=1.11
+ $X2=0 $Y2=0
cc_869 N_A_1378_125#_c_1203_n N_A_1278_102#_c_1564_n 0.00566357f $X=6.865
+ $Y=1.115 $X2=0 $Y2=0
cc_870 N_A_1378_125#_M1016_g N_A_1278_102#_c_1579_n 0.0135751f $X=8.97 $Y=2.34
+ $X2=0 $Y2=0
cc_871 N_A_1378_125#_c_1130_n N_A_1278_102#_c_1579_n 8.09836e-19 $X=8.88
+ $Y=1.485 $X2=0 $Y2=0
cc_872 N_A_1378_125#_c_1145_n N_A_1278_102#_c_1579_n 0.00449246f $X=8.545
+ $Y=2.99 $X2=0 $Y2=0
cc_873 N_A_1378_125#_c_1230_p N_A_1278_102#_c_1579_n 0.00195716f $X=8.71
+ $Y=1.485 $X2=0 $Y2=0
cc_874 N_A_1378_125#_c_1146_n N_A_1278_102#_c_1579_n 0.203328f $X=12.295
+ $Y=2.695 $X2=0 $Y2=0
cc_875 N_A_1378_125#_c_1147_n N_A_1278_102#_c_1579_n 0.0153023f $X=12.505
+ $Y=2.61 $X2=0 $Y2=0
cc_876 N_A_1378_125#_c_1150_n N_A_1278_102#_c_1579_n 0.0104146f $X=8.63 $Y=2.695
+ $X2=0 $Y2=0
cc_877 N_A_1378_125#_c_1129_n N_A_1278_102#_c_1566_n 0.0045789f $X=9.425 $Y=1.32
+ $X2=0 $Y2=0
cc_878 N_A_1378_125#_c_1129_n N_A_1278_102#_c_1568_n 0.00449284f $X=9.425
+ $Y=1.32 $X2=0 $Y2=0
cc_879 N_A_1378_125#_c_1129_n N_A_1278_102#_c_1615_n 0.00118926f $X=9.425
+ $Y=1.32 $X2=0 $Y2=0
cc_880 N_A_1378_125#_c_1135_n N_A_1278_102#_c_1569_n 0.013906f $X=12.465
+ $Y=1.095 $X2=0 $Y2=0
cc_881 N_A_1378_125#_c_1138_n N_A_1278_102#_c_1569_n 0.0836101f $X=12.505
+ $Y=1.95 $X2=0 $Y2=0
cc_882 N_A_1378_125#_M1017_s N_A_1278_102#_c_1570_n 0.00739309f $X=12.545 $Y=0.6
+ $X2=0 $Y2=0
cc_883 N_A_1378_125#_c_1135_n N_A_1278_102#_c_1570_n 0.0143583f $X=12.465
+ $Y=1.095 $X2=0 $Y2=0
cc_884 N_A_1378_125#_c_1136_n N_A_1278_102#_c_1570_n 0.0242074f $X=12.69
+ $Y=1.095 $X2=0 $Y2=0
cc_885 N_A_1378_125#_c_1136_n N_A_1278_102#_c_1571_n 0.00727261f $X=12.69
+ $Y=1.095 $X2=0 $Y2=0
cc_886 N_A_1378_125#_c_1156_n N_A_1278_102#_c_1573_n 0.00381013f $X=6.485
+ $Y=1.13 $X2=0 $Y2=0
cc_887 N_A_1378_125#_c_1203_n N_A_1278_102#_c_1573_n 0.0130965f $X=6.865
+ $Y=1.115 $X2=0 $Y2=0
cc_888 N_A_1378_125#_M1016_g N_A_1278_102#_c_1582_n 0.00143184f $X=8.97 $Y=2.34
+ $X2=0 $Y2=0
cc_889 N_A_1378_125#_c_1133_n N_A_1278_102#_c_1582_n 0.0481667f $X=7.79 $Y=2.725
+ $X2=0 $Y2=0
cc_890 N_A_1378_125#_c_1145_n N_A_1278_102#_c_1582_n 0.020353f $X=8.545 $Y=2.99
+ $X2=0 $Y2=0
cc_891 N_A_1378_125#_c_1149_n N_A_1278_102#_c_1582_n 8.51637e-19 $X=7.79 $Y=2.9
+ $X2=0 $Y2=0
cc_892 N_A_1378_125#_c_1137_n N_A_1278_102#_c_1582_n 0.00796748f $X=8.205
+ $Y=1.485 $X2=0 $Y2=0
cc_893 N_A_1378_125#_c_1146_n N_VPWR_M1016_d 0.0146946f $X=12.295 $Y=2.695 $X2=0
+ $Y2=0
cc_894 N_A_1378_125#_c_1146_n N_VPWR_M1024_s 0.00748622f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_895 N_A_1378_125#_c_1146_n N_VPWR_M1039_s 0.017084f $X=12.295 $Y=2.695 $X2=0
+ $Y2=0
cc_896 N_A_1378_125#_c_1155_n N_VPWR_c_1778_n 0.00291357f $X=6.365 $Y=2.99 $X2=0
+ $Y2=0
cc_897 N_A_1378_125#_c_1147_n N_VPWR_c_1779_n 0.00954883f $X=12.505 $Y=2.61
+ $X2=0 $Y2=0
cc_898 N_A_1378_125#_c_1146_n N_VPWR_c_1783_n 0.0241314f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_899 N_A_1378_125#_c_1146_n N_VPWR_c_1784_n 0.0132992f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_900 N_A_1378_125#_c_1146_n N_VPWR_c_1785_n 0.00373225f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_901 N_A_1378_125#_c_1147_n N_VPWR_c_1785_n 0.0125009f $X=12.505 $Y=2.61 $X2=0
+ $Y2=0
cc_902 N_A_1378_125#_M1016_g N_VPWR_c_1795_n 0.00446568f $X=8.97 $Y=2.34 $X2=0
+ $Y2=0
cc_903 N_A_1378_125#_c_1155_n N_VPWR_c_1795_n 0.0115566f $X=6.365 $Y=2.99 $X2=0
+ $Y2=0
cc_904 N_A_1378_125#_c_1145_n N_VPWR_c_1795_n 0.0426071f $X=8.545 $Y=2.99 $X2=0
+ $Y2=0
cc_905 N_A_1378_125#_c_1146_n N_VPWR_c_1795_n 0.00728235f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_906 N_A_1378_125#_c_1148_n N_VPWR_c_1795_n 0.0880113f $X=6.99 $Y=2.9 $X2=0
+ $Y2=0
cc_907 N_A_1378_125#_c_1149_n N_VPWR_c_1795_n 0.0121505f $X=7.79 $Y=2.9 $X2=0
+ $Y2=0
cc_908 N_A_1378_125#_c_1150_n N_VPWR_c_1795_n 0.0117055f $X=8.63 $Y=2.695 $X2=0
+ $Y2=0
cc_909 N_A_1378_125#_M1016_g N_VPWR_c_1796_n 3.19911e-19 $X=8.97 $Y=2.34 $X2=0
+ $Y2=0
cc_910 N_A_1378_125#_c_1146_n N_VPWR_c_1796_n 0.0417827f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_911 N_A_1378_125#_c_1150_n N_VPWR_c_1796_n 0.00569084f $X=8.63 $Y=2.695 $X2=0
+ $Y2=0
cc_912 N_A_1378_125#_c_1146_n N_VPWR_c_1797_n 0.0132992f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_913 N_A_1378_125#_c_1146_n N_VPWR_c_1798_n 0.0462415f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_914 N_A_1378_125#_M1016_g N_VPWR_c_1776_n 0.00610055f $X=8.97 $Y=2.34 $X2=0
+ $Y2=0
cc_915 N_A_1378_125#_c_1155_n N_VPWR_c_1776_n 0.00579705f $X=6.365 $Y=2.99 $X2=0
+ $Y2=0
cc_916 N_A_1378_125#_c_1145_n N_VPWR_c_1776_n 0.0243674f $X=8.545 $Y=2.99 $X2=0
+ $Y2=0
cc_917 N_A_1378_125#_c_1146_n N_VPWR_c_1776_n 0.0669606f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_918 N_A_1378_125#_c_1147_n N_VPWR_c_1776_n 0.01431f $X=12.505 $Y=2.61 $X2=0
+ $Y2=0
cc_919 N_A_1378_125#_c_1148_n N_VPWR_c_1776_n 0.0458466f $X=6.99 $Y=2.9 $X2=0
+ $Y2=0
cc_920 N_A_1378_125#_c_1149_n N_VPWR_c_1776_n 0.00660393f $X=7.79 $Y=2.9 $X2=0
+ $Y2=0
cc_921 N_A_1378_125#_c_1150_n N_VPWR_c_1776_n 0.00646822f $X=8.63 $Y=2.695 $X2=0
+ $Y2=0
cc_922 N_A_1378_125#_c_1146_n N_A_1183_102#_M1001_d 0.0032498f $X=12.295
+ $Y=2.695 $X2=0 $Y2=0
cc_923 N_A_1378_125#_c_1150_n N_A_1183_102#_M1001_d 0.00454018f $X=8.63 $Y=2.695
+ $X2=0 $Y2=0
cc_924 N_A_1378_125#_c_1132_n N_A_1183_102#_c_2137_n 0.0232953f $X=6.4 $Y=1.98
+ $X2=0 $Y2=0
cc_925 N_A_1378_125#_c_1156_n N_A_1183_102#_c_2137_n 0.0134469f $X=6.485 $Y=1.13
+ $X2=0 $Y2=0
cc_926 N_A_1378_125#_M1016_g N_A_1183_102#_c_2145_n 0.007755f $X=8.97 $Y=2.34
+ $X2=0 $Y2=0
cc_927 N_A_1378_125#_c_1130_n N_A_1183_102#_c_2145_n 0.00452406f $X=8.88
+ $Y=1.485 $X2=0 $Y2=0
cc_928 N_A_1378_125#_c_1230_p N_A_1183_102#_c_2145_n 0.0108693f $X=8.71 $Y=1.485
+ $X2=0 $Y2=0
cc_929 N_A_1378_125#_c_1128_n N_A_1183_102#_c_2138_n 0.0119665f $X=9.35 $Y=1.395
+ $X2=0 $Y2=0
cc_930 N_A_1378_125#_c_1129_n N_A_1183_102#_c_2138_n 0.00824624f $X=9.425
+ $Y=1.32 $X2=0 $Y2=0
cc_931 N_A_1378_125#_c_1131_n N_A_1183_102#_c_2138_n 0.00481137f $X=8.97
+ $Y=1.485 $X2=0 $Y2=0
cc_932 N_A_1378_125#_c_1230_p N_A_1183_102#_c_2138_n 0.017395f $X=8.71 $Y=1.485
+ $X2=0 $Y2=0
cc_933 N_A_1378_125#_M1016_g N_A_1183_102#_c_2140_n 0.00282711f $X=8.97 $Y=2.34
+ $X2=0 $Y2=0
cc_934 N_A_1378_125#_c_1130_n N_A_1183_102#_c_2140_n 0.00351064f $X=8.88
+ $Y=1.485 $X2=0 $Y2=0
cc_935 N_A_1378_125#_c_1131_n N_A_1183_102#_c_2140_n 0.00601054f $X=8.97
+ $Y=1.485 $X2=0 $Y2=0
cc_936 N_A_1378_125#_c_1132_n N_A_1183_102#_c_2140_n 0.0149711f $X=6.4 $Y=1.98
+ $X2=0 $Y2=0
cc_937 N_A_1378_125#_c_1133_n N_A_1183_102#_c_2140_n 0.013647f $X=7.79 $Y=2.725
+ $X2=0 $Y2=0
cc_938 N_A_1378_125#_c_1192_n N_A_1183_102#_c_2140_n 0.00433015f $X=7.875
+ $Y=1.565 $X2=0 $Y2=0
cc_939 N_A_1378_125#_c_1134_n N_A_1183_102#_c_2140_n 0.00551874f $X=8.37
+ $Y=1.485 $X2=0 $Y2=0
cc_940 N_A_1378_125#_c_1230_p N_A_1183_102#_c_2140_n 0.0166872f $X=8.71 $Y=1.485
+ $X2=0 $Y2=0
cc_941 N_A_1378_125#_c_1157_n N_A_1183_102#_c_2140_n 0.00172569f $X=6.4 $Y=2.065
+ $X2=0 $Y2=0
cc_942 N_A_1378_125#_c_1172_n N_A_1183_102#_c_2140_n 0.00433712f $X=7.03 $Y=1.11
+ $X2=0 $Y2=0
cc_943 N_A_1378_125#_c_1203_n N_A_1183_102#_c_2140_n 0.00826032f $X=6.865
+ $Y=1.115 $X2=0 $Y2=0
cc_944 N_A_1378_125#_c_1137_n N_A_1183_102#_c_2140_n 0.0121484f $X=8.205
+ $Y=1.485 $X2=0 $Y2=0
cc_945 N_A_1378_125#_c_1132_n N_A_1183_102#_c_2141_n 6.25769e-19 $X=6.4 $Y=1.98
+ $X2=0 $Y2=0
cc_946 N_A_1378_125#_c_1128_n N_A_1183_102#_c_2142_n 7.80307e-19 $X=9.35
+ $Y=1.395 $X2=0 $Y2=0
cc_947 N_A_1378_125#_c_1230_p N_A_1183_102#_c_2142_n 2.3631e-19 $X=8.71 $Y=1.485
+ $X2=0 $Y2=0
cc_948 N_A_1378_125#_M1016_g N_A_1183_102#_c_2143_n 0.0156462f $X=8.97 $Y=2.34
+ $X2=0 $Y2=0
cc_949 N_A_1378_125#_c_1128_n N_A_1183_102#_c_2143_n 0.00906648f $X=9.35
+ $Y=1.395 $X2=0 $Y2=0
cc_950 N_A_1378_125#_c_1131_n N_A_1183_102#_c_2143_n 0.00300299f $X=8.97
+ $Y=1.485 $X2=0 $Y2=0
cc_951 N_A_1378_125#_c_1230_p N_A_1183_102#_c_2143_n 0.00703936f $X=8.71
+ $Y=1.485 $X2=0 $Y2=0
cc_952 N_A_1378_125#_c_1132_n N_A_1183_102#_c_2144_n 0.0152081f $X=6.4 $Y=1.98
+ $X2=0 $Y2=0
cc_953 N_A_1378_125#_c_1146_n N_COUT_M1008_d 0.00410409f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_954 N_A_1378_125#_c_1146_n N_COUT_M1036_d 0.00410409f $X=12.295 $Y=2.695
+ $X2=0 $Y2=0
cc_955 N_A_1268_379#_M1041_d N_A_1278_102#_c_1564_n 0.00240242f $X=7.32 $Y=0.625
+ $X2=0 $Y2=0
cc_956 N_A_1268_379#_c_1353_n N_A_1278_102#_c_1564_n 0.0591356f $X=8.705 $Y=1.02
+ $X2=0 $Y2=0
cc_957 N_A_1268_379#_c_1356_n N_A_1278_102#_c_1564_n 0.0159286f $X=8.875 $Y=0.68
+ $X2=0 $Y2=0
cc_958 N_A_1268_379#_c_1358_n N_A_1278_102#_c_1564_n 0.0197937f $X=7.525 $Y=1.02
+ $X2=0 $Y2=0
cc_959 N_A_1268_379#_M1008_g N_A_1278_102#_c_1579_n 0.0158493f $X=9.83 $Y=2.4
+ $X2=0 $Y2=0
cc_960 N_A_1268_379#_M1024_g N_A_1278_102#_c_1579_n 0.0125275f $X=10.28 $Y=2.4
+ $X2=0 $Y2=0
cc_961 N_A_1268_379#_M1036_g N_A_1278_102#_c_1579_n 0.0125126f $X=10.9 $Y=2.4
+ $X2=0 $Y2=0
cc_962 N_A_1268_379#_M1039_g N_A_1278_102#_c_1579_n 0.0150609f $X=11.35 $Y=2.4
+ $X2=0 $Y2=0
cc_963 N_A_1268_379#_c_1357_n N_A_1278_102#_c_1579_n 0.00298542f $X=9.865
+ $Y=1.35 $X2=0 $Y2=0
cc_964 N_A_1268_379#_c_1359_n N_A_1278_102#_c_1579_n 0.0120464f $X=11.405
+ $Y=1.517 $X2=0 $Y2=0
cc_965 N_A_1268_379#_c_1353_n N_A_1278_102#_c_1566_n 0.0059494f $X=8.705 $Y=1.02
+ $X2=0 $Y2=0
cc_966 N_A_1268_379#_c_1355_n N_A_1278_102#_c_1566_n 0.0487789f $X=9.385 $Y=0.68
+ $X2=0 $Y2=0
cc_967 N_A_1268_379#_c_1356_n N_A_1278_102#_c_1566_n 0.0131348f $X=8.875 $Y=0.68
+ $X2=0 $Y2=0
cc_968 N_A_1268_379#_c_1438_p N_A_1278_102#_c_1566_n 0.00512258f $X=9.78
+ $Y=1.095 $X2=0 $Y2=0
cc_969 N_A_1268_379#_c_1348_n N_A_1278_102#_c_1568_n 0.00439367f $X=10.425
+ $Y=1.35 $X2=0 $Y2=0
cc_970 N_A_1268_379#_c_1355_n N_A_1278_102#_c_1568_n 0.00289242f $X=9.385
+ $Y=0.68 $X2=0 $Y2=0
cc_971 N_A_1268_379#_c_1348_n N_A_1278_102#_c_1645_n 0.0149351f $X=10.425
+ $Y=1.35 $X2=0 $Y2=0
cc_972 N_A_1268_379#_c_1349_n N_A_1278_102#_c_1645_n 0.0122214f $X=10.855
+ $Y=1.35 $X2=0 $Y2=0
cc_973 N_A_1268_379#_c_1350_n N_A_1278_102#_c_1645_n 0.0122187f $X=11.405
+ $Y=1.35 $X2=0 $Y2=0
cc_974 N_A_1268_379#_c_1351_n N_A_1278_102#_c_1645_n 0.0174474f $X=11.835
+ $Y=1.35 $X2=0 $Y2=0
cc_975 N_A_1268_379#_c_1438_p N_A_1278_102#_c_1645_n 0.00443282f $X=9.78
+ $Y=1.095 $X2=0 $Y2=0
cc_976 N_A_1268_379#_c_1446_p N_A_1278_102#_c_1645_n 0.0152617f $X=10.585
+ $Y=1.515 $X2=0 $Y2=0
cc_977 N_A_1268_379#_c_1359_n N_A_1278_102#_c_1645_n 0.00853237f $X=11.405
+ $Y=1.517 $X2=0 $Y2=0
cc_978 N_A_1268_379#_c_1438_p N_A_1278_102#_c_1615_n 0.0145386f $X=9.78 $Y=1.095
+ $X2=0 $Y2=0
cc_979 N_A_1268_379#_c_1359_n N_A_1278_102#_c_1615_n 4.2528e-19 $X=11.405
+ $Y=1.517 $X2=0 $Y2=0
cc_980 N_A_1268_379#_M1039_g N_A_1278_102#_c_1569_n 0.0106204f $X=11.35 $Y=2.4
+ $X2=0 $Y2=0
cc_981 N_A_1268_379#_c_1351_n N_A_1278_102#_c_1569_n 0.0225461f $X=11.835
+ $Y=1.35 $X2=0 $Y2=0
cc_982 N_A_1268_379#_M1024_g N_VPWR_c_1783_n 0.00382756f $X=10.28 $Y=2.4 $X2=0
+ $Y2=0
cc_983 N_A_1268_379#_M1036_g N_VPWR_c_1783_n 0.00382756f $X=10.9 $Y=2.4 $X2=0
+ $Y2=0
cc_984 N_A_1268_379#_M1008_g N_VPWR_c_1784_n 0.00380045f $X=9.83 $Y=2.4 $X2=0
+ $Y2=0
cc_985 N_A_1268_379#_M1024_g N_VPWR_c_1784_n 0.00380045f $X=10.28 $Y=2.4 $X2=0
+ $Y2=0
cc_986 N_A_1268_379#_M1008_g N_VPWR_c_1796_n 0.00587695f $X=9.83 $Y=2.4 $X2=0
+ $Y2=0
cc_987 N_A_1268_379#_M1036_g N_VPWR_c_1797_n 0.00380045f $X=10.9 $Y=2.4 $X2=0
+ $Y2=0
cc_988 N_A_1268_379#_M1039_g N_VPWR_c_1797_n 0.00380045f $X=11.35 $Y=2.4 $X2=0
+ $Y2=0
cc_989 N_A_1268_379#_M1039_g N_VPWR_c_1798_n 0.00616041f $X=11.35 $Y=2.4 $X2=0
+ $Y2=0
cc_990 N_A_1268_379#_M1008_g N_VPWR_c_1776_n 0.00475386f $X=9.83 $Y=2.4 $X2=0
+ $Y2=0
cc_991 N_A_1268_379#_M1024_g N_VPWR_c_1776_n 0.00471761f $X=10.28 $Y=2.4 $X2=0
+ $Y2=0
cc_992 N_A_1268_379#_M1036_g N_VPWR_c_1776_n 0.00471761f $X=10.9 $Y=2.4 $X2=0
+ $Y2=0
cc_993 N_A_1268_379#_M1039_g N_VPWR_c_1776_n 0.00475386f $X=11.35 $Y=2.4 $X2=0
+ $Y2=0
cc_994 N_A_1268_379#_c_1355_n N_A_1183_102#_M1020_s 0.00555428f $X=9.385 $Y=0.68
+ $X2=0 $Y2=0
cc_995 N_A_1268_379#_c_1353_n N_A_1183_102#_c_2138_n 0.0141318f $X=8.705 $Y=1.02
+ $X2=0 $Y2=0
cc_996 N_A_1268_379#_c_1355_n N_A_1183_102#_c_2138_n 0.0136682f $X=9.385 $Y=0.68
+ $X2=0 $Y2=0
cc_997 N_A_1268_379#_c_1418_n N_A_1183_102#_c_2138_n 0.00523147f $X=9.47 $Y=1.01
+ $X2=0 $Y2=0
cc_998 N_A_1268_379#_c_1419_n N_A_1183_102#_c_2138_n 0.0131627f $X=9.555
+ $Y=1.095 $X2=0 $Y2=0
cc_999 N_A_1268_379#_c_1357_n N_A_1183_102#_c_2138_n 0.0111278f $X=9.865 $Y=1.35
+ $X2=0 $Y2=0
cc_1000 N_A_1268_379#_c_1359_n N_A_1183_102#_c_2138_n 0.00103954f $X=11.405
+ $Y=1.517 $X2=0 $Y2=0
cc_1001 N_A_1268_379#_c_1368_n N_A_1183_102#_c_2140_n 0.00736532f $X=7.365
+ $Y=2.405 $X2=0 $Y2=0
cc_1002 N_A_1268_379#_c_1352_n N_A_1183_102#_c_2140_n 0.0206767f $X=7.45 $Y=2.32
+ $X2=0 $Y2=0
cc_1003 N_A_1268_379#_c_1353_n N_A_1183_102#_c_2140_n 0.00634108f $X=8.705
+ $Y=1.02 $X2=0 $Y2=0
cc_1004 N_A_1268_379#_c_1358_n N_A_1183_102#_c_2140_n 0.00613882f $X=7.525
+ $Y=1.02 $X2=0 $Y2=0
cc_1005 N_A_1268_379#_c_1419_n N_A_1183_102#_c_2142_n 0.00187797f $X=9.555
+ $Y=1.095 $X2=0 $Y2=0
cc_1006 N_A_1268_379#_c_1357_n N_A_1183_102#_c_2142_n 0.00396076f $X=9.865
+ $Y=1.35 $X2=0 $Y2=0
cc_1007 N_A_1268_379#_c_1359_n N_A_1183_102#_c_2142_n 0.00476444f $X=11.405
+ $Y=1.517 $X2=0 $Y2=0
cc_1008 N_A_1268_379#_M1008_g N_A_1183_102#_c_2143_n 0.00344561f $X=9.83 $Y=2.4
+ $X2=0 $Y2=0
cc_1009 N_A_1268_379#_c_1419_n N_A_1183_102#_c_2143_n 0.00274373f $X=9.555
+ $Y=1.095 $X2=0 $Y2=0
cc_1010 N_A_1268_379#_c_1357_n N_A_1183_102#_c_2143_n 0.00493762f $X=9.865
+ $Y=1.35 $X2=0 $Y2=0
cc_1011 N_A_1268_379#_c_1359_n N_A_1183_102#_c_2143_n 0.00324543f $X=11.405
+ $Y=1.517 $X2=0 $Y2=0
cc_1012 N_A_1268_379#_M1008_g N_COUT_c_2249_n 0.00663761f $X=9.83 $Y=2.4 $X2=0
+ $Y2=0
cc_1013 N_A_1268_379#_M1024_g N_COUT_c_2249_n 0.0133089f $X=10.28 $Y=2.4 $X2=0
+ $Y2=0
cc_1014 N_A_1268_379#_M1036_g N_COUT_c_2249_n 0.013935f $X=10.9 $Y=2.4 $X2=0
+ $Y2=0
cc_1015 N_A_1268_379#_c_1357_n N_COUT_c_2249_n 0.00356953f $X=9.865 $Y=1.35
+ $X2=0 $Y2=0
cc_1016 N_A_1268_379#_c_1446_p N_COUT_c_2249_n 0.0518067f $X=10.585 $Y=1.515
+ $X2=0 $Y2=0
cc_1017 N_A_1268_379#_c_1359_n N_COUT_c_2249_n 0.00860274f $X=11.405 $Y=1.517
+ $X2=0 $Y2=0
cc_1018 N_A_1268_379#_c_1348_n N_COUT_c_2255_n 0.0039161f $X=10.425 $Y=1.35
+ $X2=0 $Y2=0
cc_1019 N_A_1268_379#_c_1349_n N_COUT_c_2255_n 0.0112714f $X=10.855 $Y=1.35
+ $X2=0 $Y2=0
cc_1020 N_A_1268_379#_c_1438_p N_COUT_c_2255_n 0.00597892f $X=9.78 $Y=1.095
+ $X2=0 $Y2=0
cc_1021 N_A_1268_379#_c_1446_p N_COUT_c_2255_n 0.0151874f $X=10.585 $Y=1.515
+ $X2=0 $Y2=0
cc_1022 N_A_1268_379#_c_1359_n N_COUT_c_2255_n 0.00224206f $X=11.405 $Y=1.517
+ $X2=0 $Y2=0
cc_1023 N_A_1268_379#_c_1350_n N_COUT_c_2244_n 0.0070657f $X=11.405 $Y=1.35
+ $X2=0 $Y2=0
cc_1024 N_A_1268_379#_c_1351_n N_COUT_c_2244_n 0.00427856f $X=11.835 $Y=1.35
+ $X2=0 $Y2=0
cc_1025 N_A_1268_379#_c_1359_n N_COUT_c_2244_n 0.00428146f $X=11.405 $Y=1.517
+ $X2=0 $Y2=0
cc_1026 N_A_1268_379#_c_1349_n N_COUT_c_2245_n 0.00101776f $X=10.855 $Y=1.35
+ $X2=0 $Y2=0
cc_1027 N_A_1268_379#_c_1350_n N_COUT_c_2245_n 0.00625608f $X=11.405 $Y=1.35
+ $X2=0 $Y2=0
cc_1028 N_A_1268_379#_M1036_g N_COUT_c_2265_n 0.00108858f $X=10.9 $Y=2.4 $X2=0
+ $Y2=0
cc_1029 N_A_1268_379#_M1039_g N_COUT_c_2265_n 0.00903001f $X=11.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1030 N_A_1268_379#_M1024_g COUT 7.45537e-19 $X=10.28 $Y=2.4 $X2=0 $Y2=0
cc_1031 N_A_1268_379#_c_1349_n COUT 0.00276711f $X=10.855 $Y=1.35 $X2=0 $Y2=0
cc_1032 N_A_1268_379#_M1036_g COUT 0.00558626f $X=10.9 $Y=2.4 $X2=0 $Y2=0
cc_1033 N_A_1268_379#_M1039_g COUT 0.00640851f $X=11.35 $Y=2.4 $X2=0 $Y2=0
cc_1034 N_A_1268_379#_c_1350_n COUT 0.00304543f $X=11.405 $Y=1.35 $X2=0 $Y2=0
cc_1035 N_A_1268_379#_c_1351_n COUT 2.86206e-19 $X=11.835 $Y=1.35 $X2=0 $Y2=0
cc_1036 N_A_1268_379#_c_1446_p COUT 0.0196019f $X=10.585 $Y=1.515 $X2=0 $Y2=0
cc_1037 N_A_1268_379#_c_1359_n COUT 0.0338604f $X=11.405 $Y=1.517 $X2=0 $Y2=0
cc_1038 N_A_1268_379#_c_1438_p N_VGND_M1020_d 0.0181521f $X=9.78 $Y=1.095 $X2=0
+ $Y2=0
cc_1039 N_A_1268_379#_c_1357_n N_VGND_M1020_d 0.00168778f $X=9.865 $Y=1.35 $X2=0
+ $Y2=0
cc_1040 N_A_1268_379#_c_1348_n N_VGND_c_2356_n 0.0038192f $X=10.425 $Y=1.35
+ $X2=0 $Y2=0
cc_1041 N_A_1268_379#_c_1349_n N_VGND_c_2357_n 0.00213129f $X=10.855 $Y=1.35
+ $X2=0 $Y2=0
cc_1042 N_A_1268_379#_c_1350_n N_VGND_c_2357_n 0.00216156f $X=11.405 $Y=1.35
+ $X2=0 $Y2=0
cc_1043 N_A_1268_379#_c_1351_n N_VGND_c_2358_n 0.00382573f $X=11.835 $Y=1.35
+ $X2=0 $Y2=0
cc_1044 N_A_1268_379#_c_1348_n N_VGND_c_2369_n 0.00377304f $X=10.425 $Y=1.35
+ $X2=0 $Y2=0
cc_1045 N_A_1268_379#_c_1349_n N_VGND_c_2369_n 0.00377304f $X=10.855 $Y=1.35
+ $X2=0 $Y2=0
cc_1046 N_A_1268_379#_c_1350_n N_VGND_c_2371_n 0.00377304f $X=11.405 $Y=1.35
+ $X2=0 $Y2=0
cc_1047 N_A_1268_379#_c_1351_n N_VGND_c_2371_n 0.00377304f $X=11.835 $Y=1.35
+ $X2=0 $Y2=0
cc_1048 N_A_1268_379#_c_1348_n N_VGND_c_2380_n 0.00505379f $X=10.425 $Y=1.35
+ $X2=0 $Y2=0
cc_1049 N_A_1268_379#_c_1349_n N_VGND_c_2380_n 0.00505379f $X=10.855 $Y=1.35
+ $X2=0 $Y2=0
cc_1050 N_A_1268_379#_c_1350_n N_VGND_c_2380_n 0.00505379f $X=11.405 $Y=1.35
+ $X2=0 $Y2=0
cc_1051 N_A_1268_379#_c_1351_n N_VGND_c_2380_n 0.00505379f $X=11.835 $Y=1.35
+ $X2=0 $Y2=0
cc_1052 N_CI_M1034_g N_A_1278_102#_M1012_g 0.0169807f $X=12.775 $Y=2.34 $X2=0
+ $Y2=0
cc_1053 N_CI_c_1523_n N_A_1278_102#_M1012_g 0.0021753f $X=12.815 $Y=1.515 $X2=0
+ $Y2=0
cc_1054 N_CI_c_1524_n N_A_1278_102#_c_1560_n 0.017705f $X=12.815 $Y=1.35 $X2=0
+ $Y2=0
cc_1055 N_CI_c_1523_n N_A_1278_102#_c_1570_n 0.00369733f $X=12.815 $Y=1.515
+ $X2=0 $Y2=0
cc_1056 N_CI_c_1524_n N_A_1278_102#_c_1570_n 0.0153141f $X=12.815 $Y=1.35 $X2=0
+ $Y2=0
cc_1057 N_CI_c_1524_n N_A_1278_102#_c_1571_n 0.00840455f $X=12.815 $Y=1.35 $X2=0
+ $Y2=0
cc_1058 N_CI_c_1522_n N_A_1278_102#_c_1572_n 0.00239698f $X=12.815 $Y=1.515
+ $X2=0 $Y2=0
cc_1059 N_CI_c_1523_n N_A_1278_102#_c_1572_n 0.0219159f $X=12.815 $Y=1.515 $X2=0
+ $Y2=0
cc_1060 N_CI_c_1522_n N_A_1278_102#_c_1574_n 0.0138012f $X=12.815 $Y=1.515 $X2=0
+ $Y2=0
cc_1061 N_CI_c_1523_n N_A_1278_102#_c_1574_n 3.82865e-19 $X=12.815 $Y=1.515
+ $X2=0 $Y2=0
cc_1062 N_CI_M1034_g N_VPWR_c_1779_n 0.00873271f $X=12.775 $Y=2.34 $X2=0 $Y2=0
cc_1063 N_CI_c_1522_n N_VPWR_c_1779_n 3.50127e-19 $X=12.815 $Y=1.515 $X2=0 $Y2=0
cc_1064 N_CI_c_1523_n N_VPWR_c_1779_n 0.00510587f $X=12.815 $Y=1.515 $X2=0 $Y2=0
cc_1065 N_CI_M1034_g N_VPWR_c_1785_n 0.00567028f $X=12.775 $Y=2.34 $X2=0 $Y2=0
cc_1066 N_CI_M1034_g N_VPWR_c_1798_n 5.20033e-19 $X=12.775 $Y=2.34 $X2=0 $Y2=0
cc_1067 N_CI_M1034_g N_VPWR_c_1776_n 0.00610055f $X=12.775 $Y=2.34 $X2=0 $Y2=0
cc_1068 N_CI_M1034_g N_SUM_c_2296_n 4.61105e-19 $X=12.775 $Y=2.34 $X2=0 $Y2=0
cc_1069 N_CI_c_1524_n N_SUM_c_2290_n 9.14912e-19 $X=12.815 $Y=1.35 $X2=0 $Y2=0
cc_1070 N_CI_c_1524_n N_VGND_c_2358_n 7.59991e-19 $X=12.815 $Y=1.35 $X2=0 $Y2=0
cc_1071 N_CI_c_1524_n N_VGND_c_2359_n 8.80616e-19 $X=12.815 $Y=1.35 $X2=0 $Y2=0
cc_1072 N_CI_c_1524_n N_VGND_c_2374_n 0.00333058f $X=12.815 $Y=1.35 $X2=0 $Y2=0
cc_1073 N_CI_c_1524_n N_VGND_c_2380_n 0.00476395f $X=12.815 $Y=1.35 $X2=0 $Y2=0
cc_1074 N_A_1278_102#_c_1579_n N_VPWR_M1016_d 0.0217932f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1075 N_A_1278_102#_c_1579_n N_VPWR_M1024_s 0.00744798f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1076 N_A_1278_102#_c_1579_n N_VPWR_M1039_s 0.0195586f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1077 N_A_1278_102#_c_1569_n N_VPWR_M1039_s 0.0103656f $X=12.04 $Y=2.27 $X2=0
+ $Y2=0
cc_1078 N_A_1278_102#_M1012_g N_VPWR_c_1779_n 0.00383792f $X=13.36 $Y=2.4 $X2=0
+ $Y2=0
cc_1079 N_A_1278_102#_M1013_g N_VPWR_c_1780_n 0.00243252f $X=13.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1080 N_A_1278_102#_M1015_g N_VPWR_c_1780_n 0.00388538f $X=14.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1081 N_A_1278_102#_M1032_g N_VPWR_c_1782_n 0.00649214f $X=14.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1082 N_A_1278_102#_M1012_g N_VPWR_c_1790_n 0.005209f $X=13.36 $Y=2.4 $X2=0
+ $Y2=0
cc_1083 N_A_1278_102#_M1013_g N_VPWR_c_1790_n 0.005209f $X=13.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1084 N_A_1278_102#_M1015_g N_VPWR_c_1791_n 0.0053223f $X=14.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1085 N_A_1278_102#_M1032_g N_VPWR_c_1791_n 0.00515235f $X=14.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1086 N_A_1278_102#_M1012_g N_VPWR_c_1776_n 0.00986727f $X=13.36 $Y=2.4 $X2=0
+ $Y2=0
cc_1087 N_A_1278_102#_M1013_g N_VPWR_c_1776_n 0.0098244f $X=13.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1088 N_A_1278_102#_M1015_g N_VPWR_c_1776_n 0.01019f $X=14.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1089 N_A_1278_102#_M1032_g N_VPWR_c_1776_n 0.00967912f $X=14.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1090 N_A_1278_102#_c_1579_n N_A_1183_102#_M1001_d 0.00486963f $X=11.955
+ $Y=2.355 $X2=0 $Y2=0
cc_1091 N_A_1278_102#_c_1579_n N_A_1183_102#_c_2145_n 0.0281851f $X=11.955
+ $Y=2.355 $X2=0 $Y2=0
cc_1092 N_A_1278_102#_c_1579_n N_A_1183_102#_c_2140_n 0.00537584f $X=11.955
+ $Y=2.355 $X2=0 $Y2=0
cc_1093 N_A_1278_102#_c_1582_n N_A_1183_102#_c_2140_n 0.00814434f $X=8.21
+ $Y=2.26 $X2=0 $Y2=0
cc_1094 N_A_1278_102#_c_1579_n N_A_1183_102#_c_2142_n 0.00688913f $X=11.955
+ $Y=2.355 $X2=0 $Y2=0
cc_1095 N_A_1278_102#_c_1579_n N_A_1183_102#_c_2143_n 0.0143996f $X=11.955
+ $Y=2.355 $X2=0 $Y2=0
cc_1096 N_A_1278_102#_c_1645_n N_COUT_M1009_d 0.00465974f $X=11.955 $Y=0.755
+ $X2=-0.19 $Y2=-0.245
cc_1097 N_A_1278_102#_c_1645_n N_COUT_M1014_d 0.00465974f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1098 N_A_1278_102#_c_1579_n N_COUT_M1008_d 0.00324035f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1099 N_A_1278_102#_c_1579_n N_COUT_M1036_d 0.00323662f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1100 N_A_1278_102#_c_1579_n N_COUT_c_2249_n 0.0610881f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1101 N_A_1278_102#_c_1645_n N_COUT_c_2255_n 0.0238509f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1102 N_A_1278_102#_c_1645_n N_COUT_c_2244_n 0.0199912f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1103 N_A_1278_102#_c_1569_n N_COUT_c_2244_n 0.0111269f $X=12.04 $Y=2.27 $X2=0
+ $Y2=0
cc_1104 N_A_1278_102#_c_1645_n N_COUT_c_2245_n 0.0282199f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1105 N_A_1278_102#_c_1579_n N_COUT_c_2265_n 0.0250924f $X=11.955 $Y=2.355
+ $X2=0 $Y2=0
cc_1106 N_A_1278_102#_c_1569_n N_COUT_c_2265_n 0.00768039f $X=12.04 $Y=2.27
+ $X2=0 $Y2=0
cc_1107 N_A_1278_102#_c_1569_n COUT 0.0182058f $X=12.04 $Y=2.27 $X2=0 $Y2=0
cc_1108 N_A_1278_102#_M1012_g N_SUM_c_2296_n 0.00350401f $X=13.36 $Y=2.4 $X2=0
+ $Y2=0
cc_1109 N_A_1278_102#_M1013_g N_SUM_c_2296_n 8.84614e-19 $X=13.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1110 N_A_1278_102#_c_1702_p N_SUM_c_2296_n 0.0218858f $X=14.16 $Y=1.515 $X2=0
+ $Y2=0
cc_1111 N_A_1278_102#_c_1574_n N_SUM_c_2296_n 0.00245159f $X=14.795 $Y=1.515
+ $X2=0 $Y2=0
cc_1112 N_A_1278_102#_M1012_g N_SUM_c_2293_n 0.0116697f $X=13.36 $Y=2.4 $X2=0
+ $Y2=0
cc_1113 N_A_1278_102#_M1013_g N_SUM_c_2293_n 0.0132668f $X=13.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1114 N_A_1278_102#_M1015_g N_SUM_c_2293_n 6.25485e-19 $X=14.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1115 N_A_1278_102#_c_1560_n N_SUM_c_2290_n 0.00762192f $X=13.505 $Y=1.35
+ $X2=0 $Y2=0
cc_1116 N_A_1278_102#_M1013_g N_SUM_c_2306_n 0.0134371f $X=13.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1117 N_A_1278_102#_M1015_g N_SUM_c_2306_n 0.0155601f $X=14.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1118 N_A_1278_102#_c_1702_p N_SUM_c_2306_n 0.0377615f $X=14.16 $Y=1.515 $X2=0
+ $Y2=0
cc_1119 N_A_1278_102#_c_1574_n N_SUM_c_2306_n 0.00446909f $X=14.795 $Y=1.515
+ $X2=0 $Y2=0
cc_1120 N_A_1278_102#_c_1561_n N_SUM_c_2310_n 0.0120151f $X=13.935 $Y=1.35 $X2=0
+ $Y2=0
cc_1121 N_A_1278_102#_c_1562_n N_SUM_c_2310_n 0.01375f $X=14.365 $Y=1.35 $X2=0
+ $Y2=0
cc_1122 N_A_1278_102#_c_1702_p N_SUM_c_2310_n 0.0317758f $X=14.16 $Y=1.515 $X2=0
+ $Y2=0
cc_1123 N_A_1278_102#_c_1574_n N_SUM_c_2310_n 0.00236025f $X=14.795 $Y=1.515
+ $X2=0 $Y2=0
cc_1124 N_A_1278_102#_c_1560_n N_SUM_c_2314_n 0.00210071f $X=13.505 $Y=1.35
+ $X2=0 $Y2=0
cc_1125 N_A_1278_102#_c_1702_p N_SUM_c_2314_n 0.0179227f $X=14.16 $Y=1.515 $X2=0
+ $Y2=0
cc_1126 N_A_1278_102#_c_1574_n N_SUM_c_2314_n 0.00272203f $X=14.795 $Y=1.515
+ $X2=0 $Y2=0
cc_1127 N_A_1278_102#_c_1562_n N_SUM_c_2291_n 3.97481e-19 $X=14.365 $Y=1.35
+ $X2=0 $Y2=0
cc_1128 N_A_1278_102#_c_1563_n N_SUM_c_2291_n 0.00666962f $X=14.795 $Y=1.35
+ $X2=0 $Y2=0
cc_1129 N_A_1278_102#_M1015_g N_SUM_c_2292_n 0.00411339f $X=14.35 $Y=2.4 $X2=0
+ $Y2=0
cc_1130 N_A_1278_102#_c_1562_n N_SUM_c_2292_n 0.00280039f $X=14.365 $Y=1.35
+ $X2=0 $Y2=0
cc_1131 N_A_1278_102#_c_1563_n N_SUM_c_2292_n 0.00556993f $X=14.795 $Y=1.35
+ $X2=0 $Y2=0
cc_1132 N_A_1278_102#_M1032_g N_SUM_c_2292_n 0.00769591f $X=14.81 $Y=2.4 $X2=0
+ $Y2=0
cc_1133 N_A_1278_102#_c_1702_p N_SUM_c_2292_n 0.0256674f $X=14.16 $Y=1.515 $X2=0
+ $Y2=0
cc_1134 N_A_1278_102#_c_1574_n N_SUM_c_2292_n 0.0304506f $X=14.795 $Y=1.515
+ $X2=0 $Y2=0
cc_1135 N_A_1278_102#_c_1563_n N_SUM_c_2325_n 0.00181823f $X=14.795 $Y=1.35
+ $X2=0 $Y2=0
cc_1136 N_A_1278_102#_M1015_g SUM 8.43868e-19 $X=14.35 $Y=2.4 $X2=0 $Y2=0
cc_1137 N_A_1278_102#_M1032_g SUM 0.00269271f $X=14.81 $Y=2.4 $X2=0 $Y2=0
cc_1138 N_A_1278_102#_M1013_g SUM 6.12982e-19 $X=13.81 $Y=2.4 $X2=0 $Y2=0
cc_1139 N_A_1278_102#_M1015_g SUM 0.0125129f $X=14.35 $Y=2.4 $X2=0 $Y2=0
cc_1140 N_A_1278_102#_M1032_g SUM 0.0130241f $X=14.81 $Y=2.4 $X2=0 $Y2=0
cc_1141 N_A_1278_102#_c_1568_n N_VGND_M1020_d 0.00225064f $X=9.81 $Y=0.67 $X2=0
+ $Y2=0
cc_1142 N_A_1278_102#_c_1645_n N_VGND_M1020_d 0.0137386f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1143 N_A_1278_102#_c_1615_n N_VGND_M1020_d 0.00476653f $X=9.895 $Y=0.755
+ $X2=0 $Y2=0
cc_1144 N_A_1278_102#_c_1645_n N_VGND_M1011_s 0.00609924f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1145 N_A_1278_102#_c_1569_n N_VGND_M1022_s 0.0111503f $X=12.04 $Y=2.27 $X2=0
+ $Y2=0
cc_1146 N_A_1278_102#_c_1570_n N_VGND_M1022_s 0.00860261f $X=13.215 $Y=0.755
+ $X2=0 $Y2=0
cc_1147 N_A_1278_102#_c_1739_p N_VGND_M1022_s 0.00202028f $X=12.04 $Y=0.755
+ $X2=0 $Y2=0
cc_1148 N_A_1278_102#_c_1570_n N_VGND_M1017_d 0.0122531f $X=13.215 $Y=0.755
+ $X2=0 $Y2=0
cc_1149 N_A_1278_102#_c_1571_n N_VGND_M1017_d 0.00763515f $X=13.3 $Y=1.35 $X2=0
+ $Y2=0
cc_1150 N_A_1278_102#_c_1566_n N_VGND_c_2356_n 0.0145006f $X=9.725 $Y=0.34 $X2=0
+ $Y2=0
cc_1151 N_A_1278_102#_c_1568_n N_VGND_c_2356_n 0.00567177f $X=9.81 $Y=0.67 $X2=0
+ $Y2=0
cc_1152 N_A_1278_102#_c_1645_n N_VGND_c_2356_n 0.0184124f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1153 N_A_1278_102#_c_1645_n N_VGND_c_2357_n 0.0238802f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1154 N_A_1278_102#_c_1570_n N_VGND_c_2358_n 0.0130442f $X=13.215 $Y=0.755
+ $X2=0 $Y2=0
cc_1155 N_A_1278_102#_c_1739_p N_VGND_c_2358_n 0.0134917f $X=12.04 $Y=0.755
+ $X2=0 $Y2=0
cc_1156 N_A_1278_102#_c_1560_n N_VGND_c_2359_n 0.00323466f $X=13.505 $Y=1.35
+ $X2=0 $Y2=0
cc_1157 N_A_1278_102#_c_1570_n N_VGND_c_2359_n 0.0272503f $X=13.215 $Y=0.755
+ $X2=0 $Y2=0
cc_1158 N_A_1278_102#_c_1560_n N_VGND_c_2360_n 4.50936e-19 $X=13.505 $Y=1.35
+ $X2=0 $Y2=0
cc_1159 N_A_1278_102#_c_1561_n N_VGND_c_2360_n 0.00826597f $X=13.935 $Y=1.35
+ $X2=0 $Y2=0
cc_1160 N_A_1278_102#_c_1562_n N_VGND_c_2360_n 0.00824964f $X=14.365 $Y=1.35
+ $X2=0 $Y2=0
cc_1161 N_A_1278_102#_c_1563_n N_VGND_c_2360_n 4.4964e-19 $X=14.795 $Y=1.35
+ $X2=0 $Y2=0
cc_1162 N_A_1278_102#_c_1563_n N_VGND_c_2362_n 0.018424f $X=14.795 $Y=1.35 $X2=0
+ $Y2=0
cc_1163 N_A_1278_102#_c_1564_n N_VGND_c_2367_n 0.0033734f $X=8.365 $Y=0.68 $X2=0
+ $Y2=0
cc_1164 N_A_1278_102#_c_1566_n N_VGND_c_2367_n 0.0886485f $X=9.725 $Y=0.34 $X2=0
+ $Y2=0
cc_1165 N_A_1278_102#_c_1567_n N_VGND_c_2367_n 0.0119262f $X=8.535 $Y=0.34 $X2=0
+ $Y2=0
cc_1166 N_A_1278_102#_c_1645_n N_VGND_c_2367_n 0.00273597f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1167 N_A_1278_102#_c_1645_n N_VGND_c_2369_n 0.00883547f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1168 N_A_1278_102#_c_1645_n N_VGND_c_2371_n 0.00893371f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1169 N_A_1278_102#_c_1570_n N_VGND_c_2374_n 0.011173f $X=13.215 $Y=0.755
+ $X2=0 $Y2=0
cc_1170 N_A_1278_102#_c_1560_n N_VGND_c_2375_n 0.00467453f $X=13.505 $Y=1.35
+ $X2=0 $Y2=0
cc_1171 N_A_1278_102#_c_1561_n N_VGND_c_2375_n 0.00405273f $X=13.935 $Y=1.35
+ $X2=0 $Y2=0
cc_1172 N_A_1278_102#_c_1562_n N_VGND_c_2376_n 0.00405273f $X=14.365 $Y=1.35
+ $X2=0 $Y2=0
cc_1173 N_A_1278_102#_c_1563_n N_VGND_c_2376_n 0.00467453f $X=14.795 $Y=1.35
+ $X2=0 $Y2=0
cc_1174 N_A_1278_102#_c_1560_n N_VGND_c_2380_n 0.00505379f $X=13.505 $Y=1.35
+ $X2=0 $Y2=0
cc_1175 N_A_1278_102#_c_1561_n N_VGND_c_2380_n 0.00424518f $X=13.935 $Y=1.35
+ $X2=0 $Y2=0
cc_1176 N_A_1278_102#_c_1562_n N_VGND_c_2380_n 0.00424518f $X=14.365 $Y=1.35
+ $X2=0 $Y2=0
cc_1177 N_A_1278_102#_c_1563_n N_VGND_c_2380_n 0.00505379f $X=14.795 $Y=1.35
+ $X2=0 $Y2=0
cc_1178 N_A_1278_102#_c_1566_n N_VGND_c_2380_n 0.0513167f $X=9.725 $Y=0.34 $X2=0
+ $Y2=0
cc_1179 N_A_1278_102#_c_1567_n N_VGND_c_2380_n 0.00656035f $X=8.535 $Y=0.34
+ $X2=0 $Y2=0
cc_1180 N_A_1278_102#_c_1645_n N_VGND_c_2380_n 0.0430717f $X=11.955 $Y=0.755
+ $X2=0 $Y2=0
cc_1181 N_A_1278_102#_c_1570_n N_VGND_c_2380_n 0.0230552f $X=13.215 $Y=0.755
+ $X2=0 $Y2=0
cc_1182 N_A_1278_102#_c_1573_n N_VGND_c_2380_n 0.00870196f $X=6.705 $Y=0.72
+ $X2=0 $Y2=0
cc_1183 N_A_1278_102#_c_1739_p N_VGND_c_2380_n 0.00110116f $X=12.04 $Y=0.755
+ $X2=0 $Y2=0
cc_1184 N_VPWR_c_1777_n N_A_200_74#_c_1951_n 0.0129208f $X=0.73 $Y=2.135 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1788_n N_A_200_74#_c_1951_n 0.0146352f $X=1.575 $Y=3.33 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1793_n N_A_200_74#_c_1951_n 6.78065e-19 $X=1.745 $Y=3.055 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1776_n N_A_200_74#_c_1951_n 0.0120433f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1188 N_VPWR_M1003_s N_A_200_74#_c_1953_n 0.0133162f $X=1.595 $Y=1.81 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1788_n N_A_200_74#_c_1953_n 0.00532338f $X=1.575 $Y=3.33 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1793_n N_A_200_74#_c_1953_n 0.0190466f $X=1.745 $Y=3.055 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1776_n N_A_200_74#_c_1953_n 0.00859395f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1192 N_VPWR_M1003_s N_A_200_74#_c_1946_n 0.0169372f $X=1.595 $Y=1.81 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1789_n N_A_200_74#_c_1955_n 0.0254748f $X=5.325 $Y=3.33 $X2=0
+ $Y2=0
cc_1194 N_VPWR_c_1776_n N_A_200_74#_c_1955_n 0.032839f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1195 N_VPWR_M1003_s N_A_200_74#_c_1981_n 7.99406e-19 $X=1.595 $Y=1.81 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1789_n N_A_200_74#_c_1981_n 0.00151778f $X=5.325 $Y=3.33 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1793_n N_A_200_74#_c_1981_n 0.00635899f $X=1.745 $Y=3.055 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1776_n N_A_200_74#_c_1981_n 0.00344617f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1789_n N_A_200_74#_c_1956_n 0.0128589f $X=5.325 $Y=3.33 $X2=0
+ $Y2=0
cc_1200 N_VPWR_c_1776_n N_A_200_74#_c_1956_n 0.0103646f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1201 N_VPWR_c_1789_n N_A_430_362#_c_2058_n 0.00524178f $X=5.325 $Y=3.33 $X2=0
+ $Y2=0
cc_1202 N_VPWR_c_1776_n N_A_430_362#_c_2058_n 0.00706341f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1203 N_VPWR_M1016_d N_A_1183_102#_c_2143_n 0.00575862f $X=9.06 $Y=1.84 $X2=0
+ $Y2=0
cc_1204 N_VPWR_M1024_s N_COUT_c_2249_n 0.00785282f $X=10.37 $Y=1.84 $X2=0 $Y2=0
cc_1205 N_VPWR_c_1779_n N_SUM_c_2293_n 0.0367744f $X=13.085 $Y=2.035 $X2=0 $Y2=0
cc_1206 N_VPWR_c_1780_n N_SUM_c_2293_n 0.0304332f $X=14.085 $Y=2.355 $X2=0 $Y2=0
cc_1207 N_VPWR_c_1790_n N_SUM_c_2293_n 0.0144623f $X=13.92 $Y=3.33 $X2=0 $Y2=0
cc_1208 N_VPWR_c_1776_n N_SUM_c_2293_n 0.0118344f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1209 N_VPWR_M1013_s N_SUM_c_2306_n 0.00482477f $X=13.9 $Y=1.84 $X2=0 $Y2=0
cc_1210 N_VPWR_c_1780_n N_SUM_c_2306_n 0.0200142f $X=14.085 $Y=2.355 $X2=0 $Y2=0
cc_1211 N_VPWR_c_1782_n N_SUM_c_2292_n 0.0015622f $X=15.035 $Y=1.985 $X2=0 $Y2=0
cc_1212 N_VPWR_c_1780_n SUM 0.0305015f $X=14.085 $Y=2.355 $X2=0 $Y2=0
cc_1213 N_VPWR_c_1782_n SUM 0.0330024f $X=15.035 $Y=1.985 $X2=0 $Y2=0
cc_1214 N_VPWR_c_1791_n SUM 0.0147003f $X=14.95 $Y=3.33 $X2=0 $Y2=0
cc_1215 N_VPWR_c_1776_n SUM 0.0120432f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1216 N_VPWR_c_1782_n N_VGND_c_2362_n 0.0101049f $X=15.035 $Y=1.985 $X2=0
+ $Y2=0
cc_1217 N_A_200_74#_c_1955_n N_A_430_362#_M1003_d 0.0051819f $X=3.165 $Y=2.715
+ $X2=0 $Y2=0
cc_1218 N_A_200_74#_c_1946_n N_A_430_362#_c_2056_n 0.0177356f $X=1.92 $Y=2.63
+ $X2=0 $Y2=0
cc_1219 N_A_200_74#_c_1946_n N_A_430_362#_c_2053_n 0.0325438f $X=1.92 $Y=2.63
+ $X2=0 $Y2=0
cc_1220 N_A_200_74#_c_1947_n N_A_430_362#_c_2053_n 0.0115498f $X=2.05 $Y=0.79
+ $X2=0 $Y2=0
cc_1221 N_A_200_74#_c_1948_n N_A_430_362#_c_2053_n 0.0113185f $X=3.155 $Y=0.34
+ $X2=0 $Y2=0
cc_1222 N_A_200_74#_c_1980_n N_A_430_362#_c_2053_n 0.0133617f $X=1.92 $Y=0.895
+ $X2=0 $Y2=0
cc_1223 N_A_200_74#_M1019_d N_A_430_362#_c_2058_n 0.00899348f $X=3.11 $Y=1.81
+ $X2=0 $Y2=0
cc_1224 N_A_200_74#_c_1955_n N_A_430_362#_c_2058_n 0.0340276f $X=3.165 $Y=2.715
+ $X2=0 $Y2=0
cc_1225 N_A_200_74#_c_1956_n N_A_430_362#_c_2058_n 0.0249199f $X=3.33 $Y=2.715
+ $X2=0 $Y2=0
cc_1226 N_A_200_74#_c_1955_n N_A_430_362#_c_2086_n 0.0193975f $X=3.165 $Y=2.715
+ $X2=0 $Y2=0
cc_1227 N_A_200_74#_c_1944_n N_VGND_M1007_s 0.00976727f $X=1.835 $Y=0.895 $X2=0
+ $Y2=0
cc_1228 N_A_200_74#_c_1946_n N_VGND_M1007_s 0.00716393f $X=1.92 $Y=2.63 $X2=0
+ $Y2=0
cc_1229 N_A_200_74#_c_1947_n N_VGND_M1007_s 0.00495363f $X=2.05 $Y=0.79 $X2=0
+ $Y2=0
cc_1230 N_A_200_74#_c_1980_n N_VGND_M1007_s 0.00341922f $X=1.92 $Y=0.895 $X2=0
+ $Y2=0
cc_1231 N_A_200_74#_c_1943_n N_VGND_c_2353_n 0.0164623f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_1232 N_A_200_74#_c_1943_n N_VGND_c_2354_n 0.0178806f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_1233 N_A_200_74#_c_1944_n N_VGND_c_2354_n 0.0208409f $X=1.835 $Y=0.895 $X2=0
+ $Y2=0
cc_1234 N_A_200_74#_c_1947_n N_VGND_c_2354_n 0.014651f $X=2.05 $Y=0.79 $X2=0
+ $Y2=0
cc_1235 N_A_200_74#_c_1949_n N_VGND_c_2354_n 0.0146193f $X=2.135 $Y=0.34 $X2=0
+ $Y2=0
cc_1236 N_A_200_74#_c_1948_n N_VGND_c_2365_n 0.0827822f $X=3.155 $Y=0.34 $X2=0
+ $Y2=0
cc_1237 N_A_200_74#_c_1949_n N_VGND_c_2365_n 0.0122124f $X=2.135 $Y=0.34 $X2=0
+ $Y2=0
cc_1238 N_A_200_74#_c_1943_n N_VGND_c_2373_n 0.0145162f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_1239 N_A_200_74#_c_1943_n N_VGND_c_2380_n 0.0119798f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_1240 N_A_200_74#_c_1944_n N_VGND_c_2380_n 0.0108847f $X=1.835 $Y=0.895 $X2=0
+ $Y2=0
cc_1241 N_A_200_74#_c_1948_n N_VGND_c_2380_n 0.0463404f $X=3.155 $Y=0.34 $X2=0
+ $Y2=0
cc_1242 N_A_200_74#_c_1949_n N_VGND_c_2380_n 0.00661405f $X=2.135 $Y=0.34 $X2=0
+ $Y2=0
cc_1243 N_A_200_74#_c_1980_n N_VGND_c_2380_n 0.00535727f $X=1.92 $Y=0.895 $X2=0
+ $Y2=0
cc_1244 N_A_1183_102#_c_2143_n N_COUT_c_2249_n 0.0070394f $X=9.36 $Y=1.665 $X2=0
+ $Y2=0
cc_1245 N_COUT_c_2245_n N_VGND_M1011_s 0.00352697f $X=11.177 $Y=1.135 $X2=0
+ $Y2=0
cc_1246 N_SUM_c_2310_n N_VGND_M1028_d 0.00330483f $X=14.495 $Y=1.095 $X2=0 $Y2=0
cc_1247 N_SUM_c_2290_n N_VGND_c_2359_n 0.00148977f $X=13.72 $Y=0.645 $X2=0 $Y2=0
cc_1248 N_SUM_c_2290_n N_VGND_c_2360_n 0.0136308f $X=13.72 $Y=0.645 $X2=0 $Y2=0
cc_1249 N_SUM_c_2310_n N_VGND_c_2360_n 0.0170777f $X=14.495 $Y=1.095 $X2=0 $Y2=0
cc_1250 N_SUM_c_2291_n N_VGND_c_2360_n 0.0136308f $X=14.58 $Y=0.645 $X2=0 $Y2=0
cc_1251 N_SUM_c_2291_n N_VGND_c_2362_n 0.019813f $X=14.58 $Y=0.645 $X2=0 $Y2=0
cc_1252 N_SUM_c_2292_n N_VGND_c_2362_n 0.0036313f $X=14.62 $Y=1.85 $X2=0 $Y2=0
cc_1253 N_SUM_c_2290_n N_VGND_c_2375_n 0.00718756f $X=13.72 $Y=0.645 $X2=0 $Y2=0
cc_1254 N_SUM_c_2291_n N_VGND_c_2376_n 0.00717249f $X=14.58 $Y=0.645 $X2=0 $Y2=0
cc_1255 N_SUM_c_2290_n N_VGND_c_2380_n 0.0083989f $X=13.72 $Y=0.645 $X2=0 $Y2=0
cc_1256 N_SUM_c_2291_n N_VGND_c_2380_n 0.00838881f $X=14.58 $Y=0.645 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o2bb2ai_1.spice
* Created: Wed Sep  2 12:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2bb2ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o2bb2ai_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1009 A_114_74# N_A1_N_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1004 N_A_134_383#_M1004_d N_A2_N_M1004_g A_114_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_397_74#_M1008_d N_A_134_383#_M1008_g N_Y_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_B2_M1007_g N_A_397_74#_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1000 N_A_397_74#_M1000_d N_B1_M1000_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_134_383#_M1005_d N_A1_N_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2772 PD=1.11 PS=2.34 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.2 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1006 N_VPWR_M1006_d N_A2_N_M1006_g N_A_134_383#_M1005_d VPB PSHORT L=0.18
+ W=0.84 AD=0.305411 AS=0.1134 PD=1.57286 PS=1.11 NRD=39.0848 NRS=0 M=1
+ R=4.66667 SA=90000.7 SB=90002 A=0.1512 P=2.04 MULT=1
MM1001 N_Y_M1001_d N_A_134_383#_M1001_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.407214 PD=1.39 PS=2.09714 NRD=0 NRS=26.9693 M=1 R=6.22222
+ SA=90001.3 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1003 A_493_368# N_B2_M1003_g N_Y_M1001_d VPB PSHORT L=0.18 W=1.12 AD=0.168
+ AS=0.1512 PD=1.42 PS=1.39 NRD=16.7056 NRS=0 M=1 R=6.22222 SA=90001.7
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g A_493_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.168 PD=2.8 PS=1.42 NRD=0 NRS=16.7056 M=1 R=6.22222 SA=90002.2 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__o2bb2ai_1.pxi.spice"
*
.ends
*
*

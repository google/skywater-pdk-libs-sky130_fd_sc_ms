* NGSPICE file created from sky130_fd_sc_ms__o2bb2a_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_270_48# A2_N VPWR VPB pshort w=840000u l=180000u
+  ad=3.024e+11p pd=2.4e+06u as=1.68435e+12p ps=1.199e+07u
M1001 X a_204_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=7.087e+11p ps=6.4e+06u
M1002 VPWR A1_N a_270_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_500_74# A2_N a_270_48# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1004 VPWR a_270_48# a_204_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1005 a_204_392# a_270_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=4.699e+11p ps=4.23e+06u
M1006 a_120_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND A1_N a_500_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_204_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 VGND B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_204_392# B2 a_120_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_204_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_204_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


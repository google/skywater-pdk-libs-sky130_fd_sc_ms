* File: sky130_fd_sc_ms__a222o_2.pxi.spice
* Created: Fri Aug 28 17:02:03 2020
* 
x_PM_SKY130_FD_SC_MS__A222O_2%C1 N_C1_c_98_n N_C1_M1001_g N_C1_M1004_g
+ N_C1_c_95_n C1 N_C1_c_96_n N_C1_c_97_n PM_SKY130_FD_SC_MS__A222O_2%C1
x_PM_SKY130_FD_SC_MS__A222O_2%C2 N_C2_M1015_g N_C2_M1002_g C2 N_C2_c_128_n
+ N_C2_c_129_n PM_SKY130_FD_SC_MS__A222O_2%C2
x_PM_SKY130_FD_SC_MS__A222O_2%A_27_82# N_A_27_82#_M1004_s N_A_27_82#_M1007_d
+ N_A_27_82#_M1001_s N_A_27_82#_M1002_d N_A_27_82#_c_161_n N_A_27_82#_M1005_g
+ N_A_27_82#_c_162_n N_A_27_82#_c_163_n N_A_27_82#_M1006_g N_A_27_82#_c_165_n
+ N_A_27_82#_M1010_g N_A_27_82#_M1008_g N_A_27_82#_c_166_n N_A_27_82#_c_178_n
+ N_A_27_82#_c_179_n N_A_27_82#_c_167_n N_A_27_82#_c_168_n N_A_27_82#_c_180_n
+ N_A_27_82#_c_203_n N_A_27_82#_c_169_n N_A_27_82#_c_170_n N_A_27_82#_c_262_p
+ N_A_27_82#_c_247_p N_A_27_82#_c_171_n N_A_27_82#_c_172_n N_A_27_82#_c_173_n
+ N_A_27_82#_c_263_p N_A_27_82#_c_174_n N_A_27_82#_c_175_n
+ PM_SKY130_FD_SC_MS__A222O_2%A_27_82#
x_PM_SKY130_FD_SC_MS__A222O_2%A1 N_A1_M1003_g N_A1_M1007_g A1 A1 N_A1_c_293_n
+ N_A1_c_294_n PM_SKY130_FD_SC_MS__A222O_2%A1
x_PM_SKY130_FD_SC_MS__A222O_2%B1 N_B1_M1013_g N_B1_M1011_g B1 N_B1_c_335_n
+ N_B1_c_336_n PM_SKY130_FD_SC_MS__A222O_2%B1
x_PM_SKY130_FD_SC_MS__A222O_2%B2 N_B2_M1012_g N_B2_M1014_g B2 N_B2_c_371_n
+ N_B2_c_372_n PM_SKY130_FD_SC_MS__A222O_2%B2
x_PM_SKY130_FD_SC_MS__A222O_2%A2 N_A2_M1000_g N_A2_M1009_g A2 N_A2_c_411_n
+ PM_SKY130_FD_SC_MS__A222O_2%A2
x_PM_SKY130_FD_SC_MS__A222O_2%A_119_392# N_A_119_392#_M1001_d
+ N_A_119_392#_M1013_d N_A_119_392#_c_436_n N_A_119_392#_c_451_n
+ N_A_119_392#_c_437_n PM_SKY130_FD_SC_MS__A222O_2%A_119_392#
x_PM_SKY130_FD_SC_MS__A222O_2%VPWR N_VPWR_M1006_s N_VPWR_M1008_s N_VPWR_M1009_d
+ N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n
+ N_VPWR_c_477_n VPWR N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n
+ N_VPWR_c_471_n PM_SKY130_FD_SC_MS__A222O_2%VPWR
x_PM_SKY130_FD_SC_MS__A222O_2%X N_X_M1005_d N_X_M1006_d N_X_c_522_n X
+ N_X_c_524_n PM_SKY130_FD_SC_MS__A222O_2%X
x_PM_SKY130_FD_SC_MS__A222O_2%A_642_368# N_A_642_368#_M1003_d
+ N_A_642_368#_M1014_d N_A_642_368#_c_550_n N_A_642_368#_c_551_n
+ N_A_642_368#_c_552_n PM_SKY130_FD_SC_MS__A222O_2%A_642_368#
x_PM_SKY130_FD_SC_MS__A222O_2%VGND N_VGND_M1015_d N_VGND_M1010_s N_VGND_M1012_d
+ N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n
+ N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n VGND N_VGND_c_581_n
+ N_VGND_c_582_n PM_SKY130_FD_SC_MS__A222O_2%VGND
x_PM_SKY130_FD_SC_MS__A222O_2%A_557_74# N_A_557_74#_M1007_s N_A_557_74#_M1000_d
+ N_A_557_74#_c_636_n N_A_557_74#_c_673_p N_A_557_74#_c_637_n
+ N_A_557_74#_c_638_n N_A_557_74#_c_639_n N_A_557_74#_c_640_n
+ PM_SKY130_FD_SC_MS__A222O_2%A_557_74#
cc_1 VNB N_C1_M1004_g 0.0329894f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_C1_c_95_n 0.00186909f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.83
cc_3 VNB N_C1_c_96_n 0.00453376f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_C1_c_97_n 0.0575289f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_5 VNB N_C2_M1015_g 0.0237179f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.92
cc_6 VNB N_C2_M1002_g 0.00425652f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_7 VNB N_C2_c_128_n 0.03207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_C2_c_129_n 0.00834647f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_9 VNB N_A_27_82#_c_161_n 0.0182542f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_A_27_82#_c_162_n 0.013455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_82#_c_163_n 0.013716f $X=-0.19 $Y=-0.245 $X2=0.492 $Y2=1.465
cc_12 VNB N_A_27_82#_M1006_g 0.00447002f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_13 VNB N_A_27_82#_c_165_n 0.0165924f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_14 VNB N_A_27_82#_c_166_n 0.0220451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_82#_c_167_n 0.0109097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_82#_c_168_n 0.00886217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_82#_c_169_n 0.0102068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_82#_c_170_n 0.0021754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_82#_c_171_n 0.00257009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_82#_c_172_n 0.0538084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_82#_c_173_n 0.0255526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_82#_c_174_n 0.00378718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_82#_c_175_n 0.0103491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_M1007_g 0.0367638f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_25 VNB N_A1_c_293_n 0.028052f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_26 VNB N_A1_c_294_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_27 VNB N_B1_M1011_g 0.0313709f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_28 VNB N_B1_c_335_n 0.0315864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_336_n 0.00240839f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_30 VNB N_B2_M1012_g 0.0290869f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.92
cc_31 VNB N_B2_c_371_n 0.0224753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B2_c_372_n 0.0054107f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_33 VNB N_A2_M1000_g 0.0411723f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.92
cc_34 VNB A2 0.0159538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_411_n 0.0276826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_471_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_522_n 0.00209829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_573_n 0.00881119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_574_n 0.00671846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_575_n 0.0301057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_576_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_42 VNB N_VGND_c_577_n 0.0168493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_578_n 0.0282128f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_44 VNB N_VGND_c_579_n 0.0443678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_580_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_581_n 0.0215382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_582_n 0.330142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_557_74#_c_636_n 0.00610588f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_49 VNB N_A_557_74#_c_637_n 0.0269419f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_50 VNB N_A_557_74#_c_638_n 0.00403445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_557_74#_c_639_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_52 VNB N_A_557_74#_c_640_n 0.00917671f $X=-0.19 $Y=-0.245 $X2=0.492 $Y2=1.465
cc_53 VPB N_C1_c_98_n 0.0287202f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.92
cc_54 VPB N_C1_c_95_n 0.0118236f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.83
cc_55 VPB N_C1_c_96_n 0.00761937f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_56 VPB N_C2_M1002_g 0.0333956f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.73
cc_57 VPB N_C2_c_129_n 0.00530202f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_58 VPB N_A_27_82#_M1006_g 0.0251695f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_59 VPB N_A_27_82#_M1008_g 0.0232164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_82#_c_178_n 0.0120621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_27_82#_c_179_n 0.031021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_82#_c_180_n 0.0167668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_82#_c_169_n 0.00644725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_82#_c_172_n 0.00114409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A1_M1003_g 0.0229618f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.92
cc_66 VPB N_A1_c_293_n 0.00569525f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_67 VPB N_A1_c_294_n 0.0033873f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_68 VPB N_B1_M1013_g 0.0220617f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.92
cc_69 VPB N_B1_c_335_n 0.00810167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_B1_c_336_n 0.00419737f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_71 VPB N_B2_M1014_g 0.0206455f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.73
cc_72 VPB N_B2_c_371_n 0.00545172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_B2_c_372_n 0.00495473f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_74 VPB N_A2_M1009_g 0.0258337f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.73
cc_75 VPB A2 0.00822096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A2_c_411_n 0.00579252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_119_392#_c_436_n 0.015467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_119_392#_c_437_n 0.00231152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_472_n 0.0149882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_473_n 0.0106611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_474_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_82 VPB N_VPWR_c_475_n 0.0513304f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_83 VPB N_VPWR_c_476_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_477_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_478_n 0.0477633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_479_n 0.0459735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_480_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_471_n 0.0822233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_X_c_522_n 0.00248928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_X_c_524_n 0.0089111f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_91 VPB N_A_642_368#_c_550_n 0.0140479f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.73
cc_92 VPB N_A_642_368#_c_551_n 0.00136426f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_93 VPB N_A_642_368#_c_552_n 0.00618782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 N_C1_M1004_g N_C2_M1015_g 0.0346947f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_95 N_C1_c_98_n N_C2_M1002_g 0.0281221f $X=0.505 $Y=1.92 $X2=0 $Y2=0
cc_96 N_C1_c_97_n N_C2_M1002_g 0.00962598f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_97 N_C1_c_96_n N_C2_c_128_n 2.1027e-19 $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_98 N_C1_c_97_n N_C2_c_128_n 0.0346947f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_99 N_C1_M1004_g N_C2_c_129_n 0.00533482f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_100 N_C1_c_96_n N_C2_c_129_n 0.0395606f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_101 N_C1_M1004_g N_A_27_82#_c_166_n 5.45389e-19 $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_102 N_C1_c_96_n N_A_27_82#_c_178_n 0.0228254f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_103 N_C1_c_97_n N_A_27_82#_c_178_n 0.00137994f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_104 N_C1_c_98_n N_A_27_82#_c_179_n 4.69176e-19 $X=0.505 $Y=1.92 $X2=0 $Y2=0
cc_105 N_C1_M1004_g N_A_27_82#_c_167_n 0.0174317f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_106 N_C1_c_96_n N_A_27_82#_c_167_n 0.00448606f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_107 N_C1_c_97_n N_A_27_82#_c_167_n 3.67789e-19 $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_108 N_C1_c_96_n N_A_27_82#_c_168_n 0.0185799f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_109 N_C1_c_97_n N_A_27_82#_c_168_n 0.00192177f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_110 N_C1_c_98_n N_A_27_82#_c_180_n 0.0220105f $X=0.505 $Y=1.92 $X2=0 $Y2=0
cc_111 N_C1_c_96_n N_A_27_82#_c_180_n 0.00562319f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_112 N_C1_c_97_n N_A_27_82#_c_180_n 2.49658e-19 $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_113 N_C1_c_98_n N_A_119_392#_c_437_n 0.00848316f $X=0.505 $Y=1.92 $X2=0 $Y2=0
cc_114 N_C1_c_98_n N_VPWR_c_478_n 0.005209f $X=0.505 $Y=1.92 $X2=0 $Y2=0
cc_115 N_C1_c_98_n N_VPWR_c_471_n 0.00987216f $X=0.505 $Y=1.92 $X2=0 $Y2=0
cc_116 N_C1_M1004_g N_VGND_c_573_n 0.00160827f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_117 N_C1_M1004_g N_VGND_c_575_n 0.00548708f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_118 N_C1_M1004_g N_VGND_c_582_n 0.00533081f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_119 N_C2_M1015_g N_A_27_82#_c_161_n 0.009666f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_120 N_C2_c_128_n N_A_27_82#_c_163_n 0.00361438f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_121 N_C2_M1015_g N_A_27_82#_c_167_n 0.0150237f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_122 N_C2_c_128_n N_A_27_82#_c_167_n 0.00437059f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_123 N_C2_c_129_n N_A_27_82#_c_167_n 0.0419923f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_124 N_C2_M1002_g N_A_27_82#_c_180_n 0.0121686f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_125 N_C2_c_128_n N_A_27_82#_c_180_n 6.93298e-19 $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_126 N_C2_c_129_n N_A_27_82#_c_180_n 0.0437162f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_127 N_C2_M1015_g N_A_27_82#_c_203_n 0.00296638f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_128 N_C2_M1015_g N_A_27_82#_c_169_n 0.00304065f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_129 N_C2_M1002_g N_A_27_82#_c_169_n 0.00615715f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_130 N_C2_c_128_n N_A_27_82#_c_169_n 0.001751f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_131 N_C2_c_129_n N_A_27_82#_c_169_n 0.0348642f $X=0.975 $Y=1.425 $X2=0 $Y2=0
cc_132 N_C2_M1002_g N_A_119_392#_c_436_n 0.0117345f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_133 N_C2_M1002_g N_A_119_392#_c_437_n 0.0207448f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_134 N_C2_M1002_g N_VPWR_c_472_n 0.00980832f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_135 N_C2_M1002_g N_VPWR_c_478_n 0.005209f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_136 N_C2_M1002_g N_VPWR_c_471_n 0.00526773f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_137 N_C2_M1002_g N_X_c_524_n 5.12846e-19 $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_138 N_C2_M1015_g N_VGND_c_573_n 0.0110632f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_139 N_C2_M1015_g N_VGND_c_575_n 0.00455951f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_140 N_C2_M1015_g N_VGND_c_582_n 0.00447788f $X=0.885 $Y=0.73 $X2=0 $Y2=0
cc_141 N_A_27_82#_M1008_g N_A1_M1003_g 0.0326016f $X=2.5 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_27_82#_c_171_n N_A1_M1007_g 0.00245637f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_143 N_A_27_82#_c_172_n N_A1_M1007_g 0.00233427f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_144 N_A_27_82#_c_173_n N_A1_M1007_g 0.0132844f $X=3.265 $Y=1.095 $X2=0 $Y2=0
cc_145 N_A_27_82#_c_175_n N_A1_M1007_g 0.00113123f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_146 N_A_27_82#_c_171_n N_A1_c_293_n 9.97553e-19 $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_147 N_A_27_82#_c_172_n N_A1_c_293_n 0.0114142f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_148 N_A_27_82#_c_173_n N_A1_c_293_n 0.00125479f $X=3.265 $Y=1.095 $X2=0 $Y2=0
cc_149 N_A_27_82#_M1008_g N_A1_c_294_n 0.00573829f $X=2.5 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_27_82#_c_171_n N_A1_c_294_n 0.00975019f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_151 N_A_27_82#_c_172_n N_A1_c_294_n 0.00168361f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_152 N_A_27_82#_c_173_n N_A1_c_294_n 0.0256551f $X=3.265 $Y=1.095 $X2=0 $Y2=0
cc_153 N_A_27_82#_c_175_n N_B1_M1011_g 0.0132613f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_154 N_A_27_82#_c_175_n N_B1_c_335_n 0.0019768f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_155 N_A_27_82#_c_175_n N_B1_c_336_n 0.0236445f $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_156 N_A_27_82#_c_175_n N_B2_M1012_g 2.25597e-19 $X=3.505 $Y=0.865 $X2=0 $Y2=0
cc_157 N_A_27_82#_c_180_n N_A_119_392#_M1001_d 0.00167813f $X=1.355 $Y=2.075
+ $X2=-0.19 $Y2=-0.245
cc_158 N_A_27_82#_M1002_d N_A_119_392#_c_436_n 0.0075965f $X=1.045 $Y=1.96 $X2=0
+ $Y2=0
cc_159 N_A_27_82#_M1006_g N_A_119_392#_c_436_n 0.0152738f $X=2.05 $Y=2.4 $X2=0
+ $Y2=0
cc_160 N_A_27_82#_M1008_g N_A_119_392#_c_436_n 0.0185309f $X=2.5 $Y=2.4 $X2=0
+ $Y2=0
cc_161 N_A_27_82#_c_180_n N_A_119_392#_c_436_n 0.0436386f $X=1.355 $Y=2.075
+ $X2=0 $Y2=0
cc_162 N_A_27_82#_c_179_n N_A_119_392#_c_437_n 0.015139f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_27_82#_c_180_n N_A_119_392#_c_437_n 0.0174907f $X=1.355 $Y=2.075
+ $X2=0 $Y2=0
cc_164 N_A_27_82#_M1006_g N_VPWR_c_472_n 0.0105025f $X=2.05 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A_27_82#_M1008_g N_VPWR_c_473_n 0.00698686f $X=2.5 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_27_82#_M1006_g N_VPWR_c_476_n 0.00553757f $X=2.05 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A_27_82#_M1008_g N_VPWR_c_476_n 0.00553757f $X=2.5 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A_27_82#_c_179_n N_VPWR_c_478_n 0.011066f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_27_82#_M1006_g N_VPWR_c_471_n 0.00545239f $X=2.05 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A_27_82#_M1008_g N_VPWR_c_471_n 0.00545239f $X=2.5 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_27_82#_c_179_n N_VPWR_c_471_n 0.00915947f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_27_82#_c_170_n N_X_M1005_d 0.00435233f $X=2.23 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_27_82#_c_161_n N_X_c_522_n 0.0052405f $X=1.645 $Y=1.26 $X2=0 $Y2=0
cc_174 N_A_27_82#_c_162_n N_X_c_522_n 0.0105762f $X=1.96 $Y=1.335 $X2=0 $Y2=0
cc_175 N_A_27_82#_c_163_n N_X_c_522_n 0.00207346f $X=1.72 $Y=1.335 $X2=0 $Y2=0
cc_176 N_A_27_82#_M1006_g N_X_c_522_n 0.00966798f $X=2.05 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_27_82#_c_165_n N_X_c_522_n 0.00554882f $X=2.075 $Y=1.26 $X2=0 $Y2=0
cc_178 N_A_27_82#_c_169_n N_X_c_522_n 0.0542206f $X=1.44 $Y=1.95 $X2=0 $Y2=0
cc_179 N_A_27_82#_c_170_n N_X_c_522_n 0.0170777f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_180 N_A_27_82#_c_247_p N_X_c_522_n 0.00572056f $X=2.315 $Y=1.01 $X2=0 $Y2=0
cc_181 N_A_27_82#_c_171_n N_X_c_522_n 0.0267529f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_182 N_A_27_82#_c_172_n N_X_c_522_n 0.0117993f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_183 N_A_27_82#_c_174_n N_X_c_522_n 0.012203f $X=2.395 $Y=1.095 $X2=0 $Y2=0
cc_184 N_A_27_82#_c_163_n N_X_c_524_n 7.04168e-19 $X=1.72 $Y=1.335 $X2=0 $Y2=0
cc_185 N_A_27_82#_M1006_g N_X_c_524_n 0.022345f $X=2.05 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A_27_82#_M1008_g N_X_c_524_n 0.0083454f $X=2.5 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_27_82#_c_180_n N_X_c_524_n 0.0233303f $X=1.355 $Y=2.075 $X2=0 $Y2=0
cc_188 N_A_27_82#_c_169_n N_X_c_524_n 0.0108574f $X=1.44 $Y=1.95 $X2=0 $Y2=0
cc_189 N_A_27_82#_c_171_n N_X_c_524_n 0.0139616f $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_190 N_A_27_82#_c_172_n N_X_c_524_n 6.34955e-19 $X=2.395 $Y=1.425 $X2=0 $Y2=0
cc_191 N_A_27_82#_c_167_n A_114_82# 0.0048076f $X=1.355 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_27_82#_c_167_n N_VGND_M1015_d 0.0111604f $X=1.355 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_27_82#_c_203_n N_VGND_M1015_d 0.00267073f $X=1.44 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_27_82#_c_169_n N_VGND_M1015_d 0.00133961f $X=1.44 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_27_82#_c_262_p N_VGND_M1015_d 0.00463907f $X=1.525 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_27_82#_c_263_p N_VGND_M1015_d 0.00142544f $X=1.44 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_27_82#_c_170_n N_VGND_M1010_s 0.00562426f $X=2.23 $Y=0.665 $X2=0
+ $Y2=0
cc_198 N_A_27_82#_c_247_p N_VGND_M1010_s 0.011885f $X=2.315 $Y=1.01 $X2=0 $Y2=0
cc_199 N_A_27_82#_c_174_n N_VGND_M1010_s 0.00193901f $X=2.395 $Y=1.095 $X2=0
+ $Y2=0
cc_200 N_A_27_82#_c_161_n N_VGND_c_573_n 0.0062784f $X=1.645 $Y=1.26 $X2=0 $Y2=0
cc_201 N_A_27_82#_c_166_n N_VGND_c_573_n 0.00509935f $X=0.28 $Y=0.555 $X2=0
+ $Y2=0
cc_202 N_A_27_82#_c_167_n N_VGND_c_573_n 0.015373f $X=1.355 $Y=1.005 $X2=0 $Y2=0
cc_203 N_A_27_82#_c_262_p N_VGND_c_573_n 0.0141996f $X=1.525 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_27_82#_c_166_n N_VGND_c_575_n 0.00955085f $X=0.28 $Y=0.555 $X2=0
+ $Y2=0
cc_205 N_A_27_82#_c_165_n N_VGND_c_577_n 0.00546687f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_206 N_A_27_82#_c_170_n N_VGND_c_577_n 0.0157799f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_27_82#_c_174_n N_VGND_c_577_n 0.00480154f $X=2.395 $Y=1.095 $X2=0
+ $Y2=0
cc_208 N_A_27_82#_c_161_n N_VGND_c_578_n 0.00414982f $X=1.645 $Y=1.26 $X2=0
+ $Y2=0
cc_209 N_A_27_82#_c_165_n N_VGND_c_578_n 0.00414982f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_210 N_A_27_82#_c_170_n N_VGND_c_578_n 0.0113015f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_211 N_A_27_82#_c_262_p N_VGND_c_578_n 0.00358211f $X=1.525 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_27_82#_c_161_n N_VGND_c_582_n 0.00533081f $X=1.645 $Y=1.26 $X2=0
+ $Y2=0
cc_213 N_A_27_82#_c_165_n N_VGND_c_582_n 0.00533081f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_214 N_A_27_82#_c_166_n N_VGND_c_582_n 0.00894475f $X=0.28 $Y=0.555 $X2=0
+ $Y2=0
cc_215 N_A_27_82#_c_170_n N_VGND_c_582_n 0.0210788f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_216 N_A_27_82#_c_262_p N_VGND_c_582_n 0.00537088f $X=1.525 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_27_82#_M1007_d N_A_557_74#_c_636_n 0.00478343f $X=3.255 $Y=0.37 $X2=0
+ $Y2=0
cc_218 N_A_27_82#_c_173_n N_A_557_74#_c_636_n 0.00462336f $X=3.265 $Y=1.095
+ $X2=0 $Y2=0
cc_219 N_A_27_82#_c_175_n N_A_557_74#_c_636_n 0.0272186f $X=3.505 $Y=0.865 $X2=0
+ $Y2=0
cc_220 N_A_27_82#_c_175_n N_A_557_74#_c_638_n 0.0146766f $X=3.505 $Y=0.865 $X2=0
+ $Y2=0
cc_221 N_A_27_82#_c_165_n N_A_557_74#_c_640_n 0.00501373f $X=2.075 $Y=1.26 $X2=0
+ $Y2=0
cc_222 N_A_27_82#_c_170_n N_A_557_74#_c_640_n 0.00852177f $X=2.23 $Y=0.665 $X2=0
+ $Y2=0
cc_223 N_A_27_82#_c_247_p N_A_557_74#_c_640_n 0.00405254f $X=2.315 $Y=1.01 $X2=0
+ $Y2=0
cc_224 N_A_27_82#_c_173_n N_A_557_74#_c_640_n 0.0244887f $X=3.265 $Y=1.095 $X2=0
+ $Y2=0
cc_225 N_A1_M1003_g N_B1_M1013_g 0.0283061f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_226 N_A1_c_294_n N_B1_M1013_g 0.00243977f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A1_M1007_g N_B1_M1011_g 0.0259476f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_228 N_A1_c_293_n N_B1_c_335_n 0.0204459f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A1_c_294_n N_B1_c_335_n 0.00119705f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_230 N_A1_M1003_g N_B1_c_336_n 3.74161e-19 $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_231 N_A1_c_293_n N_B1_c_336_n 0.00114936f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_232 N_A1_c_294_n N_B1_c_336_n 0.0280926f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_233 N_A1_M1003_g N_A_119_392#_c_436_n 0.0158932f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_234 N_A1_c_293_n N_A_119_392#_c_436_n 2.26286e-19 $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_235 N_A1_c_294_n N_A_119_392#_c_436_n 0.0143022f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_236 N_A1_M1003_g N_A_119_392#_c_451_n 0.00114348f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_237 N_A1_c_294_n N_VPWR_M1008_s 0.00501169f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A1_M1003_g N_VPWR_c_473_n 0.00234955f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_239 N_A1_M1003_g N_VPWR_c_479_n 0.0059286f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_240 N_A1_M1003_g N_VPWR_c_471_n 0.00610055f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_241 N_A1_M1003_g N_X_c_524_n 5.08955e-19 $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_242 N_A1_c_294_n N_X_c_524_n 0.0119982f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_243 N_A1_M1003_g N_A_642_368#_c_552_n 0.00247266f $X=3.12 $Y=2.34 $X2=0 $Y2=0
cc_244 N_A1_M1007_g N_VGND_c_577_n 0.00265086f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_245 N_A1_M1007_g N_VGND_c_579_n 0.00291649f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_246 N_A1_M1007_g N_VGND_c_582_n 0.00365718f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_247 N_A1_M1007_g N_A_557_74#_c_636_n 0.0115929f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_248 N_A1_M1007_g N_A_557_74#_c_640_n 0.00168345f $X=3.18 $Y=0.69 $X2=0 $Y2=0
cc_249 N_B1_M1011_g N_B2_M1012_g 0.0355648f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_250 N_B1_M1013_g N_B2_M1014_g 0.0242598f $X=3.775 $Y=2.34 $X2=0 $Y2=0
cc_251 N_B1_c_335_n N_B2_c_371_n 0.0355648f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_252 N_B1_c_336_n N_B2_c_371_n 2.7993e-19 $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_253 N_B1_M1013_g N_B2_c_372_n 6.9747e-19 $X=3.775 $Y=2.34 $X2=0 $Y2=0
cc_254 N_B1_c_335_n N_B2_c_372_n 0.00249096f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_255 N_B1_c_336_n N_B2_c_372_n 0.0350349f $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_256 N_B1_M1013_g N_A_119_392#_c_436_n 0.0180423f $X=3.775 $Y=2.34 $X2=0 $Y2=0
cc_257 N_B1_c_335_n N_A_119_392#_c_436_n 8.0354e-19 $X=3.63 $Y=1.515 $X2=0 $Y2=0
cc_258 N_B1_c_336_n N_A_119_392#_c_436_n 0.00918305f $X=3.63 $Y=1.515 $X2=0
+ $Y2=0
cc_259 N_B1_M1013_g N_A_119_392#_c_451_n 0.0110441f $X=3.775 $Y=2.34 $X2=0 $Y2=0
cc_260 N_B1_M1013_g N_VPWR_c_479_n 8.71493e-19 $X=3.775 $Y=2.34 $X2=0 $Y2=0
cc_261 N_B1_M1013_g N_A_642_368#_c_550_n 0.00882386f $X=3.775 $Y=2.34 $X2=0
+ $Y2=0
cc_262 N_B1_M1013_g N_A_642_368#_c_552_n 0.00306464f $X=3.775 $Y=2.34 $X2=0
+ $Y2=0
cc_263 N_B1_M1011_g N_VGND_c_574_n 7.59698e-19 $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_264 N_B1_M1011_g N_VGND_c_579_n 0.00291649f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_265 N_B1_M1011_g N_VGND_c_582_n 0.00360429f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_266 N_B1_M1011_g N_A_557_74#_c_636_n 0.0139417f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_267 N_B1_M1011_g N_A_557_74#_c_638_n 0.00130469f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_268 N_B2_M1012_g N_A2_M1000_g 0.0231299f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_269 N_B2_M1014_g N_A2_M1009_g 0.0088376f $X=4.225 $Y=2.34 $X2=0 $Y2=0
cc_270 N_B2_c_372_n N_A2_M1009_g 4.22075e-19 $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_271 N_B2_c_371_n A2 4.19559e-19 $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_272 N_B2_c_372_n A2 0.0263802f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_273 N_B2_c_371_n N_A2_c_411_n 0.0181621f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_274 N_B2_c_372_n N_A2_c_411_n 4.19449e-19 $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_275 N_B2_M1014_g N_A_119_392#_c_436_n 0.00462888f $X=4.225 $Y=2.34 $X2=0
+ $Y2=0
cc_276 N_B2_M1014_g N_A_119_392#_c_451_n 0.00583417f $X=4.225 $Y=2.34 $X2=0
+ $Y2=0
cc_277 N_B2_c_372_n N_A_119_392#_c_451_n 0.0147873f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_278 N_B2_M1014_g N_VPWR_c_475_n 2.45511e-19 $X=4.225 $Y=2.34 $X2=0 $Y2=0
cc_279 N_B2_M1014_g N_VPWR_c_479_n 8.71493e-19 $X=4.225 $Y=2.34 $X2=0 $Y2=0
cc_280 N_B2_M1014_g N_A_642_368#_c_550_n 0.0126323f $X=4.225 $Y=2.34 $X2=0 $Y2=0
cc_281 N_B2_M1014_g N_A_642_368#_c_551_n 0.00188914f $X=4.225 $Y=2.34 $X2=0
+ $Y2=0
cc_282 N_B2_c_371_n N_A_642_368#_c_551_n 5.81599e-19 $X=4.28 $Y=1.515 $X2=0
+ $Y2=0
cc_283 N_B2_c_372_n N_A_642_368#_c_551_n 0.00801953f $X=4.28 $Y=1.515 $X2=0
+ $Y2=0
cc_284 N_B2_M1012_g N_VGND_c_574_n 0.00890008f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_285 N_B2_M1012_g N_VGND_c_579_n 0.00444681f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_286 N_B2_M1012_g N_VGND_c_582_n 0.00877228f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_287 N_B2_M1012_g N_A_557_74#_c_636_n 7.44093e-19 $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_288 N_B2_M1012_g N_A_557_74#_c_637_n 0.0147396f $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_289 N_B2_c_371_n N_A_557_74#_c_637_n 0.00423269f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_290 N_B2_c_372_n N_A_557_74#_c_637_n 0.0267388f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_291 N_B2_c_372_n N_A_557_74#_c_638_n 0.011271f $X=4.28 $Y=1.515 $X2=0 $Y2=0
cc_292 N_B2_M1012_g N_A_557_74#_c_639_n 9.43881e-19 $X=4.19 $Y=0.69 $X2=0 $Y2=0
cc_293 N_A2_M1009_g N_VPWR_c_475_n 0.0190509f $X=4.775 $Y=2.34 $X2=0 $Y2=0
cc_294 A2 N_VPWR_c_475_n 0.0254126f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_295 N_A2_c_411_n N_VPWR_c_475_n 7.81657e-19 $X=4.85 $Y=1.515 $X2=0 $Y2=0
cc_296 N_A2_M1009_g N_VPWR_c_479_n 0.00492916f $X=4.775 $Y=2.34 $X2=0 $Y2=0
cc_297 N_A2_M1009_g N_VPWR_c_471_n 0.00511769f $X=4.775 $Y=2.34 $X2=0 $Y2=0
cc_298 N_A2_M1009_g N_A_642_368#_c_550_n 6.61023e-19 $X=4.775 $Y=2.34 $X2=0
+ $Y2=0
cc_299 N_A2_M1009_g N_A_642_368#_c_551_n 6.09564e-19 $X=4.775 $Y=2.34 $X2=0
+ $Y2=0
cc_300 N_A2_M1000_g N_VGND_c_574_n 0.00752319f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_301 N_A2_M1000_g N_VGND_c_581_n 0.00434272f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_302 N_A2_M1000_g N_VGND_c_582_n 0.00826173f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_303 N_A2_M1000_g N_A_557_74#_c_637_n 0.0159753f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_304 A2 N_A_557_74#_c_637_n 0.0378526f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_305 N_A2_c_411_n N_A_557_74#_c_637_n 0.00431154f $X=4.85 $Y=1.515 $X2=0 $Y2=0
cc_306 N_A2_M1000_g N_A_557_74#_c_639_n 0.00970393f $X=4.76 $Y=0.69 $X2=0 $Y2=0
cc_307 N_A_119_392#_c_436_n N_VPWR_M1006_s 0.00472277f $X=3.835 $Y=2.455
+ $X2=-0.19 $Y2=1.66
cc_308 N_A_119_392#_c_436_n N_VPWR_M1008_s 0.0153124f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_309 N_A_119_392#_c_436_n N_VPWR_c_472_n 0.0263858f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_310 N_A_119_392#_c_436_n N_VPWR_c_473_n 0.0258995f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_311 N_A_119_392#_c_437_n N_VPWR_c_478_n 0.0143496f $X=0.73 $Y=2.455 $X2=0
+ $Y2=0
cc_312 N_A_119_392#_c_436_n N_VPWR_c_471_n 0.0609947f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_313 N_A_119_392#_c_437_n N_VPWR_c_471_n 0.01179f $X=0.73 $Y=2.455 $X2=0 $Y2=0
cc_314 N_A_119_392#_c_436_n N_X_M1006_d 0.00466364f $X=3.835 $Y=2.455 $X2=0
+ $Y2=0
cc_315 N_A_119_392#_c_436_n N_X_c_524_n 0.043221f $X=3.835 $Y=2.455 $X2=0 $Y2=0
cc_316 N_A_119_392#_c_436_n N_A_642_368#_M1003_d 0.0152695f $X=3.835 $Y=2.455
+ $X2=-0.19 $Y2=1.66
cc_317 N_A_119_392#_c_436_n N_A_642_368#_c_550_n 0.0265678f $X=3.835 $Y=2.455
+ $X2=0 $Y2=0
cc_318 N_A_119_392#_c_436_n N_A_642_368#_c_552_n 0.0271648f $X=3.835 $Y=2.455
+ $X2=0 $Y2=0
cc_319 N_VPWR_M1006_s N_X_c_524_n 0.00349912f $X=1.595 $Y=2.73 $X2=0 $Y2=0
cc_320 N_VPWR_c_475_n N_A_642_368#_c_550_n 0.0147692f $X=5 $Y=2.115 $X2=0 $Y2=0
cc_321 N_VPWR_c_479_n N_A_642_368#_c_550_n 0.0690424f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_471_n N_A_642_368#_c_550_n 0.0393321f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_475_n N_A_642_368#_c_551_n 0.0384549f $X=5 $Y=2.115 $X2=0 $Y2=0
cc_324 N_VPWR_c_473_n N_A_642_368#_c_552_n 0.0135358f $X=2.81 $Y=2.875 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_479_n N_A_642_368#_c_552_n 0.0248486f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_471_n N_A_642_368#_c_552_n 0.0138941f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_327 N_VGND_c_574_n N_A_557_74#_c_636_n 0.00729485f $X=4.425 $Y=0.635 $X2=0
+ $Y2=0
cc_328 N_VGND_c_579_n N_A_557_74#_c_636_n 0.0401161f $X=4.26 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_582_n N_A_557_74#_c_636_n 0.0340164f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_574_n N_A_557_74#_c_637_n 0.0245379f $X=4.425 $Y=0.635 $X2=0
+ $Y2=0
cc_331 N_VGND_c_574_n N_A_557_74#_c_639_n 0.0312316f $X=4.425 $Y=0.635 $X2=0
+ $Y2=0
cc_332 N_VGND_c_581_n N_A_557_74#_c_639_n 0.0145639f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_582_n N_A_557_74#_c_639_n 0.0119984f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_c_577_n N_A_557_74#_c_640_n 0.00404517f $X=2.37 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_579_n N_A_557_74#_c_640_n 0.0142934f $X=4.26 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_c_582_n N_A_557_74#_c_640_n 0.0119825f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_337 N_A_557_74#_c_673_p A_775_74# 9.797e-19 $X=4.005 $Y=1.01 $X2=-0.19
+ $Y2=-0.245

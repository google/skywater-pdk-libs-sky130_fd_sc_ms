* File: sky130_fd_sc_ms__a32oi_4.pex.spice
* Created: Wed Sep  2 11:56:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A32OI_4%B2 3 7 11 15 19 23 27 31 33 34 35 36 55
c79 31 0 8.12065e-20 $X=1.92 $Y=0.74
r80 54 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.905 $Y=1.515
+ $X2=1.92 $Y2=1.515
r81 52 54 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=1.605 $Y=1.515
+ $X2=1.905 $Y2=1.515
r82 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.605
+ $Y=1.515 $X2=1.605 $Y2=1.515
r83 50 52 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.455 $Y=1.515
+ $X2=1.605 $Y2=1.515
r84 49 50 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.455 $Y2=1.515
r85 48 49 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.005 $Y=1.515
+ $X2=1.425 $Y2=1.515
r86 47 48 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.515
+ $X2=1.005 $Y2=1.515
r87 45 47 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.995 $Y2=1.515
r88 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r89 43 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.515
+ $X2=0.585 $Y2=1.515
r90 41 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.51 $Y2=1.515
r91 36 53 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.605 $Y2=1.565
r92 35 53 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.605 $Y2=1.565
r93 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r94 34 46 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r95 33 46 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r96 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.35
+ $X2=1.92 $Y2=1.515
r97 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.92 $Y=1.35
+ $X2=1.92 $Y2=0.74
r98 25 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=1.515
r99 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=2.4
r100 21 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.515
r101 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r102 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.515
r103 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r104 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r105 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r106 9 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=1.515
r107 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=2.4
r108 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.68
+ $X2=0.51 $Y2=1.515
r109 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.51 $Y=1.68 $X2=0.51
+ $Y2=2.4
r110 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r111 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 37 57
c89 31 0 1.67277e-19 $X=3.905 $Y=2.4
c90 19 0 8.60869e-20 $X=3.28 $Y=0.74
c91 3 0 7.59056e-20 $X=2.35 $Y=0.74
r92 55 57 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=3.8 $Y=1.515
+ $X2=3.905 $Y2=1.515
r93 55 56 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.8
+ $Y=1.515 $X2=3.8 $Y2=1.515
r94 53 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.71 $Y=1.515 $X2=3.8
+ $Y2=1.515
r95 52 53 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=3.405 $Y=1.515
+ $X2=3.71 $Y2=1.515
r96 51 52 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.28 $Y=1.515
+ $X2=3.405 $Y2=1.515
r97 50 51 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.905 $Y=1.515
+ $X2=3.28 $Y2=1.515
r98 49 50 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.78 $Y=1.515
+ $X2=2.905 $Y2=1.515
r99 47 49 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.44 $Y=1.515
+ $X2=2.78 $Y2=1.515
r100 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.44
+ $Y=1.515 $X2=2.44 $Y2=1.515
r101 45 47 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.405 $Y=1.515
+ $X2=2.44 $Y2=1.515
r102 43 45 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.35 $Y=1.515
+ $X2=2.405 $Y2=1.515
r103 37 56 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.8 $Y2=1.565
r104 36 56 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.8
+ $Y2=1.565
r105 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r106 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r107 34 48 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.44
+ $Y2=1.565
r108 33 48 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.44 $Y2=1.565
r109 29 57 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=1.68
+ $X2=3.905 $Y2=1.515
r110 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.905 $Y=1.68
+ $X2=3.905 $Y2=2.4
r111 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.515
r112 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=0.74
r113 21 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.68
+ $X2=3.405 $Y2=1.515
r114 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.405 $Y=1.68
+ $X2=3.405 $Y2=2.4
r115 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=1.35
+ $X2=3.28 $Y2=1.515
r116 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.28 $Y=1.35
+ $X2=3.28 $Y2=0.74
r117 13 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.68
+ $X2=2.905 $Y2=1.515
r118 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.905 $Y=1.68
+ $X2=2.905 $Y2=2.4
r119 9 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.35
+ $X2=2.78 $Y2=1.515
r120 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.78 $Y=1.35
+ $X2=2.78 $Y2=0.74
r121 5 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=1.515
r122 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=2.4
r123 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.35
+ $X2=2.35 $Y2=1.515
r124 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.35 $Y=1.35 $X2=2.35
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A1 3 7 11 15 19 23 27 31 33 34 35 51 53
r80 52 53 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.045 $Y=1.515
+ $X2=6.06 $Y2=1.515
r81 50 52 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=5.64 $Y=1.515
+ $X2=6.045 $Y2=1.515
r82 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.64
+ $Y=1.515 $X2=5.64 $Y2=1.515
r83 48 50 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.63 $Y=1.515 $X2=5.64
+ $Y2=1.515
r84 47 48 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.495 $Y=1.515
+ $X2=5.63 $Y2=1.515
r85 46 47 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=5.2 $Y=1.515
+ $X2=5.495 $Y2=1.515
r86 45 46 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.045 $Y=1.515
+ $X2=5.2 $Y2=1.515
r87 44 45 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=4.7 $Y=1.515
+ $X2=5.045 $Y2=1.515
r88 42 44 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.62 $Y=1.515 $X2=4.7
+ $Y2=1.515
r89 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.62
+ $Y=1.515 $X2=4.62 $Y2=1.515
r90 39 42 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=1.515
+ $X2=4.62 $Y2=1.515
r91 35 51 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.64 $Y2=1.565
r92 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r93 34 43 11.2564 $w=4.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.62 $Y2=1.565
r94 33 43 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=4.56 $Y=1.565 $X2=4.62
+ $Y2=1.565
r95 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.06 $Y=1.35
+ $X2=6.06 $Y2=1.515
r96 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.06 $Y=1.35
+ $X2=6.06 $Y2=0.74
r97 25 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.68
+ $X2=6.045 $Y2=1.515
r98 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.045 $Y=1.68
+ $X2=6.045 $Y2=2.4
r99 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.35
+ $X2=5.63 $Y2=1.515
r100 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.63 $Y=1.35
+ $X2=5.63 $Y2=0.74
r101 17 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.495 $Y=1.68
+ $X2=5.495 $Y2=1.515
r102 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.495 $Y=1.68
+ $X2=5.495 $Y2=2.4
r103 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.35
+ $X2=5.2 $Y2=1.515
r104 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.2 $Y=1.35 $X2=5.2
+ $Y2=0.74
r105 9 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.045 $Y=1.68
+ $X2=5.045 $Y2=1.515
r106 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.045 $Y=1.68
+ $X2=5.045 $Y2=2.4
r107 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.7 $Y=1.35 $X2=4.7
+ $Y2=1.515
r108 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.7 $Y=1.35 $X2=4.7
+ $Y2=0.74
r109 1 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.68
+ $X2=4.545 $Y2=1.515
r110 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.545 $Y=1.68
+ $X2=4.545 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A2 3 7 11 15 19 23 27 31 33 34 35 36 55
c88 55 0 1.89024e-19 $X=7.995 $Y=1.515
c89 36 0 9.24776e-20 $X=8.4 $Y=1.665
c90 31 0 3.04851e-19 $X=7.995 $Y=2.4
r91 53 55 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.92 $Y=1.515
+ $X2=7.995 $Y2=1.515
r92 51 53 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.785 $Y=1.515
+ $X2=7.92 $Y2=1.515
r93 50 51 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=7.495 $Y=1.515
+ $X2=7.785 $Y2=1.515
r94 49 50 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=7.355 $Y=1.515
+ $X2=7.495 $Y2=1.515
r95 48 49 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=7.045 $Y=1.515
+ $X2=7.355 $Y2=1.515
r96 47 48 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.92 $Y=1.515
+ $X2=7.045 $Y2=1.515
r97 45 47 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.9 $Y=1.515 $X2=6.92
+ $Y2=1.515
r98 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.9
+ $Y=1.515 $X2=6.9 $Y2=1.515
r99 43 45 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=6.505 $Y=1.515
+ $X2=6.9 $Y2=1.515
r100 41 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.49 $Y=1.515
+ $X2=6.505 $Y2=1.515
r101 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r102 35 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.92
+ $Y=1.515 $X2=7.92 $Y2=1.515
r103 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r104 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r105 33 46 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.565 $X2=6.9
+ $Y2=1.565
r106 29 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.68
+ $X2=7.995 $Y2=1.515
r107 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.995 $Y=1.68
+ $X2=7.995 $Y2=2.4
r108 25 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.785 $Y=1.35
+ $X2=7.785 $Y2=1.515
r109 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.785 $Y=1.35
+ $X2=7.785 $Y2=0.74
r110 21 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.495 $Y=1.68
+ $X2=7.495 $Y2=1.515
r111 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.495 $Y=1.68
+ $X2=7.495 $Y2=2.4
r112 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.355 $Y=1.35
+ $X2=7.355 $Y2=1.515
r113 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.355 $Y=1.35
+ $X2=7.355 $Y2=0.74
r114 13 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.045 $Y=1.68
+ $X2=7.045 $Y2=1.515
r115 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.045 $Y=1.68
+ $X2=7.045 $Y2=2.4
r116 9 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.92 $Y=1.35
+ $X2=6.92 $Y2=1.515
r117 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.92 $Y=1.35
+ $X2=6.92 $Y2=0.74
r118 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=1.68
+ $X2=6.505 $Y2=1.515
r119 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.505 $Y=1.68
+ $X2=6.505 $Y2=2.4
r120 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.49 $Y=1.35
+ $X2=6.49 $Y2=1.515
r121 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.49 $Y=1.35 $X2=6.49
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 53
c83 36 0 1.89024e-19 $X=10.32 $Y=1.665
c84 11 0 2.64775e-19 $X=8.995 $Y=2.4
r85 53 54 2.41806 $w=2.99e-07 $l=1.5e-08 $layer=POLY_cond $X=10.05 $Y=1.515
+ $X2=10.065 $Y2=1.515
r86 51 53 16.1204 $w=2.99e-07 $l=1e-07 $layer=POLY_cond $X=9.95 $Y=1.515
+ $X2=10.05 $Y2=1.515
r87 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.95
+ $Y=1.515 $X2=9.95 $Y2=1.515
r88 49 51 50.7793 $w=2.99e-07 $l=3.15e-07 $layer=POLY_cond $X=9.635 $Y=1.515
+ $X2=9.95 $Y2=1.515
r89 48 49 22.5686 $w=2.99e-07 $l=1.4e-07 $layer=POLY_cond $X=9.495 $Y=1.515
+ $X2=9.635 $Y2=1.515
r90 46 48 36.2709 $w=2.99e-07 $l=2.25e-07 $layer=POLY_cond $X=9.27 $Y=1.515
+ $X2=9.495 $Y2=1.515
r91 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.27
+ $Y=1.515 $X2=9.27 $Y2=1.515
r92 44 46 10.4783 $w=2.99e-07 $l=6.5e-08 $layer=POLY_cond $X=9.205 $Y=1.515
+ $X2=9.27 $Y2=1.515
r93 43 44 33.8528 $w=2.99e-07 $l=2.1e-07 $layer=POLY_cond $X=8.995 $Y=1.515
+ $X2=9.205 $Y2=1.515
r94 42 43 35.4649 $w=2.99e-07 $l=2.2e-07 $layer=POLY_cond $X=8.775 $Y=1.515
+ $X2=8.995 $Y2=1.515
r95 36 52 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=9.95 $Y2=1.565
r96 35 52 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.95 $Y2=1.565
r97 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r98 34 47 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.27
+ $Y2=1.565
r99 33 47 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.27 $Y2=1.565
r100 29 54 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=1.515
r101 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=0.74
r102 25 53 14.6425 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.05 $Y=1.68
+ $X2=10.05 $Y2=1.515
r103 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.05 $Y=1.68
+ $X2=10.05 $Y2=2.4
r104 21 49 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.635 $Y=1.35
+ $X2=9.635 $Y2=1.515
r105 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.635 $Y=1.35
+ $X2=9.635 $Y2=0.74
r106 17 48 14.6425 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.495 $Y=1.68
+ $X2=9.495 $Y2=1.515
r107 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.495 $Y=1.68
+ $X2=9.495 $Y2=2.4
r108 13 44 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.205 $Y=1.35
+ $X2=9.205 $Y2=1.515
r109 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.205 $Y=1.35
+ $X2=9.205 $Y2=0.74
r110 9 43 14.6425 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.995 $Y=1.68
+ $X2=8.995 $Y2=1.515
r111 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.995 $Y=1.68
+ $X2=8.995 $Y2=2.4
r112 5 42 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.775 $Y=1.35
+ $X2=8.775 $Y2=1.515
r113 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.775 $Y=1.35
+ $X2=8.775 $Y2=0.74
r114 1 42 45.1371 $w=2.99e-07 $l=3.52987e-07 $layer=POLY_cond $X=8.495 $Y=1.68
+ $X2=8.775 $Y2=1.515
r115 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.495 $Y=1.68
+ $X2=8.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A_27_368# 1 2 3 4 5 6 7 8 9 10 11 36 40 41
+ 44 46 50 52 56 58 60 61 62 66 70 72 73 76 78 82 84 88 90 92 94 96 97 98 102
+ 104 107 109 111
c168 88 0 1.72297e-19 $X=9.27 $Y=2.815
c169 82 0 1.72297e-19 $X=8.27 $Y=2.815
c170 76 0 1.32554e-19 $X=7.27 $Y=2.815
r171 92 113 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=2.12
+ $X2=10.275 $Y2=2.035
r172 92 94 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=10.275 $Y=2.12
+ $X2=10.275 $Y2=2.815
r173 91 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=2.035
+ $X2=9.27 $Y2=2.035
r174 90 113 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.11 $Y=2.035
+ $X2=10.275 $Y2=2.035
r175 90 91 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=10.11 $Y=2.035
+ $X2=9.435 $Y2=2.035
r176 86 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.27 $Y=2.12
+ $X2=9.27 $Y2=2.035
r177 86 88 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.27 $Y=2.12
+ $X2=9.27 $Y2=2.815
r178 85 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.435 $Y=2.035
+ $X2=8.27 $Y2=2.035
r179 84 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=2.035
+ $X2=9.27 $Y2=2.035
r180 84 85 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.105 $Y=2.035
+ $X2=8.435 $Y2=2.035
r181 80 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=2.12
+ $X2=8.27 $Y2=2.035
r182 80 82 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.27 $Y=2.12
+ $X2=8.27 $Y2=2.815
r183 79 106 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=2.035
+ $X2=7.27 $Y2=2.035
r184 78 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=2.035
+ $X2=8.27 $Y2=2.035
r185 78 79 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.105 $Y=2.035
+ $X2=7.435 $Y2=2.035
r186 74 107 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=2.46
+ $X2=7.27 $Y2=2.375
r187 74 76 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.27 $Y=2.46
+ $X2=7.27 $Y2=2.815
r188 73 107 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=2.29
+ $X2=7.27 $Y2=2.375
r189 72 106 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.27 $Y=2.12
+ $X2=7.27 $Y2=2.035
r190 72 73 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.27 $Y=2.12
+ $X2=7.27 $Y2=2.29
r191 71 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=2.375
+ $X2=6.27 $Y2=2.375
r192 70 107 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=2.375
+ $X2=7.27 $Y2=2.375
r193 70 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.105 $Y=2.375
+ $X2=6.435 $Y2=2.375
r194 67 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=2.375
+ $X2=5.27 $Y2=2.375
r195 66 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=2.375
+ $X2=6.27 $Y2=2.375
r196 66 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.105 $Y=2.375
+ $X2=5.435 $Y2=2.375
r197 63 100 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=2.375
+ $X2=4.18 $Y2=2.375
r198 62 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=2.375
+ $X2=5.27 $Y2=2.375
r199 62 63 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.105 $Y=2.375
+ $X2=4.345 $Y2=2.375
r200 60 100 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=2.46
+ $X2=4.18 $Y2=2.375
r201 60 61 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.18 $Y=2.46
+ $X2=4.18 $Y2=2.905
r202 59 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=3.18 $Y2=2.99
r203 58 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=4.18 $Y2=2.905
r204 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=3.345 $Y2=2.99
r205 54 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=2.905
+ $X2=3.18 $Y2=2.99
r206 54 56 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.18 $Y=2.905
+ $X2=3.18 $Y2=2.455
r207 53 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.99
+ $X2=2.18 $Y2=2.99
r208 52 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.99
+ $X2=3.18 $Y2=2.99
r209 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.015 $Y=2.99
+ $X2=2.345 $Y2=2.99
r210 48 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.905
+ $X2=2.18 $Y2=2.99
r211 48 50 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.18 $Y=2.905
+ $X2=2.18 $Y2=2.455
r212 47 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.99
+ $X2=1.23 $Y2=2.99
r213 46 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=2.18 $Y2=2.99
r214 46 47 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=1.315 $Y2=2.99
r215 42 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.99
r216 42 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.23 $Y=2.905
+ $X2=1.23 $Y2=2.455
r217 40 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.23 $Y2=2.99
r218 40 41 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.445 $Y2=2.99
r219 36 39 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r220 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r221 34 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r222 11 113 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.84 $X2=10.275 $Y2=2.115
r223 11 94 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.84 $X2=10.275 $Y2=2.815
r224 10 111 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=9.085
+ $Y=1.84 $X2=9.27 $Y2=2.115
r225 10 88 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=9.085
+ $Y=1.84 $X2=9.27 $Y2=2.815
r226 9 109 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.84 $X2=8.27 $Y2=2.115
r227 9 82 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.84 $X2=8.27 $Y2=2.815
r228 8 106 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.135
+ $Y=1.84 $X2=7.27 $Y2=2.115
r229 8 76 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.135
+ $Y=1.84 $X2=7.27 $Y2=2.815
r230 7 104 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.135
+ $Y=1.84 $X2=6.27 $Y2=2.455
r231 6 102 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.135
+ $Y=1.84 $X2=5.27 $Y2=2.455
r232 5 100 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=3.995
+ $Y=1.84 $X2=4.18 $Y2=2.455
r233 4 56 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.84 $X2=3.18 $Y2=2.455
r234 3 50 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.84 $X2=2.18 $Y2=2.455
r235 2 44 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.455
r236 1 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r237 1 36 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%Y 1 2 3 4 5 6 7 8 27 31 35 39 45 48 50 52 54
+ 59 60 62 63 64 65 66 79 81
c121 54 0 8.12065e-20 $X=2.565 $Y=0.86
c122 35 0 7.59056e-20 $X=3.51 $Y=1.03
r123 66 74 4.96191 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=6 $Y=0.95
+ $X2=5.845 $Y2=0.95
r124 65 74 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=0.95
+ $X2=5.845 $Y2=0.95
r125 65 81 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=0.95
+ $X2=5.15 $Y2=0.95
r126 64 81 4.83878 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=0.975
+ $X2=5.15 $Y2=0.975
r127 64 79 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=0.975
+ $X2=4.82 $Y2=0.975
r128 63 66 5.76222 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=6.18 $Y=0.95 $X2=6
+ $Y2=0.95
r129 60 79 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.66 $Y=1.095
+ $X2=4.82 $Y2=1.095
r130 54 56 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.565 $Y=0.86
+ $X2=2.565 $Y2=1.03
r131 47 63 8.02311 $w=3.6e-07 $l=2.18403e-07 $layer=LI1_cond $X=6.265 $Y=1.13
+ $X2=6.18 $Y2=0.95
r132 47 48 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.265 $Y=1.13
+ $X2=6.265 $Y2=1.95
r133 46 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=2.035
+ $X2=3.68 $Y2=2.035
r134 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.18 $Y=2.035
+ $X2=6.265 $Y2=1.95
r135 45 46 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=6.18 $Y=2.035
+ $X2=3.845 $Y2=2.035
r136 40 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=2.035
+ $X2=2.68 $Y2=2.035
r137 39 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=2.035
+ $X2=3.68 $Y2=2.035
r138 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.515 $Y=2.035
+ $X2=2.845 $Y2=2.035
r139 36 56 1.29116 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=1.03
+ $X2=2.565 $Y2=1.03
r140 36 38 29.3873 $w=2.98e-07 $l=7.65e-07 $layer=LI1_cond $X=2.73 $Y=1.03
+ $X2=3.495 $Y2=1.03
r141 35 60 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.51 $Y=1.03
+ $X2=3.66 $Y2=1.03
r142 35 38 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.51 $Y=1.03
+ $X2=3.495 $Y2=1.03
r143 32 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.035
+ $X2=1.68 $Y2=2.035
r144 31 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=2.68 $Y2=2.035
r145 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=1.845 $Y2=2.035
r146 28 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r147 27 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=1.68 $Y2=2.035
r148 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.515 $Y=2.035
+ $X2=0.945 $Y2=2.035
r149 8 62 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=3.495
+ $Y=1.84 $X2=3.68 $Y2=2.115
r150 7 59 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=2.68 $Y2=2.115
r151 6 52 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.115
r152 5 50 300 $w=1.7e-07 $l=3.5373e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.84 $X2=0.78 $Y2=2.115
r153 4 74 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.37 $X2=5.845 $Y2=0.95
r154 3 64 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.37 $X2=4.985 $Y2=0.95
r155 2 38 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.37 $X2=3.495 $Y2=0.965
r156 1 54 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.37 $X2=2.565 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 53 54 56 57 58 79 85 86 89
c130 21 0 1.67277e-19 $X=4.77 $Y=2.805
r131 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r132 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r133 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r134 83 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.935 $Y=3.33
+ $X2=9.77 $Y2=3.33
r135 83 85 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.935 $Y=3.33
+ $X2=10.32 $Y2=3.33
r136 82 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r137 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 79 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.77 $Y2=3.33
r139 79 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.36 $Y2=3.33
r140 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r142 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r143 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r144 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r146 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r147 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r148 65 66 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r149 62 66 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r150 61 65 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 61 62 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r152 58 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r153 58 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 56 77 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.605 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=3.33
+ $X2=8.77 $Y2=3.33
r156 55 81 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.935 $Y=3.33
+ $X2=9.36 $Y2=3.33
r157 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=3.33
+ $X2=8.77 $Y2=3.33
r158 53 74 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.44 $Y2=3.33
r159 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=3.33
+ $X2=7.77 $Y2=3.33
r160 52 77 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.935 $Y=3.33
+ $X2=8.4 $Y2=3.33
r161 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.935 $Y=3.33
+ $X2=7.77 $Y2=3.33
r162 50 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.605 $Y=3.33
+ $X2=6.48 $Y2=3.33
r163 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=3.33
+ $X2=6.77 $Y2=3.33
r164 49 74 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.935 $Y=3.33
+ $X2=7.44 $Y2=3.33
r165 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.935 $Y=3.33
+ $X2=6.77 $Y2=3.33
r166 47 68 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.77 $Y2=3.33
r168 46 71 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.935 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=3.33
+ $X2=5.77 $Y2=3.33
r170 44 65 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.77 $Y2=3.33
r172 43 68 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=5.52 $Y2=3.33
r173 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=4.77 $Y2=3.33
r174 39 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.77 $Y=3.245
+ $X2=9.77 $Y2=3.33
r175 39 41 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=9.77 $Y=3.245
+ $X2=9.77 $Y2=2.455
r176 35 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.77 $Y=3.245
+ $X2=8.77 $Y2=3.33
r177 35 37 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=8.77 $Y=3.245
+ $X2=8.77 $Y2=2.455
r178 31 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=3.33
r179 31 33 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=2.455
r180 27 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.77 $Y=3.245
+ $X2=6.77 $Y2=3.33
r181 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=6.77 $Y=3.245
+ $X2=6.77 $Y2=2.805
r182 23 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=3.245
+ $X2=5.77 $Y2=3.33
r183 23 25 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=5.77 $Y=3.245
+ $X2=5.77 $Y2=2.805
r184 19 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=3.33
r185 19 21 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=2.805
r186 6 41 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=9.585
+ $Y=1.84 $X2=9.77 $Y2=2.455
r187 5 37 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=8.585
+ $Y=1.84 $X2=8.77 $Y2=2.455
r188 4 33 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=7.585
+ $Y=1.84 $X2=7.77 $Y2=2.455
r189 3 29 600 $w=1.7e-07 $l=1.04886e-06 $layer=licon1_PDIFF $count=1 $X=6.595
+ $Y=1.84 $X2=6.77 $Y2=2.805
r190 2 25 600 $w=1.7e-07 $l=1.05345e-06 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.84 $X2=5.77 $Y2=2.805
r191 1 21 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=4.635
+ $Y=1.84 $X2=4.77 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 32 33 34
+ 36 37 42
c74 32 0 8.60869e-20 $X=2.9 $Y=0.34
r75 42 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.925 $Y=0.34
+ $X2=3.925 $Y2=0.53
r76 37 40 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.065 $Y=0.34
+ $X2=3.065 $Y2=0.53
r77 35 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=0.34
+ $X2=3.065 $Y2=0.34
r78 34 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0.34
+ $X2=3.925 $Y2=0.34
r79 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.76 $Y=0.34
+ $X2=3.23 $Y2=0.34
r80 32 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=0.34
+ $X2=3.065 $Y2=0.34
r81 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.9 $Y=0.34 $X2=2.22
+ $Y2=0.34
r82 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.135 $Y=1.01
+ $X2=2.135 $Y2=0.515
r83 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=0.425
+ $X2=2.22 $Y2=0.34
r84 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.135 $Y=0.425
+ $X2=2.135 $Y2=0.515
r85 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=1.095
+ $X2=1.21 $Y2=1.095
r86 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=1.095
+ $X2=2.135 $Y2=1.01
r87 26 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.05 $Y=1.095
+ $X2=1.295 $Y2=1.095
r88 22 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=1.01 $X2=1.21
+ $Y2=1.095
r89 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.21 $Y=1.01
+ $X2=1.21 $Y2=0.515
r90 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=1.21 $Y2=1.095
r91 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.095
+ $X2=0.445 $Y2=1.095
r92 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r93 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r94 5 45 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.37 $X2=3.925 $Y2=0.53
r95 4 40 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.37 $X2=3.065 $Y2=0.53
r96 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.995
+ $Y=0.37 $X2=2.135 $Y2=0.515
r97 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r98 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 53 58 64 67 70 73 77
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r113 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r114 70 71 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r115 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r118 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r119 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r120 59 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.585 $Y=0 $X2=9.42
+ $Y2=0
r121 59 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.585 $Y=0
+ $X2=9.84 $Y2=0
r122 58 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.337 $Y2=0
r123 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r124 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r125 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r126 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r127 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=0 $X2=8.56
+ $Y2=0
r128 54 56 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.725 $Y=0
+ $X2=8.88 $Y2=0
r129 53 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=0 $X2=9.42
+ $Y2=0
r130 53 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.255 $Y=0
+ $X2=8.88 $Y2=0
r131 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r132 51 52 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r133 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.64
+ $Y2=0
r134 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=2.16 $Y2=0
r135 48 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.395 $Y=0 $X2=8.56
+ $Y2=0
r136 48 51 406.775 $w=1.68e-07 $l=6.235e-06 $layer=LI1_cond $X=8.395 $Y=0
+ $X2=2.16 $Y2=0
r137 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r138 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r139 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r140 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r141 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r142 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.64
+ $Y2=0
r143 43 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r144 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r146 38 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r147 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r148 36 71 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=8.4
+ $Y2=0
r149 36 52 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=2.16 $Y2=0
r150 32 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.337 $Y2=0
r151 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.515
r152 28 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.42 $Y=0.085
+ $X2=9.42 $Y2=0
r153 28 30 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=9.42 $Y=0.085
+ $X2=9.42 $Y2=0.595
r154 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=0.085
+ $X2=8.56 $Y2=0
r155 24 26 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.56 $Y=0.085
+ $X2=8.56 $Y2=0.595
r156 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0
r157 20 22 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0.595
r158 16 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r159 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.595
r160 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.14
+ $Y=0.37 $X2=10.28 $Y2=0.515
r161 4 30 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=9.28
+ $Y=0.37 $X2=9.42 $Y2=0.595
r162 3 26 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=8.415
+ $Y=0.37 $X2=8.56 $Y2=0.595
r163 2 22 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.595
r164 1 18 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A_868_74# 1 2 3 4 5 24 30 31
r40 30 31 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8 $Y=0.515
+ $X2=7.835 $Y2=0.515
r41 24 27 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.485 $Y=0.475
+ $X2=4.485 $Y2=0.595
r42 23 31 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=7.135 $Y=0.475
+ $X2=7.835 $Y2=0.475
r43 21 23 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=6.275 $Y=0.475
+ $X2=7.135 $Y2=0.475
r44 19 21 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=5.415 $Y=0.475
+ $X2=6.275 $Y2=0.475
r45 17 24 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=0.475
+ $X2=4.485 $Y2=0.475
r46 17 19 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=4.65 $Y=0.475
+ $X2=5.415 $Y2=0.475
r47 5 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.86
+ $Y=0.37 $X2=8 $Y2=0.515
r48 4 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.995
+ $Y=0.37 $X2=7.135 $Y2=0.515
r49 3 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.135
+ $Y=0.37 $X2=6.275 $Y2=0.515
r50 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.275
+ $Y=0.37 $X2=5.415 $Y2=0.515
r51 1 27 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.37 $X2=4.485 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_4%A_1313_74# 1 2 3 4 15 19 21 25 30 32 33 34
r57 32 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=1.015
+ $X2=7.735 $Y2=1.015
r58 30 32 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=6.87 $Y=1.015 $X2=7.57
+ $Y2=1.015
r59 28 30 5.11015 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.705 $Y=0.975
+ $X2=6.87 $Y2=0.975
r60 23 25 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.85 $Y=1.01
+ $X2=9.85 $Y2=0.515
r61 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=1.095
+ $X2=8.99 $Y2=1.095
r62 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.765 $Y=1.095
+ $X2=9.85 $Y2=1.01
r63 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.765 $Y=1.095
+ $X2=9.075 $Y2=1.095
r64 17 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.99 $Y=1.01 $X2=8.99
+ $Y2=1.095
r65 17 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.99 $Y=1.01
+ $X2=8.99 $Y2=0.515
r66 15 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=1.095
+ $X2=8.99 $Y2=1.095
r67 15 33 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=8.905 $Y=1.095
+ $X2=7.735 $Y2=1.095
r68 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.71
+ $Y=0.37 $X2=9.85 $Y2=0.515
r69 3 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.85
+ $Y=0.37 $X2=8.99 $Y2=0.515
r70 2 32 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.43
+ $Y=0.37 $X2=7.57 $Y2=0.95
r71 1 28 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.37 $X2=6.705 $Y2=0.95
.ends


* File: sky130_fd_sc_ms__xnor2_2.pxi.spice
* Created: Wed Sep  2 12:33:24 2020
* 
x_PM_SKY130_FD_SC_MS__XNOR2_2%A N_A_M1011_g N_A_M1014_g N_A_M1002_g N_A_M1006_g
+ N_A_M1008_g N_A_M1007_g N_A_c_98_n N_A_c_114_n N_A_c_115_n A N_A_c_100_n
+ N_A_c_101_n N_A_c_102_n N_A_c_103_n N_A_c_104_n N_A_c_105_n N_A_c_106_n
+ N_A_c_107_n N_A_c_108_n N_A_c_109_n PM_SKY130_FD_SC_MS__XNOR2_2%A
x_PM_SKY130_FD_SC_MS__XNOR2_2%B N_B_M1013_g N_B_M1012_g N_B_c_246_n N_B_M1001_g
+ N_B_M1000_g N_B_c_248_n N_B_M1005_g N_B_M1003_g N_B_c_250_n N_B_c_251_n
+ N_B_c_252_n N_B_c_264_n N_B_c_265_n N_B_c_289_n N_B_c_266_n N_B_c_344_p
+ N_B_c_253_n N_B_c_254_n N_B_c_255_n B N_B_c_257_n
+ PM_SKY130_FD_SC_MS__XNOR2_2%B
x_PM_SKY130_FD_SC_MS__XNOR2_2%A_136_368# N_A_136_368#_M1013_d
+ N_A_136_368#_M1011_d N_A_136_368#_M1009_g N_A_136_368#_c_402_n
+ N_A_136_368#_M1004_g N_A_136_368#_M1010_g N_A_136_368#_c_404_n
+ N_A_136_368#_M1015_g N_A_136_368#_c_412_n N_A_136_368#_c_405_n
+ N_A_136_368#_c_406_n N_A_136_368#_c_407_n N_A_136_368#_c_408_n
+ N_A_136_368#_c_409_n PM_SKY130_FD_SC_MS__XNOR2_2%A_136_368#
x_PM_SKY130_FD_SC_MS__XNOR2_2%VPWR N_VPWR_M1011_s N_VPWR_M1012_d N_VPWR_M1010_s
+ N_VPWR_M1008_d N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ N_VPWR_c_506_n N_VPWR_c_507_n VPWR N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_501_n PM_SKY130_FD_SC_MS__XNOR2_2%VPWR
x_PM_SKY130_FD_SC_MS__XNOR2_2%Y N_Y_M1004_d N_Y_M1009_d N_Y_M1000_d N_Y_c_568_n
+ N_Y_c_569_n N_Y_c_570_n N_Y_c_587_n N_Y_c_575_n N_Y_c_588_n N_Y_c_571_n
+ N_Y_c_590_n N_Y_c_572_n N_Y_c_573_n N_Y_c_591_n Y Y N_Y_c_592_n
+ PM_SKY130_FD_SC_MS__XNOR2_2%Y
x_PM_SKY130_FD_SC_MS__XNOR2_2%A_641_368# N_A_641_368#_M1002_s
+ N_A_641_368#_M1003_s N_A_641_368#_c_670_n N_A_641_368#_c_677_n
+ N_A_641_368#_c_671_n PM_SKY130_FD_SC_MS__XNOR2_2%A_641_368#
x_PM_SKY130_FD_SC_MS__XNOR2_2%VGND N_VGND_M1014_s N_VGND_M1006_d N_VGND_M1005_s
+ N_VGND_c_697_n N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n
+ N_VGND_c_702_n VGND N_VGND_c_703_n N_VGND_c_704_n N_VGND_c_705_n
+ N_VGND_c_706_n PM_SKY130_FD_SC_MS__XNOR2_2%VGND
x_PM_SKY130_FD_SC_MS__XNOR2_2%A_340_107# N_A_340_107#_M1004_s
+ N_A_340_107#_M1015_s N_A_340_107#_M1001_d N_A_340_107#_M1007_s
+ N_A_340_107#_c_765_n N_A_340_107#_c_766_n N_A_340_107#_c_762_n
+ N_A_340_107#_c_763_n N_A_340_107#_c_772_n N_A_340_107#_c_776_n
+ N_A_340_107#_c_764_n PM_SKY130_FD_SC_MS__XNOR2_2%A_340_107#
cc_1 VNB N_A_M1011_g 0.00690535f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.34
cc_2 VNB N_A_M1002_g 0.00685807f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=2.4
cc_3 VNB N_A_M1007_g 0.031366f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.74
cc_4 VNB N_A_c_98_n 0.00126095f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_5 VNB A 0.00491569f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_6 VNB N_A_c_100_n 0.0212635f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.295
cc_7 VNB N_A_c_101_n 0.00284076f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.295
cc_8 VNB N_A_c_102_n 0.00311998f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_9 VNB N_A_c_103_n 0.00526995f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_10 VNB N_A_c_104_n 0.0358441f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_11 VNB N_A_c_105_n 0.00770753f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_12 VNB N_A_c_106_n 0.017864f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.22
cc_13 VNB N_A_c_107_n 0.0327682f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.385
cc_14 VNB N_A_c_108_n 0.0186645f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.22
cc_15 VNB N_A_c_109_n 0.0276459f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=1.515
cc_16 VNB N_B_M1013_g 0.0267022f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.34
cc_17 VNB N_B_c_246_n 0.0190023f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=2.4
cc_18 VNB N_B_M1000_g 0.00663087f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=0.74
cc_19 VNB N_B_c_248_n 0.0181813f $X=-0.19 $Y=-0.245 $X2=4.695 $Y2=2.4
cc_20 VNB N_B_M1003_g 0.00101917f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.74
cc_21 VNB N_B_c_250_n 0.0126261f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_22 VNB N_B_c_251_n 0.00111425f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_23 VNB N_B_c_252_n 0.0372654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_253_n 0.0198025f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_25 VNB N_B_c_254_n 7.72606e-19 $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_26 VNB N_B_c_255_n 0.0227111f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_27 VNB B 0.00119299f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_28 VNB N_B_c_257_n 0.0467984f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=1.515
cc_29 VNB N_A_136_368#_M1009_g 0.00602318f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=2.4
cc_30 VNB N_A_136_368#_c_402_n 0.0206891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_136_368#_M1010_g 0.00662457f $X=-0.19 $Y=-0.245 $X2=4.695 $Y2=2.4
cc_32 VNB N_A_136_368#_c_404_n 0.0190849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_136_368#_c_405_n 0.00311207f $X=-0.19 $Y=-0.245 $X2=3.355
+ $Y2=1.805
cc_34 VNB N_A_136_368#_c_406_n 0.00644617f $X=-0.19 $Y=-0.245 $X2=0.865
+ $Y2=1.295
cc_35 VNB N_A_136_368#_c_407_n 0.0075666f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_36 VNB N_A_136_368#_c_408_n 0.00974138f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_37 VNB N_A_136_368#_c_409_n 0.0577931f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.22
cc_38 VNB N_VPWR_c_501_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_568_n 0.0311889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_569_n 0.00487916f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.22
cc_41 VNB N_Y_c_570_n 0.00986386f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=0.74
cc_42 VNB N_Y_c_571_n 5.82374e-19 $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=1.35
cc_43 VNB N_Y_c_572_n 0.00409335f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.55
cc_44 VNB N_Y_c_573_n 0.0148451f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_45 VNB N_VGND_c_697_n 0.0131748f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=2.4
cc_46 VNB N_VGND_c_698_n 0.0273582f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.22
cc_47 VNB N_VGND_c_699_n 0.00800128f $X=-0.19 $Y=-0.245 $X2=4.695 $Y2=2.4
cc_48 VNB N_VGND_c_700_n 0.00812389f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.74
cc_49 VNB N_VGND_c_701_n 0.0656586f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.55
cc_50 VNB N_VGND_c_702_n 0.0064126f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_51 VNB N_VGND_c_703_n 0.0190098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_704_n 0.0193317f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_53 VNB N_VGND_c_705_n 0.291439f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_54 VNB N_VGND_c_706_n 0.0066048f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.55
cc_55 VNB N_A_340_107#_c_762_n 0.00274459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_340_107#_c_763_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_57 VNB N_A_340_107#_c_764_n 0.0136683f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_58 VPB N_A_M1011_g 0.0242784f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.34
cc_59 VPB N_A_M1002_g 0.025329f $X=-0.19 $Y=1.66 $X2=3.115 $Y2=2.4
cc_60 VPB N_A_M1008_g 0.0226149f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=2.4
cc_61 VPB N_A_c_98_n 6.82535e-19 $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.72
cc_62 VPB N_A_c_114_n 0.0175175f $X=-0.19 $Y=1.66 $X2=4.445 $Y2=1.805
cc_63 VPB N_A_c_115_n 9.52429e-19 $X=-0.19 $Y=1.66 $X2=3.355 $Y2=1.805
cc_64 VPB A 0.00150831f $X=-0.19 $Y=1.66 $X2=4.475 $Y2=1.58
cc_65 VPB N_A_c_109_n 0.00586232f $X=-0.19 $Y=1.66 $X2=4.69 $Y2=1.515
cc_66 VPB N_B_M1012_g 0.0228871f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_67 VPB N_B_M1000_g 0.0224945f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=0.74
cc_68 VPB N_B_M1003_g 0.0211869f $X=-0.19 $Y=1.66 $X2=4.785 $Y2=0.74
cc_69 VPB N_B_c_250_n 8.0996e-19 $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.72
cc_70 VPB N_B_c_251_n 6.80183e-19 $X=-0.19 $Y=1.66 $X2=4.475 $Y2=1.58
cc_71 VPB N_B_c_252_n 0.0165375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_B_c_264_n 0.00699785f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.295
cc_73 VPB N_B_c_265_n 7.3043e-19 $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.295
cc_74 VPB N_B_c_266_n 0.0100484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_B_c_255_n 0.0168007f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_76 VPB N_A_136_368#_M1009_g 0.0243047f $X=-0.19 $Y=1.66 $X2=3.115 $Y2=2.4
cc_77 VPB N_A_136_368#_M1010_g 0.0234569f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=2.4
cc_78 VPB N_A_136_368#_c_412_n 0.00404678f $X=-0.19 $Y=1.66 $X2=4.785 $Y2=0.74
cc_79 VPB N_VPWR_c_502_n 0.0121909f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=0.74
cc_80 VPB N_VPWR_c_503_n 0.0293007f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=1.68
cc_81 VPB N_VPWR_c_504_n 0.020562f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=2.4
cc_82 VPB N_VPWR_c_505_n 0.00861433f $X=-0.19 $Y=1.66 $X2=4.785 $Y2=0.74
cc_83 VPB N_VPWR_c_506_n 0.0131441f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.55
cc_84 VPB N_VPWR_c_507_n 0.0342994f $X=-0.19 $Y=1.66 $X2=4.445 $Y2=1.805
cc_85 VPB N_VPWR_c_508_n 0.0249485f $X=-0.19 $Y=1.66 $X2=2.975 $Y2=1.295
cc_86 VPB N_VPWR_c_509_n 0.0439986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_510_n 0.0303963f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.22
cc_88 VPB N_VPWR_c_511_n 0.00632133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_501_n 0.0696905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_Y_c_568_n 0.0263982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_Y_c_575_n 0.00801979f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=1.68
cc_92 VPB Y 0.00231613f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.295
cc_93 VPB N_A_641_368#_c_670_n 0.00487134f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_94 VPB N_A_641_368#_c_671_n 0.00370087f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=0.74
cc_95 N_A_c_100_n N_B_M1013_g 0.00113884f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_96 N_A_c_101_n N_B_M1013_g 6.92697e-19 $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_97 N_A_c_105_n N_B_M1013_g 0.00207268f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A_c_106_n N_B_M1013_g 0.0342458f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_99 N_A_c_103_n N_B_c_246_n 3.87669e-19 $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_100 N_A_c_108_n N_B_c_246_n 0.0238678f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A_M1002_g N_B_M1000_g 0.0386952f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_c_98_n N_B_M1000_g 0.00365154f $X=3.19 $Y=1.72 $X2=0 $Y2=0
cc_103 N_A_c_114_n N_B_M1000_g 0.0179849f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_104 N_A_M1007_g N_B_c_248_n 0.0266017f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_M1008_g N_B_M1003_g 0.0299197f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_c_114_n N_B_M1003_g 0.0120373f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_107 N_A_M1011_g N_B_c_250_n 0.0453172f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_108 N_A_c_100_n N_B_c_250_n 2.10602e-19 $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_109 N_A_c_101_n N_B_c_250_n 7.45074e-19 $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_110 N_A_c_104_n N_B_c_250_n 0.0342458f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_c_100_n N_B_c_251_n 0.0190018f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_112 N_A_c_100_n N_B_c_252_n 0.0113639f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_113 N_A_M1002_g N_B_c_264_n 8.12181e-19 $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_c_115_n N_B_c_264_n 0.0112446f $X=3.355 $Y=1.805 $X2=0 $Y2=0
cc_115 N_A_c_100_n N_B_c_264_n 0.0164056f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_116 N_A_M1002_g N_B_c_289_n 0.00342789f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_M1002_g N_B_c_266_n 0.013108f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_M1008_g N_B_c_266_n 0.0190348f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_c_114_n N_B_c_266_n 0.0607902f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_120 N_A_c_115_n N_B_c_266_n 0.0213544f $X=3.355 $Y=1.805 $X2=0 $Y2=0
cc_121 A N_B_c_266_n 0.0192216f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A_c_107_n N_B_c_266_n 4.40757e-19 $X=3.19 $Y=1.385 $X2=0 $Y2=0
cc_123 N_A_c_109_n N_B_c_266_n 6.63683e-19 $X=4.69 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_M1007_g N_B_c_253_n 0.01286f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_c_114_n N_B_c_253_n 0.00627445f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_126 A N_B_c_253_n 0.0314518f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A_c_109_n N_B_c_253_n 0.00129427f $X=4.69 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_M1008_g N_B_c_255_n 0.00967964f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_M1007_g N_B_c_255_n 0.0132787f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_130 A N_B_c_255_n 0.0348497f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A_M1007_g B 9.31443e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_c_114_n B 0.0251802f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_133 A B 0.0148825f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A_c_103_n B 0.0105933f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_135 N_A_c_107_n B 8.71298e-19 $X=3.19 $Y=1.385 $X2=0 $Y2=0
cc_136 N_A_c_109_n B 2.21532e-19 $X=4.69 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A_c_114_n N_B_c_257_n 6.27403e-19 $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_138 A N_B_c_257_n 0.00553545f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_c_103_n N_B_c_257_n 0.00162562f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_140 N_A_c_107_n N_B_c_257_n 0.0145025f $X=3.19 $Y=1.385 $X2=0 $Y2=0
cc_141 N_A_c_109_n N_B_c_257_n 0.0160078f $X=4.69 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_A_136_368#_M1010_g 0.0203132f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_c_98_n N_A_136_368#_M1010_g 9.63074e-19 $X=3.19 $Y=1.72 $X2=0 $Y2=0
cc_144 N_A_c_102_n N_A_136_368#_c_404_n 6.76195e-19 $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_145 N_A_c_103_n N_A_136_368#_c_404_n 0.00119559f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_146 N_A_c_108_n N_A_136_368#_c_404_n 0.0132146f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_147 N_A_M1011_g N_A_136_368#_c_412_n 0.00691986f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_148 N_A_c_100_n N_A_136_368#_c_412_n 0.00506714f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_149 N_A_c_101_n N_A_136_368#_c_412_n 0.00227899f $X=0.865 $Y=1.295 $X2=0
+ $Y2=0
cc_150 N_A_c_104_n N_A_136_368#_c_412_n 0.00186935f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_151 N_A_c_105_n N_A_136_368#_c_412_n 0.00943479f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A_M1011_g N_A_136_368#_c_405_n 0.00165132f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_153 N_A_c_100_n N_A_136_368#_c_405_n 0.0262593f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_154 N_A_c_101_n N_A_136_368#_c_405_n 0.0026151f $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_155 N_A_c_105_n N_A_136_368#_c_405_n 0.0261005f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A_c_106_n N_A_136_368#_c_405_n 4.6081e-19 $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A_c_100_n N_A_136_368#_c_406_n 0.0130897f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_158 N_A_c_106_n N_A_136_368#_c_406_n 0.00147911f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A_c_100_n N_A_136_368#_c_407_n 0.0361112f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_160 N_A_c_102_n N_A_136_368#_c_407_n 0.00234524f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_161 N_A_c_103_n N_A_136_368#_c_407_n 0.0119148f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_162 N_A_c_107_n N_A_136_368#_c_407_n 4.75044e-19 $X=3.19 $Y=1.385 $X2=0 $Y2=0
cc_163 N_A_c_100_n N_A_136_368#_c_408_n 0.0150674f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_164 N_A_c_100_n N_A_136_368#_c_409_n 0.0077648f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_165 N_A_c_103_n N_A_136_368#_c_409_n 7.12902e-19 $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_166 N_A_c_107_n N_A_136_368#_c_409_n 0.0288976f $X=3.19 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A_M1011_g N_VPWR_c_503_n 0.00914406f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_168 N_A_M1002_g N_VPWR_c_505_n 0.00316613f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_M1008_g N_VPWR_c_507_n 0.00341401f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A_M1011_g N_VPWR_c_508_n 0.0059286f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_171 N_A_M1002_g N_VPWR_c_509_n 0.00406853f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_M1008_g N_VPWR_c_509_n 0.00517089f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A_M1011_g N_VPWR_c_501_n 0.00610055f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_174 N_A_M1002_g N_VPWR_c_501_n 0.00534175f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_M1008_g N_VPWR_c_501_n 0.00981361f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A_c_114_n N_Y_M1000_d 0.00166235f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_177 N_A_M1011_g N_Y_c_568_n 0.0208745f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A_c_101_n N_Y_c_568_n 0.00117441f $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_179 N_A_c_104_n N_Y_c_568_n 0.00231928f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_180 N_A_c_105_n N_Y_c_568_n 0.0273196f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_181 N_A_c_106_n N_Y_c_568_n 0.00499812f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_182 N_A_c_101_n N_Y_c_569_n 0.00665349f $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_183 N_A_c_104_n N_Y_c_569_n 0.00101244f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_184 N_A_c_105_n N_Y_c_569_n 0.0252708f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_185 N_A_c_106_n N_Y_c_569_n 0.0103528f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_186 N_A_M1011_g N_Y_c_587_n 0.0197723f $X=0.59 $Y=2.34 $X2=0 $Y2=0
cc_187 N_A_c_106_n N_Y_c_588_n 0.0132561f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_188 N_A_c_106_n N_Y_c_571_n 0.00474295f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_189 N_A_M1002_g N_Y_c_590_n 0.015388f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_M1002_g N_Y_c_591_n 8.05545e-19 $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_M1002_g N_Y_c_592_n 0.00174165f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_c_114_n N_A_641_368#_M1002_s 0.00282287f $X=4.445 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_c_115_n N_A_641_368#_M1002_s 0.00102194f $X=3.355 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_c_114_n N_A_641_368#_M1003_s 0.00108692f $X=4.445 $Y=1.805 $X2=0
+ $Y2=0
cc_195 A N_A_641_368#_M1003_s 0.00113462f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A_M1008_g N_A_641_368#_c_670_n 0.00364476f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_M1008_g N_A_641_368#_c_677_n 0.00632425f $X=4.695 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_M1002_g N_A_641_368#_c_671_n 0.00279882f $X=3.115 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_c_106_n N_VGND_c_698_n 0.00928014f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_200 N_A_c_108_n N_VGND_c_699_n 0.00418692f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_201 N_A_M1007_g N_VGND_c_700_n 0.00460763f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_c_106_n N_VGND_c_701_n 0.00351461f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_203 N_A_c_108_n N_VGND_c_701_n 0.00324657f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_204 N_A_M1007_g N_VGND_c_704_n 0.00327532f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_M1007_g N_VGND_c_705_n 0.00418429f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_c_106_n N_VGND_c_705_n 0.00401739f $X=0.59 $Y=1.22 $X2=0 $Y2=0
cc_207 N_A_c_108_n N_VGND_c_705_n 0.00411282f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_208 N_A_c_100_n N_A_340_107#_c_765_n 0.00521727f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_209 N_A_M1007_g N_A_340_107#_c_766_n 0.00984289f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_c_100_n N_A_340_107#_c_762_n 0.00314462f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_211 N_A_c_100_n N_A_340_107#_c_763_n 0.0107331f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_212 N_A_c_102_n N_A_340_107#_c_763_n 0.00234562f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_213 N_A_c_103_n N_A_340_107#_c_763_n 0.00358921f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_214 N_A_c_108_n N_A_340_107#_c_763_n 0.0103404f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A_c_102_n N_A_340_107#_c_772_n 0.00116104f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_216 N_A_c_103_n N_A_340_107#_c_772_n 0.00891553f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_217 N_A_c_107_n N_A_340_107#_c_772_n 6.51786e-19 $X=3.19 $Y=1.385 $X2=0 $Y2=0
cc_218 N_A_c_108_n N_A_340_107#_c_772_n 0.0104775f $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A_M1007_g N_A_340_107#_c_776_n 7.40195e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_c_108_n N_A_340_107#_c_776_n 7.68469e-19 $X=3.19 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A_M1007_g N_A_340_107#_c_764_n 0.00520058f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B_c_251_n N_A_136_368#_M1009_g 0.00215345f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_223 N_B_c_252_n N_A_136_368#_M1009_g 0.0066709f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_224 N_B_c_264_n N_A_136_368#_M1009_g 0.0143657f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_225 N_B_c_264_n N_A_136_368#_M1010_g 0.0133067f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_226 N_B_M1012_g N_A_136_368#_c_412_n 0.0122231f $X=1.085 $Y=2.34 $X2=0 $Y2=0
cc_227 N_B_c_265_n N_A_136_368#_c_412_n 0.00604058f $X=1.675 $Y=1.805 $X2=0
+ $Y2=0
cc_228 N_B_M1013_g N_A_136_368#_c_405_n 0.00491928f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B_M1012_g N_A_136_368#_c_405_n 0.00467603f $X=1.085 $Y=2.34 $X2=0 $Y2=0
cc_230 N_B_c_250_n N_A_136_368#_c_405_n 0.012913f $X=1.085 $Y=1.515 $X2=0 $Y2=0
cc_231 N_B_c_251_n N_A_136_368#_c_405_n 0.0262874f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B_c_265_n N_A_136_368#_c_405_n 0.00803434f $X=1.675 $Y=1.805 $X2=0
+ $Y2=0
cc_233 N_B_M1013_g N_A_136_368#_c_406_n 0.0171185f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B_c_251_n N_A_136_368#_c_406_n 0.00706196f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_235 N_B_c_252_n N_A_136_368#_c_406_n 0.00720307f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_236 N_B_c_251_n N_A_136_368#_c_407_n 0.0117923f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_237 N_B_c_252_n N_A_136_368#_c_407_n 8.33861e-19 $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_238 N_B_c_264_n N_A_136_368#_c_407_n 0.0482043f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_239 N_B_M1013_g N_A_136_368#_c_408_n 5.78457e-19 $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B_c_251_n N_A_136_368#_c_408_n 0.0139809f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_241 N_B_c_252_n N_A_136_368#_c_408_n 0.00157908f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_242 N_B_c_264_n N_A_136_368#_c_408_n 0.00353018f $X=2.605 $Y=1.805 $X2=0
+ $Y2=0
cc_243 N_B_c_251_n N_A_136_368#_c_409_n 2.6341e-19 $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B_c_252_n N_A_136_368#_c_409_n 0.0113656f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_245 N_B_c_264_n N_A_136_368#_c_409_n 0.010121f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_246 N_B_c_264_n N_VPWR_M1012_d 0.00385927f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_247 N_B_c_265_n N_VPWR_M1012_d 0.00664243f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_248 N_B_c_264_n N_VPWR_M1010_s 5.51361e-19 $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_249 N_B_c_289_n N_VPWR_M1010_s 0.00215336f $X=2.69 $Y=2.06 $X2=0 $Y2=0
cc_250 N_B_c_266_n N_VPWR_M1010_s 0.00986084f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_251 N_B_c_344_p N_VPWR_M1010_s 0.00259146f $X=2.775 $Y=2.145 $X2=0 $Y2=0
cc_252 N_B_c_266_n N_VPWR_M1008_d 0.0108078f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_253 N_B_c_255_n N_VPWR_M1008_d 0.0037127f $X=5.11 $Y=2.06 $X2=0 $Y2=0
cc_254 N_B_c_266_n N_VPWR_c_507_n 0.0247019f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_255 N_B_M1012_g N_VPWR_c_508_n 0.0059286f $X=1.085 $Y=2.34 $X2=0 $Y2=0
cc_256 N_B_M1000_g N_VPWR_c_509_n 0.00333926f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B_M1003_g N_VPWR_c_509_n 0.00333926f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B_M1012_g N_VPWR_c_510_n 0.0096343f $X=1.085 $Y=2.34 $X2=0 $Y2=0
cc_259 N_B_M1012_g N_VPWR_c_501_n 0.00610055f $X=1.085 $Y=2.34 $X2=0 $Y2=0
cc_260 N_B_M1000_g N_VPWR_c_501_n 0.00423353f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B_M1003_g N_VPWR_c_501_n 0.00423254f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B_c_264_n N_Y_M1009_d 0.00165831f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_263 N_B_c_266_n N_Y_M1000_d 0.00321778f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_264 N_B_M1013_g N_Y_c_569_n 0.00103342f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_265 N_B_M1012_g N_Y_c_587_n 0.0155615f $X=1.085 $Y=2.34 $X2=0 $Y2=0
cc_266 N_B_c_252_n N_Y_c_587_n 0.00464167f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_267 N_B_c_264_n N_Y_c_587_n 0.011036f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_268 N_B_c_265_n N_Y_c_587_n 0.0132626f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_269 N_B_M1013_g N_Y_c_588_n 0.00535018f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B_M1000_g N_Y_c_590_n 0.0111198f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_271 N_B_c_264_n N_Y_c_590_n 0.00414614f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_272 N_B_c_266_n N_Y_c_590_n 0.0607542f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_273 N_B_c_344_p N_Y_c_590_n 0.0105714f $X=2.775 $Y=2.145 $X2=0 $Y2=0
cc_274 N_B_M1013_g N_Y_c_573_n 0.0114851f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_275 N_B_M1000_g N_Y_c_591_n 0.00536651f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_276 N_B_M1003_g N_Y_c_591_n 0.00455641f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_277 N_B_c_266_n N_Y_c_591_n 0.016087f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_278 N_B_c_264_n N_Y_c_592_n 0.0215964f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_279 N_B_c_266_n N_A_641_368#_M1002_s 0.0078788f $X=5.025 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_280 N_B_c_266_n N_A_641_368#_M1003_s 0.00434617f $X=5.025 $Y=2.145 $X2=0
+ $Y2=0
cc_281 N_B_M1000_g N_A_641_368#_c_670_n 0.0104179f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_282 N_B_M1003_g N_A_641_368#_c_670_n 0.0118633f $X=4.195 $Y=2.4 $X2=0 $Y2=0
cc_283 N_B_c_266_n N_A_641_368#_c_670_n 0.00323991f $X=5.025 $Y=2.145 $X2=0
+ $Y2=0
cc_284 N_B_c_266_n N_A_641_368#_c_677_n 0.0189154f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_285 N_B_M1000_g N_A_641_368#_c_671_n 4.93815e-19 $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_286 N_B_c_253_n N_VGND_M1005_s 0.0041543f $X=5.025 $Y=1.095 $X2=0 $Y2=0
cc_287 N_B_c_246_n N_VGND_c_699_n 0.00455846f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_288 N_B_c_248_n N_VGND_c_700_n 0.00460763f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_289 N_B_M1013_g N_VGND_c_701_n 0.00278271f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_290 N_B_c_246_n N_VGND_c_703_n 0.00326539f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_291 N_B_c_248_n N_VGND_c_703_n 0.00329249f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_292 N_B_M1013_g N_VGND_c_705_n 0.00358137f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_293 N_B_c_246_n N_VGND_c_705_n 0.00416026f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_294 N_B_c_248_n N_VGND_c_705_n 0.00421564f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_295 N_B_c_254_n N_A_340_107#_M1001_d 0.00267476f $X=4.255 $Y=1.095 $X2=0
+ $Y2=0
cc_296 N_B_c_253_n N_A_340_107#_M1007_s 0.00246551f $X=5.025 $Y=1.095 $X2=0
+ $Y2=0
cc_297 N_B_c_248_n N_A_340_107#_c_766_n 0.0102985f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_298 N_B_c_253_n N_A_340_107#_c_766_n 0.0332405f $X=5.025 $Y=1.095 $X2=0 $Y2=0
cc_299 N_B_M1013_g N_A_340_107#_c_762_n 6.43207e-19 $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B_c_246_n N_A_340_107#_c_763_n 0.00164705f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_301 N_B_c_246_n N_A_340_107#_c_772_n 0.0130102f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_302 N_B_c_246_n N_A_340_107#_c_776_n 0.00555908f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_303 N_B_c_248_n N_A_340_107#_c_776_n 0.00346836f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_304 N_B_c_254_n N_A_340_107#_c_776_n 0.0214926f $X=4.255 $Y=1.095 $X2=0 $Y2=0
cc_305 N_B_c_257_n N_A_340_107#_c_776_n 0.00149766f $X=4.18 $Y=1.43 $X2=0 $Y2=0
cc_306 N_B_c_248_n N_A_340_107#_c_764_n 8.44873e-19 $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_307 N_B_c_253_n N_A_340_107#_c_764_n 0.022058f $X=5.025 $Y=1.095 $X2=0 $Y2=0
cc_308 N_A_136_368#_M1009_g N_VPWR_c_504_n 0.00452919f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_309 N_A_136_368#_M1010_g N_VPWR_c_504_n 0.0039848f $X=2.495 $Y=2.4 $X2=0
+ $Y2=0
cc_310 N_A_136_368#_M1010_g N_VPWR_c_505_n 0.00481925f $X=2.495 $Y=2.4 $X2=0
+ $Y2=0
cc_311 N_A_136_368#_M1009_g N_VPWR_c_510_n 0.0064765f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_312 N_A_136_368#_M1009_g N_VPWR_c_501_n 0.00496497f $X=2.045 $Y=2.4 $X2=0
+ $Y2=0
cc_313 N_A_136_368#_M1010_g N_VPWR_c_501_n 0.00514539f $X=2.495 $Y=2.4 $X2=0
+ $Y2=0
cc_314 N_A_136_368#_c_407_n N_Y_M1004_d 0.00456646f $X=2.42 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_136_368#_c_412_n N_Y_c_568_n 0.013159f $X=1.005 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_136_368#_c_406_n N_Y_c_569_n 0.0143386f $X=1.285 $Y=0.8 $X2=0 $Y2=0
cc_317 N_A_136_368#_M1011_d N_Y_c_587_n 0.00618296f $X=0.68 $Y=1.84 $X2=0 $Y2=0
cc_318 N_A_136_368#_M1009_g N_Y_c_587_n 0.0103539f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_319 N_A_136_368#_c_412_n N_Y_c_587_n 0.0309362f $X=1.005 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_136_368#_c_406_n N_Y_c_588_n 0.0154603f $X=1.285 $Y=0.8 $X2=0 $Y2=0
cc_321 N_A_136_368#_M1010_g N_Y_c_590_n 0.0133886f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_322 N_A_136_368#_c_404_n N_Y_c_572_n 0.00431131f $X=2.705 $Y=1.22 $X2=0 $Y2=0
cc_323 N_A_136_368#_M1013_d N_Y_c_573_n 0.00245749f $X=1.145 $Y=0.37 $X2=0 $Y2=0
cc_324 N_A_136_368#_c_402_n N_Y_c_573_n 0.0123292f $X=2.06 $Y=1.22 $X2=0 $Y2=0
cc_325 N_A_136_368#_c_406_n N_Y_c_573_n 0.0236434f $X=1.285 $Y=0.8 $X2=0 $Y2=0
cc_326 N_A_136_368#_c_408_n N_Y_c_573_n 0.00734058f $X=1.915 $Y=1.28 $X2=0 $Y2=0
cc_327 N_A_136_368#_M1009_g Y 0.0106001f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_328 N_A_136_368#_M1010_g Y 0.00717846f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_329 N_A_136_368#_M1009_g N_Y_c_592_n 0.0202297f $X=2.045 $Y=2.4 $X2=0 $Y2=0
cc_330 N_A_136_368#_M1010_g N_Y_c_592_n 0.00705991f $X=2.495 $Y=2.4 $X2=0 $Y2=0
cc_331 N_A_136_368#_c_402_n N_VGND_c_701_n 0.00278271f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_332 N_A_136_368#_c_404_n N_VGND_c_701_n 0.00324657f $X=2.705 $Y=1.22 $X2=0
+ $Y2=0
cc_333 N_A_136_368#_c_402_n N_VGND_c_705_n 0.00360197f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_334 N_A_136_368#_c_404_n N_VGND_c_705_n 0.00412609f $X=2.705 $Y=1.22 $X2=0
+ $Y2=0
cc_335 N_A_136_368#_c_408_n N_A_340_107#_M1004_s 0.0020198f $X=1.915 $Y=1.28
+ $X2=-0.19 $Y2=-0.245
cc_336 N_A_136_368#_c_402_n N_A_340_107#_c_765_n 0.00868583f $X=2.06 $Y=1.22
+ $X2=0 $Y2=0
cc_337 N_A_136_368#_c_404_n N_A_340_107#_c_765_n 0.0106562f $X=2.705 $Y=1.22
+ $X2=0 $Y2=0
cc_338 N_A_136_368#_c_407_n N_A_340_107#_c_765_n 0.0285439f $X=2.42 $Y=1.385
+ $X2=0 $Y2=0
cc_339 N_A_136_368#_c_409_n N_A_340_107#_c_765_n 0.00135058f $X=2.495 $Y=1.385
+ $X2=0 $Y2=0
cc_340 N_A_136_368#_c_402_n N_A_340_107#_c_762_n 0.00263714f $X=2.06 $Y=1.22
+ $X2=0 $Y2=0
cc_341 N_A_136_368#_c_404_n N_A_340_107#_c_762_n 3.24573e-19 $X=2.705 $Y=1.22
+ $X2=0 $Y2=0
cc_342 N_A_136_368#_c_406_n N_A_340_107#_c_762_n 0.0147768f $X=1.285 $Y=0.8
+ $X2=0 $Y2=0
cc_343 N_A_136_368#_c_408_n N_A_340_107#_c_762_n 0.0285439f $X=1.915 $Y=1.28
+ $X2=0 $Y2=0
cc_344 N_A_136_368#_c_409_n N_A_340_107#_c_762_n 2.18933e-19 $X=2.495 $Y=1.385
+ $X2=0 $Y2=0
cc_345 N_A_136_368#_c_402_n N_A_340_107#_c_763_n 0.00164025f $X=2.06 $Y=1.22
+ $X2=0 $Y2=0
cc_346 N_A_136_368#_c_404_n N_A_340_107#_c_763_n 0.0106998f $X=2.705 $Y=1.22
+ $X2=0 $Y2=0
cc_347 N_VPWR_M1011_s N_Y_c_568_n 0.00902214f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_348 N_VPWR_M1011_s N_Y_c_587_n 0.00969112f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_349 N_VPWR_M1012_d N_Y_c_587_n 0.0216743f $X=1.175 $Y=1.84 $X2=0 $Y2=0
cc_350 N_VPWR_c_503_n N_Y_c_587_n 0.0149256f $X=0.28 $Y=2.825 $X2=0 $Y2=0
cc_351 N_VPWR_c_510_n N_Y_c_587_n 0.0510878f $X=1.79 $Y=2.825 $X2=0 $Y2=0
cc_352 N_VPWR_c_501_n N_Y_c_587_n 0.0338979f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_353 N_VPWR_M1011_s N_Y_c_575_n 0.00242814f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_354 N_VPWR_c_503_n N_Y_c_575_n 0.0122531f $X=0.28 $Y=2.825 $X2=0 $Y2=0
cc_355 N_VPWR_c_501_n N_Y_c_575_n 0.00170605f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_356 N_VPWR_M1010_s N_Y_c_590_n 0.00760776f $X=2.585 $Y=1.84 $X2=0 $Y2=0
cc_357 N_VPWR_c_504_n N_Y_c_590_n 0.00224454f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_358 N_VPWR_c_505_n N_Y_c_590_n 0.0257224f $X=2.805 $Y=2.905 $X2=0 $Y2=0
cc_359 N_VPWR_c_509_n N_Y_c_590_n 0.00302133f $X=4.805 $Y=3.33 $X2=0 $Y2=0
cc_360 N_VPWR_c_501_n N_Y_c_590_n 0.0135637f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_361 N_VPWR_c_504_n Y 0.0169602f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_362 N_VPWR_c_505_n Y 0.00864627f $X=2.805 $Y=2.905 $X2=0 $Y2=0
cc_363 N_VPWR_c_510_n Y 0.0265326f $X=1.79 $Y=2.825 $X2=0 $Y2=0
cc_364 N_VPWR_c_501_n Y 0.013761f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_365 N_VPWR_c_507_n N_A_641_368#_c_670_n 0.0119238f $X=4.97 $Y=2.485 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_509_n N_A_641_368#_c_670_n 0.0678759f $X=4.805 $Y=3.33 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_501_n N_A_641_368#_c_670_n 0.0375541f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_505_n N_A_641_368#_c_671_n 0.0065515f $X=2.805 $Y=2.905 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_509_n N_A_641_368#_c_671_n 0.0229944f $X=4.805 $Y=3.33 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_501_n N_A_641_368#_c_671_n 0.012911f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_371 N_Y_c_590_n N_A_641_368#_M1002_s 0.00791485f $X=3.805 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_372 N_Y_M1000_d N_A_641_368#_c_670_n 0.00165831f $X=3.835 $Y=1.84 $X2=0 $Y2=0
cc_373 N_Y_c_590_n N_A_641_368#_c_670_n 0.00516104f $X=3.805 $Y=2.485 $X2=0
+ $Y2=0
cc_374 N_Y_c_591_n N_A_641_368#_c_670_n 0.0151027f $X=3.97 $Y=2.485 $X2=0 $Y2=0
cc_375 N_Y_c_590_n N_A_641_368#_c_671_n 0.0250247f $X=3.805 $Y=2.485 $X2=0 $Y2=0
cc_376 N_Y_c_569_n N_VGND_M1014_s 0.00690923f $X=0.665 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_377 N_Y_c_569_n N_VGND_c_698_n 0.0192864f $X=0.665 $Y=0.925 $X2=0 $Y2=0
cc_378 N_Y_c_570_n N_VGND_c_698_n 0.0127101f $X=0.255 $Y=0.925 $X2=0 $Y2=0
cc_379 N_Y_c_588_n N_VGND_c_698_n 0.0183033f $X=0.75 $Y=0.84 $X2=0 $Y2=0
cc_380 N_Y_c_571_n N_VGND_c_698_n 0.0143324f $X=0.835 $Y=0.34 $X2=0 $Y2=0
cc_381 N_Y_c_571_n N_VGND_c_701_n 0.0118705f $X=0.835 $Y=0.34 $X2=0 $Y2=0
cc_382 N_Y_c_573_n N_VGND_c_701_n 0.111797f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_383 N_Y_c_569_n N_VGND_c_705_n 0.00623186f $X=0.665 $Y=0.925 $X2=0 $Y2=0
cc_384 N_Y_c_570_n N_VGND_c_705_n 0.00172823f $X=0.255 $Y=0.925 $X2=0 $Y2=0
cc_385 N_Y_c_571_n N_VGND_c_705_n 0.0061974f $X=0.835 $Y=0.34 $X2=0 $Y2=0
cc_386 N_Y_c_573_n N_VGND_c_705_n 0.0641627f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_387 N_Y_c_569_n A_151_74# 0.00170774f $X=0.665 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_388 N_Y_c_588_n A_151_74# 0.00411005f $X=0.75 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_389 N_Y_c_573_n A_151_74# 0.00389187f $X=2.19 $Y=0.377 $X2=-0.19 $Y2=-0.245
cc_390 N_Y_c_573_n N_A_340_107#_M1004_s 0.00226585f $X=2.19 $Y=0.377 $X2=-0.19
+ $Y2=-0.245
cc_391 N_Y_M1004_d N_A_340_107#_c_765_n 0.00860281f $X=2.135 $Y=0.37 $X2=0 $Y2=0
cc_392 N_Y_c_572_n N_A_340_107#_c_765_n 0.0271762f $X=2.38 $Y=0.415 $X2=0 $Y2=0
cc_393 N_Y_c_573_n N_A_340_107#_c_765_n 0.00570513f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_394 N_Y_c_573_n N_A_340_107#_c_762_n 0.0191024f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_395 N_Y_c_572_n N_A_340_107#_c_763_n 0.00621476f $X=2.38 $Y=0.415 $X2=0 $Y2=0
cc_396 N_VGND_c_701_n N_A_340_107#_c_765_n 0.00237563f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_705_n N_A_340_107#_c_765_n 0.00549522f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_398 N_VGND_M1005_s N_A_340_107#_c_766_n 0.00787506f $X=4.255 $Y=0.37 $X2=0
+ $Y2=0
cc_399 N_VGND_c_700_n N_A_340_107#_c_766_n 0.0262746f $X=4.48 $Y=0.335 $X2=0
+ $Y2=0
cc_400 N_VGND_c_703_n N_A_340_107#_c_766_n 0.00266206f $X=4.31 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_704_n N_A_340_107#_c_766_n 0.0023667f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_705_n N_A_340_107#_c_766_n 0.0107342f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_c_699_n N_A_340_107#_c_763_n 0.00613715f $X=3.43 $Y=0.335 $X2=0
+ $Y2=0
cc_404 N_VGND_c_701_n N_A_340_107#_c_763_n 0.0144609f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_c_705_n N_A_340_107#_c_763_n 0.0118703f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_406 N_VGND_M1006_d N_A_340_107#_c_772_n 0.0145608f $X=3.21 $Y=0.37 $X2=0
+ $Y2=0
cc_407 N_VGND_c_699_n N_A_340_107#_c_772_n 0.0255041f $X=3.43 $Y=0.335 $X2=0
+ $Y2=0
cc_408 N_VGND_c_701_n N_A_340_107#_c_772_n 0.0023667f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_703_n N_A_340_107#_c_772_n 0.00236055f $X=4.31 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_705_n N_A_340_107#_c_772_n 0.0102361f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_703_n N_A_340_107#_c_776_n 0.00723046f $X=4.31 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_705_n N_A_340_107#_c_776_n 0.0106441f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_704_n N_A_340_107#_c_764_n 0.00789542f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_705_n N_A_340_107#_c_764_n 0.0106304f $X=5.04 $Y=0 $X2=0 $Y2=0

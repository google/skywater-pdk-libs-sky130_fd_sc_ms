* File: sky130_fd_sc_ms__nand3_1.pxi.spice
* Created: Fri Aug 28 17:43:03 2020
* 
x_PM_SKY130_FD_SC_MS__NAND3_1%C N_C_M1003_g N_C_c_39_n N_C_M1002_g C C
+ N_C_c_41_n PM_SKY130_FD_SC_MS__NAND3_1%C
x_PM_SKY130_FD_SC_MS__NAND3_1%B N_B_M1001_g N_B_M1005_g B B B N_B_c_65_n
+ N_B_c_66_n PM_SKY130_FD_SC_MS__NAND3_1%B
x_PM_SKY130_FD_SC_MS__NAND3_1%A N_A_M1000_g N_A_M1004_g A N_A_c_103_n
+ N_A_c_104_n PM_SKY130_FD_SC_MS__NAND3_1%A
x_PM_SKY130_FD_SC_MS__NAND3_1%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_c_134_n
+ N_VPWR_c_135_n N_VPWR_c_136_n N_VPWR_c_137_n N_VPWR_c_138_n VPWR
+ N_VPWR_c_139_n N_VPWR_c_133_n PM_SKY130_FD_SC_MS__NAND3_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND3_1%Y N_Y_M1000_d N_Y_M1003_d N_Y_M1004_d N_Y_c_165_n
+ N_Y_c_166_n N_Y_c_162_n N_Y_c_167_n N_Y_c_163_n N_Y_c_164_n N_Y_c_169_n Y Y Y
+ N_Y_c_170_n PM_SKY130_FD_SC_MS__NAND3_1%Y
x_PM_SKY130_FD_SC_MS__NAND3_1%VGND N_VGND_M1002_s N_VGND_c_213_n N_VGND_c_214_n
+ N_VGND_c_215_n VGND N_VGND_c_216_n N_VGND_c_217_n
+ PM_SKY130_FD_SC_MS__NAND3_1%VGND
cc_1 VNB N_C_M1003_g 0.00936933f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.4
cc_2 VNB N_C_c_39_n 0.0208066f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_3 VNB C 0.0311109f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C_c_41_n 0.0694136f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_5 VNB N_B_M1005_g 0.00667073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB B 0.00244094f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_7 VNB N_B_c_65_n 0.0326751f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_8 VNB N_B_c_66_n 0.0180991f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_9 VNB N_A_M1004_g 0.00735656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A 0.00684394f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_11 VNB N_A_c_103_n 0.0327357f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A_c_104_n 0.0229091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_133_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_162_n 0.02133f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.385
cc_15 VNB N_Y_c_163_n 0.0320047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_164_n 0.0146427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_213_n 0.0344107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_214_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_19 VNB N_VGND_c_215_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_VGND_c_216_n 0.0529515f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_21 VNB N_VGND_c_217_n 0.18517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_C_M1003_g 0.0280487f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.4
cc_23 VPB N_B_M1005_g 0.0233482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_24 VPB N_A_M1004_g 0.0290507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_134_n 0.012885f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_26 VPB N_VPWR_c_135_n 0.0563013f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_27 VPB N_VPWR_c_136_n 0.00976275f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_28 VPB N_VPWR_c_137_n 0.0213359f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_29 VPB N_VPWR_c_138_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_30 VPB N_VPWR_c_139_n 0.0253045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_133_n 0.0630422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_Y_c_165_n 0.00881636f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_33 VPB N_Y_c_166_n 0.00807857f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_34 VPB N_Y_c_167_n 0.055594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_Y_c_163_n 0.00301672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_Y_c_169_n 0.0165104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_Y_c_170_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 N_C_M1003_g N_B_M1005_g 0.0231643f $X=0.655 $Y=2.4 $X2=0 $Y2=0
cc_39 N_C_c_39_n B 0.0034981f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_40 C B 0.0296912f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_41 N_C_c_41_n N_B_c_65_n 0.0329663f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_42 N_C_c_39_n N_B_c_66_n 0.0329663f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_43 C N_B_c_66_n 0.00239222f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_44 N_C_M1003_g N_VPWR_c_135_n 0.0285123f $X=0.655 $Y=2.4 $X2=0 $Y2=0
cc_45 C N_VPWR_c_135_n 0.0149317f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_46 N_C_c_41_n N_VPWR_c_135_n 0.00546342f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_47 N_C_M1003_g N_VPWR_c_137_n 0.00396269f $X=0.655 $Y=2.4 $X2=0 $Y2=0
cc_48 N_C_M1003_g N_VPWR_c_133_n 0.00584081f $X=0.655 $Y=2.4 $X2=0 $Y2=0
cc_49 N_C_M1003_g N_Y_c_166_n 0.0103944f $X=0.655 $Y=2.4 $X2=0 $Y2=0
cc_50 C N_Y_c_166_n 0.0191701f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_51 N_C_c_41_n N_Y_c_166_n 8.17195e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_52 N_C_M1003_g N_Y_c_170_n 0.0229299f $X=0.655 $Y=2.4 $X2=0 $Y2=0
cc_53 N_C_c_39_n N_VGND_c_213_n 0.0151342f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_54 C N_VGND_c_213_n 0.0259403f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_55 N_C_c_41_n N_VGND_c_213_n 0.00199349f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_56 N_C_c_39_n N_VGND_c_216_n 0.00383152f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_57 N_C_c_39_n N_VGND_c_217_n 0.0075725f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_58 N_B_M1005_g N_A_M1004_g 0.0274726f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_59 B A 0.0244362f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_60 N_B_c_65_n A 0.00202352f $X=1.18 $Y=1.385 $X2=0 $Y2=0
cc_61 B N_A_c_103_n 4.06701e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_62 N_B_c_65_n N_A_c_103_n 0.0175474f $X=1.18 $Y=1.385 $X2=0 $Y2=0
cc_63 B N_A_c_104_n 0.00897929f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_64 N_B_c_66_n N_A_c_104_n 0.0246919f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_65 N_B_M1005_g N_VPWR_c_136_n 0.00347203f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_66 N_B_M1005_g N_VPWR_c_137_n 0.005209f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_67 N_B_M1005_g N_VPWR_c_133_n 0.00982843f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_68 N_B_M1005_g N_Y_c_165_n 0.0135147f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_69 B N_Y_c_165_n 0.0232997f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_70 N_B_c_65_n N_Y_c_165_n 0.00105037f $X=1.18 $Y=1.385 $X2=0 $Y2=0
cc_71 N_B_M1005_g N_Y_c_166_n 0.00224432f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_72 B N_Y_c_166_n 0.00245488f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_73 B N_Y_c_162_n 0.0172672f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_B_c_66_n N_Y_c_162_n 7.56255e-19 $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_75 N_B_M1005_g N_Y_c_167_n 7.0357e-19 $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_76 B N_Y_c_164_n 0.00754251f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_77 N_B_M1005_g N_Y_c_170_n 0.015174f $X=1.105 $Y=2.4 $X2=0 $Y2=0
cc_78 B N_VGND_c_213_n 0.023155f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_79 N_B_c_66_n N_VGND_c_213_n 0.00251629f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_80 B N_VGND_c_216_n 0.00930091f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_81 N_B_c_66_n N_VGND_c_216_n 0.00304348f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_82 B N_VGND_c_217_n 0.0106938f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_83 N_B_c_66_n N_VGND_c_217_n 0.00371612f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_84 B A_233_74# 0.00988329f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_85 N_A_M1004_g N_VPWR_c_136_n 0.00879843f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VPWR_c_139_n 0.005209f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_VPWR_c_133_n 0.00987481f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_Y_c_165_n 0.0135147f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_89 A N_Y_c_165_n 0.0123606f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A_c_104_n N_Y_c_162_n 0.00846119f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_91 N_A_M1004_g N_Y_c_167_n 0.0164413f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_M1004_g N_Y_c_163_n 0.00503397f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_93 A N_Y_c_163_n 0.0280999f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A_c_103_n N_Y_c_163_n 0.00739878f $X=1.75 $Y=1.385 $X2=0 $Y2=0
cc_95 N_A_c_104_n N_Y_c_163_n 0.00394268f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_96 A N_Y_c_164_n 0.0138478f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A_c_103_n N_Y_c_164_n 0.001011f $X=1.75 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A_c_104_n N_Y_c_164_n 0.00296171f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_99 N_A_M1004_g N_Y_c_169_n 0.00357848f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_100 A N_Y_c_169_n 0.0151534f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A_c_103_n N_Y_c_169_n 0.0011793f $X=1.75 $Y=1.385 $X2=0 $Y2=0
cc_102 N_A_M1004_g N_Y_c_170_n 9.51264e-19 $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_c_104_n N_VGND_c_216_n 0.00434272f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_104 N_A_c_104_n N_VGND_c_217_n 0.00822158f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_105 N_VPWR_M1005_d N_Y_c_165_n 0.0030153f $X=1.195 $Y=1.84 $X2=0 $Y2=0
cc_106 N_VPWR_c_136_n N_Y_c_165_n 0.022455f $X=1.38 $Y=2.145 $X2=0 $Y2=0
cc_107 N_VPWR_c_135_n N_Y_c_166_n 0.0056822f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_108 N_VPWR_c_136_n N_Y_c_167_n 0.0345826f $X=1.38 $Y=2.145 $X2=0 $Y2=0
cc_109 N_VPWR_c_139_n N_Y_c_167_n 0.0230269f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_110 N_VPWR_c_133_n N_Y_c_167_n 0.0189916f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_111 N_VPWR_c_135_n N_Y_c_170_n 0.0846655f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_112 N_VPWR_c_136_n N_Y_c_170_n 0.0368642f $X=1.38 $Y=2.145 $X2=0 $Y2=0
cc_113 N_VPWR_c_137_n N_Y_c_170_n 0.0190418f $X=1.215 $Y=3.33 $X2=0 $Y2=0
cc_114 N_VPWR_c_133_n N_Y_c_170_n 0.0153665f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_115 N_Y_c_162_n N_VGND_c_216_n 0.0142249f $X=1.875 $Y=0.515 $X2=0 $Y2=0
cc_116 N_Y_c_162_n N_VGND_c_217_n 0.011867f $X=1.875 $Y=0.515 $X2=0 $Y2=0
cc_117 N_Y_c_164_n N_VGND_c_217_n 0.00749433f $X=2.17 $Y=0.925 $X2=0 $Y2=0

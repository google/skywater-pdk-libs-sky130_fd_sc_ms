* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 Y B1 a_351_74# VNB nlowvt w=740000u l=150000u
+  ad=8.695e+11p pd=5.31e+06u as=1.554e+11p ps=1.9e+06u
M1001 a_121_368# B2 a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=5.936e+11p pd=5.54e+06u as=9.184e+11p ps=8.36e+06u
M1002 VPWR A1 a_263_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.032e+11p pd=2.96e+06u as=0p ps=0u
M1003 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=0p ps=0u
M1004 a_263_368# B1 a_121_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_263_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_567_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1007 VGND A2 a_567_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_351_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_121_368# C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
.ends

* File: sky130_fd_sc_ms__or2_1.pex.spice
* Created: Fri Aug 28 18:06:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR2_1%B 5 7 9 10 13 14
r27 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r28 10 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r29 7 13 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.7 $Y=1.22
+ $X2=0.685 $Y2=1.385
r30 7 9 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.7 $Y=1.22 $X2=0.7
+ $Y2=0.835
r31 3 13 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.685 $Y=1.55
+ $X2=0.685 $Y2=1.385
r32 3 5 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=0.685 $Y=1.55
+ $X2=0.685 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_1%A 3 7 9 13 14
c40 13 0 6.83128e-20 $X=1.21 $Y=1.515
c41 7 0 7.78164e-20 $X=1.325 $Y=0.835
r42 13 15 17.5968 $w=3.15e-07 $l=1.15e-07 $layer=POLY_cond $X=1.21 $Y=1.515
+ $X2=1.325 $Y2=1.515
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.515 $X2=1.21 $Y2=1.515
r44 11 13 16.0667 $w=3.15e-07 $l=1.05e-07 $layer=POLY_cond $X=1.105 $Y=1.515
+ $X2=1.21 $Y2=1.515
r45 9 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.21 $Y=1.665
+ $X2=1.21 $Y2=1.515
r46 5 15 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.35
+ $X2=1.325 $Y2=1.515
r47 5 7 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.325 $Y=1.35
+ $X2=1.325 $Y2=0.835
r48 1 11 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.68
+ $X2=1.105 $Y2=1.515
r49 1 3 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.105 $Y=1.68
+ $X2=1.105 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_1%A_63_368# 1 2 9 13 17 21 23 24 25 26 28 32
c72 23 0 6.83128e-20 $X=1.615 $Y=1.095
r73 32 35 40.7387 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.812 $Y=1.465
+ $X2=1.812 $Y2=1.63
r74 32 34 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.812 $Y=1.465
+ $X2=1.812 $Y2=1.3
r75 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.805
+ $Y=1.465 $X2=1.805 $Y2=1.465
r76 25 31 9.13575 $w=2.68e-07 $l=2.05925e-07 $layer=LI1_cond $X=1.7 $Y=1.63
+ $X2=1.792 $Y2=1.465
r77 25 26 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.7 $Y=1.63 $X2=1.7
+ $Y2=1.95
r78 23 31 16.8433 $w=2.68e-07 $l=4.49878e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=1.792 $Y2=1.465
r79 23 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.615 $Y=1.095
+ $X2=1.24 $Y2=1.095
r80 19 24 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.092 $Y=1.01
+ $X2=1.24 $Y2=1.095
r81 19 21 7.42251 $w=2.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.092 $Y=1.01
+ $X2=1.092 $Y2=0.82
r82 18 28 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.625 $Y=2.035
+ $X2=0.46 $Y2=1.97
r83 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=1.7 $Y2=1.95
r84 17 18 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=0.625 $Y2=2.035
r85 13 34 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.905 $Y=0.74
+ $X2=1.905 $Y2=1.3
r86 9 35 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.895 $Y=2.4
+ $X2=1.895 $Y2=1.63
r87 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.315
+ $Y=1.84 $X2=0.46 $Y2=1.985
r88 1 21 182 $w=1.7e-07 $l=4.09878e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.56 $X2=1.075 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_1%VPWR 1 6 8 10 17 18 21
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 15 21 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.475 $Y2=3.33
r29 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=1.475 $Y2=3.33
r32 10 12 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r34 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r35 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 4 21 2.59604 $w=6.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=3.33
r37 4 6 15.2404 $w=6.18e-07 $l=7.9e-07 $layer=LI1_cond $X=1.475 $Y=3.245
+ $X2=1.475 $Y2=2.455
r38 1 6 200 $w=1.7e-07 $l=8.18749e-07 $layer=licon1_PDIFF $count=3 $X=1.195
+ $Y=1.84 $X2=1.67 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_1%X 1 2 9 13 14 15 16 23 32
c25 13 0 7.78164e-20 $X=2.132 $Y=1.13
r26 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=2.132 $Y=1.997
+ $X2=2.132 $Y2=2.035
r27 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.132 $Y=2.405
+ $X2=2.132 $Y2=2.775
r28 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=2.132 $Y=1.973
+ $X2=2.132 $Y2=1.997
r29 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=2.132 $Y=1.973
+ $X2=2.132 $Y2=1.82
r30 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=2.132 $Y=2.058
+ $X2=2.132 $Y2=2.405
r31 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=2.132 $Y=2.058
+ $X2=2.132 $Y2=2.035
r32 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.225 $Y=1.13
+ $X2=2.225 $Y2=1.82
r33 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=2.132 $Y=0.953
+ $X2=2.132 $Y2=1.13
r34 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=2.132 $Y=0.953
+ $X2=2.132 $Y2=0.515
r35 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=1.985
r36 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.37 $X2=2.12 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2_1%VGND 1 2 9 13 16 17 18 23 29 30 33
r32 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r33 30 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r34 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 27 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r36 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.16
+ $Y2=0
r37 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r38 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.2
+ $Y2=0
r39 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 18 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r41 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r42 18 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 16 21 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.24
+ $Y2=0
r44 16 17 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.472
+ $Y2=0
r45 15 25 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=1.2
+ $Y2=0
r46 15 17 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.472
+ $Y2=0
r47 11 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r48 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.675
r49 7 17 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.472 $Y=0.085
+ $X2=0.472 $Y2=0
r50 7 9 24.1851 $w=3.53e-07 $l=7.45e-07 $layer=LI1_cond $X=0.472 $Y=0.085
+ $X2=0.472 $Y2=0.83
r51 2 13 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.56 $X2=1.62 $Y2=0.675
r52 1 9 182 $w=1.7e-07 $l=4.65833e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.485 $Y2=0.83
.ends


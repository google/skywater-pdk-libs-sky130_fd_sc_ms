* File: sky130_fd_sc_ms__o221ai_4.pxi.spice
* Created: Wed Sep  2 12:23:22 2020
* 
x_PM_SKY130_FD_SC_MS__O221AI_4%C1 N_C1_M1013_g N_C1_M1000_g N_C1_M1002_g
+ N_C1_M1014_g N_C1_M1004_g N_C1_M1024_g N_C1_M1018_g N_C1_M1035_g C1 C1 C1
+ N_C1_c_151_n N_C1_c_152_n PM_SKY130_FD_SC_MS__O221AI_4%C1
x_PM_SKY130_FD_SC_MS__O221AI_4%B1 N_B1_M1003_g N_B1_M1009_g N_B1_M1020_g
+ N_B1_c_232_n N_B1_M1011_g N_B1_M1022_g N_B1_c_233_n N_B1_M1030_g N_B1_M1037_g
+ N_B1_M1028_g N_B1_c_249_n N_B1_c_243_n N_B1_c_235_n B1 N_B1_c_236_n
+ N_B1_c_237_n N_B1_c_238_n PM_SKY130_FD_SC_MS__O221AI_4%B1
x_PM_SKY130_FD_SC_MS__O221AI_4%B2 N_B2_c_366_n N_B2_M1005_g N_B2_c_358_n
+ N_B2_M1006_g N_B2_c_367_n N_B2_M1025_g N_B2_c_359_n N_B2_M1015_g N_B2_M1032_g
+ N_B2_c_361_n N_B2_M1016_g N_B2_c_362_n N_B2_M1036_g N_B2_c_364_n N_B2_M1026_g
+ B2 B2 PM_SKY130_FD_SC_MS__O221AI_4%B2
x_PM_SKY130_FD_SC_MS__O221AI_4%A1 N_A1_M1008_g N_A1_M1001_g N_A1_M1027_g
+ N_A1_M1010_g N_A1_M1038_g N_A1_M1031_g N_A1_M1039_g N_A1_M1034_g N_A1_c_450_n
+ N_A1_c_451_n A1 A1 A1 A1 N_A1_c_453_n N_A1_c_454_n A1 N_A1_c_455_n
+ PM_SKY130_FD_SC_MS__O221AI_4%A1
x_PM_SKY130_FD_SC_MS__O221AI_4%A2 N_A2_M1007_g N_A2_M1021_g N_A2_M1012_g
+ N_A2_M1023_g N_A2_M1029_g N_A2_M1017_g N_A2_M1033_g N_A2_M1019_g A2 A2 A2
+ N_A2_c_568_n PM_SKY130_FD_SC_MS__O221AI_4%A2
x_PM_SKY130_FD_SC_MS__O221AI_4%VPWR N_VPWR_M1013_s N_VPWR_M1014_s N_VPWR_M1035_s
+ N_VPWR_M1020_d N_VPWR_M1028_d N_VPWR_M1010_s N_VPWR_M1039_s N_VPWR_c_649_n
+ N_VPWR_c_650_n N_VPWR_c_651_n N_VPWR_c_652_n N_VPWR_c_653_n N_VPWR_c_654_n
+ N_VPWR_c_655_n N_VPWR_c_656_n N_VPWR_c_657_n VPWR N_VPWR_c_658_n
+ N_VPWR_c_659_n N_VPWR_c_660_n N_VPWR_c_661_n N_VPWR_c_662_n N_VPWR_c_663_n
+ N_VPWR_c_664_n N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n
+ N_VPWR_c_648_n PM_SKY130_FD_SC_MS__O221AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O221AI_4%Y N_Y_M1000_s N_Y_M1004_s N_Y_M1013_d N_Y_M1024_d
+ N_Y_M1005_s N_Y_M1032_s N_Y_M1021_d N_Y_M1029_d N_Y_c_784_n N_Y_c_787_n
+ N_Y_c_780_n N_Y_c_776_n N_Y_c_777_n N_Y_c_802_n N_Y_c_806_n N_Y_c_781_n
+ N_Y_c_811_n N_Y_c_890_p N_Y_c_833_n N_Y_c_834_n N_Y_c_835_n N_Y_c_854_n
+ N_Y_c_778_n N_Y_c_782_n N_Y_c_779_n N_Y_c_840_n N_Y_c_841_n N_Y_c_858_n Y
+ PM_SKY130_FD_SC_MS__O221AI_4%Y
x_PM_SKY130_FD_SC_MS__O221AI_4%A_511_368# N_A_511_368#_M1003_s
+ N_A_511_368#_M1022_s N_A_511_368#_M1025_d N_A_511_368#_M1036_d
+ N_A_511_368#_c_924_n N_A_511_368#_c_926_n N_A_511_368#_c_927_n
+ N_A_511_368#_c_915_n N_A_511_368#_c_916_n N_A_511_368#_c_941_n
+ N_A_511_368#_c_917_n N_A_511_368#_c_931_n N_A_511_368#_c_918_n
+ N_A_511_368#_c_919_n PM_SKY130_FD_SC_MS__O221AI_4%A_511_368#
x_PM_SKY130_FD_SC_MS__O221AI_4%A_1291_368# N_A_1291_368#_M1001_d
+ N_A_1291_368#_M1023_s N_A_1291_368#_M1033_s N_A_1291_368#_M1038_d
+ N_A_1291_368#_c_979_n N_A_1291_368#_c_1022_n N_A_1291_368#_c_980_n
+ N_A_1291_368#_c_985_n N_A_1291_368#_c_986_n N_A_1291_368#_c_990_n
+ N_A_1291_368#_c_981_n N_A_1291_368#_c_982_n N_A_1291_368#_c_983_n
+ PM_SKY130_FD_SC_MS__O221AI_4%A_1291_368#
x_PM_SKY130_FD_SC_MS__O221AI_4%A_27_84# N_A_27_84#_M1000_d N_A_27_84#_M1002_d
+ N_A_27_84#_M1018_d N_A_27_84#_M1009_d N_A_27_84#_M1030_d N_A_27_84#_M1015_s
+ N_A_27_84#_M1026_s N_A_27_84#_c_1027_n N_A_27_84#_c_1028_n N_A_27_84#_c_1029_n
+ N_A_27_84#_c_1078_n N_A_27_84#_c_1030_n N_A_27_84#_c_1031_n
+ N_A_27_84#_c_1032_n N_A_27_84#_c_1033_n N_A_27_84#_c_1034_n
+ N_A_27_84#_c_1035_n N_A_27_84#_c_1036_n N_A_27_84#_c_1037_n
+ N_A_27_84#_c_1061_n N_A_27_84#_c_1067_n PM_SKY130_FD_SC_MS__O221AI_4%A_27_84#
x_PM_SKY130_FD_SC_MS__O221AI_4%A_483_74# N_A_483_74#_M1009_s N_A_483_74#_M1011_s
+ N_A_483_74#_M1006_d N_A_483_74#_M1016_d N_A_483_74#_M1037_s
+ N_A_483_74#_M1007_s N_A_483_74#_M1017_s N_A_483_74#_M1027_d
+ N_A_483_74#_M1034_d N_A_483_74#_c_1107_n N_A_483_74#_c_1108_n
+ N_A_483_74#_c_1129_n N_A_483_74#_c_1109_n N_A_483_74#_c_1134_n
+ N_A_483_74#_c_1110_n N_A_483_74#_c_1135_n N_A_483_74#_c_1111_n
+ N_A_483_74#_c_1112_n N_A_483_74#_c_1113_n N_A_483_74#_c_1114_n
+ N_A_483_74#_c_1147_n N_A_483_74#_c_1148_n N_A_483_74#_c_1149_n
+ PM_SKY130_FD_SC_MS__O221AI_4%A_483_74#
x_PM_SKY130_FD_SC_MS__O221AI_4%VGND N_VGND_M1008_s N_VGND_M1012_d N_VGND_M1019_d
+ N_VGND_M1031_s N_VGND_c_1217_n N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n
+ VGND N_VGND_c_1221_n N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n
+ N_VGND_c_1225_n N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n
+ N_VGND_c_1229_n N_VGND_c_1230_n PM_SKY130_FD_SC_MS__O221AI_4%VGND
cc_1 VNB N_C1_M1000_g 0.0263359f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_2 VNB N_C1_M1002_g 0.0191476f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_3 VNB N_C1_M1004_g 0.0191247f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.79
cc_4 VNB N_C1_M1018_g 0.0256157f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_5 VNB N_C1_c_151_n 0.0167416f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.515
cc_6 VNB N_C1_c_152_n 0.0837029f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.515
cc_7 VNB N_B1_M1009_g 0.0308588f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_8 VNB N_B1_c_232_n 0.0146162f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_9 VNB N_B1_c_233_n 0.0147307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1037_g 0.0257119f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_11 VNB N_B1_c_235_n 0.0037594f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_12 VNB N_B1_c_236_n 0.0862693f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.515
cc_13 VNB N_B1_c_237_n 0.0250033f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_14 VNB N_B1_c_238_n 0.00725477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_358_n 0.0169363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B2_c_359_n 0.0166753f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_17 VNB N_B2_M1032_g 0.00601454f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_18 VNB N_B2_c_361_n 0.0166979f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_19 VNB N_B2_c_362_n 0.094423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_M1036_g 0.0061634f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.4
cc_21 VNB N_B2_c_364_n 0.017373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B2 0.00745009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_M1008_g 0.021903f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_24 VNB N_A1_M1001_g 0.00405989f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_25 VNB N_A1_M1027_g 0.0196218f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_26 VNB N_A1_M1010_g 0.00309826f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_27 VNB N_A1_M1038_g 0.00309312f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.79
cc_28 VNB N_A1_M1031_g 0.0192941f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.4
cc_29 VNB N_A1_M1039_g 0.00418093f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_30 VNB N_A1_M1034_g 0.0262473f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_31 VNB N_A1_c_450_n 0.0104553f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_A1_c_451_n 0.0286608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB A1 0.0222352f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_34 VNB N_A1_c_453_n 0.063562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A1_c_454_n 0.0147594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A1_c_455_n 0.0016599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A2_M1007_g 0.0238876f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_38 VNB N_A2_M1012_g 0.0227944f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.79
cc_39 VNB N_A2_M1017_g 0.0233499f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.4
cc_40 VNB N_A2_M1019_g 0.0216231f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_41 VNB N_A2_c_568_n 0.0694159f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.515
cc_42 VNB N_VPWR_c_648_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_776_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_44 VNB N_Y_c_777_n 0.00229834f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_45 VNB N_Y_c_778_n 0.00421298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_779_n 0.00159633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_84#_c_1027_n 0.0307564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_84#_c_1028_n 0.00475623f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_49 VNB N_A_27_84#_c_1029_n 0.00958293f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_50 VNB N_A_27_84#_c_1030_n 0.00952739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_84#_c_1031_n 0.00400018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_84#_c_1032_n 0.0199341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_84#_c_1033_n 0.00690962f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_54 VNB N_A_27_84#_c_1034_n 0.00225825f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_55 VNB N_A_27_84#_c_1035_n 0.00136506f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.515
cc_56 VNB N_A_27_84#_c_1036_n 0.00138842f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.515
cc_57 VNB N_A_27_84#_c_1037_n 0.00348266f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=1.515
cc_58 VNB N_A_483_74#_c_1107_n 0.00940936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_483_74#_c_1108_n 0.0127258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_483_74#_c_1109_n 0.00206045f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_61 VNB N_A_483_74#_c_1110_n 0.00206045f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.515
cc_62 VNB N_A_483_74#_c_1111_n 0.00252795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_483_74#_c_1112_n 0.0075506f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_64 VNB N_A_483_74#_c_1113_n 0.0233055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_483_74#_c_1114_n 0.0026414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1217_n 0.00886652f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_67 VNB N_VGND_c_1218_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.79
cc_68 VNB N_VGND_c_1219_n 0.00269659f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=2.4
cc_69 VNB N_VGND_c_1220_n 0.00333063f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.79
cc_70 VNB N_VGND_c_1221_n 0.156139f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_71 VNB N_VGND_c_1222_n 0.0156795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1223_n 0.0156795f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.515
cc_73 VNB N_VGND_c_1224_n 0.0161665f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.515
cc_74 VNB N_VGND_c_1225_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_75 VNB N_VGND_c_1226_n 0.523727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1227_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1228_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1229_n 0.00619876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1230_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VPB N_C1_M1013_g 0.0246442f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_81 VPB N_C1_M1014_g 0.0214289f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_82 VPB N_C1_M1024_g 0.0214468f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=2.4
cc_83 VPB N_C1_M1035_g 0.0218077f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_84 VPB N_C1_c_151_n 0.0152619f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=1.515
cc_85 VPB N_C1_c_152_n 0.015808f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.515
cc_86 VPB N_B1_M1003_g 0.0216803f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_87 VPB N_B1_M1020_g 0.0210122f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.79
cc_88 VPB N_B1_M1022_g 0.0206593f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.79
cc_89 VPB N_B1_M1028_g 0.0214186f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.68
cc_90 VPB N_B1_c_243_n 0.00897985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_B1_c_235_n 6.0265e-19 $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.515
cc_92 VPB N_B1_c_236_n 0.0111879f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.515
cc_93 VPB N_B1_c_237_n 0.0056017f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_94 VPB N_B1_c_238_n 0.00271992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_B2_c_366_n 0.0170979f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.68
cc_96 VPB N_B2_c_367_n 0.0170611f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.79
cc_97 VPB N_B2_M1032_g 0.0210656f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_98 VPB N_B2_c_362_n 0.00911485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_B2_M1036_g 0.0217462f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=2.4
cc_100 VPB N_A1_M1001_g 0.0245657f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.79
cc_101 VPB N_A1_M1010_g 0.0211602f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_102 VPB N_A1_M1038_g 0.0214394f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.79
cc_103 VPB N_A1_M1039_g 0.0259175f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.79
cc_104 VPB A1 0.015855f $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.515
cc_105 VPB N_A1_c_455_n 0.00293155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A2_M1021_g 0.0209767f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.79
cc_107 VPB N_A2_M1023_g 0.0196385f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_108 VPB N_A2_M1029_g 0.0196385f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.79
cc_109 VPB N_A2_M1033_g 0.0201709f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.79
cc_110 VPB A2 0.00731208f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_111 VPB N_A2_c_568_n 0.0116455f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.515
cc_112 VPB N_VPWR_c_649_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=2.4
cc_113 VPB N_VPWR_c_650_n 0.0498587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_651_n 0.00898286f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_115 VPB N_VPWR_c_652_n 0.00506286f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_116 VPB N_VPWR_c_653_n 0.00858545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_654_n 0.00885887f $X=-0.19 $Y=1.66 $X2=0.9 $Y2=1.515
cc_118 VPB N_VPWR_c_655_n 0.00554449f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=1.515
cc_119 VPB N_VPWR_c_656_n 0.0107598f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=1.515
cc_120 VPB N_VPWR_c_657_n 0.0495391f $X=-0.19 $Y=1.66 $X2=1.49 $Y2=1.515
cc_121 VPB N_VPWR_c_658_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_122 VPB N_VPWR_c_659_n 0.0178177f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=1.565
cc_123 VPB N_VPWR_c_660_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_661_n 0.0599347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_662_n 0.0580859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_663_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_664_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_665_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_666_n 0.00631813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_667_n 0.00631418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_668_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_648_n 0.0879003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_Y_c_780_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_134 VPB N_Y_c_781_n 0.00225649f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.515
cc_135 VPB N_Y_c_782_n 0.00221543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_Y_c_779_n 0.00130166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_511_368#_c_915_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.79
cc_138 VPB N_A_511_368#_c_916_n 0.00196576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_511_368#_c_917_n 0.00458349f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.35
cc_140 VPB N_A_511_368#_c_918_n 0.0023101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_511_368#_c_919_n 0.00196576f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_142 VPB N_A_1291_368#_c_979_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_143 VPB N_A_1291_368#_c_980_n 0.00473643f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.79
cc_144 VPB N_A_1291_368#_c_981_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.68
cc_145 VPB N_A_1291_368#_c_982_n 0.00220034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_1291_368#_c_983_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_147 N_C1_M1035_g N_B1_M1003_g 0.017418f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_148 N_C1_c_152_n N_B1_c_249_n 0.00258062f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_149 N_C1_c_152_n N_B1_c_236_n 0.0219622f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_150 N_C1_M1013_g N_VPWR_c_650_n 0.00501904f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_151 N_C1_c_151_n N_VPWR_c_650_n 0.0208754f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_152 N_C1_M1014_g N_VPWR_c_651_n 0.00341061f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_153 N_C1_M1024_g N_VPWR_c_651_n 0.00202538f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_154 N_C1_M1024_g N_VPWR_c_652_n 5.27444e-19 $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_155 N_C1_M1035_g N_VPWR_c_652_n 0.0117033f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_156 N_C1_M1013_g N_VPWR_c_658_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_157 N_C1_M1014_g N_VPWR_c_658_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_158 N_C1_M1024_g N_VPWR_c_659_n 0.00549225f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_159 N_C1_M1035_g N_VPWR_c_659_n 0.00460063f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_160 N_C1_M1013_g N_VPWR_c_648_n 0.00986008f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_161 N_C1_M1014_g N_VPWR_c_648_n 0.00982397f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_162 N_C1_M1024_g N_VPWR_c_648_n 0.0107024f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_163 N_C1_M1035_g N_VPWR_c_648_n 0.00908804f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_164 N_C1_M1000_g N_Y_c_784_n 0.00473639f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_165 N_C1_M1002_g N_Y_c_784_n 0.00575058f $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_166 N_C1_M1004_g N_Y_c_784_n 5.36571e-19 $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_167 N_C1_M1013_g N_Y_c_787_n 0.0025567f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_168 N_C1_M1014_g N_Y_c_787_n 8.84614e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_169 N_C1_c_151_n N_Y_c_787_n 0.0235495f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_170 N_C1_c_152_n N_Y_c_787_n 5.53716e-19 $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_171 N_C1_M1013_g N_Y_c_780_n 0.0112644f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_172 N_C1_M1014_g N_Y_c_780_n 0.0117613f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_173 N_C1_M1024_g N_Y_c_780_n 8.62186e-19 $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_174 N_C1_M1002_g N_Y_c_776_n 0.00900535f $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_175 N_C1_M1004_g N_Y_c_776_n 0.00900535f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_176 N_C1_c_151_n N_Y_c_776_n 0.039654f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_177 N_C1_c_152_n N_Y_c_776_n 0.00241935f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_178 N_C1_M1000_g N_Y_c_777_n 0.0023927f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_179 N_C1_M1002_g N_Y_c_777_n 9.58661e-19 $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_180 N_C1_c_151_n N_Y_c_777_n 0.0277843f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_181 N_C1_c_152_n N_Y_c_777_n 0.00241407f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_182 N_C1_M1014_g N_Y_c_802_n 0.013412f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_183 N_C1_M1024_g N_Y_c_802_n 0.0212056f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_184 N_C1_c_151_n N_Y_c_802_n 0.0354114f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_185 N_C1_c_152_n N_Y_c_802_n 9.45805e-19 $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_186 N_C1_M1002_g N_Y_c_806_n 5.3642e-19 $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_187 N_C1_M1004_g N_Y_c_806_n 0.00575058f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_188 N_C1_M1018_g N_Y_c_806_n 0.0051579f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_189 N_C1_M1024_g N_Y_c_781_n 0.00843542f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_190 N_C1_M1035_g N_Y_c_781_n 2.76437e-19 $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_191 N_C1_M1035_g N_Y_c_811_n 0.0196821f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_192 N_C1_M1004_g N_Y_c_778_n 0.00183768f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_193 N_C1_M1018_g N_Y_c_778_n 0.0021587f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_194 N_C1_c_152_n N_Y_c_778_n 0.00259964f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_195 N_C1_M1014_g N_Y_c_782_n 9.08817e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_196 N_C1_M1024_g N_Y_c_782_n 0.00516064f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_197 N_C1_M1035_g N_Y_c_782_n 5.03246e-19 $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_198 N_C1_c_152_n N_Y_c_782_n 0.00199936f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_199 N_C1_M1014_g N_Y_c_779_n 8.222e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_200 N_C1_M1004_g N_Y_c_779_n 0.00360365f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_201 N_C1_M1024_g N_Y_c_779_n 0.00312689f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_202 N_C1_M1018_g N_Y_c_779_n 0.00809756f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_203 N_C1_M1035_g N_Y_c_779_n 0.00306551f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_204 N_C1_c_151_n N_Y_c_779_n 0.0325268f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_205 N_C1_c_152_n N_Y_c_779_n 0.0187585f $X=1.785 $Y=1.515 $X2=0 $Y2=0
cc_206 N_C1_M1000_g N_A_27_84#_c_1027_n 0.00160853f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_207 N_C1_c_151_n N_A_27_84#_c_1027_n 0.0224519f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_208 N_C1_M1000_g N_A_27_84#_c_1028_n 0.0141481f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_209 N_C1_M1002_g N_A_27_84#_c_1028_n 0.0109808f $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_210 N_C1_M1004_g N_A_27_84#_c_1030_n 0.0109808f $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_211 N_C1_M1018_g N_A_27_84#_c_1030_n 0.0138423f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_212 N_C1_M1018_g N_A_27_84#_c_1033_n 0.00141527f $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_213 N_C1_c_152_n N_A_27_84#_c_1033_n 0.00559349f $X=1.785 $Y=1.515 $X2=0
+ $Y2=0
cc_214 N_C1_M1018_g N_A_483_74#_c_1107_n 3.01901e-19 $X=1.785 $Y=0.79 $X2=0
+ $Y2=0
cc_215 N_C1_M1000_g N_VGND_c_1221_n 8.76084e-19 $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_216 N_C1_M1002_g N_VGND_c_1221_n 8.76084e-19 $X=0.925 $Y=0.79 $X2=0 $Y2=0
cc_217 N_C1_M1004_g N_VGND_c_1221_n 8.76084e-19 $X=1.355 $Y=0.79 $X2=0 $Y2=0
cc_218 N_C1_M1018_g N_VGND_c_1221_n 8.76084e-19 $X=1.785 $Y=0.79 $X2=0 $Y2=0
cc_219 N_B1_M1022_g N_B2_c_366_n 0.0204691f $X=3.465 $Y=2.4 $X2=-0.19 $Y2=-0.245
cc_220 N_B1_c_243_n N_B2_c_366_n 0.008563f $X=5.405 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_221 N_B1_c_233_n N_B2_c_358_n 0.0179023f $X=3.635 $Y=1.185 $X2=0 $Y2=0
cc_222 N_B1_c_243_n N_B2_c_367_n 0.00859825f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_223 N_B1_c_243_n N_B2_M1032_g 0.0119597f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_224 N_B1_c_243_n N_B2_c_362_n 0.0234439f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_225 N_B1_c_235_n N_B2_c_362_n 0.00219148f $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_226 N_B1_c_236_n N_B2_c_362_n 0.0448508f $X=3.465 $Y=1.432 $X2=0 $Y2=0
cc_227 N_B1_c_237_n N_B2_c_362_n 0.0110451f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_228 N_B1_c_238_n N_B2_c_362_n 0.00710875f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_229 N_B1_M1028_g N_B2_M1036_g 0.0292422f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_230 N_B1_c_243_n N_B2_M1036_g 0.0155118f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_231 N_B1_c_237_n N_B2_M1036_g 0.00565698f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B1_c_238_n N_B2_M1036_g 0.00762987f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_233 N_B1_M1037_g N_B2_c_364_n 0.0347442f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B1_M1037_g B2 5.14568e-19 $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B1_c_243_n B2 0.0747366f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_236 N_B1_c_235_n B2 0.00532239f $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_237 N_B1_c_236_n B2 8.13044e-19 $X=3.465 $Y=1.432 $X2=0 $Y2=0
cc_238 N_B1_c_238_n B2 0.0132957f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_239 N_B1_M1037_g N_A1_M1008_g 0.0237178f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1028_g N_A1_M1001_g 0.0234927f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B1_c_237_n N_A1_M1001_g 0.00439601f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_242 N_B1_c_238_n N_A1_M1001_g 0.00543157f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_243 N_B1_M1037_g N_A1_c_450_n 5.32822e-19 $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B1_c_237_n N_A1_c_450_n 8.36735e-19 $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_245 N_B1_c_238_n N_A1_c_450_n 0.0161127f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_246 N_B1_c_237_n N_A1_c_451_n 0.0150967f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_247 N_B1_c_238_n N_A1_c_451_n 3.00906e-19 $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_248 N_B1_c_249_n N_VPWR_M1020_d 0.00250498f $X=3.29 $Y=1.615 $X2=0 $Y2=0
cc_249 N_B1_c_235_n N_VPWR_M1020_d 3.08984e-19 $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_250 N_B1_c_238_n N_VPWR_M1028_d 9.92712e-19 $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_251 N_B1_M1003_g N_VPWR_c_652_n 0.00194999f $X=2.465 $Y=2.4 $X2=0 $Y2=0
cc_252 N_B1_M1020_g N_VPWR_c_653_n 0.00203999f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_253 N_B1_M1022_g N_VPWR_c_653_n 0.00150551f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_254 N_B1_M1028_g N_VPWR_c_654_n 0.00150551f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_255 N_B1_M1003_g N_VPWR_c_660_n 0.005209f $X=2.465 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B1_M1020_g N_VPWR_c_660_n 0.005209f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B1_M1022_g N_VPWR_c_661_n 0.00517089f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B1_M1028_g N_VPWR_c_661_n 0.00517089f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_259 N_B1_M1003_g N_VPWR_c_648_n 0.0098216f $X=2.465 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B1_M1020_g N_VPWR_c_648_n 0.00515684f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B1_M1022_g N_VPWR_c_648_n 0.00515622f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B1_M1028_g N_VPWR_c_648_n 0.00978354f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_263 N_B1_c_243_n N_Y_M1005_s 0.00165831f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_264 N_B1_c_243_n N_Y_M1032_s 0.00218982f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_265 N_B1_M1003_g N_Y_c_811_n 0.0216828f $X=2.465 $Y=2.4 $X2=0 $Y2=0
cc_266 N_B1_M1020_g N_Y_c_811_n 0.0122174f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_267 N_B1_M1022_g N_Y_c_811_n 0.0121787f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_268 N_B1_c_249_n N_Y_c_811_n 0.0836148f $X=3.29 $Y=1.615 $X2=0 $Y2=0
cc_269 N_B1_c_236_n N_Y_c_811_n 0.00122287f $X=3.465 $Y=1.432 $X2=0 $Y2=0
cc_270 N_B1_c_243_n N_Y_c_833_n 0.0356639f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_271 N_B1_M1028_g N_Y_c_834_n 5.42618e-19 $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_272 N_B1_M1028_g N_Y_c_835_n 0.0170123f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_273 N_B1_c_243_n N_Y_c_835_n 0.0101332f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_274 N_B1_c_237_n N_Y_c_835_n 3.2897e-19 $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_275 N_B1_c_238_n N_Y_c_835_n 0.0328037f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_276 N_B1_c_236_n N_Y_c_779_n 0.00163472f $X=3.465 $Y=1.432 $X2=0 $Y2=0
cc_277 N_B1_c_243_n N_Y_c_840_n 0.0126995f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_278 N_B1_c_243_n N_Y_c_841_n 0.0190144f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_279 N_B1_c_249_n N_A_511_368#_M1003_s 0.00172148f $X=3.29 $Y=1.615 $X2=-0.19
+ $Y2=-0.245
cc_280 N_B1_c_243_n N_A_511_368#_M1022_s 0.00166235f $X=5.405 $Y=1.795 $X2=0
+ $Y2=0
cc_281 N_B1_c_243_n N_A_511_368#_M1025_d 0.00166235f $X=5.405 $Y=1.795 $X2=0
+ $Y2=0
cc_282 N_B1_c_238_n N_A_511_368#_M1036_d 0.00226794f $X=5.835 $Y=1.515 $X2=0
+ $Y2=0
cc_283 N_B1_M1020_g N_A_511_368#_c_924_n 0.0100971f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_284 N_B1_M1022_g N_A_511_368#_c_924_n 0.0100971f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_285 N_B1_M1022_g N_A_511_368#_c_926_n 8.84747e-19 $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_286 N_B1_M1020_g N_A_511_368#_c_927_n 3.0069e-19 $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_287 N_B1_M1022_g N_A_511_368#_c_927_n 0.00555833f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_288 N_B1_M1022_g N_A_511_368#_c_916_n 0.00338824f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_289 N_B1_M1028_g N_A_511_368#_c_917_n 0.00357739f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_290 N_B1_M1028_g N_A_511_368#_c_931_n 0.00623735f $X=5.815 $Y=2.4 $X2=0 $Y2=0
cc_291 N_B1_M1003_g N_A_511_368#_c_918_n 0.00755618f $X=2.465 $Y=2.4 $X2=0 $Y2=0
cc_292 N_B1_M1020_g N_A_511_368#_c_918_n 0.0077957f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_293 N_B1_M1022_g N_A_511_368#_c_918_n 3.16734e-19 $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_294 N_B1_M1009_g N_A_27_84#_c_1030_n 0.00288917f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_295 N_B1_M1009_g N_A_27_84#_c_1031_n 0.00289242f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_296 N_B1_M1009_g N_A_27_84#_c_1032_n 0.0206145f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_c_249_n N_A_27_84#_c_1032_n 0.040357f $X=3.29 $Y=1.615 $X2=0 $Y2=0
cc_298 N_B1_c_236_n N_A_27_84#_c_1032_n 0.0143454f $X=3.465 $Y=1.432 $X2=0 $Y2=0
cc_299 N_B1_c_232_n N_A_27_84#_c_1034_n 0.00841735f $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_300 N_B1_c_233_n N_A_27_84#_c_1034_n 0.00950816f $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_301 N_B1_c_243_n N_A_27_84#_c_1034_n 0.00395856f $X=5.405 $Y=1.795 $X2=0
+ $Y2=0
cc_302 N_B1_c_236_n N_A_27_84#_c_1034_n 0.00320458f $X=3.465 $Y=1.432 $X2=0
+ $Y2=0
cc_303 N_B1_c_232_n N_A_27_84#_c_1036_n 0.00558702f $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_304 N_B1_c_233_n N_A_27_84#_c_1036_n 5.18778e-19 $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_305 N_B1_c_235_n N_A_27_84#_c_1036_n 0.040357f $X=3.555 $Y=1.615 $X2=0 $Y2=0
cc_306 N_B1_c_232_n N_A_27_84#_c_1037_n 6.02585e-19 $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_307 N_B1_c_233_n N_A_27_84#_c_1037_n 0.00612157f $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_308 N_B1_c_243_n N_A_27_84#_c_1037_n 0.0111311f $X=5.405 $Y=1.795 $X2=0 $Y2=0
cc_309 N_B1_M1037_g N_A_27_84#_c_1061_n 0.00364331f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B1_c_238_n N_A_27_84#_c_1061_n 0.0149317f $X=5.835 $Y=1.515 $X2=0 $Y2=0
cc_311 N_B1_M1009_g N_A_483_74#_c_1107_n 0.0102979f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_312 N_B1_c_232_n N_A_483_74#_c_1107_n 0.0113119f $X=3.205 $Y=1.185 $X2=0
+ $Y2=0
cc_313 N_B1_c_233_n N_A_483_74#_c_1108_n 0.0112282f $X=3.635 $Y=1.185 $X2=0
+ $Y2=0
cc_314 N_B1_M1037_g N_A_483_74#_c_1108_n 0.0154814f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_315 N_B1_M1037_g N_A_483_74#_c_1114_n 6.56207e-19 $X=5.785 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_B1_c_237_n N_A_483_74#_c_1114_n 6.57592e-19 $X=5.835 $Y=1.515 $X2=0
+ $Y2=0
cc_317 N_B1_c_238_n N_A_483_74#_c_1114_n 0.00538446f $X=5.835 $Y=1.515 $X2=0
+ $Y2=0
cc_318 N_B1_M1009_g N_VGND_c_1221_n 0.00291649f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_319 N_B1_c_232_n N_VGND_c_1221_n 0.00291649f $X=3.205 $Y=1.185 $X2=0 $Y2=0
cc_320 N_B1_c_233_n N_VGND_c_1221_n 0.00291649f $X=3.635 $Y=1.185 $X2=0 $Y2=0
cc_321 N_B1_M1037_g N_VGND_c_1221_n 0.00291649f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_322 N_B1_M1009_g N_VGND_c_1226_n 0.0036412f $X=2.775 $Y=0.74 $X2=0 $Y2=0
cc_323 N_B1_c_232_n N_VGND_c_1226_n 0.00359121f $X=3.205 $Y=1.185 $X2=0 $Y2=0
cc_324 N_B1_c_233_n N_VGND_c_1226_n 0.00359219f $X=3.635 $Y=1.185 $X2=0 $Y2=0
cc_325 N_B1_M1037_g N_VGND_c_1226_n 0.0035993f $X=5.785 $Y=0.74 $X2=0 $Y2=0
cc_326 N_B2_c_366_n N_VPWR_c_661_n 0.00333896f $X=3.915 $Y=1.725 $X2=0 $Y2=0
cc_327 N_B2_c_367_n N_VPWR_c_661_n 0.00333896f $X=4.365 $Y=1.725 $X2=0 $Y2=0
cc_328 N_B2_M1032_g N_VPWR_c_661_n 0.00333896f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_329 N_B2_M1036_g N_VPWR_c_661_n 0.00333926f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_330 N_B2_c_366_n N_VPWR_c_648_n 0.00422796f $X=3.915 $Y=1.725 $X2=0 $Y2=0
cc_331 N_B2_c_367_n N_VPWR_c_648_n 0.00422685f $X=4.365 $Y=1.725 $X2=0 $Y2=0
cc_332 N_B2_M1032_g N_VPWR_c_648_n 0.00423173f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_333 N_B2_M1036_g N_VPWR_c_648_n 0.00423742f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_334 N_B2_c_366_n N_Y_c_811_n 0.0141869f $X=3.915 $Y=1.725 $X2=0 $Y2=0
cc_335 N_B2_c_367_n N_Y_c_833_n 0.0142562f $X=4.365 $Y=1.725 $X2=0 $Y2=0
cc_336 N_B2_M1032_g N_Y_c_833_n 0.0142562f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_337 N_B2_M1036_g N_Y_c_834_n 0.00815121f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_338 N_B2_M1036_g N_Y_c_835_n 0.0131783f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_339 N_B2_c_362_n N_Y_c_840_n 4.84876e-19 $X=5.315 $Y=1.55 $X2=0 $Y2=0
cc_340 N_B2_M1036_g N_Y_c_841_n 8.70246e-19 $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_341 N_B2_c_366_n N_A_511_368#_c_926_n 0.00244711f $X=3.915 $Y=1.725 $X2=0
+ $Y2=0
cc_342 N_B2_c_366_n N_A_511_368#_c_927_n 0.00530339f $X=3.915 $Y=1.725 $X2=0
+ $Y2=0
cc_343 N_B2_c_367_n N_A_511_368#_c_927_n 4.87357e-19 $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_344 N_B2_c_366_n N_A_511_368#_c_915_n 0.0116345f $X=3.915 $Y=1.725 $X2=0
+ $Y2=0
cc_345 N_B2_c_367_n N_A_511_368#_c_915_n 0.0116345f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_346 N_B2_c_366_n N_A_511_368#_c_916_n 0.001916f $X=3.915 $Y=1.725 $X2=0 $Y2=0
cc_347 N_B2_c_366_n N_A_511_368#_c_941_n 5.41427e-19 $X=3.915 $Y=1.725 $X2=0
+ $Y2=0
cc_348 N_B2_c_367_n N_A_511_368#_c_941_n 0.00773996f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_349 N_B2_M1032_g N_A_511_368#_c_941_n 0.00782866f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_350 N_B2_M1036_g N_A_511_368#_c_941_n 4.54422e-19 $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_351 N_B2_M1032_g N_A_511_368#_c_917_n 0.0119307f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_352 N_B2_M1036_g N_A_511_368#_c_917_n 0.0144846f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_353 N_B2_c_367_n N_A_511_368#_c_919_n 0.00193733f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_354 N_B2_M1032_g N_A_511_368#_c_919_n 0.00193733f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_355 N_B2_c_358_n N_A_27_84#_c_1037_n 0.00612289f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_356 N_B2_c_359_n N_A_27_84#_c_1037_n 9.42328e-19 $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_357 N_B2_c_362_n N_A_27_84#_c_1037_n 0.00394764f $X=5.315 $Y=1.55 $X2=0 $Y2=0
cc_358 N_B2_c_364_n N_A_27_84#_c_1061_n 0.00202711f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_359 N_B2_c_358_n N_A_27_84#_c_1067_n 0.0138321f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_360 N_B2_c_359_n N_A_27_84#_c_1067_n 0.0103131f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_361 N_B2_c_361_n N_A_27_84#_c_1067_n 0.0103131f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_362 N_B2_c_362_n N_A_27_84#_c_1067_n 0.00192366f $X=5.315 $Y=1.55 $X2=0 $Y2=0
cc_363 N_B2_c_364_n N_A_27_84#_c_1067_n 0.0130444f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_364 B2 N_A_27_84#_c_1067_n 0.0699825f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_365 N_B2_c_358_n N_A_483_74#_c_1108_n 0.0101343f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_366 N_B2_c_359_n N_A_483_74#_c_1108_n 0.010218f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_367 N_B2_c_361_n N_A_483_74#_c_1108_n 0.010218f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_368 N_B2_c_364_n N_A_483_74#_c_1108_n 0.0101492f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_369 N_B2_c_358_n N_VGND_c_1221_n 0.00291649f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_370 N_B2_c_359_n N_VGND_c_1221_n 0.00291649f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_371 N_B2_c_361_n N_VGND_c_1221_n 0.00291649f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_372 N_B2_c_364_n N_VGND_c_1221_n 0.00291649f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_373 N_B2_c_358_n N_VGND_c_1226_n 0.00358272f $X=4.065 $Y=1.22 $X2=0 $Y2=0
cc_374 N_B2_c_359_n N_VGND_c_1226_n 0.00359121f $X=4.495 $Y=1.22 $X2=0 $Y2=0
cc_375 N_B2_c_361_n N_VGND_c_1226_n 0.00359121f $X=4.925 $Y=1.22 $X2=0 $Y2=0
cc_376 N_B2_c_364_n N_VGND_c_1226_n 0.00359219f $X=5.355 $Y=1.22 $X2=0 $Y2=0
cc_377 N_A1_M1008_g N_A2_M1007_g 0.0240526f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A1_c_450_n N_A2_M1007_g 0.00517694f $X=6.575 $Y=1.175 $X2=0 $Y2=0
cc_379 N_A1_c_451_n N_A2_M1007_g 0.0179795f $X=6.375 $Y=1.425 $X2=0 $Y2=0
cc_380 N_A1_c_454_n N_A2_M1007_g 0.0128792f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_381 N_A1_c_454_n N_A2_M1012_g 0.0108858f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_382 N_A1_c_454_n N_A2_M1017_g 0.0108382f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_383 N_A1_c_455_n N_A2_M1017_g 4.14448e-19 $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_384 N_A1_M1010_g N_A2_M1033_g 0.0125152f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_385 N_A1_c_455_n N_A2_M1033_g 0.00366435f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_386 N_A1_M1027_g N_A2_M1019_g 0.0206073f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A1_c_454_n N_A2_M1019_g 0.0104992f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_388 N_A1_c_455_n N_A2_M1019_g 0.00421415f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_389 N_A1_M1001_g A2 0.00101517f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_390 N_A1_c_450_n A2 0.00953035f $X=6.575 $Y=1.175 $X2=0 $Y2=0
cc_391 N_A1_c_454_n A2 0.0884035f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_392 N_A1_c_455_n A2 0.0220095f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_393 N_A1_M1001_g N_A2_c_568_n 0.0458106f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_394 N_A1_c_453_n N_A2_c_568_n 0.0331225f $X=9.585 $Y=1.425 $X2=0 $Y2=0
cc_395 N_A1_c_454_n N_A2_c_568_n 0.00988025f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_396 N_A1_c_455_n N_A2_c_568_n 0.0134688f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_397 N_A1_M1001_g N_VPWR_c_654_n 0.00150551f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A1_M1010_g N_VPWR_c_655_n 0.0117336f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_399 N_A1_M1038_g N_VPWR_c_655_n 0.002979f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_400 N_A1_M1039_g N_VPWR_c_657_n 0.00501904f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_401 A1 N_VPWR_c_657_n 0.0216354f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_402 N_A1_M1001_g N_VPWR_c_662_n 0.00517089f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_403 N_A1_M1010_g N_VPWR_c_662_n 0.00460063f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_404 N_A1_M1038_g N_VPWR_c_663_n 0.005209f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_405 N_A1_M1039_g N_VPWR_c_663_n 0.005209f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A1_M1001_g N_VPWR_c_648_n 0.00978398f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_407 N_A1_M1010_g N_VPWR_c_648_n 0.00908665f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_408 N_A1_M1038_g N_VPWR_c_648_n 0.00982266f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_409 N_A1_M1039_g N_VPWR_c_648_n 0.00986025f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_410 N_A1_M1001_g N_Y_c_835_n 0.0190785f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A1_c_450_n N_Y_c_835_n 0.010431f $X=6.575 $Y=1.175 $X2=0 $Y2=0
cc_412 N_A1_c_451_n N_Y_c_835_n 4.77286e-19 $X=6.375 $Y=1.425 $X2=0 $Y2=0
cc_413 N_A1_M1001_g Y 0.00225758f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A1_M1010_g N_A_1291_368#_c_980_n 0.00101073f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_415 N_A1_c_455_n N_A_1291_368#_c_985_n 0.0147553f $X=8.455 $Y=1.435 $X2=0
+ $Y2=0
cc_416 N_A1_M1010_g N_A_1291_368#_c_986_n 0.0142562f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_417 N_A1_M1038_g N_A_1291_368#_c_986_n 0.0128923f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_418 A1 N_A_1291_368#_c_986_n 0.0443262f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_419 N_A1_c_453_n N_A_1291_368#_c_986_n 4.05102e-19 $X=9.585 $Y=1.425 $X2=0
+ $Y2=0
cc_420 N_A1_M1038_g N_A_1291_368#_c_990_n 8.84614e-19 $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_421 N_A1_M1039_g N_A_1291_368#_c_990_n 0.0025567f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_422 A1 N_A_1291_368#_c_990_n 0.0239609f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_423 N_A1_c_453_n N_A_1291_368#_c_990_n 4.57942e-19 $X=9.585 $Y=1.425 $X2=0
+ $Y2=0
cc_424 N_A1_M1010_g N_A_1291_368#_c_981_n 6.74232e-19 $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_425 N_A1_M1038_g N_A_1291_368#_c_981_n 0.0121366f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_426 N_A1_M1039_g N_A_1291_368#_c_981_n 0.0112644f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_427 N_A1_M1001_g N_A_1291_368#_c_982_n 0.0071932f $X=6.365 $Y=2.4 $X2=0 $Y2=0
cc_428 N_A1_c_454_n N_A_483_74#_M1007_s 0.00176461f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_429 N_A1_c_454_n N_A_483_74#_M1017_s 0.00176461f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_430 N_A1_M1008_g N_A_483_74#_c_1129_n 0.0107566f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A1_c_450_n N_A_483_74#_c_1129_n 0.0186469f $X=6.575 $Y=1.175 $X2=0
+ $Y2=0
cc_432 N_A1_c_451_n N_A_483_74#_c_1129_n 6.09656e-19 $X=6.375 $Y=1.425 $X2=0
+ $Y2=0
cc_433 N_A1_c_454_n N_A_483_74#_c_1129_n 0.0195621f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_434 N_A1_M1008_g N_A_483_74#_c_1109_n 5.78282e-19 $X=6.285 $Y=0.74 $X2=0
+ $Y2=0
cc_435 N_A1_c_454_n N_A_483_74#_c_1134_n 0.0357472f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_436 N_A1_M1027_g N_A_483_74#_c_1135_n 0.0118367f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_437 A1 N_A_483_74#_c_1135_n 0.0123244f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_438 N_A1_c_454_n N_A_483_74#_c_1135_n 0.019324f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_439 N_A1_M1027_g N_A_483_74#_c_1111_n 0.00214936f $X=8.655 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A1_M1031_g N_A_483_74#_c_1111_n 2.6509e-19 $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_441 N_A1_M1031_g N_A_483_74#_c_1112_n 0.0122595f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_442 N_A1_M1034_g N_A_483_74#_c_1112_n 0.0122129f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_443 A1 N_A_483_74#_c_1112_n 0.0655704f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_444 N_A1_c_453_n N_A_483_74#_c_1112_n 0.00236025f $X=9.585 $Y=1.425 $X2=0
+ $Y2=0
cc_445 N_A1_M1034_g N_A_483_74#_c_1113_n 8.26992e-19 $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_446 N_A1_M1008_g N_A_483_74#_c_1114_n 0.0112264f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_447 N_A1_c_450_n N_A_483_74#_c_1114_n 0.00188346f $X=6.575 $Y=1.175 $X2=0
+ $Y2=0
cc_448 N_A1_c_454_n N_A_483_74#_c_1147_n 0.0151907f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_449 N_A1_c_454_n N_A_483_74#_c_1148_n 0.0151907f $X=8.285 $Y=1.435 $X2=0
+ $Y2=0
cc_450 A1 N_A_483_74#_c_1149_n 0.0206148f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_451 N_A1_c_453_n N_A_483_74#_c_1149_n 0.0042758f $X=9.585 $Y=1.425 $X2=0
+ $Y2=0
cc_452 N_A1_c_450_n N_VGND_M1008_s 0.0017364f $X=6.575 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_453 N_A1_c_454_n N_VGND_M1008_s 0.00158921f $X=8.285 $Y=1.435 $X2=-0.19
+ $Y2=-0.245
cc_454 N_A1_c_454_n N_VGND_M1012_d 0.00251484f $X=8.285 $Y=1.435 $X2=0 $Y2=0
cc_455 N_A1_c_455_n N_VGND_M1019_d 0.00145497f $X=8.455 $Y=1.435 $X2=0 $Y2=0
cc_456 N_A1_M1008_g N_VGND_c_1217_n 0.00464693f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_457 N_A1_M1027_g N_VGND_c_1219_n 0.00679571f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A1_M1031_g N_VGND_c_1219_n 3.92591e-19 $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A1_M1027_g N_VGND_c_1220_n 4.37937e-19 $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_460 N_A1_M1031_g N_VGND_c_1220_n 0.00869262f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_461 N_A1_M1034_g N_VGND_c_1220_n 0.0114756f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A1_M1008_g N_VGND_c_1221_n 0.00331438f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A1_M1027_g N_VGND_c_1224_n 0.00281141f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_464 N_A1_M1031_g N_VGND_c_1224_n 0.00383152f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_465 N_A1_M1034_g N_VGND_c_1225_n 0.00383152f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_466 N_A1_M1008_g N_VGND_c_1226_n 0.0042805f $X=6.285 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A1_M1027_g N_VGND_c_1226_n 0.00365724f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_468 N_A1_M1031_g N_VGND_c_1226_n 0.00758198f $X=9.155 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A1_M1034_g N_VGND_c_1226_n 0.00761198f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A2_M1021_g N_VPWR_c_662_n 0.00333926f $X=6.87 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A2_M1023_g N_VPWR_c_662_n 0.00333926f $X=7.32 $Y=2.4 $X2=0 $Y2=0
cc_472 N_A2_M1029_g N_VPWR_c_662_n 0.00333926f $X=7.77 $Y=2.4 $X2=0 $Y2=0
cc_473 N_A2_M1033_g N_VPWR_c_662_n 0.00333926f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_474 N_A2_M1021_g N_VPWR_c_648_n 0.00423297f $X=6.87 $Y=2.4 $X2=0 $Y2=0
cc_475 N_A2_M1023_g N_VPWR_c_648_n 0.00422687f $X=7.32 $Y=2.4 $X2=0 $Y2=0
cc_476 N_A2_M1029_g N_VPWR_c_648_n 0.00422687f $X=7.77 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A2_M1033_g N_VPWR_c_648_n 0.00422798f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_478 N_A2_M1021_g N_Y_c_835_n 0.00889187f $X=6.87 $Y=2.4 $X2=0 $Y2=0
cc_479 N_A2_M1023_g N_Y_c_854_n 0.012931f $X=7.32 $Y=2.4 $X2=0 $Y2=0
cc_480 N_A2_M1029_g N_Y_c_854_n 0.012931f $X=7.77 $Y=2.4 $X2=0 $Y2=0
cc_481 A2 N_Y_c_854_n 0.0384651f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_482 N_A2_c_568_n N_Y_c_854_n 4.90767e-19 $X=8.215 $Y=1.515 $X2=0 $Y2=0
cc_483 N_A2_M1023_g N_Y_c_858_n 5.72851e-19 $X=7.32 $Y=2.4 $X2=0 $Y2=0
cc_484 N_A2_M1029_g N_Y_c_858_n 0.0105614f $X=7.77 $Y=2.4 $X2=0 $Y2=0
cc_485 N_A2_M1033_g N_Y_c_858_n 0.0119589f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_486 A2 N_Y_c_858_n 0.0150408f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A2_c_568_n N_Y_c_858_n 7.23585e-19 $X=8.215 $Y=1.515 $X2=0 $Y2=0
cc_488 N_A2_M1021_g Y 0.021025f $X=6.87 $Y=2.4 $X2=0 $Y2=0
cc_489 N_A2_M1023_g Y 0.0106272f $X=7.32 $Y=2.4 $X2=0 $Y2=0
cc_490 N_A2_M1029_g Y 5.71911e-19 $X=7.77 $Y=2.4 $X2=0 $Y2=0
cc_491 A2 Y 0.0298358f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_492 N_A2_c_568_n Y 5.53363e-19 $X=8.215 $Y=1.515 $X2=0 $Y2=0
cc_493 N_A2_M1021_g N_A_1291_368#_c_979_n 0.0122346f $X=6.87 $Y=2.4 $X2=0 $Y2=0
cc_494 N_A2_M1023_g N_A_1291_368#_c_979_n 0.0139915f $X=7.32 $Y=2.4 $X2=0 $Y2=0
cc_495 N_A2_M1029_g N_A_1291_368#_c_980_n 0.0139834f $X=7.77 $Y=2.4 $X2=0 $Y2=0
cc_496 N_A2_M1033_g N_A_1291_368#_c_980_n 0.0137017f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_497 N_A2_M1007_g N_A_483_74#_c_1129_n 0.00941575f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A2_M1007_g N_A_483_74#_c_1109_n 0.00687331f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A2_M1012_g N_A_483_74#_c_1109_n 4.39567e-19 $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A2_M1012_g N_A_483_74#_c_1134_n 0.0113092f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A2_M1017_g N_A_483_74#_c_1134_n 0.00916065f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_A2_M1012_g N_A_483_74#_c_1110_n 6.09957e-19 $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_503 N_A2_M1017_g N_A_483_74#_c_1110_n 0.00657942f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_504 N_A2_M1019_g N_A_483_74#_c_1110_n 4.39567e-19 $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A2_M1019_g N_A_483_74#_c_1135_n 0.0109279f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_506 N_A2_M1007_g N_A_483_74#_c_1114_n 0.00144055f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A2_M1007_g N_A_483_74#_c_1147_n 0.00181289f $X=6.855 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A2_M1017_g N_A_483_74#_c_1148_n 0.00181289f $X=7.785 $Y=0.74 $X2=0
+ $Y2=0
cc_509 N_A2_M1007_g N_VGND_c_1217_n 0.00317556f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_510 N_A2_M1007_g N_VGND_c_1218_n 4.44774e-19 $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_511 N_A2_M1012_g N_VGND_c_1218_n 0.00678063f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_512 N_A2_M1017_g N_VGND_c_1218_n 0.0028836f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_513 N_A2_M1017_g N_VGND_c_1219_n 4.44681e-19 $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_514 N_A2_M1019_g N_VGND_c_1219_n 0.00678207f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_515 N_A2_M1007_g N_VGND_c_1222_n 0.00331438f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_516 N_A2_M1012_g N_VGND_c_1222_n 0.00281141f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_517 N_A2_M1017_g N_VGND_c_1223_n 0.00331438f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_518 N_A2_M1019_g N_VGND_c_1223_n 0.00281141f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_519 N_A2_M1007_g N_VGND_c_1226_n 0.00427339f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A2_M1012_g N_VGND_c_1226_n 0.00365066f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A2_M1017_g N_VGND_c_1226_n 0.00426745f $X=7.785 $Y=0.74 $X2=0 $Y2=0
cc_522 N_A2_M1019_g N_VGND_c_1226_n 0.00365066f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_523 N_VPWR_c_650_n N_Y_c_780_n 0.0289761f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_524 N_VPWR_c_651_n N_Y_c_780_n 0.0266809f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_525 N_VPWR_c_658_n N_Y_c_780_n 0.0144623f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_648_n N_Y_c_780_n 0.0118344f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_M1014_s N_Y_c_802_n 0.00478602f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_528 N_VPWR_c_651_n N_Y_c_802_n 0.0196074f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_529 N_VPWR_c_651_n N_Y_c_781_n 0.0244596f $X=1.23 $Y=2.455 $X2=0 $Y2=0
cc_530 N_VPWR_c_652_n N_Y_c_781_n 0.0201138f $X=2.19 $Y=2.475 $X2=0 $Y2=0
cc_531 N_VPWR_c_659_n N_Y_c_781_n 0.011054f $X=2.025 $Y=3.33 $X2=0 $Y2=0
cc_532 N_VPWR_c_648_n N_Y_c_781_n 0.00914017f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_533 N_VPWR_M1035_s N_Y_c_811_n 0.0100499f $X=2.055 $Y=1.84 $X2=0 $Y2=0
cc_534 N_VPWR_M1020_d N_Y_c_811_n 0.00524267f $X=3.005 $Y=1.84 $X2=0 $Y2=0
cc_535 N_VPWR_c_652_n N_Y_c_811_n 0.0189268f $X=2.19 $Y=2.475 $X2=0 $Y2=0
cc_536 N_VPWR_M1028_d N_Y_c_835_n 0.0113144f $X=5.905 $Y=1.84 $X2=0 $Y2=0
cc_537 N_VPWR_c_654_n N_Y_c_835_n 0.0208278f $X=6.09 $Y=2.475 $X2=0 $Y2=0
cc_538 N_VPWR_M1020_d N_A_511_368#_c_924_n 0.00548861f $X=3.005 $Y=1.84 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_653_n N_A_511_368#_c_924_n 0.0202465f $X=3.19 $Y=2.815 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_648_n N_A_511_368#_c_924_n 0.0115311f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_661_n N_A_511_368#_c_915_n 0.0357927f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_648_n N_A_511_368#_c_915_n 0.0200586f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_653_n N_A_511_368#_c_916_n 0.0119238f $X=3.19 $Y=2.815 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_661_n N_A_511_368#_c_916_n 0.0234587f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_648_n N_A_511_368#_c_916_n 0.0125576f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_654_n N_A_511_368#_c_917_n 0.0119238f $X=6.09 $Y=2.475 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_661_n N_A_511_368#_c_917_n 0.0656793f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_648_n N_A_511_368#_c_917_n 0.0363721f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_652_n N_A_511_368#_c_918_n 0.0165124f $X=2.19 $Y=2.475 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_653_n N_A_511_368#_c_918_n 0.0101711f $X=3.19 $Y=2.815 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_660_n N_A_511_368#_c_918_n 0.0143153f $X=3.025 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_648_n N_A_511_368#_c_918_n 0.0117766f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_661_n N_A_511_368#_c_919_n 0.0234587f $X=5.925 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_648_n N_A_511_368#_c_919_n 0.0125576f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_662_n N_A_1291_368#_c_979_n 0.0439866f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_648_n N_A_1291_368#_c_979_n 0.0246722f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_655_n N_A_1291_368#_c_980_n 0.010126f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_662_n N_A_1291_368#_c_980_n 0.0581059f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_648_n N_A_1291_368#_c_980_n 0.0324093f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_M1010_s N_A_1291_368#_c_986_n 0.00317244f $X=8.76 $Y=1.84 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_655_n N_A_1291_368#_c_986_n 0.0148589f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_655_n N_A_1291_368#_c_981_n 0.0234083f $X=8.895 $Y=2.455 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_657_n N_A_1291_368#_c_981_n 0.0289761f $X=9.795 $Y=2.115 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_663_n N_A_1291_368#_c_981_n 0.0144623f $X=9.71 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_648_n N_A_1291_368#_c_981_n 0.0118344f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_654_n N_A_1291_368#_c_982_n 0.0214366f $X=6.09 $Y=2.475 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_662_n N_A_1291_368#_c_982_n 0.023f $X=8.73 $Y=3.33 $X2=0 $Y2=0
cc_568 N_VPWR_c_648_n N_A_1291_368#_c_982_n 0.0127161f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_662_n N_A_1291_368#_c_983_n 0.0121867f $X=8.73 $Y=3.33 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_648_n N_A_1291_368#_c_983_n 0.00660921f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_Y_c_811_n N_A_511_368#_M1003_s 0.0031756f $X=4.055 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_572 N_Y_c_811_n N_A_511_368#_M1022_s 0.00332066f $X=4.055 $Y=2.135 $X2=0
+ $Y2=0
cc_573 N_Y_c_833_n N_A_511_368#_M1025_d 0.00321395f $X=4.925 $Y=2.135 $X2=0
+ $Y2=0
cc_574 N_Y_c_835_n N_A_511_368#_M1036_d 0.00437964f $X=6.845 $Y=2.135 $X2=0
+ $Y2=0
cc_575 N_Y_c_811_n N_A_511_368#_c_924_n 0.0388605f $X=4.055 $Y=2.135 $X2=0 $Y2=0
cc_576 N_Y_c_811_n N_A_511_368#_c_926_n 0.0171885f $X=4.055 $Y=2.135 $X2=0 $Y2=0
cc_577 N_Y_M1005_s N_A_511_368#_c_915_n 0.00165831f $X=4.005 $Y=1.84 $X2=0 $Y2=0
cc_578 N_Y_c_890_p N_A_511_368#_c_915_n 0.0118804f $X=4.14 $Y=2.57 $X2=0 $Y2=0
cc_579 N_Y_c_833_n N_A_511_368#_c_941_n 0.0170361f $X=4.925 $Y=2.135 $X2=0 $Y2=0
cc_580 N_Y_M1032_s N_A_511_368#_c_917_n 0.00218982f $X=4.905 $Y=1.84 $X2=0 $Y2=0
cc_581 N_Y_c_834_n N_A_511_368#_c_917_n 0.0177184f $X=5.09 $Y=2.57 $X2=0 $Y2=0
cc_582 N_Y_c_835_n N_A_511_368#_c_931_n 0.0189382f $X=6.845 $Y=2.135 $X2=0 $Y2=0
cc_583 N_Y_c_811_n N_A_511_368#_c_918_n 0.0169819f $X=4.055 $Y=2.135 $X2=0 $Y2=0
cc_584 N_Y_c_835_n N_A_1291_368#_M1001_d 0.0102437f $X=6.845 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_585 N_Y_c_854_n N_A_1291_368#_M1023_s 0.00314376f $X=7.83 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_Y_M1021_d N_A_1291_368#_c_979_n 0.00165831f $X=6.96 $Y=1.84 $X2=0 $Y2=0
cc_587 Y N_A_1291_368#_c_979_n 0.0188729f $X=6.875 $Y=2.32 $X2=0 $Y2=0
cc_588 N_Y_c_854_n N_A_1291_368#_c_1022_n 0.0126919f $X=7.83 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_Y_M1029_d N_A_1291_368#_c_980_n 0.00165831f $X=7.86 $Y=1.84 $X2=0 $Y2=0
cc_590 N_Y_c_858_n N_A_1291_368#_c_980_n 0.0159318f $X=7.995 $Y=2.115 $X2=0
+ $Y2=0
cc_591 N_Y_c_835_n N_A_1291_368#_c_982_n 0.00907667f $X=6.845 $Y=2.135 $X2=0
+ $Y2=0
cc_592 Y N_A_1291_368#_c_982_n 0.00448535f $X=6.875 $Y=2.32 $X2=0 $Y2=0
cc_593 N_Y_c_776_n N_A_27_84#_M1002_d 0.00176461f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_594 N_Y_c_777_n N_A_27_84#_c_1027_n 0.00792678f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_595 N_Y_M1000_s N_A_27_84#_c_1028_n 0.00176461f $X=0.57 $Y=0.42 $X2=0 $Y2=0
cc_596 N_Y_c_784_n N_A_27_84#_c_1028_n 0.0157965f $X=0.71 $Y=0.68 $X2=0 $Y2=0
cc_597 N_Y_c_776_n N_A_27_84#_c_1028_n 0.00304353f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_598 N_Y_c_776_n N_A_27_84#_c_1078_n 0.0133411f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_599 N_Y_M1004_s N_A_27_84#_c_1030_n 0.00176461f $X=1.43 $Y=0.42 $X2=0 $Y2=0
cc_600 N_Y_c_776_n N_A_27_84#_c_1030_n 0.00304353f $X=1.405 $Y=1.095 $X2=0 $Y2=0
cc_601 N_Y_c_806_n N_A_27_84#_c_1030_n 0.0165966f $X=1.57 $Y=0.68 $X2=0 $Y2=0
cc_602 N_Y_c_778_n N_A_27_84#_c_1033_n 0.00808484f $X=1.575 $Y=1.095 $X2=0 $Y2=0
cc_603 N_A_27_84#_c_1032_n N_A_483_74#_M1009_s 0.00441709f $X=2.95 $Y=0.975
+ $X2=-0.19 $Y2=-0.245
cc_604 N_A_27_84#_c_1034_n N_A_483_74#_M1011_s 0.00176461f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_605 N_A_27_84#_c_1067_n N_A_483_74#_M1006_d 0.00332127f $X=5.405 $Y=0.91
+ $X2=0 $Y2=0
cc_606 N_A_27_84#_c_1067_n N_A_483_74#_M1016_d 0.00413357f $X=5.405 $Y=0.91
+ $X2=0 $Y2=0
cc_607 N_A_27_84#_M1009_d N_A_483_74#_c_1107_n 0.00179007f $X=2.85 $Y=0.37 $X2=0
+ $Y2=0
cc_608 N_A_27_84#_c_1030_n N_A_483_74#_c_1107_n 0.00560069f $X=1.915 $Y=0.34
+ $X2=0 $Y2=0
cc_609 N_A_27_84#_c_1031_n N_A_483_74#_c_1107_n 0.0121732f $X=2 $Y=0.565 $X2=0
+ $Y2=0
cc_610 N_A_27_84#_c_1032_n N_A_483_74#_c_1107_n 0.0445249f $X=2.95 $Y=0.975
+ $X2=0 $Y2=0
cc_611 N_A_27_84#_c_1034_n N_A_483_74#_c_1107_n 0.0174102f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_612 N_A_27_84#_M1030_d N_A_483_74#_c_1108_n 0.00178571f $X=3.71 $Y=0.37 $X2=0
+ $Y2=0
cc_613 N_A_27_84#_M1015_s N_A_483_74#_c_1108_n 0.00170263f $X=4.57 $Y=0.37 $X2=0
+ $Y2=0
cc_614 N_A_27_84#_M1026_s N_A_483_74#_c_1108_n 0.00179007f $X=5.43 $Y=0.37 $X2=0
+ $Y2=0
cc_615 N_A_27_84#_c_1034_n N_A_483_74#_c_1108_n 0.00427478f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_616 N_A_27_84#_c_1037_n N_A_483_74#_c_1108_n 0.0162997f $X=3.85 $Y=0.89 $X2=0
+ $Y2=0
cc_617 N_A_27_84#_c_1067_n N_A_483_74#_c_1108_n 0.0907973f $X=5.405 $Y=0.91
+ $X2=0 $Y2=0
cc_618 N_A_27_84#_c_1028_n N_VGND_c_1221_n 0.043102f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_27_84#_c_1029_n N_VGND_c_1221_n 0.0186386f $X=0.375 $Y=0.34 $X2=0
+ $Y2=0
cc_620 N_A_27_84#_c_1030_n N_VGND_c_1221_n 0.0616678f $X=1.915 $Y=0.34 $X2=0
+ $Y2=0
cc_621 N_A_27_84#_c_1035_n N_VGND_c_1221_n 0.0134682f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_27_84#_c_1028_n N_VGND_c_1226_n 0.0251825f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_623 N_A_27_84#_c_1029_n N_VGND_c_1226_n 0.0101082f $X=0.375 $Y=0.34 $X2=0
+ $Y2=0
cc_624 N_A_27_84#_c_1030_n N_VGND_c_1226_n 0.0352779f $X=1.915 $Y=0.34 $X2=0
+ $Y2=0
cc_625 N_A_27_84#_c_1032_n N_VGND_c_1226_n 0.0105008f $X=2.95 $Y=0.975 $X2=0
+ $Y2=0
cc_626 N_A_27_84#_c_1035_n N_VGND_c_1226_n 0.00735812f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_483_74#_c_1129_n N_VGND_M1008_s 0.00678566f $X=6.905 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_628 N_A_483_74#_c_1134_n N_VGND_M1012_d 0.00472947f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_629 N_A_483_74#_c_1135_n N_VGND_M1019_d 0.00398331f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_630 N_A_483_74#_c_1112_n N_VGND_M1031_s 0.00330483f $X=9.715 $Y=1.005 $X2=0
+ $Y2=0
cc_631 N_A_483_74#_c_1129_n N_VGND_c_1217_n 0.0240865f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_632 N_A_483_74#_c_1109_n N_VGND_c_1217_n 0.00906117f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_633 N_A_483_74#_c_1114_n N_VGND_c_1217_n 0.00942064f $X=6.07 $Y=0.475 $X2=0
+ $Y2=0
cc_634 N_A_483_74#_c_1109_n N_VGND_c_1218_n 0.00897147f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_635 N_A_483_74#_c_1134_n N_VGND_c_1218_n 0.0203034f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_636 N_A_483_74#_c_1110_n N_VGND_c_1218_n 0.00906117f $X=8 $Y=0.635 $X2=0
+ $Y2=0
cc_637 N_A_483_74#_c_1110_n N_VGND_c_1219_n 0.00900923f $X=8 $Y=0.635 $X2=0
+ $Y2=0
cc_638 N_A_483_74#_c_1135_n N_VGND_c_1219_n 0.0173074f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_639 N_A_483_74#_c_1111_n N_VGND_c_1219_n 0.00942763f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_640 N_A_483_74#_c_1111_n N_VGND_c_1220_n 0.0150645f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_483_74#_c_1112_n N_VGND_c_1220_n 0.0171619f $X=9.715 $Y=1.005 $X2=0
+ $Y2=0
cc_642 N_A_483_74#_c_1113_n N_VGND_c_1220_n 0.0150645f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_643 N_A_483_74#_c_1107_n N_VGND_c_1221_n 0.0454606f $X=3.335 $Y=0.475 $X2=0
+ $Y2=0
cc_644 N_A_483_74#_c_1108_n N_VGND_c_1221_n 0.0970299f $X=5.905 $Y=0.475 $X2=0
+ $Y2=0
cc_645 N_A_483_74#_c_1129_n N_VGND_c_1221_n 0.00190416f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_646 N_A_483_74#_c_1114_n N_VGND_c_1221_n 0.0145639f $X=6.07 $Y=0.475 $X2=0
+ $Y2=0
cc_647 N_A_483_74#_c_1129_n N_VGND_c_1222_n 0.00189877f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_648 N_A_483_74#_c_1109_n N_VGND_c_1222_n 0.0108551f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_649 N_A_483_74#_c_1134_n N_VGND_c_1222_n 0.00197156f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_650 N_A_483_74#_c_1134_n N_VGND_c_1223_n 0.00189877f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_651 N_A_483_74#_c_1110_n N_VGND_c_1223_n 0.0108551f $X=8 $Y=0.635 $X2=0 $Y2=0
cc_652 N_A_483_74#_c_1135_n N_VGND_c_1223_n 0.00197156f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_653 N_A_483_74#_c_1135_n N_VGND_c_1224_n 0.00190416f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_654 N_A_483_74#_c_1111_n N_VGND_c_1224_n 0.011066f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_483_74#_c_1113_n N_VGND_c_1225_n 0.011066f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_656 N_A_483_74#_c_1107_n N_VGND_c_1226_n 0.0383078f $X=3.335 $Y=0.475 $X2=0
+ $Y2=0
cc_657 N_A_483_74#_c_1108_n N_VGND_c_1226_n 0.0814955f $X=5.905 $Y=0.475 $X2=0
+ $Y2=0
cc_658 N_A_483_74#_c_1129_n N_VGND_c_1226_n 0.00891641f $X=6.905 $Y=0.835 $X2=0
+ $Y2=0
cc_659 N_A_483_74#_c_1109_n N_VGND_c_1226_n 0.00898945f $X=7.07 $Y=0.635 $X2=0
+ $Y2=0
cc_660 N_A_483_74#_c_1134_n N_VGND_c_1226_n 0.00914714f $X=7.835 $Y=0.835 $X2=0
+ $Y2=0
cc_661 N_A_483_74#_c_1110_n N_VGND_c_1226_n 0.00898945f $X=8 $Y=0.635 $X2=0
+ $Y2=0
cc_662 N_A_483_74#_c_1135_n N_VGND_c_1226_n 0.00917295f $X=8.775 $Y=0.835 $X2=0
+ $Y2=0
cc_663 N_A_483_74#_c_1111_n N_VGND_c_1226_n 0.00915947f $X=8.94 $Y=0.515 $X2=0
+ $Y2=0
cc_664 N_A_483_74#_c_1113_n N_VGND_c_1226_n 0.00915947f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_665 N_A_483_74#_c_1114_n N_VGND_c_1226_n 0.0119984f $X=6.07 $Y=0.475 $X2=0
+ $Y2=0

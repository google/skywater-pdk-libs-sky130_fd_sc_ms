* File: sky130_fd_sc_ms__o22ai_2.pxi.spice
* Created: Fri Aug 28 17:58:49 2020
* 
x_PM_SKY130_FD_SC_MS__O22AI_2%B1 N_B1_M1007_g N_B1_M1001_g N_B1_M1015_g
+ N_B1_M1013_g B1 B1 B1 N_B1_c_83_n PM_SKY130_FD_SC_MS__O22AI_2%B1
x_PM_SKY130_FD_SC_MS__O22AI_2%B2 N_B2_M1000_g N_B2_M1004_g N_B2_M1002_g
+ N_B2_M1006_g B2 N_B2_c_128_n N_B2_c_129_n PM_SKY130_FD_SC_MS__O22AI_2%B2
x_PM_SKY130_FD_SC_MS__O22AI_2%A2 N_A2_M1010_g N_A2_M1008_g N_A2_M1009_g
+ N_A2_M1014_g A2 N_A2_c_185_n N_A2_c_186_n PM_SKY130_FD_SC_MS__O22AI_2%A2
x_PM_SKY130_FD_SC_MS__O22AI_2%A1 N_A1_M1003_g N_A1_M1011_g N_A1_M1012_g
+ N_A1_M1005_g A1 A1 N_A1_c_243_n PM_SKY130_FD_SC_MS__O22AI_2%A1
x_PM_SKY130_FD_SC_MS__O22AI_2%A_28_368# N_A_28_368#_M1001_s N_A_28_368#_M1015_s
+ N_A_28_368#_M1002_s N_A_28_368#_c_287_n N_A_28_368#_c_288_n
+ N_A_28_368#_c_294_n N_A_28_368#_c_298_n N_A_28_368#_c_300_n
+ N_A_28_368#_c_289_n N_A_28_368#_c_290_n N_A_28_368#_c_291_n
+ PM_SKY130_FD_SC_MS__O22AI_2%A_28_368#
x_PM_SKY130_FD_SC_MS__O22AI_2%VPWR N_VPWR_M1001_d N_VPWR_M1011_d N_VPWR_c_333_n
+ N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n VPWR N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_332_n N_VPWR_c_340_n PM_SKY130_FD_SC_MS__O22AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O22AI_2%Y N_Y_M1007_s N_Y_M1004_s N_Y_M1000_d N_Y_M1008_d
+ N_Y_c_435_p N_Y_c_381_n N_Y_c_382_n N_Y_c_396_n N_Y_c_397_n N_Y_c_385_n
+ N_Y_c_412_n N_Y_c_398_n N_Y_c_383_n N_Y_c_386_n Y
+ PM_SKY130_FD_SC_MS__O22AI_2%Y
x_PM_SKY130_FD_SC_MS__O22AI_2%A_510_368# N_A_510_368#_M1008_s
+ N_A_510_368#_M1009_s N_A_510_368#_M1012_s N_A_510_368#_c_444_n
+ N_A_510_368#_c_445_n N_A_510_368#_c_446_n N_A_510_368#_c_456_n
+ N_A_510_368#_c_458_n N_A_510_368#_c_447_n N_A_510_368#_c_448_n
+ PM_SKY130_FD_SC_MS__O22AI_2%A_510_368#
x_PM_SKY130_FD_SC_MS__O22AI_2%A_27_74# N_A_27_74#_M1007_d N_A_27_74#_M1013_d
+ N_A_27_74#_M1006_d N_A_27_74#_M1014_d N_A_27_74#_M1005_d N_A_27_74#_c_483_n
+ N_A_27_74#_c_484_n N_A_27_74#_c_485_n N_A_27_74#_c_500_n N_A_27_74#_c_486_n
+ N_A_27_74#_c_487_n N_A_27_74#_c_488_n N_A_27_74#_c_489_n N_A_27_74#_c_490_n
+ N_A_27_74#_c_491_n N_A_27_74#_c_492_n N_A_27_74#_c_493_n
+ PM_SKY130_FD_SC_MS__O22AI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O22AI_2%VGND N_VGND_M1010_s N_VGND_M1003_s N_VGND_c_561_n
+ N_VGND_c_562_n VGND N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n
+ N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n PM_SKY130_FD_SC_MS__O22AI_2%VGND
cc_1 VNB N_B1_M1007_g 0.033015f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_M1013_g 0.0244807f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_3 VNB B1 0.0210388f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B1_c_83_n 0.040125f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.515
cc_5 VNB N_B2_M1004_g 0.0240538f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_6 VNB N_B2_M1006_g 0.0279479f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_7 VNB N_B2_c_128_n 0.00143484f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_8 VNB N_B2_c_129_n 0.0439761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_M1010_g 0.0239562f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A2_M1008_g 0.00191348f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_11 VNB N_A2_M1009_g 0.00158639f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_12 VNB N_A2_M1014_g 0.0219989f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_13 VNB A2 0.00672635f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_14 VNB N_A2_c_185_n 0.00345565f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_15 VNB N_A2_c_186_n 0.0542117f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_16 VNB N_A1_M1003_g 0.0244981f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_17 VNB N_A1_M1005_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_18 VNB A1 0.0134698f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB N_A1_c_243_n 0.0518765f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_20 VNB N_VPWR_c_332_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_381_n 0.00474786f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_Y_c_382_n 0.00340221f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_Y_c_383_n 0.00615473f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.565
cc_24 VNB Y 0.00712626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_483_n 0.0302158f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_26 VNB N_A_27_74#_c_484_n 0.00288965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_485_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_486_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_29 VNB N_A_27_74#_c_487_n 0.00329829f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_30 VNB N_A_27_74#_c_488_n 0.00207407f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_31 VNB N_A_27_74#_c_489_n 0.0132237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_490_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_33 VNB N_A_27_74#_c_491_n 0.00220733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_492_n 0.012391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_493_n 0.00327131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_561_n 0.00572435f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.68
cc_37 VNB N_VGND_c_562_n 0.00566037f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.35
cc_38 VNB N_VGND_c_563_n 0.0703081f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_39 VNB N_VGND_c_564_n 0.0183651f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_40 VNB N_VGND_c_565_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_41 VNB N_VGND_c_566_n 0.276858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_567_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_568_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_B1_M1001_g 0.0273599f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_45 VPB N_B1_M1015_g 0.0208199f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_46 VPB B1 0.0139021f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_47 VPB N_B1_c_83_n 0.0062744f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.515
cc_48 VPB N_B2_M1000_g 0.020326f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_49 VPB N_B2_M1002_g 0.0233473f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_50 VPB N_B2_c_128_n 0.00368074f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_51 VPB N_B2_c_129_n 0.00478561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A2_M1008_g 0.0258129f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_53 VPB N_A2_M1009_g 0.0216939f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_54 VPB A2 0.00500544f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_55 VPB N_A1_M1011_g 0.0207639f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_56 VPB N_A1_M1012_g 0.027583f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_57 VPB A1 0.0107393f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_58 VPB N_A1_c_243_n 0.0116224f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_59 VPB N_A_28_368#_c_287_n 0.00739392f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_60 VPB N_A_28_368#_c_288_n 0.0339247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_28_368#_c_289_n 0.00605183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_28_368#_c_290_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_28_368#_c_291_n 0.0056491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_333_n 0.0059449f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.68
cc_65 VPB N_VPWR_c_334_n 0.00554449f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.35
cc_66 VPB N_VPWR_c_335_n 0.0715147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_336_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_68 VPB N_VPWR_c_337_n 0.0181665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_338_n 0.0209017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_332_n 0.0795606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_340_n 0.0061237f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.565
cc_72 VPB N_Y_c_385_n 0.023148f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_73 VPB N_Y_c_386_n 5.97342e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB Y 0.00377136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_510_368#_c_444_n 0.00784838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_510_368#_c_445_n 0.00438754f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=0.74
cc_77 VPB N_A_510_368#_c_446_n 0.0041294f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=0.74
cc_78 VPB N_A_510_368#_c_447_n 0.00723723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_510_368#_c_448_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 N_B1_M1015_g N_B2_M1000_g 0.0167407f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_81 N_B1_M1013_g N_B2_M1004_g 0.0279646f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_82 B1 N_B2_c_128_n 0.0360516f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_83 N_B1_c_83_n N_B2_c_128_n 3.19042e-19 $X=1.025 $Y=1.515 $X2=0 $Y2=0
cc_84 B1 N_B2_c_129_n 0.0039539f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_85 N_B1_c_83_n N_B2_c_129_n 0.0167407f $X=1.025 $Y=1.515 $X2=0 $Y2=0
cc_86 B1 N_A_28_368#_c_287_n 0.0213698f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_87 N_B1_M1001_g N_A_28_368#_c_288_n 4.69176e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_88 N_B1_M1001_g N_A_28_368#_c_294_n 0.0145524f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_89 N_B1_M1015_g N_A_28_368#_c_294_n 0.0132272f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_90 B1 N_A_28_368#_c_294_n 0.047525f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_91 N_B1_c_83_n N_A_28_368#_c_294_n 7.63416e-19 $X=1.025 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B1_M1015_g N_A_28_368#_c_298_n 8.84614e-19 $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_93 B1 N_A_28_368#_c_298_n 0.0187568f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_94 N_B1_M1001_g N_A_28_368#_c_300_n 7.24402e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_95 N_B1_M1015_g N_A_28_368#_c_300_n 0.0102703f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_96 N_B1_M1015_g N_A_28_368#_c_290_n 0.00337536f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_97 N_B1_M1001_g N_VPWR_c_333_n 0.0158556f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_98 N_B1_M1015_g N_VPWR_c_333_n 0.00141551f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_99 N_B1_M1015_g N_VPWR_c_335_n 0.00517089f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_100 N_B1_M1001_g N_VPWR_c_337_n 0.00460063f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_101 N_B1_M1001_g N_VPWR_c_332_n 0.00912313f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_102 N_B1_M1015_g N_VPWR_c_332_n 0.00977404f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_103 N_B1_M1013_g N_Y_c_381_n 0.012846f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_104 B1 N_Y_c_381_n 0.0287022f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_105 N_B1_M1007_g N_Y_c_382_n 0.00241337f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_106 B1 N_Y_c_382_n 0.0280045f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B1_c_83_n N_Y_c_382_n 0.00486759f $X=1.025 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_M1007_g N_A_27_74#_c_483_n 0.0108851f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B1_M1013_g N_A_27_74#_c_483_n 6.35781e-19 $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_110 B1 N_A_27_74#_c_483_n 0.023775f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B1_M1007_g N_A_27_74#_c_484_n 0.0106115f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B1_M1013_g N_A_27_74#_c_484_n 0.0118932f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B1_M1007_g N_A_27_74#_c_485_n 0.00282152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_M1007_g N_VGND_c_563_n 0.00278247f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B1_M1013_g N_VGND_c_563_n 0.00278271f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_116 N_B1_M1007_g N_VGND_c_566_n 0.00357999f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_117 N_B1_M1013_g N_VGND_c_566_n 0.00354801f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B2_M1006_g N_A2_c_186_n 0.00279892f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_119 N_B2_c_129_n N_A2_c_186_n 0.00143843f $X=1.91 $Y=1.515 $X2=0 $Y2=0
cc_120 N_B2_M1000_g N_A_28_368#_c_298_n 0.00332483f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_121 N_B2_M1000_g N_A_28_368#_c_300_n 0.0101035f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B2_M1002_g N_A_28_368#_c_300_n 5.99195e-19 $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B2_M1000_g N_A_28_368#_c_289_n 0.0116345f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B2_M1002_g N_A_28_368#_c_289_n 0.014552f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B2_M1000_g N_A_28_368#_c_290_n 0.001916f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_126 N_B2_M1000_g N_A_28_368#_c_291_n 5.53268e-19 $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B2_M1002_g N_A_28_368#_c_291_n 0.00962971f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_128 N_B2_M1000_g N_VPWR_c_335_n 0.00333896f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B2_M1002_g N_VPWR_c_335_n 0.00333896f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_130 N_B2_M1000_g N_VPWR_c_332_n 0.00422796f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_131 N_B2_M1002_g N_VPWR_c_332_n 0.00427818f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_132 N_B2_M1004_g N_Y_c_381_n 0.014657f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_133 N_B2_c_128_n N_Y_c_381_n 0.0249311f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_134 N_B2_c_129_n N_Y_c_381_n 0.00207531f $X=1.91 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B2_M1006_g N_Y_c_396_n 0.0068998f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_136 N_B2_M1002_g N_Y_c_397_n 0.0202664f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_137 N_B2_c_128_n N_Y_c_398_n 0.0170903f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B2_c_129_n N_Y_c_398_n 5.52121e-19 $X=1.91 $Y=1.515 $X2=0 $Y2=0
cc_139 N_B2_M1006_g N_Y_c_383_n 0.0168118f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_140 N_B2_c_129_n N_Y_c_383_n 0.00174181f $X=1.91 $Y=1.515 $X2=0 $Y2=0
cc_141 N_B2_M1002_g N_Y_c_386_n 0.00535904f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_142 N_B2_M1004_g Y 8.02322e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_143 N_B2_M1006_g Y 0.00612352f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_144 N_B2_c_128_n Y 0.0261971f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_145 N_B2_c_129_n Y 0.0108092f $X=1.91 $Y=1.515 $X2=0 $Y2=0
cc_146 N_B2_M1002_g N_A_510_368#_c_444_n 0.00374777f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_147 N_B2_M1002_g N_A_510_368#_c_446_n 6.06861e-19 $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_148 N_B2_M1004_g N_A_27_74#_c_500_n 0.00682727f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_149 N_B2_M1006_g N_A_27_74#_c_500_n 4.62551e-19 $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_150 N_B2_M1004_g N_A_27_74#_c_486_n 0.00831967f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B2_M1006_g N_A_27_74#_c_486_n 0.0132502f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_152 N_B2_M1004_g N_A_27_74#_c_491_n 0.00272972f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_153 N_B2_M1006_g N_A_27_74#_c_492_n 0.0033343f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_154 N_B2_M1004_g N_VGND_c_563_n 0.00278247f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_155 N_B2_M1006_g N_VGND_c_563_n 0.00278271f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B2_M1004_g N_VGND_c_566_n 0.00354543f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B2_M1006_g N_VGND_c_566_n 0.00359085f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1014_g N_A1_M1003_g 0.0167769f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_159 A2 N_A1_M1003_g 3.98292e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A2_c_186_n N_A1_M1003_g 0.0173095f $X=3.375 $Y=1.465 $X2=0 $Y2=0
cc_161 A2 A1 0.0314575f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A2_c_186_n A1 2.9359e-19 $X=3.375 $Y=1.465 $X2=0 $Y2=0
cc_163 N_A2_M1009_g N_A1_c_243_n 0.0173095f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_164 A2 N_A1_c_243_n 0.0040064f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A2_M1008_g N_A_28_368#_c_289_n 6.06861e-19 $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A2_M1008_g N_A_28_368#_c_291_n 0.00133844f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A2_M1008_g N_VPWR_c_335_n 0.00333896f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A2_M1009_g N_VPWR_c_335_n 0.00333926f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A2_M1008_g N_VPWR_c_332_n 0.00427818f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A2_M1009_g N_VPWR_c_332_n 0.00422798f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_Y_c_385_n 0.0166271f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A2_M1009_g N_Y_c_385_n 0.00420946f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_173 A2 N_Y_c_385_n 0.0117309f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A2_c_185_n N_Y_c_385_n 0.0382159f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_175 N_A2_c_186_n N_Y_c_385_n 0.00548838f $X=3.375 $Y=1.465 $X2=0 $Y2=0
cc_176 N_A2_M1009_g N_Y_c_412_n 0.0111773f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A2_M1010_g N_Y_c_383_n 0.00158819f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_M1008_g N_Y_c_386_n 0.00389642f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A2_M1010_g Y 0.00283903f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A2_M1008_g Y 0.00411964f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A2_c_185_n Y 0.0143507f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_182 N_A2_c_186_n Y 0.0013782f $X=3.375 $Y=1.465 $X2=0 $Y2=0
cc_183 N_A2_M1008_g N_A_510_368#_c_444_n 0.0133315f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A2_M1009_g N_A_510_368#_c_444_n 7.17719e-19 $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A2_M1008_g N_A_510_368#_c_445_n 0.0115958f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A2_M1009_g N_A_510_368#_c_445_n 0.0137017f $X=3.37 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A2_M1008_g N_A_510_368#_c_446_n 0.00291744f $X=2.92 $Y=2.4 $X2=0 $Y2=0
cc_188 A2 N_A_510_368#_c_456_n 0.0143582f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_M1010_g N_A_27_74#_c_487_n 0.01289f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A2_M1014_g N_A_27_74#_c_487_n 0.0138493f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_191 A2 N_A_27_74#_c_487_n 0.0212066f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A2_c_185_n N_A_27_74#_c_487_n 0.0283f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_193 N_A2_c_186_n N_A_27_74#_c_487_n 0.00392092f $X=3.375 $Y=1.465 $X2=0 $Y2=0
cc_194 N_A2_M1014_g N_A_27_74#_c_488_n 4.09578e-19 $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A2_M1010_g N_A_27_74#_c_492_n 0.00384249f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A2_c_185_n N_A_27_74#_c_492_n 0.01012f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_197 N_A2_c_186_n N_A_27_74#_c_492_n 0.00279548f $X=3.375 $Y=1.465 $X2=0 $Y2=0
cc_198 N_A2_M1014_g N_A_27_74#_c_493_n 0.00158218f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_199 A2 N_A_27_74#_c_493_n 0.0162604f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A2_M1010_g N_VGND_c_561_n 0.0092302f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_M1014_g N_VGND_c_561_n 0.00222839f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A2_M1010_g N_VGND_c_563_n 0.00383152f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_M1014_g N_VGND_c_564_n 0.00461464f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A2_M1010_g N_VGND_c_566_n 0.00762539f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A2_M1014_g N_VGND_c_566_n 0.00907921f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A1_M1011_g N_VPWR_c_334_n 0.0117336f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A1_M1012_g N_VPWR_c_334_n 0.002979f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A1_M1011_g N_VPWR_c_335_n 0.00460063f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_M1012_g N_VPWR_c_338_n 0.005209f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A1_M1011_g N_VPWR_c_332_n 0.00908665f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A1_M1012_g N_VPWR_c_332_n 0.00986091f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_M1011_g N_Y_c_385_n 6.44128e-19 $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A1_M1011_g N_A_510_368#_c_445_n 0.00101073f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A1_M1011_g N_A_510_368#_c_458_n 0.0197231f $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A1_M1012_g N_A_510_368#_c_458_n 0.0128923f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_216 A1 N_A_510_368#_c_458_n 0.0282763f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A1_c_243_n N_A_510_368#_c_458_n 4.90767e-19 $X=4.415 $Y=1.515 $X2=0
+ $Y2=0
cc_218 N_A1_M1012_g N_A_510_368#_c_447_n 8.84614e-19 $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_219 A1 N_A_510_368#_c_447_n 0.0263957f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_220 N_A1_c_243_n N_A_510_368#_c_447_n 0.00121174f $X=4.415 $Y=1.515 $X2=0
+ $Y2=0
cc_221 N_A1_M1011_g N_A_510_368#_c_448_n 6.74232e-19 $X=3.82 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A1_M1012_g N_A_510_368#_c_448_n 0.0122988f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A1_M1003_g N_A_27_74#_c_488_n 0.00819795f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1005_g N_A_27_74#_c_488_n 6.73095e-19 $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_M1003_g N_A_27_74#_c_489_n 0.0153304f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1005_g N_A_27_74#_c_489_n 0.0140467f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_227 A1 N_A_27_74#_c_489_n 0.0606947f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_228 N_A1_c_243_n N_A_27_74#_c_489_n 0.00873549f $X=4.415 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A1_M1005_g N_A_27_74#_c_490_n 0.00159319f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1003_g N_A_27_74#_c_493_n 0.00340873f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1005_g N_A_27_74#_c_493_n 2.34371e-19 $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_M1003_g N_VGND_c_562_n 0.00429078f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1005_g N_VGND_c_562_n 0.0137334f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1003_g N_VGND_c_564_n 0.00434272f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1005_g N_VGND_c_565_n 0.00383152f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1003_g N_VGND_c_566_n 0.00820816f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1005_g N_VGND_c_566_n 0.00761198f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_28_368#_c_294_n N_VPWR_M1001_d 0.00410979f $X=1.07 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_239 N_A_28_368#_c_288_n N_VPWR_c_333_n 0.0234083f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_240 N_A_28_368#_c_294_n N_VPWR_c_333_n 0.0189268f $X=1.07 $Y=2.035 $X2=0
+ $Y2=0
cc_241 N_A_28_368#_c_290_n N_VPWR_c_333_n 0.0119238f $X=1.4 $Y=2.99 $X2=0 $Y2=0
cc_242 N_A_28_368#_c_289_n N_VPWR_c_335_n 0.0593439f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_243 N_A_28_368#_c_290_n N_VPWR_c_335_n 0.0234458f $X=1.4 $Y=2.99 $X2=0 $Y2=0
cc_244 N_A_28_368#_c_288_n N_VPWR_c_337_n 0.011066f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_245 N_A_28_368#_c_288_n N_VPWR_c_332_n 0.00915947f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_246 N_A_28_368#_c_289_n N_VPWR_c_332_n 0.032751f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_247 N_A_28_368#_c_290_n N_VPWR_c_332_n 0.0125551f $X=1.4 $Y=2.99 $X2=0 $Y2=0
cc_248 N_A_28_368#_c_289_n N_Y_M1000_d 0.00165831f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_249 N_A_28_368#_c_291_n N_Y_c_397_n 0.00216696f $X=2.135 $Y=2.375 $X2=0 $Y2=0
cc_250 N_A_28_368#_M1002_s N_Y_c_385_n 4.3007e-19 $X=2 $Y=1.84 $X2=0 $Y2=0
cc_251 N_A_28_368#_c_291_n N_Y_c_385_n 0.00128853f $X=2.135 $Y=2.375 $X2=0 $Y2=0
cc_252 N_A_28_368#_c_289_n N_Y_c_398_n 0.0118736f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_253 N_A_28_368#_M1002_s N_Y_c_386_n 0.00674064f $X=2 $Y=1.84 $X2=0 $Y2=0
cc_254 N_A_28_368#_c_291_n N_Y_c_386_n 0.0195651f $X=2.135 $Y=2.375 $X2=0 $Y2=0
cc_255 N_A_28_368#_c_291_n N_A_510_368#_c_444_n 0.0413949f $X=2.135 $Y=2.375
+ $X2=0 $Y2=0
cc_256 N_A_28_368#_c_289_n N_A_510_368#_c_446_n 0.0128664f $X=1.97 $Y=2.99 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_334_n N_A_510_368#_c_445_n 0.010126f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_335_n N_A_510_368#_c_445_n 0.0530426f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_332_n N_A_510_368#_c_445_n 0.0295386f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_335_n N_A_510_368#_c_446_n 0.0235512f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_332_n N_A_510_368#_c_446_n 0.0126924f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_M1011_d N_A_510_368#_c_458_n 0.00314376f $X=3.91 $Y=1.84 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_334_n N_A_510_368#_c_458_n 0.0148589f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_334_n N_A_510_368#_c_448_n 0.0234083f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_338_n N_A_510_368#_c_448_n 0.014549f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_332_n N_A_510_368#_c_448_n 0.0119743f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_Y_c_385_n N_A_510_368#_M1008_s 0.00308455f $X=3.06 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_268 N_Y_c_385_n N_A_510_368#_c_444_n 0.0219147f $X=3.06 $Y=1.885 $X2=0 $Y2=0
cc_269 N_Y_M1008_d N_A_510_368#_c_445_n 0.00165831f $X=3.01 $Y=1.84 $X2=0 $Y2=0
cc_270 N_Y_c_412_n N_A_510_368#_c_445_n 0.0139027f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_271 N_Y_c_381_n N_A_27_74#_M1013_d 0.00218982f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_272 N_Y_c_383_n N_A_27_74#_M1006_d 0.00272289f $X=2.16 $Y=1.18 $X2=0 $Y2=0
cc_273 N_Y_c_382_n N_A_27_74#_c_483_n 0.00540984f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_274 N_Y_M1007_s N_A_27_74#_c_484_n 0.00288741f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_275 N_Y_c_435_p N_A_27_74#_c_484_n 0.0200134f $X=0.78 $Y=0.76 $X2=0 $Y2=0
cc_276 N_Y_c_381_n N_A_27_74#_c_484_n 0.0036669f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_277 N_Y_c_381_n N_A_27_74#_c_500_n 0.0183199f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_278 N_Y_M1004_s N_A_27_74#_c_486_n 0.00250873f $X=1.57 $Y=0.37 $X2=0 $Y2=0
cc_279 N_Y_c_381_n N_A_27_74#_c_486_n 0.00612372f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_280 N_Y_c_396_n N_A_27_74#_c_486_n 0.018913f $X=1.78 $Y=0.76 $X2=0 $Y2=0
cc_281 N_Y_c_396_n N_A_27_74#_c_492_n 0.00573111f $X=1.78 $Y=0.76 $X2=0 $Y2=0
cc_282 N_Y_c_385_n N_A_27_74#_c_492_n 0.00678392f $X=3.06 $Y=1.885 $X2=0 $Y2=0
cc_283 N_Y_c_383_n N_A_27_74#_c_492_n 0.0222436f $X=2.16 $Y=1.18 $X2=0 $Y2=0
cc_284 N_A_27_74#_c_487_n N_VGND_M1010_s 0.00218982f $X=3.505 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_285 N_A_27_74#_c_489_n N_VGND_M1003_s 0.00250873f $X=4.435 $Y=1.095 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_487_n N_VGND_c_561_n 0.0185459f $X=3.505 $Y=1.045 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_c_488_n N_VGND_c_561_n 0.00129215f $X=3.59 $Y=0.515 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_c_492_n N_VGND_c_561_n 0.0254844f $X=2.69 $Y=0.965 $X2=0 $Y2=0
cc_289 N_A_27_74#_c_488_n N_VGND_c_562_n 0.0184106f $X=3.59 $Y=0.515 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_489_n N_VGND_c_562_n 0.0209867f $X=4.435 $Y=1.095 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_c_490_n N_VGND_c_562_n 0.0182902f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_484_n N_VGND_c_563_n 0.0423044f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_485_n N_VGND_c_563_n 0.0235688f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_486_n N_VGND_c_563_n 0.0423044f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_491_n N_VGND_c_563_n 0.0233048f $X=1.28 $Y=0.34 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_492_n N_VGND_c_563_n 0.0477547f $X=2.69 $Y=0.965 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_488_n N_VGND_c_564_n 0.0109942f $X=3.59 $Y=0.515 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_490_n N_VGND_c_565_n 0.011066f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_484_n N_VGND_c_566_n 0.0239316f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_485_n N_VGND_c_566_n 0.0127152f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_486_n N_VGND_c_566_n 0.0239316f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_488_n N_VGND_c_566_n 0.00904371f $X=3.59 $Y=0.515 $X2=0
+ $Y2=0
cc_303 N_A_27_74#_c_490_n N_VGND_c_566_n 0.00915947f $X=4.52 $Y=0.515 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_491_n N_VGND_c_566_n 0.0126653f $X=1.28 $Y=0.34 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_492_n N_VGND_c_566_n 0.0259963f $X=2.69 $Y=0.965 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dfsbp_2.pex.spice
* Created: Wed Sep  2 12:03:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFSBP_2%D 2 5 9 11 12 16 17 20
c34 17 0 1.14039e-19 $X=0.64 $Y=1.145
r35 20 22 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.825
+ $X2=0.61 $Y2=1.99
r36 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r37 16 18 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.145
+ $X2=0.61 $Y2=0.98
r38 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r39 12 21 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r40 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r41 11 17 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r42 9 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r43 5 22 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.505 $Y=2.75
+ $X2=0.505 $Y2=1.99
r44 2 20 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.795 $X2=0.61
+ $Y2=1.825
r45 1 16 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.145
r46 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%CLK 3 6 8 11 13
c39 11 0 1.39813e-19 $X=1.465 $Y=1.385
c40 6 0 1.14039e-19 $X=1.515 $Y=2.35
r41 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.55
r42 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.22
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r44 8 12 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r45 6 14 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=1.515 $Y=2.35 $X2=1.515
+ $Y2=1.55
r46 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=0.74
+ $X2=1.485 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_398_74# 1 2 7 8 11 13 17 21 24 26 29 33 35
+ 36 37 38 41 48 49 52 53 56 57 58 60 61 62 64 66 67 68 71 72 76 77 80 82 89 93
c270 80 0 2.30667e-19 $X=7.415 $Y=2.185
c271 77 0 8.86437e-20 $X=6.71 $Y=1.285
c272 62 0 1.1883e-19 $X=5.53 $Y=2.275
c273 61 0 1.74055e-19 $X=6.33 $Y=2.275
c274 26 0 1.40033e-19 $X=2.95 $Y=2.105
r275 81 93 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.415 $Y=2.185
+ $X2=7.53 $Y2=2.185
r276 80 82 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=2.185
+ $X2=7.415 $Y2=2.02
r277 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.415
+ $Y=2.185 $X2=7.415 $Y2=2.185
r278 77 89 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.71 $Y=1.285
+ $X2=6.71 $Y2=1.12
r279 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.285 $X2=6.71 $Y2=1.285
r280 73 76 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.415 $Y=1.285
+ $X2=6.71 $Y2=1.285
r281 69 82 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=7.47 $Y=0.45
+ $X2=7.47 $Y2=2.02
r282 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=0.365
+ $X2=7.47 $Y2=0.45
r283 67 68 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=7.385 $Y=0.365
+ $X2=6.5 $Y2=0.365
r284 65 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=1.45
+ $X2=6.415 $Y2=1.285
r285 65 66 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.415 $Y=1.45
+ $X2=6.415 $Y2=2.19
r286 64 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=1.12
+ $X2=6.415 $Y2=1.285
r287 63 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=0.45
+ $X2=6.5 $Y2=0.365
r288 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.415 $Y=0.45
+ $X2=6.415 $Y2=1.12
r289 61 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=2.275
+ $X2=6.415 $Y2=2.19
r290 61 62 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.33 $Y=2.275
+ $X2=5.53 $Y2=2.275
r291 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.445 $Y=2.36
+ $X2=5.53 $Y2=2.275
r292 59 60 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.445 $Y=2.36
+ $X2=5.445 $Y2=2.905
r293 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.36 $Y=2.99
+ $X2=5.445 $Y2=2.905
r294 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.36 $Y=2.99
+ $X2=4.69 $Y2=2.99
r295 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.605 $Y=2.905
+ $X2=4.69 $Y2=2.99
r296 55 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.605 $Y=2.565
+ $X2=4.605 $Y2=2.905
r297 54 72 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.845 $Y=2.48
+ $X2=3.735 $Y2=2.48
r298 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.52 $Y=2.48
+ $X2=4.605 $Y2=2.565
r299 53 54 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.52 $Y=2.48
+ $X2=3.845 $Y2=2.48
r300 51 72 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=2.565
+ $X2=3.735 $Y2=2.48
r301 51 52 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=3.735 $Y=2.565
+ $X2=3.735 $Y2=2.905
r302 49 85 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.735 $Y=1.6
+ $X2=3.58 $Y2=1.6
r303 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.735
+ $Y=1.6 $X2=3.735 $Y2=1.6
r304 46 72 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=2.395
+ $X2=3.735 $Y2=2.48
r305 46 48 41.6451 $w=2.18e-07 $l=7.95e-07 $layer=LI1_cond $X=3.735 $Y=2.395
+ $X2=3.735 $Y2=1.6
r306 44 71 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.025 $Y=0.425
+ $X2=3.025 $Y2=1.435
r307 41 71 8.30336 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.6
+ $X2=2.95 $Y2=1.435
r308 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.6 $X2=2.95 $Y2=1.6
r309 37 52 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=3.735 $Y2=2.905
r310 37 38 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=2.275 $Y2=2.99
r311 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.94 $Y=0.34
+ $X2=3.025 $Y2=0.425
r312 35 36 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.94 $Y=0.34
+ $X2=2.215 $Y2=0.34
r313 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.275 $Y2=2.99
r314 31 33 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.19 $Y2=2.665
r315 27 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.215 $Y2=0.34
r316 27 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r317 22 93 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.53 $Y=2.35
+ $X2=7.53 $Y2=2.185
r318 22 24 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=7.53 $Y=2.35 $X2=7.53
+ $Y2=2.75
r319 21 89 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.62 $Y=0.69
+ $X2=6.62 $Y2=1.12
r320 15 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.435
+ $X2=3.58 $Y2=1.6
r321 15 17 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.58 $Y=1.435
+ $X2=3.58 $Y2=0.695
r322 14 42 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.6
+ $X2=2.95 $Y2=1.6
r323 13 85 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=1.6
+ $X2=3.58 $Y2=1.6
r324 13 14 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=3.505 $Y=1.6
+ $X2=3.115 $Y2=1.6
r325 11 26 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=3.005 $Y=2.525
+ $X2=3.005 $Y2=2.105
r326 8 26 38.198 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.94
+ $X2=2.95 $Y2=2.105
r327 7 42 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.765
+ $X2=2.95 $Y2=1.6
r328 7 8 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.95 $Y=1.765
+ $X2=2.95 $Y2=1.94
r329 2 33 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.79 $X2=2.19 $Y2=2.665
r330 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_757_401# 1 2 9 11 13 14 15 16 17 20 23 24
+ 29 33 37
c88 23 0 1.10712e-19 $X=4.305 $Y=1.99
c89 9 0 9.24866e-20 $X=3.875 $Y=2.525
r90 37 43 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.37 $Y=1.825
+ $X2=4.37 $Y2=1.345
r91 33 35 16.7582 $w=2.73e-07 $l=3.75e-07 $layer=LI1_cond $X=5.025 $Y=2.14
+ $X2=5.025 $Y2=2.515
r92 32 43 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.462 $Y=1.18
+ $X2=4.462 $Y2=1.345
r93 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.465
+ $Y=1.18 $X2=4.465 $Y2=1.18
r94 29 31 18.866 $w=3.88e-07 $l=6.71714e-07 $layer=LI1_cond $X=4.617 $Y=0.58
+ $X2=4.465 $Y2=1.18
r95 24 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.99
+ $X2=4.305 $Y2=2.08
r96 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.99
+ $X2=4.305 $Y2=1.825
r97 23 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.305 $Y=1.99
+ $X2=4.305 $Y2=2.14
r98 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=1.99 $X2=4.305 $Y2=1.99
r99 21 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=2.14
+ $X2=4.305 $Y2=2.14
r100 20 33 3.50848 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=2.14
+ $X2=5.025 $Y2=2.14
r101 20 21 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.86 $Y=2.14
+ $X2=4.47 $Y2=2.14
r102 16 32 15.5026 $w=3.35e-07 $l=9e-08 $layer=POLY_cond $X=4.462 $Y=1.09
+ $X2=4.462 $Y2=1.18
r103 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.295 $Y=1.09
+ $X2=4.015 $Y2=1.09
r104 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=2.08
+ $X2=4.305 $Y2=2.08
r105 14 15 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.14 $Y=2.08
+ $X2=3.965 $Y2=2.08
r106 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.94 $Y=1.015
+ $X2=4.015 $Y2=1.09
r107 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.94 $Y=1.015
+ $X2=3.94 $Y2=0.695
r108 7 15 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.875 $Y=2.155
+ $X2=3.965 $Y2=2.08
r109 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.875 $Y=2.155
+ $X2=3.875 $Y2=2.525
r110 2 35 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.315 $X2=5.025 $Y2=2.515
r111 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.715 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_595_97# 1 2 9 13 15 19 21 23 24 27 30 32
+ 33 36 37 38 44 46 47 48 53 56 58 63
c163 56 0 8.86437e-20 $X=5.75 $Y=1.285
c164 53 0 2.29347e-19 $X=4.85 $Y=1.72
c165 46 0 1.55885e-19 $X=3.405 $Y=0.925
c166 44 0 1.40033e-19 $X=3.37 $Y=2.515
c167 32 0 9.24866e-20 $X=3.37 $Y=2.295
c168 9 0 1.1883e-19 $X=4.8 $Y=2.525
r169 57 63 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.75 $Y=1.285
+ $X2=5.75 $Y2=1.195
r170 56 58 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=1.265
+ $X2=5.585 $Y2=1.265
r171 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.75
+ $Y=1.285 $X2=5.75 $Y2=1.285
r172 53 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.72
+ $X2=4.85 $Y2=1.885
r173 53 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.72
+ $X2=4.85 $Y2=1.555
r174 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.72 $X2=4.85 $Y2=1.72
r175 42 44 3.66686 $w=4.38e-07 $l=1.4e-07 $layer=LI1_cond $X=3.23 $Y=2.515
+ $X2=3.37 $Y2=2.515
r176 40 48 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.015 $Y=1.325
+ $X2=4.882 $Y2=1.325
r177 40 58 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.015 $Y=1.325
+ $X2=5.585 $Y2=1.325
r178 37 52 5.21861 $w=2.63e-07 $l=1.2e-07 $layer=LI1_cond $X=4.882 $Y=1.6
+ $X2=4.882 $Y2=1.72
r179 37 48 11.9593 $w=2.63e-07 $l=2.75e-07 $layer=LI1_cond $X=4.882 $Y=1.6
+ $X2=4.882 $Y2=1.325
r180 37 38 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.75 $Y=1.6
+ $X2=4.185 $Y2=1.6
r181 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.1 $Y=1.515
+ $X2=4.185 $Y2=1.6
r182 35 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.1 $Y=1.265
+ $X2=4.1 $Y2=1.515
r183 34 47 2.06925 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.53 $Y=1.18
+ $X2=3.407 $Y2=1.18
r184 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=1.18
+ $X2=4.1 $Y2=1.265
r185 33 34 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.015 $Y=1.18
+ $X2=3.53 $Y2=1.18
r186 32 44 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.37 $Y=2.295
+ $X2=3.37 $Y2=2.515
r187 31 47 4.36305 $w=2.07e-07 $l=1.01833e-07 $layer=LI1_cond $X=3.37 $Y=1.265
+ $X2=3.407 $Y2=1.18
r188 31 32 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.37 $Y=1.265
+ $X2=3.37 $Y2=2.295
r189 30 47 4.36305 $w=2.07e-07 $l=8.5e-08 $layer=LI1_cond $X=3.407 $Y=1.095
+ $X2=3.407 $Y2=1.18
r190 30 46 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=3.407 $Y=1.095
+ $X2=3.407 $Y2=0.925
r191 25 46 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.405 $Y=0.8
+ $X2=3.405 $Y2=0.925
r192 25 27 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=3.405 $Y=0.8
+ $X2=3.405 $Y2=0.695
r193 21 24 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.23 $Y=1.12
+ $X2=6.215 $Y2=1.195
r194 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.23 $Y=1.12
+ $X2=6.23 $Y2=0.69
r195 17 24 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=6.215 $Y=1.27
+ $X2=6.215 $Y2=1.195
r196 17 19 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=6.215 $Y=1.27
+ $X2=6.215 $Y2=2.205
r197 16 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.195
+ $X2=5.75 $Y2=1.195
r198 15 24 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.125 $Y=1.195
+ $X2=6.215 $Y2=1.195
r199 15 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.125 $Y=1.195
+ $X2=5.915 $Y2=1.195
r200 13 61 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=4.93 $Y=0.58
+ $X2=4.93 $Y2=1.555
r201 9 62 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=4.8 $Y=2.525 $X2=4.8
+ $Y2=1.885
r202 2 42 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=2.315 $X2=3.23 $Y2=2.515
r203 1 27 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.485 $X2=3.365 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%SET_B 3 8 10 12 13 14 17 19 20 21 22 25 27
+ 30 32 34 38
c121 30 0 1.74055e-19 $X=5.39 $Y=1.855
c122 22 0 1.18634e-19 $X=5.665 $Y=1.665
r123 38 47 10.3882 $w=3.53e-07 $l=3.2e-07 $layer=LI1_cond $X=8.462 $Y=1.345
+ $X2=8.462 $Y2=1.665
r124 37 39 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.475 $Y=1.345
+ $X2=8.475 $Y2=1.51
r125 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.475
+ $Y=1.345 $X2=8.475 $Y2=1.345
r126 34 37 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.475 $Y=1.165
+ $X2=8.475 $Y2=1.345
r127 30 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.39 $Y=1.855
+ $X2=5.39 $Y2=2.02
r128 30 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.39 $Y=1.855
+ $X2=5.39 $Y2=1.69
r129 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.39
+ $Y=1.855 $X2=5.39 $Y2=1.855
r130 27 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r131 25 31 5.34059 $w=4.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=1.855
r132 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r133 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r134 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r135 21 22 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.665 $Y2=1.665
r136 20 32 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=5.3 $Y=1.015
+ $X2=5.3 $Y2=1.69
r137 19 20 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=5.295 $Y=0.865
+ $X2=5.295 $Y2=1.015
r138 17 39 482 $w=1.8e-07 $l=1.24e-06 $layer=POLY_cond $X=8.4 $Y=2.75 $X2=8.4
+ $Y2=1.51
r139 13 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.31 $Y=1.165
+ $X2=8.475 $Y2=1.165
r140 13 14 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.31 $Y=1.165
+ $X2=8.045 $Y2=1.165
r141 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.97 $Y=1.09
+ $X2=8.045 $Y2=1.165
r142 10 12 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.97 $Y=1.09
+ $X2=7.97 $Y2=0.8
r143 8 33 196.298 $w=1.8e-07 $l=5.05e-07 $layer=POLY_cond $X=5.315 $Y=2.525
+ $X2=5.315 $Y2=2.02
r144 3 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.29 $Y=0.58 $X2=5.29
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_225_74# 1 2 9 13 16 17 19 20 23 27 29 34
+ 35 36 39 42 43 46 47 49 50 51 54 58 62 65
c181 54 0 2.99812e-20 $X=1.945 $Y=1.805
c182 35 0 1.08117e-19 $X=7.115 $Y=1.735
r183 62 64 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r184 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.465 $X2=2.11 $Y2=1.465
r185 56 58 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.465
r186 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=2.11 $Y2=1.72
r187 54 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.455 $Y2=1.805
r188 51 53 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=1.87
+ $X2=1.29 $Y2=1.87
r189 50 65 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.455 $Y2=1.87
r190 50 53 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.29 $Y2=1.87
r191 49 51 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.145 $Y2=1.87
r192 49 64 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r193 46 59 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.11 $Y2=1.465
r194 43 46 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.485 $Y=1.12
+ $X2=2.485 $Y2=1.465
r195 41 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=2.11 $Y2=1.465
r196 41 42 3.90195 $w=3.3e-07 $l=1.08e-07 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=1.947 $Y2=1.465
r197 37 39 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.19 $Y=1.66
+ $X2=7.19 $Y2=0.8
r198 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.115 $Y=1.735
+ $X2=7.19 $Y2=1.66
r199 35 36 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.115 $Y=1.735
+ $X2=6.81 $Y2=1.735
r200 32 34 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=6.72 $Y=3.075
+ $X2=6.72 $Y2=2.46
r201 31 36 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.72 $Y=1.81
+ $X2=6.81 $Y2=1.735
r202 31 34 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=6.72 $Y=1.81
+ $X2=6.72 $Y2=2.46
r203 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.545 $Y=3.15
+ $X2=3.455 $Y2=3.15
r204 29 32 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.63 $Y=3.15
+ $X2=6.72 $Y2=3.075
r205 29 30 1581.88 $w=1.5e-07 $l=3.085e-06 $layer=POLY_cond $X=6.63 $Y=3.15
+ $X2=3.545 $Y2=3.15
r206 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.455 $Y=3.075
+ $X2=3.455 $Y2=3.15
r207 25 27 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.455 $Y=3.075
+ $X2=3.455 $Y2=2.525
r208 21 23 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.9 $Y=1.045
+ $X2=2.9 $Y2=0.695
r209 19 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.365 $Y=3.15
+ $X2=3.455 $Y2=3.15
r210 19 20 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.365 $Y=3.15
+ $X2=2.56 $Y2=3.15
r211 18 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.12
+ $X2=2.485 $Y2=1.12
r212 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.825 $Y=1.12
+ $X2=2.9 $Y2=1.045
r213 17 18 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.825 $Y=1.12
+ $X2=2.56 $Y2=1.12
r214 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r215 15 46 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=1.465
r216 15 16 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=3.075
r217 11 42 34.7346 $w=1.65e-07 $l=1.73767e-07 $layer=POLY_cond $X=1.965 $Y=1.63
+ $X2=1.947 $Y2=1.465
r218 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.965 $Y=1.63
+ $X2=1.965 $Y2=2.35
r219 7 42 34.7346 $w=1.65e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.947 $Y2=1.465
r220 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.915 $Y2=0.74
r221 2 53 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.79 $X2=1.29 $Y2=1.935
r222 1 62 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_1501_92# 1 2 9 13 17 18 20 21 22 24 27 28
+ 34
c99 22 0 1.4228e-19 $X=9.74 $Y=2.375
c100 18 0 2.30361e-19 $X=7.89 $Y=1.615
r101 36 37 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.27 $Y=0.925
+ $X2=9.27 $Y2=1.095
r102 34 36 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.27 $Y=0.8
+ $X2=9.27 $Y2=0.925
r103 28 31 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.18 $Y=2.375 $X2=9.18
+ $Y2=2.455
r104 26 27 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=9.825 $Y=1.18
+ $X2=9.825 $Y2=2.29
r105 25 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=1.095
+ $X2=9.27 $Y2=1.095
r106 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.74 $Y=1.095
+ $X2=9.825 $Y2=1.18
r107 24 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.74 $Y=1.095
+ $X2=9.435 $Y2=1.095
r108 23 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.345 $Y=2.375
+ $X2=9.18 $Y2=2.375
r109 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.74 $Y=2.375
+ $X2=9.825 $Y2=2.29
r110 22 23 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.74 $Y=2.375
+ $X2=9.345 $Y2=2.375
r111 20 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=0.925
+ $X2=9.27 $Y2=0.925
r112 20 21 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=9.105 $Y=0.925
+ $X2=8.055 $Y2=0.925
r113 18 41 11.2093 $w=2.58e-07 $l=6e-08 $layer=POLY_cond $X=7.89 $Y=1.615
+ $X2=7.95 $Y2=1.615
r114 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.615 $X2=7.89 $Y2=1.615
r115 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.89 $Y=1.01
+ $X2=8.055 $Y2=0.925
r116 15 17 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=7.89 $Y=1.01
+ $X2=7.89 $Y2=1.615
r117 11 41 11.2427 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.95 $Y=1.78
+ $X2=7.95 $Y2=1.615
r118 11 13 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=7.95 $Y=1.78
+ $X2=7.95 $Y2=2.75
r119 7 18 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=7.58 $Y=1.45
+ $X2=7.89 $Y2=1.615
r120 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=7.58 $Y=1.45 $X2=7.58
+ $Y2=0.8
r121 2 31 600 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=1 $X=9.035
+ $Y=1.84 $X2=9.18 $Y2=2.455
r122 1 34 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=9.05
+ $Y=0.59 $X2=9.27 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_1339_74# 1 2 3 12 14 15 18 20 24 28 32 36
+ 38 39 42 46 52 53 60 62 65 67 69 73 79 80 81 84
c185 65 0 1.07812e-19 $X=8.46 $Y=2.215
c186 52 0 8.81429e-20 $X=11.475 $Y=1.49
c187 14 0 1.4228e-19 $X=9.395 $Y=1.515
r188 83 84 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.405
+ $Y=1.515 $X2=9.405 $Y2=1.515
r189 80 81 9.81721 $w=5.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.75 $Y=2.3
+ $X2=7.92 $Y2=2.3
r190 79 80 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.47 $Y=2.565
+ $X2=7.75 $Y2=2.565
r191 78 79 9.51712 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=2.73
+ $X2=7.47 $Y2=2.73
r192 75 78 9.56863 $w=4.98e-07 $l=4e-07 $layer=LI1_cond $X=6.905 $Y=2.73
+ $X2=7.305 $Y2=2.73
r193 67 69 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.625 $Y=2.48
+ $X2=8.625 $Y2=2.75
r194 65 67 7.87997 $w=6.27e-07 $l=3.37565e-07 $layer=LI1_cond $X=8.46 $Y=2.215
+ $X2=8.625 $Y2=2.48
r195 65 83 13.6204 $w=6.27e-07 $l=9.37283e-07 $layer=LI1_cond $X=8.46 $Y=2.215
+ $X2=9.015 $Y2=1.515
r196 65 81 12.1865 $w=5.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.46 $Y=2.215
+ $X2=7.92 $Y2=2.215
r197 62 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.13 $Y=1.68
+ $X2=7.13 $Y2=1.765
r198 61 62 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.13 $Y=0.95
+ $X2=7.13 $Y2=1.68
r199 58 75 4.80115 $w=2.5e-07 $l=2.5e-07 $layer=LI1_cond $X=6.905 $Y=2.48
+ $X2=6.905 $Y2=2.73
r200 58 60 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=6.905 $Y=2.48
+ $X2=6.905 $Y2=2.135
r201 57 73 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.905 $Y=1.765
+ $X2=7.13 $Y2=1.765
r202 57 60 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.905 $Y=1.85
+ $X2=6.905 $Y2=2.135
r203 53 61 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.045 $Y=0.785
+ $X2=7.13 $Y2=0.95
r204 53 55 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.045 $Y=0.785
+ $X2=6.905 $Y2=0.785
r205 50 51 1.07119 $w=2.8e-07 $l=5e-09 $layer=POLY_cond $X=10.47 $Y=1.49
+ $X2=10.475 $Y2=1.49
r206 49 50 91.0515 $w=2.8e-07 $l=4.25e-07 $layer=POLY_cond $X=10.045 $Y=1.49
+ $X2=10.47 $Y2=1.49
r207 48 49 5.35597 $w=2.8e-07 $l=2.5e-08 $layer=POLY_cond $X=10.02 $Y=1.49
+ $X2=10.045 $Y2=1.49
r208 44 52 30.8978 $w=1.65e-07 $l=1.44914e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.475 $Y2=1.49
r209 44 46 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.465 $Y2=0.69
r210 40 52 30.8978 $w=1.65e-07 $l=1.4e-07 $layer=POLY_cond $X=11.475 $Y=1.63
+ $X2=11.475 $Y2=1.49
r211 40 42 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=11.475 $Y=1.63
+ $X2=11.475 $Y2=2.34
r212 39 51 18.2103 $w=2.8e-07 $l=8.5e-08 $layer=POLY_cond $X=10.56 $Y=1.49
+ $X2=10.475 $Y2=1.49
r213 38 52 1.86552 $w=2.8e-07 $l=9e-08 $layer=POLY_cond $X=11.385 $Y=1.49
+ $X2=11.475 $Y2=1.49
r214 38 39 176.747 $w=2.8e-07 $l=8.25e-07 $layer=POLY_cond $X=11.385 $Y=1.49
+ $X2=10.56 $Y2=1.49
r215 34 51 17.3521 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=10.475 $Y=1.35
+ $X2=10.475 $Y2=1.49
r216 34 36 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.475 $Y=1.35
+ $X2=10.475 $Y2=0.74
r217 30 50 13.127 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=10.47 $Y=1.63
+ $X2=10.47 $Y2=1.49
r218 30 32 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.47 $Y=1.63
+ $X2=10.47 $Y2=2.4
r219 26 49 17.3521 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=10.045 $Y=1.35
+ $X2=10.045 $Y2=1.49
r220 26 28 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.045 $Y=1.35
+ $X2=10.045 $Y2=0.74
r221 22 48 13.127 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=10.02 $Y=1.63
+ $X2=10.02 $Y2=1.49
r222 22 24 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.02 $Y=1.63
+ $X2=10.02 $Y2=2.4
r223 21 84 12.9058 $w=3.05e-07 $l=1.01735e-07 $layer=POLY_cond $X=9.575 $Y=1.49
+ $X2=9.485 $Y2=1.515
r224 20 48 19.2815 $w=2.8e-07 $l=9e-08 $layer=POLY_cond $X=9.93 $Y=1.49
+ $X2=10.02 $Y2=1.49
r225 20 21 76.0548 $w=2.8e-07 $l=3.55e-07 $layer=POLY_cond $X=9.93 $Y=1.49
+ $X2=9.575 $Y2=1.49
r226 16 84 13.0159 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.485 $Y=1.68
+ $X2=9.485 $Y2=1.515
r227 16 18 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.485 $Y=1.68
+ $X2=9.485 $Y2=2.05
r228 14 84 12.9058 $w=3.05e-07 $l=9e-08 $layer=POLY_cond $X=9.395 $Y=1.515
+ $X2=9.485 $Y2=1.515
r229 14 15 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=9.395 $Y=1.515
+ $X2=9.05 $Y2=1.515
r230 10 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.975 $Y=1.35
+ $X2=9.05 $Y2=1.515
r231 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.975 $Y=1.35
+ $X2=8.975 $Y2=0.8
r232 3 69 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.49
+ $Y=2.54 $X2=8.625 $Y2=2.75
r233 2 78 300 $w=1.7e-07 $l=1.07436e-06 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=1.96 $X2=7.305 $Y2=2.815
r234 2 60 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.81
+ $Y=1.96 $X2=6.945 $Y2=2.135
r235 1 55 182 $w=1.7e-07 $l=5.09289e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.37 $X2=6.905 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_2221_74# 1 2 9 13 17 21 25 29 35 38 44
r71 43 44 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=12.455 $Y=1.465
+ $X2=12.465 $Y2=1.465
r72 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.035 $Y=1.465
+ $X2=12.455 $Y2=1.465
r73 41 42 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=12.005 $Y=1.465
+ $X2=12.035 $Y2=1.465
r74 36 41 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=11.94 $Y=1.465
+ $X2=12.005 $Y2=1.465
r75 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.94
+ $Y=1.465 $X2=11.94 $Y2=1.465
r76 33 38 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.415 $Y=1.465
+ $X2=11.25 $Y2=1.465
r77 33 35 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=11.415 $Y=1.465
+ $X2=11.94 $Y2=1.465
r78 29 31 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.25 $Y=1.985
+ $X2=11.25 $Y2=2.695
r79 27 38 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.25 $Y=1.63
+ $X2=11.25 $Y2=1.465
r80 27 29 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=11.25 $Y=1.63
+ $X2=11.25 $Y2=1.985
r81 23 38 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.25 $Y=1.3
+ $X2=11.25 $Y2=1.465
r82 23 25 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=11.25 $Y=1.3
+ $X2=11.25 $Y2=0.515
r83 19 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.465 $Y=1.3
+ $X2=12.465 $Y2=1.465
r84 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.465 $Y=1.3
+ $X2=12.465 $Y2=0.74
r85 15 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.455 $Y=1.63
+ $X2=12.455 $Y2=1.465
r86 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=12.455 $Y=1.63
+ $X2=12.455 $Y2=2.4
r87 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.035 $Y=1.3
+ $X2=12.035 $Y2=1.465
r88 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.035 $Y=1.3
+ $X2=12.035 $Y2=0.74
r89 7 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.005 $Y=1.63
+ $X2=12.005 $Y2=1.465
r90 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=12.005 $Y=1.63
+ $X2=12.005 $Y2=2.4
r91 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.25 $Y2=2.695
r92 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.25 $Y2=1.985
r93 1 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=11.105
+ $Y=0.37 $X2=11.25 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%A_27_74# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 38
r69 35 38 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.53 $Y=0.76
+ $X2=2.685 $Y2=0.76
r70 31 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.71 $Y=2.145
+ $X2=1.71 $Y2=2.275
r71 27 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=0.76
r72 27 28 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=2.06
r73 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.71 $Y2=2.145
r74 25 42 13.5964 $w=3.32e-07 $l=4.63249e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.655 $Y2=2.515
r75 25 28 6.01991 $w=3.32e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.53 $Y2=2.06
r76 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=1.795 $Y2=2.145
r77 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.275
+ $X2=0.24 $Y2=2.275
r78 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=1.71 $Y2=2.275
r79 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=0.365 $Y2=2.275
r80 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.36 $X2=0.24
+ $Y2=2.275
r81 19 21 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=2.36
+ $X2=0.24 $Y2=2.75
r82 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.24 $Y2=2.275
r83 18 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.2 $Y=2.19 $X2=0.2
+ $Y2=0.81
r84 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.81
r85 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.58
r86 4 42 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.315 $X2=2.78 $Y2=2.515
r87 3 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r88 2 38 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.485 $X2=2.685 $Y2=0.76
r89 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 60 64 66 71 72 74 75 76 78 83 88 93 105 116 120 126 129 132 135 138 141 145
c144 34 0 2.99812e-20 $X=1.74 $Y=2.73
r145 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r146 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r147 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r148 135 136 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r149 132 133 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r152 124 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r153 124 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r154 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r155 121 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.865 $Y=3.33
+ $X2=11.74 $Y2=3.33
r156 121 123 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.865 $Y=3.33
+ $X2=12.24 $Y2=3.33
r157 120 144 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.595 $Y=3.33
+ $X2=12.777 $Y2=3.33
r158 120 123 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.595 $Y=3.33
+ $X2=12.24 $Y2=3.33
r159 119 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r160 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r161 116 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.615 $Y=3.33
+ $X2=11.74 $Y2=3.33
r162 116 118 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.615 $Y=3.33
+ $X2=11.28 $Y2=3.33
r163 115 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r164 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r165 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r166 112 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=9.795 $Y2=3.33
r167 112 114 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=10.32 $Y2=3.33
r168 111 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r169 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r170 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r171 107 110 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r172 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r173 105 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=3.33
+ $X2=9.795 $Y2=3.33
r174 105 110 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.63 $Y=3.33
+ $X2=9.36 $Y2=3.33
r175 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r176 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r177 101 135 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=5.885 $Y2=3.33
r178 101 103 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 100 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r180 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r181 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r182 97 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r184 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r185 94 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.185 $Y2=3.33
r186 94 96 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 93 135 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.885 $Y2=3.33
r188 93 99 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.52 $Y2=3.33
r189 92 133 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r190 92 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r191 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r192 89 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r193 89 91 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r194 88 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=4.185 $Y2=3.33
r195 88 91 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=2.16 $Y2=3.33
r196 87 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r197 87 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r198 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r199 84 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r200 84 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r201 83 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r202 83 86 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 81 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r205 78 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r206 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r207 76 104 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 76 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r209 74 114 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.32 $Y2=3.33
r210 74 75 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.732 $Y2=3.33
r211 73 118 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=11.28 $Y2=3.33
r212 73 75 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=10.732 $Y2=3.33
r213 71 103 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.09 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.09 $Y=3.33
+ $X2=8.175 $Y2=3.33
r215 70 107 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.26 $Y=3.33
+ $X2=8.4 $Y2=3.33
r216 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.26 $Y=3.33
+ $X2=8.175 $Y2=3.33
r217 66 69 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.72 $Y2=2.815
r218 64 144 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.72 $Y=3.245
+ $X2=12.777 $Y2=3.33
r219 64 69 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.72 $Y=3.245
+ $X2=12.72 $Y2=2.815
r220 60 63 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=11.74 $Y=1.985
+ $X2=11.74 $Y2=2.695
r221 58 141 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.74 $Y=3.245
+ $X2=11.74 $Y2=3.33
r222 58 63 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=11.74 $Y=3.245
+ $X2=11.74 $Y2=2.695
r223 54 57 37.059 $w=2.53e-07 $l=8.2e-07 $layer=LI1_cond $X=10.732 $Y=1.985
+ $X2=10.732 $Y2=2.805
r224 52 75 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.732 $Y=3.245
+ $X2=10.732 $Y2=3.33
r225 52 57 19.8853 $w=2.53e-07 $l=4.4e-07 $layer=LI1_cond $X=10.732 $Y=3.245
+ $X2=10.732 $Y2=2.805
r226 48 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=3.245
+ $X2=9.795 $Y2=3.33
r227 48 50 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=9.795 $Y=3.245
+ $X2=9.795 $Y2=2.805
r228 44 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.175 $Y=3.245
+ $X2=8.175 $Y2=3.33
r229 44 46 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.175 $Y=3.245
+ $X2=8.175 $Y2=2.815
r230 40 135 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=3.245
+ $X2=5.885 $Y2=3.33
r231 40 42 17.1309 $w=3.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.885 $Y=3.245
+ $X2=5.885 $Y2=2.695
r232 36 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=3.245
+ $X2=4.185 $Y2=3.33
r233 36 38 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.185 $Y=3.245
+ $X2=4.185 $Y2=2.82
r234 32 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r235 32 34 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.73
r236 28 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r237 28 30 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.755
r238 9 69 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.545
+ $Y=1.84 $X2=12.68 $Y2=2.815
r239 9 66 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.545
+ $Y=1.84 $X2=12.68 $Y2=1.985
r240 8 63 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=11.565
+ $Y=1.84 $X2=11.78 $Y2=2.695
r241 8 60 400 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=11.565
+ $Y=1.84 $X2=11.78 $Y2=1.985
r242 7 57 400 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=10.56
+ $Y=1.84 $X2=10.695 $Y2=2.805
r243 7 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.56
+ $Y=1.84 $X2=10.695 $Y2=1.985
r244 6 50 600 $w=1.7e-07 $l=1.06936e-06 $layer=licon1_PDIFF $count=1 $X=9.575
+ $Y=1.84 $X2=9.795 $Y2=2.805
r245 5 46 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.04
+ $Y=2.54 $X2=8.175 $Y2=2.815
r246 4 42 600 $w=1.7e-07 $l=6.42495e-07 $layer=licon1_PDIFF $count=1 $X=5.405
+ $Y=2.315 $X2=5.885 $Y2=2.695
r247 3 38 600 $w=1.7e-07 $l=6.05083e-07 $layer=licon1_PDIFF $count=1 $X=3.965
+ $Y=2.315 $X2=4.185 $Y2=2.82
r248 2 34 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.79 $X2=1.74 $Y2=2.73
r249 1 30 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.54 $X2=0.73 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%Q_N 1 2 7 8 9 10 11 32
r26 29 32 0.491205 $w=3.03e-07 $l=1.3e-08 $layer=LI1_cond $X=10.282 $Y=1.972
+ $X2=10.282 $Y2=1.985
r27 11 29 0.415635 $w=3.03e-07 $l=1.1e-08 $layer=LI1_cond $X=10.282 $Y=1.961
+ $X2=10.282 $Y2=1.972
r28 11 38 5.61139 $w=3.03e-07 $l=1.41e-07 $layer=LI1_cond $X=10.282 $Y=1.961
+ $X2=10.282 $Y2=1.82
r29 11 35 28.6788 $w=3.03e-07 $l=7.59e-07 $layer=LI1_cond $X=10.282 $Y=2.046
+ $X2=10.282 $Y2=2.805
r30 11 32 2.30489 $w=3.03e-07 $l=6.1e-08 $layer=LI1_cond $X=10.282 $Y=2.046
+ $X2=10.282 $Y2=1.985
r31 10 38 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=10.305 $Y=1.665
+ $X2=10.305 $Y2=1.82
r32 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=10.305 $Y=1.295
+ $X2=10.305 $Y2=1.665
r33 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=10.305 $Y=0.925
+ $X2=10.305 $Y2=1.295
r34 7 8 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=10.305 $Y=0.515
+ $X2=10.305 $Y2=0.925
r35 2 35 400 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.84 $X2=10.245 $Y2=2.805
r36 2 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.84 $X2=10.245 $Y2=1.985
r37 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.12
+ $Y=0.37 $X2=10.26 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%Q 1 2 9 14 15 16 17 28
c33 15 0 8.81429e-20 $X=12.245 $Y=1.82
r34 21 28 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=12.255 $Y=0.96
+ $X2=12.255 $Y2=0.925
r35 17 30 7.79401 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=12.255 $Y=0.985
+ $X2=12.255 $Y2=1.13
r36 17 21 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=12.255 $Y=0.985
+ $X2=12.255 $Y2=0.96
r37 17 28 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=12.255 $Y=0.9
+ $X2=12.255 $Y2=0.925
r38 16 17 13.0497 $w=3.38e-07 $l=3.85e-07 $layer=LI1_cond $X=12.255 $Y=0.515
+ $X2=12.255 $Y2=0.9
r39 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.34 $Y=1.82
+ $X2=12.34 $Y2=1.13
r40 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=1.985
+ $X2=12.245 $Y2=1.82
r41 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=12.245 $Y=2
+ $X2=12.245 $Y2=1.985
r42 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=12.245 $Y=2 $X2=12.245
+ $Y2=2.815
r43 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.095
+ $Y=1.84 $X2=12.23 $Y2=1.985
r44 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.095
+ $Y=1.84 $X2=12.23 $Y2=2.815
r45 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.11
+ $Y=0.37 $X2=12.25 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_2%VGND 1 2 3 4 5 6 7 8 9 30 32 36 40 44 48 52
+ 54 56 59 60 61 63 68 89 98 102 108 111 114 119 125 129 132 134 137 141
c142 36 0 1.39813e-19 $X=1.7 $Y=0.505
r143 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r144 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r145 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r146 131 132 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=0.292
+ $X2=8.845 $Y2=0.292
r147 127 131 4.43579 $w=7.53e-07 $l=2.8e-07 $layer=LI1_cond $X=8.4 $Y=0.292
+ $X2=8.68 $Y2=0.292
r148 127 129 13.2931 $w=7.53e-07 $l=3e-07 $layer=LI1_cond $X=8.4 $Y=0.292
+ $X2=8.1 $Y2=0.292
r149 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r150 123 125 11.1389 $w=7.63e-07 $l=1.6e-07 $layer=LI1_cond $X=6 $Y=0.297
+ $X2=6.16 $Y2=0.297
r151 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r152 121 123 0.0781751 $w=7.63e-07 $l=5e-09 $layer=LI1_cond $X=5.995 $Y=0.297
+ $X2=6 $Y2=0.297
r153 118 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r154 117 121 7.42663 $w=7.63e-07 $l=4.75e-07 $layer=LI1_cond $X=5.52 $Y=0.297
+ $X2=5.995 $Y2=0.297
r155 117 119 11.4516 $w=7.63e-07 $l=1.8e-07 $layer=LI1_cond $X=5.52 $Y=0.297
+ $X2=5.34 $Y2=0.297
r156 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r158 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r159 109 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r160 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r161 106 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r162 106 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r163 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r164 103 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=11.75 $Y2=0
r165 103 105 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=12.24 $Y2=0
r166 102 140 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.595 $Y=0
+ $X2=12.777 $Y2=0
r167 102 105 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.595 $Y=0
+ $X2=12.24 $Y2=0
r168 101 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r169 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r170 98 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.75 $Y2=0
r171 98 100 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.28 $Y2=0
r172 97 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r173 97 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r174 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r175 94 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.995 $Y=0
+ $X2=9.83 $Y2=0
r176 94 96 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.995 $Y=0
+ $X2=10.32 $Y2=0
r177 93 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r178 93 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.4
+ $Y2=0
r179 92 132 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=8.845 $Y2=0
r180 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r181 89 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.83 $Y2=0
r182 89 92 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.36 $Y2=0
r183 88 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r184 87 129 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=8.1
+ $Y2=0
r185 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r186 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r187 84 125 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.16
+ $Y2=0
r188 80 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r189 80 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.08 $Y2=0
r190 79 119 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.34
+ $Y2=0
r191 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r192 77 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=0
+ $X2=4.115 $Y2=0
r193 77 79 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=5.04
+ $Y2=0
r194 75 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r195 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r196 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r197 72 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r198 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r199 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r200 69 111 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.735 $Y2=0
r201 69 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r202 68 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=0
+ $X2=4.115 $Y2=0
r203 68 74 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.6
+ $Y2=0
r204 66 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r205 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r206 63 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.67 $Y2=0
r207 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r208 61 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r209 61 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r210 61 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r211 59 96 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=0
+ $X2=10.32 $Y2=0
r212 59 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.605 $Y=0
+ $X2=10.73 $Y2=0
r213 58 100 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.855 $Y=0
+ $X2=11.28 $Y2=0
r214 58 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.855 $Y=0
+ $X2=10.73 $Y2=0
r215 54 140 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.72 $Y=0.085
+ $X2=12.777 $Y2=0
r216 54 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.72 $Y=0.085
+ $X2=12.72 $Y2=0.515
r217 50 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.75 $Y=0.085
+ $X2=11.75 $Y2=0
r218 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.75 $Y=0.085
+ $X2=11.75 $Y2=0.515
r219 46 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0
r220 46 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0.515
r221 42 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=0.085
+ $X2=9.83 $Y2=0
r222 42 44 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.83 $Y=0.085
+ $X2=9.83 $Y2=0.675
r223 38 114 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=0.085
+ $X2=4.115 $Y2=0
r224 38 40 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=4.115 $Y=0.085
+ $X2=4.115 $Y2=0.655
r225 34 111 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r226 34 36 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.505
r227 33 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.67 $Y2=0
r228 32 111 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=1.735 $Y2=0
r229 32 33 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.795 $Y2=0
r230 28 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r231 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r232 9 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.54
+ $Y=0.37 $X2=12.68 $Y2=0.515
r233 8 52 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=11.54
+ $Y=0.37 $X2=11.75 $Y2=0.515
r234 7 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.55
+ $Y=0.37 $X2=10.69 $Y2=0.515
r235 6 44 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=9.685
+ $Y=0.37 $X2=9.83 $Y2=0.675
r236 5 131 91 $w=1.7e-07 $l=6.76166e-07 $layer=licon1_NDIFF $count=2 $X=8.045
+ $Y=0.59 $X2=8.68 $Y2=0.505
r237 4 121 91 $w=1.7e-07 $l=6.98749e-07 $layer=licon1_NDIFF $count=2 $X=5.365
+ $Y=0.37 $X2=5.995 $Y2=0.515
r238 3 40 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.485 $X2=4.155 $Y2=0.655
r239 2 36 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.505
r240 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__nor3b_2.spice
* Created: Fri Aug 28 17:48:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor3b_2.pex.spice"
.subckt sky130_fd_sc_ms__nor3b_2  VNB VPB C_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_N_M1008_g N_A_27_392#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1008_d N_A_27_392#_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157545 AS=0.10915 PD=1.24406 PS=1.035 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_27_392#_M1012_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2664 AS=0.10915 PD=1.46 PS=1.035 NRD=0 NRS=2.424 M=1 R=4.93333 SA=75001.1
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2664 PD=1.02 PS=1.46 NRD=0 NRS=0 M=1 R=4.93333 SA=75002 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1001_d N_B_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.3108 PD=1.02 PS=1.58 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.3108 PD=1.07 PS=1.58 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1002_d N_A_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.2257 PD=1.07 PS=2.09 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75003.9 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_C_N_M1003_g N_A_27_392#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.275 AS=0.275 PD=2.55 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_Y_M1005_d N_A_27_392#_M1005_g N_A_227_368#_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1005_d N_A_27_392#_M1006_g N_A_227_368#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_A_498_368#_M1007_d N_B_M1007_g N_A_227_368#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_A_498_368#_M1007_d N_B_M1010_g N_A_227_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1009 N_A_498_368#_M1009_d N_A_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_A_498_368#_M1009_d N_A_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__nor3b_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__xor3_1.pex.spice
* Created: Fri Aug 28 18:19:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_84_108# 1 2 3 4 15 19 23 24 26 27 31 36 38
+ 39 41 44 46 47 52
r114 50 52 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.15 $Y=1.1 $X2=4.31
+ $Y2=1.1
r115 46 48 19.8947 $w=6.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.06 $Y=2.07
+ $X2=4.06 $Y2=2.755
r116 46 47 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=2.07
+ $X2=4.06 $Y2=1.905
r117 42 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=1.265
+ $X2=4.31 $Y2=1.1
r118 42 47 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.31 $Y=1.265
+ $X2=4.31 $Y2=1.905
r119 41 48 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.755
r120 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=2.99
+ $X2=3.81 $Y2=2.905
r121 38 39 132.112 $w=1.68e-07 $l=2.025e-06 $layer=LI1_cond $X=3.725 $Y=2.99
+ $X2=1.7 $Y2=2.99
r122 34 44 3.70735 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=1.54 $Y=1.92
+ $X2=1.37 $Y2=1.92
r123 34 36 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.54 $Y=1.92
+ $X2=1.54 $Y2=1.165
r124 31 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.535 $Y=2.105
+ $X2=1.535 $Y2=2.815
r125 29 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.535 $Y=2.905
+ $X2=1.7 $Y2=2.99
r126 29 33 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.535 $Y=2.905
+ $X2=1.535 $Y2=2.815
r127 28 44 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=1.535 $Y=2.09
+ $X2=1.37 $Y2=1.92
r128 28 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.535 $Y=2.09
+ $X2=1.535 $Y2=2.105
r129 26 44 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.005
+ $X2=1.37 $Y2=1.92
r130 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.37 $Y=2.005
+ $X2=0.75 $Y2=2.005
r131 24 56 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.635
+ $X2=0.585 $Y2=1.8
r132 24 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.635
+ $X2=0.585 $Y2=1.47
r133 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.635 $X2=0.585 $Y2=1.635
r134 21 27 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=0.587 $Y=1.92
+ $X2=0.75 $Y2=2.005
r135 21 23 10.106 $w=3.23e-07 $l=2.85e-07 $layer=LI1_cond $X=0.587 $Y=1.92
+ $X2=0.587 $Y2=1.635
r136 19 56 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.66 $Y=2.46
+ $X2=0.66 $Y2=1.8
r137 15 55 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.99
+ $X2=0.495 $Y2=1.47
r138 4 46 300 $w=1.7e-07 $l=4.43959e-07 $layer=licon1_PDIFF $count=2 $X=3.445
+ $Y=1.895 $X2=3.81 $Y2=2.07
r139 3 33 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.4
+ $Y=1.96 $X2=1.535 $Y2=2.815
r140 3 31 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=1.96 $X2=1.535 $Y2=2.105
r141 2 50 182 $w=1.7e-07 $l=6.10635e-07 $layer=licon1_NDIFF $count=1 $X=3.84
+ $Y=0.625 $X2=4.15 $Y2=1.1
r142 1 36 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.67 $X2=1.54 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A 3 5 7 8 15
c36 3 0 1.7856e-19 $X=1.31 $Y=2.46
r37 14 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.31 $Y=1.585
+ $X2=1.325 $Y2=1.585
r38 11 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.125 $Y=1.585
+ $X2=1.31 $Y2=1.585
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.125
+ $Y=1.585 $X2=1.125 $Y2=1.585
r40 8 12 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.122 $Y=1.295
+ $X2=1.122 $Y2=1.585
r41 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.325 $Y2=1.585
r42 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.325 $Y2=0.99
r43 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.75
+ $X2=1.31 $Y2=1.585
r44 1 3 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.31 $Y=1.75 $X2=1.31
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_452_288# 1 2 9 13 15 16 19 25 30 32 33 34
+ 38 41 48 49 51 53
c109 9 0 1.75672e-19 $X=2.35 $Y=2.28
r110 52 53 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.57
+ $X2=3.69 $Y2=1.57
r111 49 52 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.89 $Y=1.57
+ $X2=3.765 $Y2=1.57
r112 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.57 $X2=3.89 $Y2=1.57
r113 45 48 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=3.81 $Y=1.585
+ $X2=3.89 $Y2=1.585
r114 41 43 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.665 $Y=1.985
+ $X2=4.665 $Y2=2.815
r115 41 51 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.665 $Y=1.985
+ $X2=4.665 $Y2=1.13
r116 36 51 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=4.692 $Y=1.018
+ $X2=4.692 $Y2=1.13
r117 36 38 8.09271 $w=2.23e-07 $l=1.58e-07 $layer=LI1_cond $X=4.692 $Y=1.018
+ $X2=4.692 $Y2=0.86
r118 35 38 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=4.692 $Y=0.765
+ $X2=4.692 $Y2=0.86
r119 33 35 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.58 $Y=0.68
+ $X2=4.692 $Y2=0.765
r120 33 34 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.58 $Y=0.68
+ $X2=3.895 $Y2=0.68
r121 32 45 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.81 $Y=1.435 $X2=3.81
+ $Y2=1.585
r122 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.765
+ $X2=3.895 $Y2=0.68
r123 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.81 $Y=0.765
+ $X2=3.81 $Y2=1.435
r124 23 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.405
+ $X2=3.765 $Y2=1.57
r125 23 25 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.765 $Y=1.405
+ $X2=3.765 $Y2=0.945
r126 22 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.445 $Y=1.515
+ $X2=3.355 $Y2=1.515
r127 22 53 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.445 $Y=1.515
+ $X2=3.69 $Y2=1.515
r128 17 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.355 $Y=1.59
+ $X2=3.355 $Y2=1.515
r129 17 19 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=3.355 $Y=1.59
+ $X2=3.355 $Y2=2.315
r130 16 29 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.515
+ $X2=2.505 $Y2=1.515
r131 15 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.265 $Y=1.515
+ $X2=3.355 $Y2=1.515
r132 15 16 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.265 $Y=1.515
+ $X2=2.58 $Y2=1.515
r133 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=1.44
+ $X2=2.505 $Y2=1.515
r134 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.505 $Y=1.44
+ $X2=2.505 $Y2=0.86
r135 7 29 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.35 $Y=1.515
+ $X2=2.505 $Y2=1.515
r136 7 9 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=2.35 $Y=1.59 $X2=2.35
+ $Y2=2.28
r137 2 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.84 $X2=4.665 $Y2=2.815
r138 2 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.84 $X2=4.665 $Y2=1.985
r139 1 38 182 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.37 $X2=4.72 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%B 3 7 9 10 11 12 15 17 21 23 26 28 33 37 39
+ 40 41 42 45 48 49
c136 21 0 1.96802e-19 $X=3.175 $Y=0.75
c137 7 0 1.59849e-19 $X=2.005 $Y=0.75
r138 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.085
+ $Y=1.515 $X2=5.085 $Y2=1.515
r139 46 48 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.935 $Y=1.515
+ $X2=5.085 $Y2=1.515
r140 44 46 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=4.89 $Y=1.515
+ $X2=4.935 $Y2=1.515
r141 44 45 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.89 $Y=1.515 $X2=4.8
+ $Y2=1.515
r142 42 49 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.085 $Y=1.665
+ $X2=5.085 $Y2=1.515
r143 35 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.35
+ $X2=4.935 $Y2=1.515
r144 35 37 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.935 $Y=1.35
+ $X2=4.935 $Y2=0.74
r145 31 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.68
+ $X2=4.89 $Y2=1.515
r146 31 33 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.89 $Y=1.68
+ $X2=4.89 $Y2=2.4
r147 30 41 5.30422 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=4.51 $Y=1.425
+ $X2=4.402 $Y2=1.425
r148 30 45 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.51 $Y=1.425
+ $X2=4.8 $Y2=1.425
r149 28 41 20.4101 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.435 $Y=1.35
+ $X2=4.402 $Y2=1.425
r150 27 28 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=4.435 $Y=0.255
+ $X2=4.435 $Y2=1.35
r151 25 41 20.4101 $w=1.5e-07 $l=8.95824e-08 $layer=POLY_cond $X=4.37 $Y=1.5
+ $X2=4.402 $Y2=1.425
r152 25 26 807.606 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=4.37 $Y=1.5
+ $X2=4.37 $Y2=3.075
r153 24 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.25 $Y=0.18
+ $X2=3.175 $Y2=0.18
r154 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.36 $Y=0.18
+ $X2=4.435 $Y2=0.255
r155 23 24 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=4.36 $Y=0.18
+ $X2=3.25 $Y2=0.18
r156 19 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.175 $Y=0.255
+ $X2=3.175 $Y2=0.18
r157 19 21 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.175 $Y=0.255
+ $X2=3.175 $Y2=0.75
r158 18 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.91 $Y=3.15 $X2=2.82
+ $Y2=3.15
r159 17 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.295 $Y=3.15
+ $X2=4.37 $Y2=3.075
r160 17 18 710.181 $w=1.5e-07 $l=1.385e-06 $layer=POLY_cond $X=4.295 $Y=3.15
+ $X2=2.91 $Y2=3.15
r161 13 39 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.82 $Y=3.075
+ $X2=2.82 $Y2=3.15
r162 13 15 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=2.82 $Y=3.075
+ $X2=2.82 $Y2=2.28
r163 11 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=0.18
+ $X2=3.175 $Y2=0.18
r164 11 12 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.1 $Y=0.18
+ $X2=2.08 $Y2=0.18
r165 9 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.73 $Y=3.15 $X2=2.82
+ $Y2=3.15
r166 9 10 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.73 $Y=3.15
+ $X2=1.935 $Y2=3.15
r167 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.08 $Y2=0.18
r168 5 7 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.005 $Y2=0.75
r169 1 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.845 $Y=3.075
+ $X2=1.935 $Y2=3.15
r170 1 3 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=1.845 $Y=3.075
+ $X2=1.845 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_1157_298# 1 2 9 13 16 17 18 20 23 26 31 37
+ 39 43
c91 23 0 1.49313e-19 $X=7.9 $Y=0.63
c92 13 0 1.40824e-19 $X=6.155 $Y=0.925
r93 42 43 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=6 $Y=1.655
+ $X2=6.155 $Y2=1.655
r94 36 37 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.65 $Y=2.36 $X2=7.9
+ $Y2=2.36
r95 33 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.52 $Y=2.36
+ $X2=7.65 $Y2=2.36
r96 29 42 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.97 $Y=1.655 $X2=6
+ $Y2=1.655
r97 28 31 5.56352 $w=2.88e-07 $l=1.4e-07 $layer=LI1_cond $X=5.97 $Y=1.675
+ $X2=6.11 $Y2=1.675
r98 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.97
+ $Y=1.655 $X2=5.97 $Y2=1.655
r99 26 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.9 $Y=2.195 $X2=7.9
+ $Y2=2.36
r100 26 39 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=7.9 $Y=2.195
+ $X2=7.9 $Y2=0.86
r101 21 39 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.94 $Y=0.735
+ $X2=7.94 $Y2=0.86
r102 21 23 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=7.94 $Y=0.735
+ $X2=7.94 $Y2=0.63
r103 19 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.52 $Y=2.525
+ $X2=7.52 $Y2=2.36
r104 19 20 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.52 $Y=2.525
+ $X2=7.52 $Y2=2.905
r105 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.435 $Y=2.99
+ $X2=7.52 $Y2=2.905
r106 17 18 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.435 $Y=2.99
+ $X2=6.195 $Y2=2.99
r107 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.11 $Y=2.905
+ $X2=6.195 $Y2=2.99
r108 15 31 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.11 $Y=1.82
+ $X2=6.11 $Y2=1.675
r109 15 16 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=6.11 $Y=1.82
+ $X2=6.11 $Y2=2.905
r110 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.49
+ $X2=6.155 $Y2=1.655
r111 11 13 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.155 $Y=1.49
+ $X2=6.155 $Y2=0.925
r112 7 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6 $Y=1.82 $X2=6
+ $Y2=1.655
r113 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6 $Y=1.82 $X2=6
+ $Y2=2.4
r114 2 36 600 $w=1.7e-07 $l=5.84423e-07 $layer=licon1_PDIFF $count=1 $X=7.455
+ $Y=1.865 $X2=7.65 $Y2=2.36
r115 1 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.755
+ $Y=0.42 $X2=7.9 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%C 3 5 7 8 9 11 14 16 18 21 23 24
r87 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.04
+ $Y=1.52 $X2=7.04 $Y2=1.52
r88 27 29 33.1577 $w=2.98e-07 $l=2.05e-07 $layer=POLY_cond $X=6.835 $Y=1.52
+ $X2=7.04 $Y2=1.52
r89 24 30 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.04 $Y=1.295
+ $X2=7.04 $Y2=1.52
r90 19 21 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=7.91 $Y=0.99
+ $X2=8.115 $Y2=0.99
r91 16 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.115 $Y=0.915
+ $X2=8.115 $Y2=0.99
r92 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.115 $Y=0.915
+ $X2=8.115 $Y2=0.63
r93 12 23 18.8402 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=7.925 $Y=1.595
+ $X2=7.835 $Y2=1.355
r94 12 14 229.339 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=7.925 $Y=1.595
+ $X2=7.925 $Y2=2.185
r95 11 23 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.91 $Y=1.355
+ $X2=7.835 $Y2=1.355
r96 10 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.91 $Y=1.065
+ $X2=7.91 $Y2=0.99
r97 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.91 $Y=1.065
+ $X2=7.91 $Y2=1.355
r98 9 29 38.561 $w=2.98e-07 $l=2.05122e-07 $layer=POLY_cond $X=7.205 $Y=1.43
+ $X2=7.04 $Y2=1.52
r99 8 23 6.66866 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.835 $Y=1.43
+ $X2=7.835 $Y2=1.355
r100 8 9 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=7.835 $Y=1.43
+ $X2=7.205 $Y2=1.43
r101 5 27 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.835 $Y=1.355
+ $X2=6.835 $Y2=1.52
r102 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.835 $Y=1.355
+ $X2=6.835 $Y2=0.925
r103 1 27 12.9396 $w=2.98e-07 $l=2.0106e-07 $layer=POLY_cond $X=6.755 $Y=1.685
+ $X2=6.835 $Y2=1.52
r104 1 3 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=6.755 $Y=1.685
+ $X2=6.755 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_1218_396# 1 2 9 13 17 21 23 24 27 30 35 36
c86 13 0 1.49313e-19 $X=8.625 $Y=0.79
r87 36 37 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.515
+ $X2=8.625 $Y2=1.515
r88 34 36 28.6555 $w=3.28e-07 $l=1.95e-07 $layer=POLY_cond $X=8.42 $Y=1.515
+ $X2=8.615 $Y2=1.515
r89 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.42
+ $Y=1.515 $X2=8.42 $Y2=1.515
r90 30 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665 $X2=8.4
+ $Y2=1.665
r91 27 42 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=6.535 $Y=1.665
+ $X2=6.535 $Y2=1.55
r92 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r93 24 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.665
+ $X2=6.48 $Y2=1.665
r94 23 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r95 23 24 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=6.625 $Y2=1.665
r96 21 42 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.62 $Y=1.1 $X2=6.62
+ $Y2=1.55
r97 15 27 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=1.665
r98 15 17 13.7276 $w=3.38e-07 $l=4.05e-07 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=2.125
r99 11 37 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=1.515
r100 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=0.79
r101 7 36 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.68
+ $X2=8.615 $Y2=1.515
r102 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.615 $Y=1.68
+ $X2=8.615 $Y2=2.4
r103 2 17 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=6.09
+ $Y=1.98 $X2=6.53 $Y2=2.125
r104 1 21 182 $w=1.7e-07 $l=6.61872e-07 $layer=licon1_NDIFF $count=1 $X=6.23
+ $Y=0.605 $X2=6.62 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_27_134# 1 2 3 4 13 14 17 20 21 22 25 29 32
+ 35 37 38 40 41
r85 37 38 9.60999 $w=5.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.342 $Y=2.425
+ $X2=0.342 $Y2=2.26
r86 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.17 $Y=1.3 $X2=0.17
+ $Y2=2.26
r87 32 40 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.675 $Y=1.26
+ $X2=2.595 $Y2=1.345
r88 32 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.675 $Y=1.26
+ $X2=2.675 $Y2=1.09
r89 27 41 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.72 $Y=0.96
+ $X2=2.72 $Y2=1.09
r90 27 29 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=2.72 $Y=0.96 $X2=2.72
+ $Y2=0.86
r91 23 40 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.43
+ $X2=2.595 $Y2=1.345
r92 23 25 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=2.595 $Y=1.43
+ $X2=2.595 $Y2=2.205
r93 21 40 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=1.345
+ $X2=2.595 $Y2=1.345
r94 21 22 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.43 $Y=1.345
+ $X2=1.965 $Y2=1.345
r95 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.88 $Y=1.26
+ $X2=1.965 $Y2=1.345
r96 19 20 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.88 $Y=0.83
+ $X2=1.88 $Y2=1.26
r97 18 34 5.39736 $w=1.7e-07 $l=1.82483e-07 $layer=LI1_cond $X=0.445 $Y=0.745
+ $X2=0.265 $Y2=0.74
r98 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=0.745
+ $X2=1.88 $Y2=0.83
r99 17 18 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=1.795 $Y=0.745
+ $X2=0.445 $Y2=0.745
r100 14 35 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1.12
+ $X2=0.265 $Y2=1.3
r101 13 34 2.62574 $w=3.6e-07 $l=9e-08 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.74
r102 13 14 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=1.12
r103 4 25 600 $w=1.7e-07 $l=3.1305e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.96 $X2=2.595 $Y2=2.205
r104 3 37 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=0.29
+ $Y=1.96 $X2=0.435 $Y2=2.425
r105 2 29 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.65 $X2=2.765 $Y2=0.86
r106 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.67 $X2=0.28 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%VPWR 1 2 3 12 16 22 27 28 29 35 42 52 53 56
+ 59
r76 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r77 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r78 53 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r79 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r80 50 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.39 $Y2=3.33
r81 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.88 $Y2=3.33
r82 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r83 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r84 46 49 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r85 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 45 48 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r87 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 43 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.075 $Y2=3.33
r89 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.2 $Y=3.33 $X2=5.52
+ $Y2=3.33
r90 42 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=3.33
+ $X2=8.39 $Y2=3.33
r91 42 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.225 $Y=3.33
+ $X2=7.92 $Y2=3.33
r92 37 40 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 37 38 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r94 35 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.95 $Y=3.33
+ $X2=5.075 $Y2=3.33
r95 35 40 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.95 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 33 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 29 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r99 29 38 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r100 29 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r101 27 32 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=3.33 $X2=0.72
+ $Y2=3.33
r102 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=3.33
+ $X2=0.935 $Y2=3.33
r103 26 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r104 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.935 $Y2=3.33
r105 22 25 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.39 $Y=2.115
+ $X2=8.39 $Y2=2.465
r106 20 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=3.245
+ $X2=8.39 $Y2=3.33
r107 20 25 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.39 $Y=3.245
+ $X2=8.39 $Y2=2.465
r108 16 19 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.075 $Y=2.115
+ $X2=5.075 $Y2=2.815
r109 14 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=3.33
r110 14 19 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=2.815
r111 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=3.33
r112 10 12 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=2.425
r113 3 25 300 $w=1.7e-07 $l=7.64853e-07 $layer=licon1_PDIFF $count=2 $X=8.015
+ $Y=1.865 $X2=8.39 $Y2=2.465
r114 3 22 600 $w=1.7e-07 $l=4.84123e-07 $layer=licon1_PDIFF $count=1 $X=8.015
+ $Y=1.865 $X2=8.39 $Y2=2.115
r115 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.84 $X2=5.115 $Y2=2.815
r116 2 16 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.84 $X2=5.115 $Y2=2.115
r117 1 12 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=0.75
+ $Y=1.96 $X2=0.935 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_387_392# 1 2 3 4 15 17 18 22 23 24 26 27 28
+ 32 33 34 37 39 40 42
c127 15 0 3.54233e-19 $X=2.095 $Y=2.105
r128 41 42 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.56 $Y=0.425
+ $X2=7.56 $Y2=1.855
r129 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=1.94
+ $X2=7.56 $Y2=1.855
r130 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.475 $Y=1.94
+ $X2=7.205 $Y2=1.94
r131 35 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.04 $Y=2.025
+ $X2=7.205 $Y2=1.94
r132 35 37 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=7.04 $Y=2.025
+ $X2=7.04 $Y2=2.125
r133 33 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=0.34
+ $X2=7.56 $Y2=0.425
r134 33 34 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=7.475 $Y=0.34
+ $X2=6.025 $Y2=0.34
r135 30 32 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=5.9 $Y=0.85 $X2=5.9
+ $Y2=0.8
r136 29 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.9 $Y=0.425
+ $X2=6.025 $Y2=0.34
r137 29 32 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=5.9 $Y=0.425
+ $X2=5.9 $Y2=0.8
r138 27 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.775 $Y=0.935
+ $X2=5.9 $Y2=0.85
r139 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.775 $Y=0.935
+ $X2=5.145 $Y2=0.935
r140 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=0.85
+ $X2=5.145 $Y2=0.935
r141 25 26 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.06 $Y=0.425
+ $X2=5.06 $Y2=0.85
r142 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=5.06 $Y2=0.425
r143 23 24 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=3.555 $Y2=0.34
r144 20 22 129.829 $w=1.68e-07 $l=1.99e-06 $layer=LI1_cond $X=3.47 $Y=2.565
+ $X2=3.47 $Y2=0.575
r145 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=0.425
+ $X2=3.555 $Y2=0.34
r146 19 22 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.47 $Y=0.425
+ $X2=3.47 $Y2=0.575
r147 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=2.65
+ $X2=3.47 $Y2=2.565
r148 17 18 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=3.385 $Y=2.65
+ $X2=2.26 $Y2=2.65
r149 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.095 $Y=2.565
+ $X2=2.26 $Y2=2.65
r150 13 15 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.095 $Y=2.565
+ $X2=2.095 $Y2=2.105
r151 4 37 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=6.845
+ $Y=1.98 $X2=7.04 $Y2=2.125
r152 3 15 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=1.935
+ $Y=1.96 $X2=2.095 $Y2=2.105
r153 2 32 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.605 $X2=5.94 $Y2=0.8
r154 1 22 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=3.25
+ $Y=0.43 $X2=3.47 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%A_416_86# 1 2 3 4 15 19 20 21 23 27 28 30 32
+ 38 41 42 44 45 48 51 52
c129 45 0 1.96802e-19 $X=3.265 $Y=1.665
c130 41 0 1.40824e-19 $X=7.095 $Y=0.76
c131 15 0 1.59849e-19 $X=2.22 $Y=0.575
r132 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r133 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r134 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r135 44 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=5.52 $Y2=1.665
r136 44 45 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=3.265 $Y2=1.665
r137 41 42 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.095 $Y=0.76
+ $X2=6.885 $Y2=0.76
r138 39 52 16.5011 $w=2.03e-07 $l=3.05e-07 $layer=LI1_cond $X=5.522 $Y=1.36
+ $X2=5.522 $Y2=1.665
r139 36 52 15.4191 $w=2.03e-07 $l=2.85e-07 $layer=LI1_cond $X=5.522 $Y=1.95
+ $X2=5.522 $Y2=1.665
r140 36 38 8.27032 $w=4.15e-07 $l=2.22542e-07 $layer=LI1_cond $X=5.522 $Y=1.95
+ $X2=5.63 $Y2=2.125
r141 35 48 68.5361 $w=1.93e-07 $l=1.205e-06 $layer=LI1_cond $X=3.117 $Y=0.46
+ $X2=3.117 $Y2=1.665
r142 34 48 11.9441 $w=1.93e-07 $l=2.1e-07 $layer=LI1_cond $X=3.117 $Y=1.875
+ $X2=3.117 $Y2=1.665
r143 32 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.365 $Y=0.68
+ $X2=6.885 $Y2=0.68
r144 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.28 $Y=0.765
+ $X2=6.365 $Y2=0.68
r145 29 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.28 $Y=0.765
+ $X2=6.28 $Y2=1.19
r146 28 39 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=5.625 $Y=1.275
+ $X2=5.522 $Y2=1.36
r147 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.195 $Y=1.275
+ $X2=6.28 $Y2=1.19
r148 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.195 $Y=1.275
+ $X2=5.625 $Y2=1.275
r149 21 34 6.35106 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=2 $X2=3.09
+ $Y2=1.875
r150 21 23 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.09 $Y=2 $X2=3.09
+ $Y2=2.135
r151 19 35 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=3.02 $Y=0.375
+ $X2=3.117 $Y2=0.46
r152 19 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.02 $Y=0.375
+ $X2=2.385 $Y2=0.375
r153 15 17 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=2.26 $Y=0.575
+ $X2=2.26 $Y2=0.925
r154 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.26 $Y=0.46
+ $X2=2.385 $Y2=0.375
r155 13 15 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.26 $Y=0.46
+ $X2=2.26 $Y2=0.575
r156 4 38 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.545
+ $Y=1.98 $X2=5.69 $Y2=2.125
r157 3 23 600 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=1.96 $X2=3.13 $Y2=2.135
r158 2 41 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.91
+ $Y=0.605 $X2=7.095 $Y2=0.76
r159 1 17 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.43 $X2=2.22 $Y2=0.925
r160 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.43 $X2=2.22 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%X 1 2 7 8 9 10 11 12 13
r12 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=2.405
+ $X2=8.88 $Y2=2.775
r13 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.405
r14 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.985
r15 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.665
r16 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=0.925 $X2=8.88
+ $Y2=1.295
r17 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=0.555 $X2=8.88
+ $Y2=0.925
r18 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.815
r19 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=1.985
r20 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7 $Y=0.42
+ $X2=8.84 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__XOR3_1%VGND 1 2 3 12 16 20 27 35 42 43 48 51 53 56
r71 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r72 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r73 50 51 12.4896 $w=5.73e-07 $l=2.85e-07 $layer=LI1_cond $X=0.91 $Y=0.202
+ $X2=1.195 $Y2=0.202
r74 46 50 3.95226 $w=5.73e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=0.202
+ $X2=0.91 $Y2=0.202
r75 46 48 8.53733 $w=5.73e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=0.202
+ $X2=0.625 $Y2=0.202
r76 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 43 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r78 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r79 40 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.575 $Y=0 $X2=8.41
+ $Y2=0
r80 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.575 $Y=0 $X2=8.88
+ $Y2=0
r81 39 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r82 39 54 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=0 $X2=5.52
+ $Y2=0
r83 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r84 36 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.44
+ $Y2=0
r85 36 38 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=7.92 $Y2=0
r86 35 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.41
+ $Y2=0
r87 35 38 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=7.92
+ $Y2=0
r88 34 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r89 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r90 31 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r91 30 33 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r92 30 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.195
+ $Y2=0
r93 30 31 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r94 27 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.44
+ $Y2=0
r95 27 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r96 25 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r97 24 48 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.625
+ $Y2=0
r98 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r99 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r100 20 31 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r101 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.41 $Y=0.565
+ $X2=8.41 $Y2=1.015
r102 14 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0
r103 14 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0.565
r104 10 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0
r105 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0.515
r106 3 18 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.42 $X2=8.41 $Y2=1.015
r107 3 16 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.42 $X2=8.41 $Y2=0.565
r108 2 12 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.37 $X2=5.4 $Y2=0.515
r109 1 50 182 $w=1.7e-07 $l=4.86133e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.67 $X2=0.91 $Y2=0.325
.ends


* File: sky130_fd_sc_ms__xnor3_2.pxi.spice
* Created: Fri Aug 28 18:18:15 2020
* 
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_83_247# N_A_83_247#_M1010_d N_A_83_247#_M1002_d
+ N_A_83_247#_M1022_d N_A_83_247#_M1001_d N_A_83_247#_M1015_g
+ N_A_83_247#_M1012_g N_A_83_247#_c_176_n N_A_83_247#_c_177_n
+ N_A_83_247#_c_178_n N_A_83_247#_c_179_n N_A_83_247#_c_189_p
+ N_A_83_247#_c_261_p N_A_83_247#_c_197_p N_A_83_247#_c_190_p
+ N_A_83_247#_c_185_n N_A_83_247#_c_180_n N_A_83_247#_c_186_n
+ N_A_83_247#_c_187_n N_A_83_247#_c_181_n N_A_83_247#_c_182_n
+ N_A_83_247#_c_188_n PM_SKY130_FD_SC_MS__XNOR3_2%A_83_247#
x_PM_SKY130_FD_SC_MS__XNOR3_2%A N_A_M1022_g N_A_M1010_g A N_A_c_306_n
+ N_A_c_307_n PM_SKY130_FD_SC_MS__XNOR3_2%A
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_397_21# N_A_397_21#_M1016_s N_A_397_21#_M1021_s
+ N_A_397_21#_M1004_g N_A_397_21#_c_351_n N_A_397_21#_M1011_g
+ N_A_397_21#_c_353_n N_A_397_21#_c_354_n N_A_397_21#_M1002_g
+ N_A_397_21#_M1001_g N_A_397_21#_c_363_n N_A_397_21#_c_356_n
+ N_A_397_21#_c_357_n N_A_397_21#_c_376_n N_A_397_21#_c_364_n
+ N_A_397_21#_c_358_n N_A_397_21#_c_359_n N_A_397_21#_c_360_n
+ PM_SKY130_FD_SC_MS__XNOR3_2%A_397_21#
x_PM_SKY130_FD_SC_MS__XNOR3_2%B N_B_M1018_g N_B_c_468_n N_B_M1000_g N_B_c_476_n
+ N_B_c_477_n N_B_M1003_g N_B_M1014_g N_B_c_479_n N_B_c_480_n N_B_M1016_g
+ N_B_M1021_g N_B_c_472_n N_B_c_482_n B N_B_c_473_n N_B_c_474_n
+ PM_SKY130_FD_SC_MS__XNOR3_2%B
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_1027_48# N_A_1027_48#_M1013_s
+ N_A_1027_48#_M1020_s N_A_1027_48#_M1023_g N_A_1027_48#_M1005_g
+ N_A_1027_48#_c_590_n N_A_1027_48#_c_591_n N_A_1027_48#_c_592_n
+ N_A_1027_48#_c_598_n N_A_1027_48#_c_593_n N_A_1027_48#_c_594_n
+ N_A_1027_48#_c_600_n PM_SKY130_FD_SC_MS__XNOR3_2%A_1027_48#
x_PM_SKY130_FD_SC_MS__XNOR3_2%C N_C_c_668_n N_C_M1019_g N_C_c_669_n N_C_c_670_n
+ N_C_c_671_n N_C_M1007_g N_C_c_673_n N_C_M1013_g N_C_M1020_g C N_C_c_674_n
+ N_C_c_675_n N_C_c_676_n PM_SKY130_FD_SC_MS__XNOR3_2%C
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_1057_74# N_A_1057_74#_M1023_d
+ N_A_1057_74#_M1005_d N_A_1057_74#_M1006_g N_A_1057_74#_c_754_n
+ N_A_1057_74#_M1009_g N_A_1057_74#_c_755_n N_A_1057_74#_M1008_g
+ N_A_1057_74#_c_757_n N_A_1057_74#_M1017_g N_A_1057_74#_c_786_n
+ N_A_1057_74#_c_758_n N_A_1057_74#_c_759_n N_A_1057_74#_c_768_n
+ N_A_1057_74#_c_760_n N_A_1057_74#_c_761_n N_A_1057_74#_c_762_n
+ N_A_1057_74#_c_857_p N_A_1057_74#_c_769_n N_A_1057_74#_c_797_n
+ N_A_1057_74#_c_799_n N_A_1057_74#_c_810_p N_A_1057_74#_c_801_n
+ N_A_1057_74#_c_770_n N_A_1057_74#_c_771_n N_A_1057_74#_c_763_n
+ N_A_1057_74#_c_764_n PM_SKY130_FD_SC_MS__XNOR3_2%A_1057_74#
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_27_373# N_A_27_373#_M1012_s N_A_27_373#_M1004_d
+ N_A_27_373#_M1015_s N_A_27_373#_M1011_d N_A_27_373#_c_879_n
+ N_A_27_373#_c_880_n N_A_27_373#_c_881_n N_A_27_373#_c_882_n
+ N_A_27_373#_c_890_n N_A_27_373#_c_891_n N_A_27_373#_c_935_n
+ N_A_27_373#_c_883_n N_A_27_373#_c_892_n N_A_27_373#_c_884_n
+ N_A_27_373#_c_885_n N_A_27_373#_c_886_n N_A_27_373#_c_887_n
+ N_A_27_373#_c_888_n PM_SKY130_FD_SC_MS__XNOR3_2%A_27_373#
x_PM_SKY130_FD_SC_MS__XNOR3_2%VPWR N_VPWR_M1015_d N_VPWR_M1021_d N_VPWR_M1020_d
+ N_VPWR_M1008_s N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n N_VPWR_c_986_n
+ N_VPWR_c_987_n VPWR N_VPWR_c_988_n N_VPWR_c_989_n N_VPWR_c_990_n
+ N_VPWR_c_991_n N_VPWR_c_992_n N_VPWR_c_993_n N_VPWR_c_982_n
+ PM_SKY130_FD_SC_MS__XNOR3_2%VPWR
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_335_373# N_A_335_373#_M1003_d
+ N_A_335_373#_M1019_d N_A_335_373#_M1000_d N_A_335_373#_M1005_s
+ N_A_335_373#_c_1077_n N_A_335_373#_c_1066_n N_A_335_373#_c_1067_n
+ N_A_335_373#_c_1068_n N_A_335_373#_c_1069_n N_A_335_373#_c_1070_n
+ N_A_335_373#_c_1071_n N_A_335_373#_c_1072_n N_A_335_373#_c_1081_n
+ N_A_335_373#_c_1073_n N_A_335_373#_c_1074_n N_A_335_373#_c_1075_n
+ N_A_335_373#_c_1076_n PM_SKY130_FD_SC_MS__XNOR3_2%A_335_373#
x_PM_SKY130_FD_SC_MS__XNOR3_2%A_329_81# N_A_329_81#_M1018_d N_A_329_81#_M1023_s
+ N_A_329_81#_M1014_d N_A_329_81#_M1007_d N_A_329_81#_c_1178_n
+ N_A_329_81#_c_1206_n N_A_329_81#_c_1184_n N_A_329_81#_c_1185_n
+ N_A_329_81#_c_1179_n N_A_329_81#_c_1180_n N_A_329_81#_c_1187_n
+ N_A_329_81#_c_1188_n N_A_329_81#_c_1181_n N_A_329_81#_c_1182_n
+ N_A_329_81#_c_1183_n N_A_329_81#_c_1241_n
+ PM_SKY130_FD_SC_MS__XNOR3_2%A_329_81#
x_PM_SKY130_FD_SC_MS__XNOR3_2%X N_X_M1009_d N_X_M1006_d N_X_c_1308_n
+ N_X_c_1309_n N_X_c_1306_n X X X PM_SKY130_FD_SC_MS__XNOR3_2%X
x_PM_SKY130_FD_SC_MS__XNOR3_2%VGND N_VGND_M1012_d N_VGND_M1016_d N_VGND_M1013_d
+ N_VGND_M1017_s N_VGND_c_1340_n N_VGND_c_1341_n N_VGND_c_1342_n N_VGND_c_1343_n
+ N_VGND_c_1344_n VGND N_VGND_c_1345_n N_VGND_c_1346_n N_VGND_c_1347_n
+ N_VGND_c_1348_n N_VGND_c_1349_n N_VGND_c_1350_n N_VGND_c_1351_n
+ PM_SKY130_FD_SC_MS__XNOR3_2%VGND
cc_1 VNB N_A_83_247#_M1015_g 0.00538716f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_2 VNB N_A_83_247#_M1012_g 0.0240792f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_3 VNB N_A_83_247#_c_176_n 0.00193372f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_4 VNB N_A_83_247#_c_177_n 6.25663e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_5 VNB N_A_83_247#_c_178_n 0.0350196f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_6 VNB N_A_83_247#_c_179_n 0.00535503f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.12
cc_7 VNB N_A_83_247#_c_180_n 0.00209465f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.34
cc_8 VNB N_A_83_247#_c_181_n 0.00538013f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.36
cc_9 VNB N_A_83_247#_c_182_n 0.0208851f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.35
cc_10 VNB N_A_M1010_g 0.0268525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_306_n 0.0232599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_307_n 0.00334759f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.565
cc_13 VNB N_A_397_21#_M1004_g 0.0385893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_397_21#_c_351_n 0.0171757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_397_21#_M1011_g 0.00877638f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.565
cc_16 VNB N_A_397_21#_c_353_n 0.0693021f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_17 VNB N_A_397_21#_c_354_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_397_21#_M1002_g 0.0373065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_397_21#_c_356_n 8.62302e-19 $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=0.55
cc_20 VNB N_A_397_21#_c_357_n 0.00521129f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.905
cc_21 VNB N_A_397_21#_c_358_n 0.00440373f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.115
cc_22 VNB N_A_397_21#_c_359_n 0.0335584f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_23 VNB N_A_397_21#_c_360_n 0.00404841f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.36
cc_24 VNB N_B_M1018_g 0.0344444f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.865
cc_25 VNB N_B_c_468_n 0.00570286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_M1000_g 0.00344654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_M1003_g 0.0212321f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.565
cc_28 VNB N_B_M1016_g 0.025787f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_29 VNB N_B_c_472_n 0.0133483f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=0.55
cc_30 VNB N_B_c_473_n 0.0030506f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.115
cc_31 VNB N_B_c_474_n 0.0515705f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_32 VNB N_A_1027_48#_M1023_g 0.0450805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1027_48#_c_590_n 0.00182968f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.365
cc_34 VNB N_A_1027_48#_c_591_n 0.0270322f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_35 VNB N_A_1027_48#_c_592_n 0.00260252f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_36 VNB N_A_1027_48#_c_593_n 0.00161761f $X=-0.19 $Y=-0.245 $X2=1.095
+ $Y2=2.035
cc_37 VNB N_A_1027_48#_c_594_n 9.42831e-19 $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.035
cc_38 VNB N_C_c_668_n 0.0175588f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.405
cc_39 VNB N_C_c_669_n 0.0115589f $X=-0.19 $Y=-0.245 $X2=3.295 $Y2=1.865
cc_40 VNB N_C_c_670_n 0.00905308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_c_671_n 0.0295931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_C_M1007_g 0.00372515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_C_c_673_n 0.0222798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_C_c_674_n 0.0409078f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_45 VNB N_C_c_675_n 0.035156f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.12
cc_46 VNB N_C_c_676_n 0.00330598f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.12
cc_47 VNB N_A_1057_74#_c_754_n 0.0170165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1057_74#_c_755_n 0.060644f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_49 VNB N_A_1057_74#_M1008_g 0.00429303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1057_74#_c_757_n 0.0188693f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_51 VNB N_A_1057_74#_c_758_n 0.0163721f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_52 VNB N_A_1057_74#_c_759_n 0.00383604f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.12
cc_53 VNB N_A_1057_74#_c_760_n 0.0104484f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.425
cc_54 VNB N_A_1057_74#_c_761_n 0.00552332f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.035
cc_55 VNB N_A_1057_74#_c_762_n 0.00315591f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.55
cc_56 VNB N_A_1057_74#_c_763_n 0.00443367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1057_74#_c_764_n 0.00228435f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.235
cc_58 VNB N_A_27_373#_c_879_n 0.0241546f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_59 VNB N_A_27_373#_c_880_n 6.56034e-19 $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_60 VNB N_A_27_373#_c_881_n 0.00263335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_373#_c_882_n 0.00475524f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_62 VNB N_A_27_373#_c_883_n 0.00770296f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=0.425
cc_63 VNB N_A_27_373#_c_884_n 0.00157907f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_64 VNB N_A_27_373#_c_885_n 0.0203735f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.12
cc_65 VNB N_A_27_373#_c_886_n 0.0033312f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.035
cc_66 VNB N_A_27_373#_c_887_n 0.029419f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.36
cc_67 VNB N_A_27_373#_c_888_n 0.00459486f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.795
cc_68 VNB N_VPWR_c_982_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_335_373#_c_1066_n 0.00562726f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=1.235
cc_70 VNB N_A_335_373#_c_1067_n 0.00249128f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.725
cc_71 VNB N_A_335_373#_c_1068_n 0.00300639f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.725
cc_72 VNB N_A_335_373#_c_1069_n 0.00255368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_335_373#_c_1070_n 0.0112843f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_74 VNB N_A_335_373#_c_1071_n 0.00652094f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_75 VNB N_A_335_373#_c_1072_n 0.00257282f $X=-0.19 $Y=-0.245 $X2=1.22
+ $Y2=1.035
cc_76 VNB N_A_335_373#_c_1073_n 0.0262647f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=2.99
cc_77 VNB N_A_335_373#_c_1074_n 0.00286242f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.12
cc_78 VNB N_A_335_373#_c_1075_n 0.00185916f $X=-0.19 $Y=-0.245 $X2=3.365
+ $Y2=0.35
cc_79 VNB N_A_335_373#_c_1076_n 0.00202343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_329_81#_c_1178_n 0.009648f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_81 VNB N_A_329_81#_c_1179_n 0.0164249f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.4
cc_82 VNB N_A_329_81#_c_1180_n 0.0153705f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_83 VNB N_A_329_81#_c_1181_n 0.00141657f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.035
cc_84 VNB N_A_329_81#_c_1182_n 0.00408737f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_85 VNB N_A_329_81#_c_1183_n 6.99046e-19 $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.34
cc_86 VNB N_X_c_1306_n 0.00115496f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_87 VNB X 0.00279061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1340_n 0.0080712f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_89 VNB N_VGND_c_1341_n 0.0123225f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.725
cc_90 VNB N_VGND_c_1342_n 0.0566416f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.36
cc_91 VNB N_VGND_c_1343_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.4
cc_92 VNB N_VGND_c_1344_n 0.0540788f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.4
cc_93 VNB N_VGND_c_1345_n 0.0184398f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.035
cc_94 VNB N_VGND_c_1346_n 0.0801099f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.12
cc_95 VNB N_VGND_c_1347_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=2.115
cc_96 VNB N_VGND_c_1348_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.795
cc_97 VNB N_VGND_c_1349_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1350_n 0.0297566f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.565
cc_99 VNB N_VGND_c_1351_n 0.466708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VPB N_A_83_247#_M1015_g 0.0277932f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_101 VPB N_A_83_247#_c_177_n 0.00167094f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_102 VPB N_A_83_247#_c_185_n 3.86242e-19 $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.905
cc_103 VPB N_A_83_247#_c_186_n 0.0342063f $X=-0.19 $Y=1.66 $X2=3.345 $Y2=2.99
cc_104 VPB N_A_83_247#_c_187_n 0.00278955f $X=-0.19 $Y=1.66 $X2=1.375 $Y2=2.99
cc_105 VPB N_A_83_247#_c_188_n 0.00876689f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=2.795
cc_106 VPB N_A_M1022_g 0.0219625f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.865
cc_107 VPB N_A_c_306_n 0.00732101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_c_307_n 0.0024708f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.565
cc_109 VPB N_A_397_21#_M1011_g 0.0224056f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.565
cc_110 VPB N_A_397_21#_M1001_g 0.0220534f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.4
cc_111 VPB N_A_397_21#_c_363_n 0.00272306f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=0.55
cc_112 VPB N_A_397_21#_c_364_n 0.00338753f $X=-0.19 $Y=1.66 $X2=1.375 $Y2=2.99
cc_113 VPB N_A_397_21#_c_358_n 0.00197208f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.115
cc_114 VPB N_A_397_21#_c_359_n 0.0122158f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_115 VPB N_B_M1000_g 0.0408459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_B_c_476_n 0.0603623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_B_c_477_n 0.014099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B_M1014_g 0.0543003f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.725
cc_119 VPB N_B_c_479_n 0.0786862f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.725
cc_120 VPB N_B_c_480_n 0.0783711f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_121 VPB N_B_M1021_g 0.0235492f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.035
cc_122 VPB N_B_c_482_n 0.00898883f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.12
cc_123 VPB N_B_c_473_n 0.00326101f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=2.115
cc_124 VPB N_B_c_474_n 0.00718655f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_125 VPB N_A_1027_48#_M1005_g 0.0270225f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.565
cc_126 VPB N_A_1027_48#_c_590_n 0.0093761f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_127 VPB N_A_1027_48#_c_591_n 0.023951f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.725
cc_128 VPB N_A_1027_48#_c_598_n 0.0116465f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_129 VPB N_A_1027_48#_c_594_n 0.00701589f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.035
cc_130 VPB N_A_1027_48#_c_600_n 0.00278791f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=0.55
cc_131 VPB N_C_M1007_g 0.0375189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_C_M1020_g 0.0248662f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.235
cc_133 VPB N_C_c_675_n 0.0104008f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.12
cc_134 VPB N_C_c_676_n 0.00456929f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.12
cc_135 VPB N_A_1057_74#_M1006_g 0.0239262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_1057_74#_c_755_n 0.00590784f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_137 VPB N_A_1057_74#_M1008_g 0.0274138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_1057_74#_c_768_n 0.0338257f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.12
cc_139 VPB N_A_1057_74#_c_769_n 0.0136763f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.34
cc_140 VPB N_A_1057_74#_c_770_n 0.00274009f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.36
cc_141 VPB N_A_1057_74#_c_771_n 0.00978494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_1057_74#_c_763_n 8.15627e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_27_373#_c_881_n 0.00137242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_27_373#_c_890_n 0.00701431f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.4
cc_145 VPB N_A_27_373#_c_891_n 3.23193e-19 $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_146 VPB N_A_27_373#_c_892_n 0.0268183f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=0.55
cc_147 VPB N_A_27_373#_c_887_n 0.0262562f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.36
cc_148 VPB N_VPWR_c_983_n 0.0138235f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.235
cc_149 VPB N_VPWR_c_984_n 0.0160348f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.36
cc_150 VPB N_VPWR_c_985_n 0.00830203f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_151 VPB N_VPWR_c_986_n 0.0104926f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.12
cc_152 VPB N_VPWR_c_987_n 0.0587358f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.035
cc_153 VPB N_VPWR_c_988_n 0.0877154f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.905
cc_154 VPB N_VPWR_c_989_n 0.0667808f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_155 VPB N_VPWR_c_990_n 0.0204869f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=2.795
cc_156 VPB N_VPWR_c_991_n 0.0257077f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.565
cc_157 VPB N_VPWR_c_992_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_993_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_982_n 0.101481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_335_373#_c_1077_n 0.00242978f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.365
cc_161 VPB N_A_335_373#_c_1066_n 0.00320013f $X=-0.19 $Y=1.66 $X2=0.535
+ $Y2=1.235
cc_162 VPB N_A_335_373#_c_1067_n 4.66474e-19 $X=-0.19 $Y=1.66 $X2=0.535
+ $Y2=0.725
cc_163 VPB N_A_335_373#_c_1069_n 0.00495167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_335_373#_c_1081_n 0.00567696f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=0.34
cc_165 VPB N_A_329_81#_c_1184_n 0.00366045f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.36
cc_166 VPB N_A_329_81#_c_1185_n 7.42911e-19 $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_167 VPB N_A_329_81#_c_1180_n 0.00366055f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_168 VPB N_A_329_81#_c_1187_n 0.0124642f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.4
cc_169 VPB N_A_329_81#_c_1188_n 0.00176765f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.035
cc_170 VPB N_X_c_1308_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_X_c_1309_n 8.15497e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_172 VPB N_X_c_1306_n 9.676e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_173 N_A_83_247#_c_189_p N_A_M1022_g 0.012575f $X=1.095 $Y=2.035 $X2=0 $Y2=0
cc_174 N_A_83_247#_c_190_p N_A_M1022_g 0.00118624f $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_175 N_A_83_247#_c_185_n N_A_M1022_g 0.0138739f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_176 N_A_83_247#_c_187_n N_A_M1022_g 0.00300855f $X=1.375 $Y=2.99 $X2=0 $Y2=0
cc_177 N_A_83_247#_M1012_g N_A_M1010_g 0.0220707f $X=0.535 $Y=0.725 $X2=0 $Y2=0
cc_178 N_A_83_247#_c_176_n N_A_M1010_g 0.00186641f $X=0.62 $Y=1.36 $X2=0 $Y2=0
cc_179 N_A_83_247#_c_178_n N_A_M1010_g 0.00862331f $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_180 N_A_83_247#_c_179_n N_A_M1010_g 0.0139401f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_181 N_A_83_247#_c_197_p N_A_M1010_g 0.00778962f $X=1.26 $Y=0.55 $X2=0 $Y2=0
cc_182 N_A_83_247#_c_180_n N_A_M1010_g 0.00383348f $X=1.345 $Y=0.34 $X2=0 $Y2=0
cc_183 N_A_83_247#_M1015_g N_A_c_306_n 0.0350998f $X=0.505 $Y=2.365 $X2=0 $Y2=0
cc_184 N_A_83_247#_c_177_n N_A_c_306_n 0.00593762f $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_185 N_A_83_247#_c_178_n N_A_c_306_n 0.0115787f $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_186 N_A_83_247#_c_179_n N_A_c_306_n 0.00140189f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_187 N_A_83_247#_c_190_p N_A_c_306_n 8.28178e-19 $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_188 N_A_83_247#_M1015_g N_A_c_307_n 2.20531e-19 $X=0.505 $Y=2.365 $X2=0 $Y2=0
cc_189 N_A_83_247#_c_177_n N_A_c_307_n 0.0260342f $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_190 N_A_83_247#_c_178_n N_A_c_307_n 6.61488e-19 $X=0.58 $Y=1.4 $X2=0 $Y2=0
cc_191 N_A_83_247#_c_179_n N_A_c_307_n 0.0225458f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_192 N_A_83_247#_c_189_p N_A_c_307_n 0.00987176f $X=1.095 $Y=2.035 $X2=0 $Y2=0
cc_193 N_A_83_247#_c_190_p N_A_c_307_n 0.0161144f $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_194 N_A_83_247#_c_182_n N_A_397_21#_M1004_g 0.012253f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_195 N_A_83_247#_c_186_n N_A_397_21#_M1011_g 5.03968e-19 $X=3.345 $Y=2.99
+ $X2=0 $Y2=0
cc_196 N_A_83_247#_c_182_n N_A_397_21#_c_353_n 0.0135339f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_197 N_A_83_247#_c_181_n N_A_397_21#_M1002_g 8.00488e-19 $X=3.365 $Y=0.36
+ $X2=0 $Y2=0
cc_198 N_A_83_247#_c_182_n N_A_397_21#_M1002_g 0.0134669f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_199 N_A_83_247#_c_186_n N_A_397_21#_M1001_g 0.0018681f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_200 N_A_83_247#_c_188_n N_A_397_21#_M1001_g 0.00367682f $X=3.51 $Y=2.795
+ $X2=0 $Y2=0
cc_201 N_A_83_247#_M1001_d N_A_397_21#_c_363_n 0.00231439f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_202 N_A_83_247#_M1002_d N_A_397_21#_c_356_n 0.00454958f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_203 N_A_83_247#_M1001_d N_A_397_21#_c_376_n 0.00639042f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_204 N_A_83_247#_M1001_d N_A_397_21#_c_364_n 0.00266017f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_205 N_A_83_247#_M1002_d N_A_397_21#_c_360_n 0.00205319f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_206 N_A_83_247#_c_179_n N_B_M1018_g 0.00412463f $X=1.095 $Y=1.12 $X2=0 $Y2=0
cc_207 N_A_83_247#_c_197_p N_B_M1018_g 0.00833237f $X=1.26 $Y=0.55 $X2=0 $Y2=0
cc_208 N_A_83_247#_c_182_n N_B_M1018_g 0.0145029f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_209 N_A_83_247#_c_190_p N_B_M1000_g 0.00138862f $X=1.235 $Y=2.12 $X2=0 $Y2=0
cc_210 N_A_83_247#_c_185_n N_B_M1000_g 0.00889795f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_211 N_A_83_247#_c_186_n N_B_M1000_g 0.0154033f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_212 N_A_83_247#_c_186_n N_B_c_476_n 0.0144886f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_213 N_A_83_247#_c_182_n N_B_M1003_g 0.00116683f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_214 N_A_83_247#_c_186_n N_B_M1014_g 0.0194072f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_215 N_A_83_247#_c_188_n N_B_M1014_g 0.00232951f $X=3.51 $Y=2.795 $X2=0 $Y2=0
cc_216 N_A_83_247#_c_186_n N_B_c_479_n 0.00881996f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_217 N_A_83_247#_c_188_n N_B_c_479_n 0.00889438f $X=3.51 $Y=2.795 $X2=0 $Y2=0
cc_218 N_A_83_247#_c_188_n N_B_c_480_n 0.0137734f $X=3.51 $Y=2.795 $X2=0 $Y2=0
cc_219 N_A_83_247#_c_181_n N_B_M1016_g 0.00356999f $X=3.365 $Y=0.36 $X2=0 $Y2=0
cc_220 N_A_83_247#_M1012_g N_A_27_373#_c_879_n 8.91276e-19 $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_221 N_A_83_247#_c_179_n N_A_27_373#_c_880_n 0.00266509f $X=1.095 $Y=1.12
+ $X2=0 $Y2=0
cc_222 N_A_83_247#_c_190_p N_A_27_373#_c_881_n 0.0134182f $X=1.235 $Y=2.12 $X2=0
+ $Y2=0
cc_223 N_A_83_247#_c_185_n N_A_27_373#_c_881_n 0.0324214f $X=1.235 $Y=2.905
+ $X2=0 $Y2=0
cc_224 N_A_83_247#_c_186_n N_A_27_373#_c_890_n 0.0654508f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_225 N_A_83_247#_c_185_n N_A_27_373#_c_891_n 0.0138427f $X=1.235 $Y=2.905
+ $X2=0 $Y2=0
cc_226 N_A_83_247#_c_186_n N_A_27_373#_c_891_n 0.0123447f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_227 N_A_83_247#_c_176_n N_A_27_373#_c_883_n 0.00205386f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_228 N_A_83_247#_M1015_g N_A_27_373#_c_892_n 0.00946157f $X=0.505 $Y=2.365
+ $X2=0 $Y2=0
cc_229 N_A_83_247#_c_185_n N_A_27_373#_c_892_n 3.65835e-19 $X=1.235 $Y=2.905
+ $X2=0 $Y2=0
cc_230 N_A_83_247#_M1012_g N_A_27_373#_c_885_n 0.00484232f $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_231 N_A_83_247#_c_176_n N_A_27_373#_c_885_n 0.0125183f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_232 N_A_83_247#_c_177_n N_A_27_373#_c_885_n 0.0133627f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_233 N_A_83_247#_c_178_n N_A_27_373#_c_885_n 0.00601258f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_234 N_A_83_247#_c_179_n N_A_27_373#_c_885_n 0.0234041f $X=1.095 $Y=1.12 $X2=0
+ $Y2=0
cc_235 N_A_83_247#_c_189_p N_A_27_373#_c_885_n 0.00660061f $X=1.095 $Y=2.035
+ $X2=0 $Y2=0
cc_236 N_A_83_247#_c_190_p N_A_27_373#_c_885_n 0.00256289f $X=1.235 $Y=2.12
+ $X2=0 $Y2=0
cc_237 N_A_83_247#_M1012_g N_A_27_373#_c_886_n 0.00113427f $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_238 N_A_83_247#_c_176_n N_A_27_373#_c_886_n 0.00131456f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_239 N_A_83_247#_c_177_n N_A_27_373#_c_886_n 0.00136538f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_240 N_A_83_247#_c_178_n N_A_27_373#_c_886_n 0.00130928f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_241 N_A_83_247#_M1012_g N_A_27_373#_c_887_n 0.00350179f $X=0.535 $Y=0.725
+ $X2=0 $Y2=0
cc_242 N_A_83_247#_c_176_n N_A_27_373#_c_887_n 0.0180374f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_243 N_A_83_247#_c_177_n N_A_27_373#_c_887_n 0.0438297f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_244 N_A_83_247#_c_178_n N_A_27_373#_c_887_n 0.0242641f $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_245 N_A_83_247#_c_261_p N_A_27_373#_c_887_n 0.0136904f $X=0.745 $Y=2.035
+ $X2=0 $Y2=0
cc_246 N_A_83_247#_c_179_n N_A_27_373#_c_888_n 6.39812e-19 $X=1.095 $Y=1.12
+ $X2=0 $Y2=0
cc_247 N_A_83_247#_c_177_n N_VPWR_M1015_d 0.0010503f $X=0.58 $Y=1.4 $X2=-0.19
+ $Y2=-0.245
cc_248 N_A_83_247#_c_189_p N_VPWR_M1015_d 0.00470439f $X=1.095 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_249 N_A_83_247#_c_261_p N_VPWR_M1015_d 0.00105545f $X=0.745 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_250 N_A_83_247#_M1015_g N_VPWR_c_983_n 0.00416111f $X=0.505 $Y=2.365 $X2=0
+ $Y2=0
cc_251 N_A_83_247#_c_189_p N_VPWR_c_983_n 0.0116514f $X=1.095 $Y=2.035 $X2=0
+ $Y2=0
cc_252 N_A_83_247#_c_261_p N_VPWR_c_983_n 0.00782629f $X=0.745 $Y=2.035 $X2=0
+ $Y2=0
cc_253 N_A_83_247#_c_185_n N_VPWR_c_983_n 0.0235f $X=1.235 $Y=2.905 $X2=0 $Y2=0
cc_254 N_A_83_247#_c_187_n N_VPWR_c_983_n 0.0144537f $X=1.375 $Y=2.99 $X2=0
+ $Y2=0
cc_255 N_A_83_247#_c_186_n N_VPWR_c_988_n 0.1258f $X=3.345 $Y=2.99 $X2=0 $Y2=0
cc_256 N_A_83_247#_c_187_n N_VPWR_c_988_n 0.0200723f $X=1.375 $Y=2.99 $X2=0
+ $Y2=0
cc_257 N_A_83_247#_c_188_n N_VPWR_c_988_n 0.0213919f $X=3.51 $Y=2.795 $X2=0
+ $Y2=0
cc_258 N_A_83_247#_M1015_g N_VPWR_c_991_n 0.00586114f $X=0.505 $Y=2.365 $X2=0
+ $Y2=0
cc_259 N_A_83_247#_M1015_g N_VPWR_c_982_n 0.00619157f $X=0.505 $Y=2.365 $X2=0
+ $Y2=0
cc_260 N_A_83_247#_c_186_n N_VPWR_c_982_n 0.0663994f $X=3.345 $Y=2.99 $X2=0
+ $Y2=0
cc_261 N_A_83_247#_c_187_n N_VPWR_c_982_n 0.0108858f $X=1.375 $Y=2.99 $X2=0
+ $Y2=0
cc_262 N_A_83_247#_c_188_n N_VPWR_c_982_n 0.0110564f $X=3.51 $Y=2.795 $X2=0
+ $Y2=0
cc_263 N_A_83_247#_M1002_d N_A_335_373#_c_1073_n 0.00275472f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_264 N_A_83_247#_c_182_n N_A_329_81#_M1018_d 0.00221108f $X=3.2 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_265 N_A_83_247#_M1002_d N_A_329_81#_c_1178_n 0.00880418f $X=3.145 $Y=0.625
+ $X2=0 $Y2=0
cc_266 N_A_83_247#_c_181_n N_A_329_81#_c_1178_n 0.022946f $X=3.365 $Y=0.36 $X2=0
+ $Y2=0
cc_267 N_A_83_247#_c_182_n N_A_329_81#_c_1178_n 0.0296435f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_268 N_A_83_247#_M1001_d N_A_329_81#_c_1184_n 0.00687526f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_269 N_A_83_247#_c_186_n N_A_329_81#_c_1184_n 0.00642816f $X=3.345 $Y=2.99
+ $X2=0 $Y2=0
cc_270 N_A_83_247#_c_188_n N_A_329_81#_c_1184_n 0.0245806f $X=3.51 $Y=2.795
+ $X2=0 $Y2=0
cc_271 N_A_83_247#_c_186_n N_A_329_81#_c_1185_n 0.0136531f $X=3.345 $Y=2.99
+ $X2=0 $Y2=0
cc_272 N_A_83_247#_c_197_p N_A_329_81#_c_1181_n 0.0207307f $X=1.26 $Y=0.55 $X2=0
+ $Y2=0
cc_273 N_A_83_247#_c_182_n N_A_329_81#_c_1181_n 0.0198438f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_274 N_A_83_247#_c_182_n N_A_329_81#_c_1182_n 0.0530595f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_275 N_A_83_247#_c_176_n N_VGND_M1012_d 8.63167e-19 $X=0.62 $Y=1.36 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_83_247#_c_179_n N_VGND_M1012_d 0.00177524f $X=1.095 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_83_247#_M1012_g N_VGND_c_1340_n 0.0146489f $X=0.535 $Y=0.725 $X2=0
+ $Y2=0
cc_278 N_A_83_247#_c_176_n N_VGND_c_1340_n 0.00852004f $X=0.62 $Y=1.36 $X2=0
+ $Y2=0
cc_279 N_A_83_247#_c_178_n N_VGND_c_1340_n 5.55578e-19 $X=0.58 $Y=1.4 $X2=0
+ $Y2=0
cc_280 N_A_83_247#_c_179_n N_VGND_c_1340_n 0.0127781f $X=1.095 $Y=1.12 $X2=0
+ $Y2=0
cc_281 N_A_83_247#_c_180_n N_VGND_c_1340_n 0.0129079f $X=1.345 $Y=0.34 $X2=0
+ $Y2=0
cc_282 N_A_83_247#_M1012_g N_VGND_c_1345_n 0.0045897f $X=0.535 $Y=0.725 $X2=0
+ $Y2=0
cc_283 N_A_83_247#_c_180_n N_VGND_c_1346_n 0.0179217f $X=1.345 $Y=0.34 $X2=0
+ $Y2=0
cc_284 N_A_83_247#_c_182_n N_VGND_c_1346_n 0.139665f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_285 N_A_83_247#_M1002_d N_VGND_c_1351_n 0.00251887f $X=3.145 $Y=0.625 $X2=0
+ $Y2=0
cc_286 N_A_83_247#_M1012_g N_VGND_c_1351_n 0.0044912f $X=0.535 $Y=0.725 $X2=0
+ $Y2=0
cc_287 N_A_83_247#_c_180_n N_VGND_c_1351_n 0.00971942f $X=1.345 $Y=0.34 $X2=0
+ $Y2=0
cc_288 N_A_83_247#_c_182_n N_VGND_c_1351_n 0.0773214f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_289 N_A_M1010_g N_B_M1018_g 0.0218506f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_290 N_A_c_306_n N_B_M1018_g 0.0196375f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_291 N_A_c_307_n N_B_M1018_g 0.00253285f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_292 N_A_M1022_g N_B_M1000_g 0.0268594f $X=1.045 $Y=2.365 $X2=0 $Y2=0
cc_293 N_A_M1010_g N_A_27_373#_c_880_n 0.00146258f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_294 N_A_c_307_n N_A_27_373#_c_880_n 2.43113e-19 $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_295 N_A_M1022_g N_A_27_373#_c_881_n 0.00122091f $X=1.045 $Y=2.365 $X2=0 $Y2=0
cc_296 N_A_c_306_n N_A_27_373#_c_881_n 3.77853e-19 $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_297 N_A_c_307_n N_A_27_373#_c_881_n 0.0238428f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_298 N_A_M1010_g N_A_27_373#_c_885_n 0.00523989f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_299 N_A_c_307_n N_A_27_373#_c_885_n 0.0103716f $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_300 N_A_c_307_n N_A_27_373#_c_888_n 8.6259e-19 $X=1.12 $Y=1.54 $X2=0 $Y2=0
cc_301 N_A_M1022_g N_VPWR_c_983_n 0.00438321f $X=1.045 $Y=2.365 $X2=0 $Y2=0
cc_302 N_A_M1022_g N_VPWR_c_988_n 0.00497021f $X=1.045 $Y=2.365 $X2=0 $Y2=0
cc_303 N_A_M1022_g N_VPWR_c_982_n 0.00481567f $X=1.045 $Y=2.365 $X2=0 $Y2=0
cc_304 N_A_M1010_g N_VGND_c_1340_n 0.00352423f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_305 N_A_M1010_g N_VGND_c_1346_n 0.0047553f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_306 N_A_M1010_g N_VGND_c_1351_n 0.00445555f $X=1.045 $Y=0.725 $X2=0 $Y2=0
cc_307 N_A_397_21#_M1004_g N_B_M1018_g 0.0348758f $X=2.06 $Y=1.055 $X2=0 $Y2=0
cc_308 N_A_397_21#_M1011_g N_B_M1018_g 2.98053e-19 $X=2.195 $Y=2.185 $X2=0 $Y2=0
cc_309 N_A_397_21#_M1011_g N_B_c_468_n 0.022065f $X=2.195 $Y=2.185 $X2=0 $Y2=0
cc_310 N_A_397_21#_M1011_g N_B_c_476_n 0.00376062f $X=2.195 $Y=2.185 $X2=0 $Y2=0
cc_311 N_A_397_21#_M1004_g N_B_M1003_g 0.022321f $X=2.06 $Y=1.055 $X2=0 $Y2=0
cc_312 N_A_397_21#_c_351_n N_B_M1003_g 0.0101362f $X=2.195 $Y=1.49 $X2=0 $Y2=0
cc_313 N_A_397_21#_c_353_n N_B_M1003_g 0.00737859f $X=2.995 $Y=0.18 $X2=0 $Y2=0
cc_314 N_A_397_21#_M1002_g N_B_M1003_g 0.0245034f $X=3.07 $Y=0.945 $X2=0 $Y2=0
cc_315 N_A_397_21#_M1011_g N_B_M1014_g 0.0150308f $X=2.195 $Y=2.185 $X2=0 $Y2=0
cc_316 N_A_397_21#_M1001_g N_B_M1014_g 0.0230488f $X=3.205 $Y=2.285 $X2=0 $Y2=0
cc_317 N_A_397_21#_M1001_g N_B_c_479_n 0.00885431f $X=3.205 $Y=2.285 $X2=0 $Y2=0
cc_318 N_A_397_21#_M1001_g N_B_c_480_n 0.0273672f $X=3.205 $Y=2.285 $X2=0 $Y2=0
cc_319 N_A_397_21#_c_364_n N_B_c_480_n 0.0147642f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_320 N_A_397_21#_c_358_n N_B_c_480_n 0.00340873f $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_321 N_A_397_21#_c_357_n N_B_M1016_g 0.00383817f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_322 N_A_397_21#_c_360_n N_B_M1016_g 0.00357912f $X=3.36 $Y=1.375 $X2=0 $Y2=0
cc_323 N_A_397_21#_c_364_n N_B_M1021_g 0.0047394f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_324 N_A_397_21#_M1011_g N_B_c_472_n 0.0101362f $X=2.195 $Y=2.185 $X2=0 $Y2=0
cc_325 N_A_397_21#_c_358_n N_B_c_472_n 2.81261e-19 $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_326 N_A_397_21#_c_359_n N_B_c_472_n 0.0109156f $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_327 N_A_397_21#_c_357_n N_B_c_473_n 0.0145936f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_328 N_A_397_21#_c_364_n N_B_c_473_n 0.0384932f $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_329 N_A_397_21#_c_359_n N_B_c_473_n 3.47661e-19 $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_330 N_A_397_21#_c_360_n N_B_c_473_n 0.0356463f $X=3.36 $Y=1.375 $X2=0 $Y2=0
cc_331 N_A_397_21#_M1002_g N_B_c_474_n 4.40661e-19 $X=3.07 $Y=0.945 $X2=0 $Y2=0
cc_332 N_A_397_21#_c_357_n N_B_c_474_n 0.00236562f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_333 N_A_397_21#_c_364_n N_B_c_474_n 9.48761e-19 $X=4.09 $Y=2.115 $X2=0 $Y2=0
cc_334 N_A_397_21#_c_359_n N_B_c_474_n 0.0181869f $X=3.32 $Y=1.54 $X2=0 $Y2=0
cc_335 N_A_397_21#_c_360_n N_B_c_474_n 0.00340873f $X=3.36 $Y=1.375 $X2=0 $Y2=0
cc_336 N_A_397_21#_c_351_n N_A_27_373#_c_881_n 0.00200088f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_337 N_A_397_21#_M1011_g N_A_27_373#_c_881_n 0.00216918f $X=2.195 $Y=2.185
+ $X2=0 $Y2=0
cc_338 N_A_397_21#_M1004_g N_A_27_373#_c_882_n 0.00808752f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_339 N_A_397_21#_c_351_n N_A_27_373#_c_882_n 0.00253261f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_340 N_A_397_21#_M1011_g N_A_27_373#_c_890_n 0.0122509f $X=2.195 $Y=2.185
+ $X2=0 $Y2=0
cc_341 N_A_397_21#_M1001_g N_A_27_373#_c_890_n 4.69481e-19 $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_342 N_A_397_21#_M1011_g N_A_27_373#_c_935_n 0.00898312f $X=2.195 $Y=2.185
+ $X2=0 $Y2=0
cc_343 N_A_397_21#_M1004_g N_A_27_373#_c_884_n 0.00115834f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_344 N_A_397_21#_c_351_n N_A_27_373#_c_884_n 0.00618395f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_345 N_A_397_21#_c_351_n N_A_27_373#_c_888_n 5.07152e-19 $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_346 N_A_397_21#_M1011_g N_A_335_373#_c_1077_n 0.00518624f $X=2.195 $Y=2.185
+ $X2=0 $Y2=0
cc_347 N_A_397_21#_M1011_g N_A_335_373#_c_1066_n 0.0146093f $X=2.195 $Y=2.185
+ $X2=0 $Y2=0
cc_348 N_A_397_21#_c_363_n N_A_335_373#_c_1066_n 4.14392e-19 $X=3.48 $Y=1.95
+ $X2=0 $Y2=0
cc_349 N_A_397_21#_c_358_n N_A_335_373#_c_1066_n 0.00626949f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_350 N_A_397_21#_c_359_n N_A_335_373#_c_1066_n 6.6902e-19 $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_351 N_A_397_21#_c_351_n N_A_335_373#_c_1067_n 0.00373139f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_352 N_A_397_21#_M1011_g N_A_335_373#_c_1067_n 0.00201423f $X=2.195 $Y=2.185
+ $X2=0 $Y2=0
cc_353 N_A_397_21#_M1002_g N_A_335_373#_c_1072_n 3.44089e-19 $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_354 N_A_397_21#_c_360_n N_A_335_373#_c_1072_n 0.00301081f $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_355 N_A_397_21#_M1002_g N_A_335_373#_c_1073_n 0.00697065f $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_356 N_A_397_21#_c_357_n N_A_335_373#_c_1073_n 0.018201f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_357 N_A_397_21#_c_364_n N_A_335_373#_c_1073_n 0.00714503f $X=4.09 $Y=2.115
+ $X2=0 $Y2=0
cc_358 N_A_397_21#_c_358_n N_A_335_373#_c_1073_n 0.00904642f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_359 N_A_397_21#_c_359_n N_A_335_373#_c_1073_n 3.48429e-19 $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_360 N_A_397_21#_c_360_n N_A_335_373#_c_1073_n 0.0193866f $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_361 N_A_397_21#_M1002_g N_A_335_373#_c_1074_n 7.21505e-19 $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_362 N_A_397_21#_c_358_n N_A_335_373#_c_1074_n 8.91892e-19 $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_363 N_A_397_21#_c_360_n N_A_335_373#_c_1074_n 4.32441e-19 $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_364 N_A_397_21#_c_351_n N_A_335_373#_c_1075_n 0.00119995f $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_365 N_A_397_21#_M1002_g N_A_335_373#_c_1075_n 0.00178826f $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_366 N_A_397_21#_c_358_n N_A_335_373#_c_1075_n 0.00645185f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_367 N_A_397_21#_c_360_n N_A_335_373#_c_1075_n 0.00139636f $X=3.36 $Y=1.375
+ $X2=0 $Y2=0
cc_368 N_A_397_21#_M1016_s N_A_329_81#_c_1178_n 0.00698754f $X=3.78 $Y=0.445
+ $X2=0 $Y2=0
cc_369 N_A_397_21#_M1002_g N_A_329_81#_c_1178_n 0.0140287f $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_370 N_A_397_21#_c_356_n N_A_329_81#_c_1178_n 0.01346f $X=3.565 $Y=1.04 $X2=0
+ $Y2=0
cc_371 N_A_397_21#_c_357_n N_A_329_81#_c_1178_n 0.0328652f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_372 N_A_397_21#_c_358_n N_A_329_81#_c_1178_n 0.00253746f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_373 N_A_397_21#_c_359_n N_A_329_81#_c_1178_n 0.00133832f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_374 N_A_397_21#_M1001_g N_A_329_81#_c_1206_n 0.00895034f $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_375 N_A_397_21#_c_363_n N_A_329_81#_c_1206_n 0.00407016f $X=3.48 $Y=1.95
+ $X2=0 $Y2=0
cc_376 N_A_397_21#_c_376_n N_A_329_81#_c_1206_n 0.0152789f $X=3.565 $Y=2.075
+ $X2=0 $Y2=0
cc_377 N_A_397_21#_c_359_n N_A_329_81#_c_1206_n 0.00442727f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_378 N_A_397_21#_M1021_s N_A_329_81#_c_1184_n 0.00639623f $X=3.95 $Y=1.84
+ $X2=0 $Y2=0
cc_379 N_A_397_21#_M1001_g N_A_329_81#_c_1184_n 0.0118459f $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_380 N_A_397_21#_c_376_n N_A_329_81#_c_1184_n 0.0137412f $X=3.565 $Y=2.075
+ $X2=0 $Y2=0
cc_381 N_A_397_21#_c_364_n N_A_329_81#_c_1184_n 0.0467965f $X=4.09 $Y=2.115
+ $X2=0 $Y2=0
cc_382 N_A_397_21#_c_358_n N_A_329_81#_c_1184_n 0.00494645f $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_383 N_A_397_21#_c_359_n N_A_329_81#_c_1184_n 5.45112e-19 $X=3.32 $Y=1.54
+ $X2=0 $Y2=0
cc_384 N_A_397_21#_M1001_g N_A_329_81#_c_1185_n 9.04191e-19 $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_385 N_A_397_21#_c_357_n N_A_329_81#_c_1179_n 3.53781e-19 $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_386 N_A_397_21#_c_357_n N_A_329_81#_c_1180_n 0.00564206f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_387 N_A_397_21#_c_364_n N_A_329_81#_c_1180_n 0.0116679f $X=4.09 $Y=2.115
+ $X2=0 $Y2=0
cc_388 N_A_397_21#_M1004_g N_A_329_81#_c_1181_n 0.0033689f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_389 N_A_397_21#_M1004_g N_A_329_81#_c_1182_n 0.0109418f $X=2.06 $Y=1.055
+ $X2=0 $Y2=0
cc_390 N_A_397_21#_c_351_n N_A_329_81#_c_1182_n 4.49044e-19 $X=2.195 $Y=1.49
+ $X2=0 $Y2=0
cc_391 N_A_397_21#_M1002_g N_A_329_81#_c_1183_n 4.77048e-19 $X=3.07 $Y=0.945
+ $X2=0 $Y2=0
cc_392 N_A_397_21#_c_354_n N_VGND_c_1346_n 0.0250991f $X=2.135 $Y=0.18 $X2=0
+ $Y2=0
cc_393 N_A_397_21#_c_353_n N_VGND_c_1351_n 0.0262914f $X=2.995 $Y=0.18 $X2=0
+ $Y2=0
cc_394 N_A_397_21#_c_354_n N_VGND_c_1351_n 0.00604517f $X=2.135 $Y=0.18 $X2=0
+ $Y2=0
cc_395 N_B_M1018_g N_A_27_373#_c_880_n 0.0126155f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_396 N_B_M1018_g N_A_27_373#_c_881_n 0.00273704f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_397 N_B_c_468_n N_A_27_373#_c_881_n 0.00300456f $X=1.585 $Y=1.595 $X2=0 $Y2=0
cc_398 N_B_M1000_g N_A_27_373#_c_881_n 0.0262378f $X=1.585 $Y=2.285 $X2=0 $Y2=0
cc_399 N_B_M1014_g N_A_27_373#_c_890_n 0.00695077f $X=2.665 $Y=2.185 $X2=0 $Y2=0
cc_400 N_B_M1000_g N_A_27_373#_c_891_n 0.00847779f $X=1.585 $Y=2.285 $X2=0 $Y2=0
cc_401 N_B_M1000_g N_A_27_373#_c_935_n 2.48102e-19 $X=1.585 $Y=2.285 $X2=0 $Y2=0
cc_402 N_B_M1014_g N_A_27_373#_c_935_n 0.0096966f $X=2.665 $Y=2.185 $X2=0 $Y2=0
cc_403 N_B_c_472_n N_A_27_373#_c_935_n 3.94564e-19 $X=2.625 $Y=1.655 $X2=0 $Y2=0
cc_404 N_B_M1003_g N_A_27_373#_c_884_n 0.00345094f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_405 N_B_M1018_g N_A_27_373#_c_885_n 0.0043171f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_406 N_B_M1018_g N_A_27_373#_c_888_n 0.00193489f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_407 N_B_M1000_g N_VPWR_c_983_n 2.89414e-19 $X=1.585 $Y=2.285 $X2=0 $Y2=0
cc_408 N_B_c_477_n N_VPWR_c_983_n 0.00242213f $X=1.675 $Y=3.15 $X2=0 $Y2=0
cc_409 N_B_c_480_n N_VPWR_c_984_n 0.00274317f $X=3.8 $Y=3.075 $X2=0 $Y2=0
cc_410 N_B_M1021_g N_VPWR_c_984_n 0.0100591f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_411 N_B_c_477_n N_VPWR_c_988_n 0.0541298f $X=1.675 $Y=3.15 $X2=0 $Y2=0
cc_412 N_B_M1021_g N_VPWR_c_988_n 0.00553757f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_413 N_B_c_476_n N_VPWR_c_982_n 0.0211783f $X=2.575 $Y=3.15 $X2=0 $Y2=0
cc_414 N_B_c_477_n N_VPWR_c_982_n 0.00678686f $X=1.675 $Y=3.15 $X2=0 $Y2=0
cc_415 N_B_c_479_n N_VPWR_c_982_n 0.0301161f $X=3.725 $Y=3.15 $X2=0 $Y2=0
cc_416 N_B_M1021_g N_VPWR_c_982_n 0.00545887f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_417 N_B_c_482_n N_VPWR_c_982_n 0.00445015f $X=2.665 $Y=3.15 $X2=0 $Y2=0
cc_418 N_B_M1000_g N_A_335_373#_c_1077_n 0.00226644f $X=1.585 $Y=2.285 $X2=0
+ $Y2=0
cc_419 N_B_M1014_g N_A_335_373#_c_1066_n 0.00990605f $X=2.665 $Y=2.185 $X2=0
+ $Y2=0
cc_420 N_B_c_472_n N_A_335_373#_c_1066_n 0.00602964f $X=2.625 $Y=1.655 $X2=0
+ $Y2=0
cc_421 N_B_c_468_n N_A_335_373#_c_1067_n 6.83818e-19 $X=1.585 $Y=1.595 $X2=0
+ $Y2=0
cc_422 N_B_M1003_g N_A_335_373#_c_1072_n 0.00588367f $X=2.57 $Y=0.945 $X2=0
+ $Y2=0
cc_423 N_B_c_472_n N_A_335_373#_c_1072_n 4.46333e-19 $X=2.625 $Y=1.655 $X2=0
+ $Y2=0
cc_424 N_B_M1016_g N_A_335_373#_c_1073_n 0.00592452f $X=4.14 $Y=0.815 $X2=0
+ $Y2=0
cc_425 N_B_c_473_n N_A_335_373#_c_1073_n 0.0255335f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_426 N_B_c_474_n N_A_335_373#_c_1073_n 0.00595754f $X=4.315 $Y=1.515 $X2=0
+ $Y2=0
cc_427 N_B_M1003_g N_A_335_373#_c_1074_n 0.00173286f $X=2.57 $Y=0.945 $X2=0
+ $Y2=0
cc_428 N_B_M1003_g N_A_335_373#_c_1075_n 0.005578f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_429 N_B_c_472_n N_A_335_373#_c_1075_n 0.00384975f $X=2.625 $Y=1.655 $X2=0
+ $Y2=0
cc_430 N_B_M1016_g N_A_329_81#_c_1178_n 0.0169621f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_431 N_B_c_473_n N_A_329_81#_c_1178_n 0.00378334f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_432 N_B_c_474_n N_A_329_81#_c_1178_n 7.94901e-19 $X=4.315 $Y=1.515 $X2=0
+ $Y2=0
cc_433 N_B_M1014_g N_A_329_81#_c_1206_n 0.00480308f $X=2.665 $Y=2.185 $X2=0
+ $Y2=0
cc_434 N_B_c_480_n N_A_329_81#_c_1206_n 9.37421e-19 $X=3.8 $Y=3.075 $X2=0 $Y2=0
cc_435 N_B_c_479_n N_A_329_81#_c_1184_n 9.48738e-19 $X=3.725 $Y=3.15 $X2=0 $Y2=0
cc_436 N_B_c_480_n N_A_329_81#_c_1184_n 0.012978f $X=3.8 $Y=3.075 $X2=0 $Y2=0
cc_437 N_B_M1021_g N_A_329_81#_c_1184_n 0.0176013f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_438 N_B_c_473_n N_A_329_81#_c_1184_n 0.0038981f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_439 N_B_M1014_g N_A_329_81#_c_1185_n 0.00241551f $X=2.665 $Y=2.185 $X2=0
+ $Y2=0
cc_440 N_B_M1016_g N_A_329_81#_c_1179_n 0.00981436f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_441 N_B_M1016_g N_A_329_81#_c_1180_n 0.00795796f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_442 N_B_c_473_n N_A_329_81#_c_1180_n 0.032345f $X=4.24 $Y=1.515 $X2=0 $Y2=0
cc_443 N_B_c_474_n N_A_329_81#_c_1180_n 0.0274616f $X=4.315 $Y=1.515 $X2=0 $Y2=0
cc_444 N_B_M1018_g N_A_329_81#_c_1181_n 0.00561682f $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_445 N_B_M1003_g N_A_329_81#_c_1182_n 0.00493879f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_446 N_B_M1003_g N_A_329_81#_c_1183_n 0.00621366f $X=2.57 $Y=0.945 $X2=0 $Y2=0
cc_447 N_B_M1021_g N_A_329_81#_c_1241_n 0.00103443f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_448 N_B_M1016_g N_VGND_c_1341_n 0.00546687f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_449 N_B_M1018_g N_VGND_c_1346_n 9.15902e-19 $X=1.57 $Y=0.725 $X2=0 $Y2=0
cc_450 N_B_M1016_g N_VGND_c_1346_n 0.00399972f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_451 N_B_M1016_g N_VGND_c_1351_n 0.0052212f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_452 N_A_1027_48#_M1023_g N_C_c_668_n 0.0203498f $X=5.21 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_453 N_A_1027_48#_c_590_n N_C_c_670_n 0.00175105f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_454 N_A_1027_48#_c_591_n N_C_c_670_n 0.0010582f $X=5.49 $Y=1.64 $X2=0 $Y2=0
cc_455 N_A_1027_48#_M1023_g N_C_c_671_n 0.00501499f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_456 N_A_1027_48#_c_590_n N_C_c_671_n 0.00706975f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_457 N_A_1027_48#_c_591_n N_C_c_671_n 0.0158957f $X=5.49 $Y=1.64 $X2=0 $Y2=0
cc_458 N_A_1027_48#_c_592_n N_C_c_671_n 0.00100186f $X=6.532 $Y=1.475 $X2=0
+ $Y2=0
cc_459 N_A_1027_48#_c_593_n N_C_c_671_n 8.39659e-19 $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_460 N_A_1027_48#_M1005_g N_C_M1007_g 0.0309953f $X=5.395 $Y=2.415 $X2=0 $Y2=0
cc_461 N_A_1027_48#_c_590_n N_C_M1007_g 0.0151199f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_462 N_A_1027_48#_c_598_n N_C_M1007_g 0.00111666f $X=6.687 $Y=2.132 $X2=0
+ $Y2=0
cc_463 N_A_1027_48#_c_600_n N_C_M1007_g 0.00467187f $X=6.687 $Y=1.95 $X2=0 $Y2=0
cc_464 N_A_1027_48#_c_592_n N_C_c_673_n 0.00373839f $X=6.532 $Y=1.475 $X2=0
+ $Y2=0
cc_465 N_A_1027_48#_c_593_n N_C_c_673_n 0.00308441f $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_466 N_A_1027_48#_c_598_n N_C_M1020_g 0.00327621f $X=6.687 $Y=2.132 $X2=0
+ $Y2=0
cc_467 N_A_1027_48#_c_594_n N_C_M1020_g 0.00161975f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_468 N_A_1027_48#_c_600_n N_C_M1020_g 0.00464426f $X=6.687 $Y=1.95 $X2=0 $Y2=0
cc_469 N_A_1027_48#_c_590_n N_C_c_674_n 0.0156516f $X=6.39 $Y=1.64 $X2=0 $Y2=0
cc_470 N_A_1027_48#_c_592_n N_C_c_674_n 0.0149313f $X=6.532 $Y=1.475 $X2=0 $Y2=0
cc_471 N_A_1027_48#_c_598_n N_C_c_674_n 6.80956e-19 $X=6.687 $Y=2.132 $X2=0
+ $Y2=0
cc_472 N_A_1027_48#_c_594_n N_C_c_674_n 0.00752536f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_473 N_A_1027_48#_c_598_n N_C_c_675_n 0.0064887f $X=6.687 $Y=2.132 $X2=0 $Y2=0
cc_474 N_A_1027_48#_c_594_n N_C_c_675_n 0.00272504f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_475 N_A_1027_48#_c_592_n N_C_c_676_n 0.00923975f $X=6.532 $Y=1.475 $X2=0
+ $Y2=0
cc_476 N_A_1027_48#_c_598_n N_C_c_676_n 0.00174839f $X=6.687 $Y=2.132 $X2=0
+ $Y2=0
cc_477 N_A_1027_48#_c_594_n N_C_c_676_n 0.0260181f $X=6.532 $Y=1.64 $X2=0 $Y2=0
cc_478 N_A_1027_48#_M1023_g N_A_1057_74#_c_759_n 0.00359689f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_479 N_A_1027_48#_c_598_n N_A_1057_74#_c_768_n 0.0140322f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_480 N_A_1027_48#_M1013_s N_A_1057_74#_c_761_n 0.0013543f $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_481 N_A_1027_48#_c_593_n N_A_1057_74#_c_761_n 0.0127928f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_482 N_A_1027_48#_M1013_s N_A_1057_74#_c_762_n 9.85725e-19 $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_483 N_A_1027_48#_c_590_n N_A_1057_74#_c_762_n 0.00180192f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_484 N_A_1027_48#_c_593_n N_A_1057_74#_c_762_n 0.00977295f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_485 N_A_1027_48#_c_598_n N_A_1057_74#_c_769_n 0.013647f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_486 N_A_1027_48#_M1005_g N_A_1057_74#_c_771_n 0.00445389f $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_487 N_A_1027_48#_M1005_g N_VPWR_c_984_n 0.00602983f $X=5.395 $Y=2.415 $X2=0
+ $Y2=0
cc_488 N_A_1027_48#_M1005_g N_VPWR_c_989_n 0.00589014f $X=5.395 $Y=2.415 $X2=0
+ $Y2=0
cc_489 N_A_1027_48#_M1005_g N_VPWR_c_982_n 0.00608252f $X=5.395 $Y=2.415 $X2=0
+ $Y2=0
cc_490 N_A_1027_48#_M1023_g N_A_335_373#_c_1068_n 0.00376703f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_491 N_A_1027_48#_M1023_g N_A_335_373#_c_1069_n 0.00796217f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_492 N_A_1027_48#_M1005_g N_A_335_373#_c_1069_n 0.00627158f $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_493 N_A_1027_48#_c_590_n N_A_335_373#_c_1069_n 0.0255168f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_494 N_A_1027_48#_c_591_n N_A_335_373#_c_1069_n 0.0115875f $X=5.49 $Y=1.64
+ $X2=0 $Y2=0
cc_495 N_A_1027_48#_M1023_g N_A_335_373#_c_1070_n 0.0134853f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_496 N_A_1027_48#_c_590_n N_A_335_373#_c_1070_n 0.0663436f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_497 N_A_1027_48#_c_591_n N_A_335_373#_c_1070_n 0.00886681f $X=5.49 $Y=1.64
+ $X2=0 $Y2=0
cc_498 N_A_1027_48#_c_593_n N_A_335_373#_c_1070_n 0.0120264f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_499 N_A_1027_48#_M1023_g N_A_335_373#_c_1071_n 2.07613e-19 $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_500 N_A_1027_48#_c_593_n N_A_335_373#_c_1071_n 0.00906723f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_501 N_A_1027_48#_M1005_g N_A_335_373#_c_1081_n 0.00693831f $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_502 N_A_1027_48#_c_590_n N_A_335_373#_c_1081_n 7.34818e-19 $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_503 N_A_1027_48#_c_591_n N_A_335_373#_c_1081_n 0.00484723f $X=5.49 $Y=1.64
+ $X2=0 $Y2=0
cc_504 N_A_1027_48#_M1023_g N_A_335_373#_c_1076_n 0.00454209f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_505 N_A_1027_48#_M1023_g N_A_329_81#_c_1179_n 0.00727684f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_506 N_A_1027_48#_M1023_g N_A_329_81#_c_1180_n 0.00688376f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_507 N_A_1027_48#_M1005_g N_A_329_81#_c_1180_n 0.00262639f $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_508 N_A_1027_48#_M1005_g N_A_329_81#_c_1187_n 0.0186224f $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_509 N_A_1027_48#_c_590_n N_A_329_81#_c_1187_n 0.019188f $X=6.39 $Y=1.64 $X2=0
+ $Y2=0
cc_510 N_A_1027_48#_c_591_n N_A_329_81#_c_1187_n 0.00257854f $X=5.49 $Y=1.64
+ $X2=0 $Y2=0
cc_511 N_A_1027_48#_c_598_n N_A_329_81#_c_1187_n 0.008622f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_512 N_A_1027_48#_M1005_g N_A_329_81#_c_1188_n 0.00187175f $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_513 N_A_1027_48#_c_590_n N_A_329_81#_c_1188_n 0.0216878f $X=6.39 $Y=1.64
+ $X2=0 $Y2=0
cc_514 N_A_1027_48#_c_598_n N_A_329_81#_c_1188_n 0.0318579f $X=6.687 $Y=2.132
+ $X2=0 $Y2=0
cc_515 N_A_1027_48#_M1005_g N_A_329_81#_c_1241_n 7.03353e-19 $X=5.395 $Y=2.415
+ $X2=0 $Y2=0
cc_516 N_A_1027_48#_M1023_g N_VGND_c_1341_n 0.00294228f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_517 N_A_1027_48#_M1023_g N_VGND_c_1342_n 0.00433139f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_518 N_A_1027_48#_M1023_g N_VGND_c_1351_n 0.00823312f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_519 N_C_M1020_g N_A_1057_74#_M1006_g 0.0132317f $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_520 N_C_c_675_n N_A_1057_74#_M1006_g 2.06203e-19 $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_521 N_C_c_675_n N_A_1057_74#_c_755_n 0.0169513f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_522 N_C_c_676_n N_A_1057_74#_c_755_n 3.96458e-19 $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_523 N_C_c_668_n N_A_1057_74#_c_786_n 0.00798135f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_524 N_C_c_668_n N_A_1057_74#_c_758_n 0.0120726f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_525 N_C_c_669_n N_A_1057_74#_c_758_n 7.03833e-19 $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_526 N_C_c_668_n N_A_1057_74#_c_759_n 0.00188363f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_527 N_C_M1007_g N_A_1057_74#_c_768_n 0.00925854f $X=6.01 $Y=2.415 $X2=0 $Y2=0
cc_528 N_C_M1020_g N_A_1057_74#_c_768_n 0.00434263f $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_529 N_C_c_668_n N_A_1057_74#_c_760_n 0.00264822f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_530 N_C_c_673_n N_A_1057_74#_c_761_n 0.0160581f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_531 N_C_c_674_n N_A_1057_74#_c_761_n 3.54962e-19 $X=6.695 $Y=1.515 $X2=0
+ $Y2=0
cc_532 N_C_c_674_n N_A_1057_74#_c_762_n 0.0014427f $X=6.695 $Y=1.515 $X2=0 $Y2=0
cc_533 N_C_M1020_g N_A_1057_74#_c_769_n 0.0165132f $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_534 N_C_c_675_n N_A_1057_74#_c_797_n 7.97692e-19 $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_535 N_C_c_676_n N_A_1057_74#_c_797_n 0.00860034f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_536 N_C_c_675_n N_A_1057_74#_c_799_n 0.00126166f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_537 N_C_c_676_n N_A_1057_74#_c_799_n 0.0135553f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_538 N_C_M1020_g N_A_1057_74#_c_801_n 0.00609446f $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_539 N_C_c_675_n N_A_1057_74#_c_801_n 3.12944e-19 $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_540 N_C_c_676_n N_A_1057_74#_c_801_n 0.0089103f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_541 N_C_M1020_g N_A_1057_74#_c_770_n 0.003601f $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_542 N_C_M1007_g N_A_1057_74#_c_771_n 0.00286409f $X=6.01 $Y=2.415 $X2=0 $Y2=0
cc_543 N_C_c_675_n N_A_1057_74#_c_763_n 0.00221788f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_544 N_C_c_676_n N_A_1057_74#_c_763_n 0.0268459f $X=7.01 $Y=1.515 $X2=0 $Y2=0
cc_545 N_C_c_673_n N_A_1057_74#_c_764_n 0.00377046f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_546 N_C_M1020_g N_VPWR_c_985_n 9.12636e-19 $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_547 N_C_M1007_g N_VPWR_c_989_n 8.60732e-19 $X=6.01 $Y=2.415 $X2=0 $Y2=0
cc_548 N_C_M1020_g N_VPWR_c_989_n 2.1643e-19 $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_549 N_C_c_669_n N_A_335_373#_c_1070_n 0.00532259f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_550 N_C_c_670_n N_A_335_373#_c_1070_n 0.0108015f $X=5.785 $Y=1.16 $X2=0 $Y2=0
cc_551 N_C_c_671_n N_A_335_373#_c_1070_n 0.00787198f $X=6.01 $Y=1.59 $X2=0 $Y2=0
cc_552 N_C_c_668_n N_A_335_373#_c_1071_n 0.0111838f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_553 N_C_c_669_n N_A_335_373#_c_1071_n 0.00410159f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_554 N_C_c_671_n N_A_335_373#_c_1071_n 0.00456415f $X=6.01 $Y=1.59 $X2=0 $Y2=0
cc_555 N_C_c_673_n N_A_335_373#_c_1071_n 0.0035702f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_556 N_C_M1007_g N_A_335_373#_c_1081_n 0.00110201f $X=6.01 $Y=2.415 $X2=0
+ $Y2=0
cc_557 N_C_M1007_g N_A_329_81#_c_1187_n 0.0165138f $X=6.01 $Y=2.415 $X2=0 $Y2=0
cc_558 N_C_M1020_g N_A_329_81#_c_1187_n 0.00295397f $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_559 N_C_M1007_g N_A_329_81#_c_1188_n 0.0103211f $X=6.01 $Y=2.415 $X2=0 $Y2=0
cc_560 N_C_c_674_n N_A_329_81#_c_1188_n 9.00942e-19 $X=6.695 $Y=1.515 $X2=0
+ $Y2=0
cc_561 N_C_M1020_g N_X_c_1309_n 3.07464e-19 $X=7.01 $Y=2.16 $X2=0 $Y2=0
cc_562 N_C_c_668_n N_VGND_c_1342_n 0.00278247f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_563 N_C_c_673_n N_VGND_c_1342_n 5.51389e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_564 N_C_c_673_n N_VGND_c_1350_n 7.18285e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_565 N_C_c_668_n N_VGND_c_1351_n 0.00359137f $X=5.71 $Y=1.085 $X2=0 $Y2=0
cc_566 N_A_1057_74#_c_769_n N_VPWR_M1020_d 0.00427178f $X=7.125 $Y=2.905 $X2=0
+ $Y2=0
cc_567 N_A_1057_74#_c_810_p N_VPWR_M1020_d 0.0182507f $X=7.41 $Y=2.035 $X2=0
+ $Y2=0
cc_568 N_A_1057_74#_c_801_n N_VPWR_M1020_d 0.00177741f $X=7.21 $Y=2.035 $X2=0
+ $Y2=0
cc_569 N_A_1057_74#_c_770_n N_VPWR_M1020_d 0.00213754f $X=7.495 $Y=1.95 $X2=0
+ $Y2=0
cc_570 N_A_1057_74#_M1006_g N_VPWR_c_985_n 0.00481633f $X=7.69 $Y=2.4 $X2=0
+ $Y2=0
cc_571 N_A_1057_74#_c_755_n N_VPWR_c_985_n 3.90858e-19 $X=8.14 $Y=1.605 $X2=0
+ $Y2=0
cc_572 N_A_1057_74#_c_768_n N_VPWR_c_985_n 0.0142846f $X=7.04 $Y=2.99 $X2=0
+ $Y2=0
cc_573 N_A_1057_74#_c_769_n N_VPWR_c_985_n 0.0451976f $X=7.125 $Y=2.905 $X2=0
+ $Y2=0
cc_574 N_A_1057_74#_c_810_p N_VPWR_c_985_n 0.0142694f $X=7.41 $Y=2.035 $X2=0
+ $Y2=0
cc_575 N_A_1057_74#_M1008_g N_VPWR_c_987_n 0.00648292f $X=8.14 $Y=2.4 $X2=0
+ $Y2=0
cc_576 N_A_1057_74#_c_768_n N_VPWR_c_989_n 0.0878491f $X=7.04 $Y=2.99 $X2=0
+ $Y2=0
cc_577 N_A_1057_74#_c_771_n N_VPWR_c_989_n 0.0223379f $X=5.7 $Y=2.82 $X2=0 $Y2=0
cc_578 N_A_1057_74#_M1006_g N_VPWR_c_990_n 0.005209f $X=7.69 $Y=2.4 $X2=0 $Y2=0
cc_579 N_A_1057_74#_M1008_g N_VPWR_c_990_n 0.00503905f $X=8.14 $Y=2.4 $X2=0
+ $Y2=0
cc_580 N_A_1057_74#_M1006_g N_VPWR_c_982_n 0.00987399f $X=7.69 $Y=2.4 $X2=0
+ $Y2=0
cc_581 N_A_1057_74#_M1008_g N_VPWR_c_982_n 0.0093096f $X=8.14 $Y=2.4 $X2=0 $Y2=0
cc_582 N_A_1057_74#_c_768_n N_VPWR_c_982_n 0.0507826f $X=7.04 $Y=2.99 $X2=0
+ $Y2=0
cc_583 N_A_1057_74#_c_771_n N_VPWR_c_982_n 0.0125334f $X=5.7 $Y=2.82 $X2=0 $Y2=0
cc_584 N_A_1057_74#_c_758_n N_A_335_373#_M1019_d 0.00349202f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_585 N_A_1057_74#_c_786_n N_A_335_373#_c_1070_n 0.0239462f $X=5.495 $Y=0.495
+ $X2=0 $Y2=0
cc_586 N_A_1057_74#_c_758_n N_A_335_373#_c_1071_n 0.0242638f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_587 N_A_1057_74#_c_760_n N_A_335_373#_c_1071_n 0.00511588f $X=6.415 $Y=0.66
+ $X2=0 $Y2=0
cc_588 N_A_1057_74#_c_762_n N_A_335_373#_c_1071_n 0.0150383f $X=6.5 $Y=0.745
+ $X2=0 $Y2=0
cc_589 N_A_1057_74#_c_759_n N_A_329_81#_c_1179_n 0.00373319f $X=5.66 $Y=0.34
+ $X2=0 $Y2=0
cc_590 N_A_1057_74#_M1005_d N_A_329_81#_c_1187_n 0.0100632f $X=5.485 $Y=1.995
+ $X2=0 $Y2=0
cc_591 N_A_1057_74#_c_768_n N_A_329_81#_c_1187_n 0.0231978f $X=7.04 $Y=2.99
+ $X2=0 $Y2=0
cc_592 N_A_1057_74#_c_771_n N_A_329_81#_c_1187_n 0.0239502f $X=5.7 $Y=2.82 $X2=0
+ $Y2=0
cc_593 N_A_1057_74#_M1006_g N_X_c_1308_n 0.0139761f $X=7.69 $Y=2.4 $X2=0 $Y2=0
cc_594 N_A_1057_74#_M1008_g N_X_c_1308_n 0.0137472f $X=8.14 $Y=2.4 $X2=0 $Y2=0
cc_595 N_A_1057_74#_c_769_n N_X_c_1308_n 0.00508689f $X=7.125 $Y=2.905 $X2=0
+ $Y2=0
cc_596 N_A_1057_74#_M1006_g N_X_c_1309_n 0.00312384f $X=7.69 $Y=2.4 $X2=0 $Y2=0
cc_597 N_A_1057_74#_c_755_n N_X_c_1309_n 0.0036149f $X=8.14 $Y=1.605 $X2=0 $Y2=0
cc_598 N_A_1057_74#_M1008_g N_X_c_1309_n 0.0022664f $X=8.14 $Y=2.4 $X2=0 $Y2=0
cc_599 N_A_1057_74#_M1006_g N_X_c_1306_n 9.4295e-19 $X=7.69 $Y=2.4 $X2=0 $Y2=0
cc_600 N_A_1057_74#_c_754_n N_X_c_1306_n 9.57805e-19 $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_601 N_A_1057_74#_c_755_n N_X_c_1306_n 0.0227709f $X=8.14 $Y=1.605 $X2=0 $Y2=0
cc_602 N_A_1057_74#_M1008_g N_X_c_1306_n 0.0112732f $X=8.14 $Y=2.4 $X2=0 $Y2=0
cc_603 N_A_1057_74#_c_757_n N_X_c_1306_n 0.00556338f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_604 N_A_1057_74#_c_770_n N_X_c_1306_n 0.00549586f $X=7.495 $Y=1.95 $X2=0
+ $Y2=0
cc_605 N_A_1057_74#_c_763_n N_X_c_1306_n 0.0238938f $X=7.59 $Y=1.505 $X2=0 $Y2=0
cc_606 N_A_1057_74#_c_764_n N_X_c_1306_n 0.00546742f $X=7.582 $Y=1.34 $X2=0
+ $Y2=0
cc_607 N_A_1057_74#_c_754_n X 0.0123221f $X=7.715 $Y=1.34 $X2=0 $Y2=0
cc_608 N_A_1057_74#_c_757_n X 0.00701411f $X=8.145 $Y=1.34 $X2=0 $Y2=0
cc_609 N_A_1057_74#_c_754_n X 0.00260923f $X=7.715 $Y=1.34 $X2=0 $Y2=0
cc_610 N_A_1057_74#_c_755_n X 0.00131295f $X=8.14 $Y=1.605 $X2=0 $Y2=0
cc_611 N_A_1057_74#_c_757_n X 0.00180034f $X=8.145 $Y=1.34 $X2=0 $Y2=0
cc_612 N_A_1057_74#_c_797_n X 0.0123899f $X=7.41 $Y=1.095 $X2=0 $Y2=0
cc_613 N_A_1057_74#_c_761_n N_VGND_M1013_d 0.00352419f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_614 N_A_1057_74#_c_857_p N_VGND_M1013_d 0.00320933f $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_615 N_A_1057_74#_c_797_n N_VGND_M1013_d 0.0227231f $X=7.41 $Y=1.095 $X2=0
+ $Y2=0
cc_616 N_A_1057_74#_c_799_n N_VGND_M1013_d 0.00276146f $X=7.06 $Y=1.095 $X2=0
+ $Y2=0
cc_617 N_A_1057_74#_c_764_n N_VGND_M1013_d 0.00133582f $X=7.582 $Y=1.34 $X2=0
+ $Y2=0
cc_618 N_A_1057_74#_c_758_n N_VGND_c_1342_n 0.0547745f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_1057_74#_c_759_n N_VGND_c_1342_n 0.0236456f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_620 N_A_1057_74#_c_761_n N_VGND_c_1342_n 0.00691154f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_621 N_A_1057_74#_c_757_n N_VGND_c_1344_n 0.00595876f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_622 N_A_1057_74#_c_754_n N_VGND_c_1347_n 0.00472938f $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_623 N_A_1057_74#_c_757_n N_VGND_c_1347_n 0.00472938f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_624 N_A_1057_74#_c_754_n N_VGND_c_1350_n 0.0115709f $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_625 N_A_1057_74#_c_755_n N_VGND_c_1350_n 6.33745e-19 $X=8.14 $Y=1.605 $X2=0
+ $Y2=0
cc_626 N_A_1057_74#_c_758_n N_VGND_c_1350_n 0.0087818f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_1057_74#_c_760_n N_VGND_c_1350_n 0.00301349f $X=6.415 $Y=0.66 $X2=0
+ $Y2=0
cc_628 N_A_1057_74#_c_761_n N_VGND_c_1350_n 0.0280097f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_629 N_A_1057_74#_c_857_p N_VGND_c_1350_n 7.35861e-19 $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_630 N_A_1057_74#_c_797_n N_VGND_c_1350_n 0.0358553f $X=7.41 $Y=1.095 $X2=0
+ $Y2=0
cc_631 N_A_1057_74#_c_754_n N_VGND_c_1351_n 0.00508379f $X=7.715 $Y=1.34 $X2=0
+ $Y2=0
cc_632 N_A_1057_74#_c_757_n N_VGND_c_1351_n 0.00508379f $X=8.145 $Y=1.34 $X2=0
+ $Y2=0
cc_633 N_A_1057_74#_c_758_n N_VGND_c_1351_n 0.0311946f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_634 N_A_1057_74#_c_759_n N_VGND_c_1351_n 0.0127298f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_635 N_A_1057_74#_c_761_n N_VGND_c_1351_n 0.0119702f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_636 N_A_27_373#_c_892_n N_VPWR_c_983_n 0.0200188f $X=0.28 $Y=2.375 $X2=0
+ $Y2=0
cc_637 N_A_27_373#_c_892_n N_VPWR_c_991_n 0.0114213f $X=0.28 $Y=2.375 $X2=0
+ $Y2=0
cc_638 N_A_27_373#_c_892_n N_VPWR_c_982_n 0.0123902f $X=0.28 $Y=2.375 $X2=0
+ $Y2=0
cc_639 N_A_27_373#_c_890_n N_A_335_373#_M1000_d 0.00688224f $X=2.275 $Y=2.65
+ $X2=0 $Y2=0
cc_640 N_A_27_373#_c_881_n N_A_335_373#_c_1077_n 0.0310633f $X=1.63 $Y=2.565
+ $X2=0 $Y2=0
cc_641 N_A_27_373#_c_890_n N_A_335_373#_c_1077_n 0.0154544f $X=2.275 $Y=2.65
+ $X2=0 $Y2=0
cc_642 N_A_27_373#_c_935_n N_A_335_373#_c_1077_n 0.0342077f $X=2.44 $Y=2.01
+ $X2=0 $Y2=0
cc_643 N_A_27_373#_c_882_n N_A_335_373#_c_1066_n 0.00203691f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_644 N_A_27_373#_c_935_n N_A_335_373#_c_1066_n 0.0217586f $X=2.44 $Y=2.01
+ $X2=0 $Y2=0
cc_645 N_A_27_373#_c_884_n N_A_335_373#_c_1066_n 0.0190342f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_646 N_A_27_373#_c_881_n N_A_335_373#_c_1067_n 0.0143553f $X=1.63 $Y=2.565
+ $X2=0 $Y2=0
cc_647 N_A_27_373#_c_882_n N_A_335_373#_c_1067_n 0.0184143f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_648 N_A_27_373#_c_884_n N_A_335_373#_c_1072_n 0.0240865f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_649 N_A_27_373#_M1004_d N_A_335_373#_c_1074_n 7.00965e-19 $X=2.135 $Y=0.845
+ $X2=0 $Y2=0
cc_650 N_A_27_373#_c_935_n N_A_335_373#_c_1074_n 3.4889e-19 $X=2.44 $Y=2.01
+ $X2=0 $Y2=0
cc_651 N_A_27_373#_c_884_n N_A_335_373#_c_1074_n 0.00607915f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_652 N_A_27_373#_c_884_n N_A_335_373#_c_1075_n 0.00608382f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_653 N_A_27_373#_c_882_n N_A_329_81#_M1018_d 0.00206654f $X=2.135 $Y=1.272
+ $X2=-0.19 $Y2=-0.245
cc_654 N_A_27_373#_c_935_n N_A_329_81#_c_1206_n 0.0293668f $X=2.44 $Y=2.01 $X2=0
+ $Y2=0
cc_655 N_A_27_373#_c_890_n N_A_329_81#_c_1185_n 0.00350811f $X=2.275 $Y=2.65
+ $X2=0 $Y2=0
cc_656 N_A_27_373#_c_935_n N_A_329_81#_c_1185_n 0.0125952f $X=2.44 $Y=2.01 $X2=0
+ $Y2=0
cc_657 N_A_27_373#_c_880_n N_A_329_81#_c_1181_n 0.00510362f $X=1.63 $Y=1.38
+ $X2=0 $Y2=0
cc_658 N_A_27_373#_c_882_n N_A_329_81#_c_1181_n 0.0160417f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_659 N_A_27_373#_c_888_n N_A_329_81#_c_1181_n 0.00154277f $X=1.68 $Y=1.295
+ $X2=0 $Y2=0
cc_660 N_A_27_373#_M1004_d N_A_329_81#_c_1182_n 0.00349911f $X=2.135 $Y=0.845
+ $X2=0 $Y2=0
cc_661 N_A_27_373#_c_882_n N_A_329_81#_c_1182_n 0.00580419f $X=2.135 $Y=1.272
+ $X2=0 $Y2=0
cc_662 N_A_27_373#_c_884_n N_A_329_81#_c_1182_n 0.0172834f $X=2.275 $Y=1.11
+ $X2=0 $Y2=0
cc_663 N_A_27_373#_c_879_n N_VGND_c_1340_n 0.0179595f $X=0.32 $Y=0.55 $X2=0
+ $Y2=0
cc_664 N_A_27_373#_c_885_n N_VGND_c_1340_n 8.78751e-19 $X=1.535 $Y=1.295 $X2=0
+ $Y2=0
cc_665 N_A_27_373#_c_879_n N_VGND_c_1345_n 0.0124374f $X=0.32 $Y=0.55 $X2=0
+ $Y2=0
cc_666 N_A_27_373#_c_879_n N_VGND_c_1351_n 0.0114937f $X=0.32 $Y=0.55 $X2=0
+ $Y2=0
cc_667 N_VPWR_M1021_d N_A_329_81#_c_1184_n 0.00600362f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_984_n N_A_329_81#_c_1184_n 0.00866046f $X=4.62 $Y=2.9 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_982_n N_A_329_81#_c_1184_n 0.0271416f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_670 N_VPWR_M1021_d N_A_329_81#_c_1180_n 0.0169398f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_984_n N_A_329_81#_c_1187_n 0.00232914f $X=4.62 $Y=2.9 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_982_n N_A_329_81#_c_1187_n 0.0283293f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_673 N_VPWR_M1021_d N_A_329_81#_c_1241_n 0.00447615f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_984_n N_A_329_81#_c_1241_n 0.0147528f $X=4.62 $Y=2.9 $X2=0 $Y2=0
cc_675 N_VPWR_c_982_n N_A_329_81#_c_1241_n 6.89689e-19 $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_985_n N_X_c_1308_n 0.0235251f $X=7.465 $Y=2.455 $X2=0 $Y2=0
cc_677 N_VPWR_c_990_n N_X_c_1308_n 0.0150868f $X=8.28 $Y=3.33 $X2=0 $Y2=0
cc_678 N_VPWR_c_982_n N_X_c_1308_n 0.012316f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_679 N_VPWR_c_987_n N_X_c_1306_n 0.0423827f $X=8.365 $Y=1.985 $X2=0 $Y2=0
cc_680 N_VPWR_c_987_n N_VGND_c_1344_n 0.00977564f $X=8.365 $Y=1.985 $X2=0 $Y2=0
cc_681 N_A_335_373#_M1003_d N_A_329_81#_c_1178_n 0.00218533f $X=2.645 $Y=0.625
+ $X2=0 $Y2=0
cc_682 N_A_335_373#_c_1073_n N_A_329_81#_c_1178_n 0.0256726f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_683 N_A_335_373#_c_1072_n N_A_329_81#_c_1206_n 0.00277093f $X=2.8 $Y=1.12
+ $X2=0 $Y2=0
cc_684 N_A_335_373#_c_1073_n N_A_329_81#_c_1206_n 0.00875291f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_685 N_A_335_373#_c_1068_n N_A_329_81#_c_1179_n 0.0169928f $X=5.04 $Y=1.305
+ $X2=0 $Y2=0
cc_686 N_A_335_373#_c_1070_n N_A_329_81#_c_1179_n 3.08288e-19 $X=5.83 $Y=1.22
+ $X2=0 $Y2=0
cc_687 N_A_335_373#_c_1073_n N_A_329_81#_c_1179_n 0.00643723f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_688 N_A_335_373#_c_1076_n N_A_329_81#_c_1179_n 0.0032994f $X=5.04 $Y=1.295
+ $X2=0 $Y2=0
cc_689 N_A_335_373#_c_1068_n N_A_329_81#_c_1180_n 0.0126364f $X=5.04 $Y=1.305
+ $X2=0 $Y2=0
cc_690 N_A_335_373#_c_1069_n N_A_329_81#_c_1180_n 0.0505384f $X=5.04 $Y=1.975
+ $X2=0 $Y2=0
cc_691 N_A_335_373#_c_1081_n N_A_329_81#_c_1180_n 0.0197685f $X=5.17 $Y=2.14
+ $X2=0 $Y2=0
cc_692 N_A_335_373#_c_1073_n N_A_329_81#_c_1180_n 0.0264059f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_693 N_A_335_373#_c_1076_n N_A_329_81#_c_1180_n 0.0026622f $X=5.04 $Y=1.295
+ $X2=0 $Y2=0
cc_694 N_A_335_373#_M1005_s N_A_329_81#_c_1187_n 0.00719868f $X=5.03 $Y=1.995
+ $X2=0 $Y2=0
cc_695 N_A_335_373#_c_1081_n N_A_329_81#_c_1187_n 0.0264695f $X=5.17 $Y=2.14
+ $X2=0 $Y2=0
cc_696 N_A_335_373#_c_1074_n N_A_329_81#_c_1182_n 0.00180844f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_697 N_A_335_373#_M1003_d N_A_329_81#_c_1183_n 2.36577e-19 $X=2.645 $Y=0.625
+ $X2=0 $Y2=0
cc_698 N_A_335_373#_c_1072_n N_A_329_81#_c_1183_n 0.0233474f $X=2.8 $Y=1.12
+ $X2=0 $Y2=0
cc_699 N_A_335_373#_c_1074_n N_A_329_81#_c_1183_n 0.00102588f $X=2.785 $Y=1.295
+ $X2=0 $Y2=0
cc_700 N_A_329_81#_c_1178_n N_VGND_M1016_d 0.00993346f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_701 N_A_329_81#_c_1178_n N_VGND_c_1341_n 0.0237317f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_702 N_A_329_81#_c_1179_n N_VGND_c_1341_n 0.00764375f $X=4.67 $Y=0.965 $X2=0
+ $Y2=0
cc_703 N_A_329_81#_c_1179_n N_VGND_c_1342_n 0.0193145f $X=4.67 $Y=0.965 $X2=0
+ $Y2=0
cc_704 N_A_329_81#_c_1178_n N_VGND_c_1346_n 0.0126356f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_705 N_A_329_81#_c_1178_n N_VGND_c_1351_n 0.0244914f $X=4.585 $Y=0.7 $X2=0
+ $Y2=0
cc_706 N_A_329_81#_c_1179_n N_VGND_c_1351_n 0.0191643f $X=4.67 $Y=0.965 $X2=0
+ $Y2=0
cc_707 X N_VGND_c_1344_n 0.0316671f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_708 X N_VGND_c_1347_n 0.0105983f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_709 X N_VGND_c_1350_n 0.0165965f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_710 X N_VGND_c_1351_n 0.0113894f $X=7.835 $Y=0.47 $X2=0 $Y2=0

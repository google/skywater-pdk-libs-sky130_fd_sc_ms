* File: sky130_fd_sc_ms__fa_2.pex.spice
* Created: Fri Aug 28 17:35:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FA_2%A 3 7 11 14 18 22 25 29 31 32 33 34 35 36 42 44
+ 47 51 52 55 56 57 60 62 65 66
c230 36 0 2.13543e-19 $X=4.225 $Y=1.665
c231 35 0 2.31284e-19 $X=6.335 $Y=1.665
c232 34 0 1.12499e-19 $X=2.785 $Y=1.665
c233 33 0 5.276e-20 $X=3.935 $Y=1.665
c234 32 0 1.73388e-19 $X=0.385 $Y=1.665
c235 25 0 1.1376e-19 $X=6.34 $Y=0.765
c236 14 0 1.67707e-19 $X=2.765 $Y=2.235
r237 65 68 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.515
+ $X2=6.43 $Y2=1.68
r238 65 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.515
+ $X2=6.43 $Y2=1.35
r239 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.515 $X2=6.43 $Y2=1.515
r240 60 63 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.41
+ $X2=4.36 $Y2=1.575
r241 60 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.41
+ $X2=4.36 $Y2=1.245
r242 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.41 $X2=4.36 $Y2=1.41
r243 55 58 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.41
+ $X2=2.84 $Y2=1.575
r244 55 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.41
+ $X2=2.84 $Y2=1.245
r245 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.41 $X2=2.84 $Y2=1.41
r246 52 53 1.50625 $w=3.2e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r247 51 72 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.465 $X2=0.27
+ $Y2=1.665
r248 50 52 33.8906 $w=3.2e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.495 $Y2=1.465
r249 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r250 47 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.665
r251 44 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r252 42 61 8.69211 $w=3.93e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.512
+ $X2=4.36 $Y2=1.512
r253 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r254 39 56 8.16535 $w=3.81e-07 $l=3.11288e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.765 $Y2=1.41
r255 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r256 36 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r257 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r258 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=4.225 $Y2=1.665
r259 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r260 33 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r261 33 34 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=2.785 $Y2=1.665
r262 32 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.665
+ $X2=0.24 $Y2=1.665
r263 31 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=2.64 $Y2=1.665
r264 31 32 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=0.385 $Y2=1.665
r265 29 68 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.355 $Y=2.34
+ $X2=6.355 $Y2=1.68
r266 25 67 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=6.34 $Y=0.765
+ $X2=6.34 $Y2=1.35
r267 22 62 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.45 $Y=0.765
+ $X2=4.45 $Y2=1.245
r268 18 63 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.435 $Y=2.235
+ $X2=4.435 $Y2=1.575
r269 14 58 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.765 $Y=2.235
+ $X2=2.765 $Y2=1.575
r270 11 57 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.75 $Y=0.765
+ $X2=2.75 $Y2=1.245
r271 5 52 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r272 5 7 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.765
r273 1 53 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r274 1 3 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%CIN 3 5 7 10 14 17 21 22 25 28 29 30 32 33 34
+ 37 38 41 42 45 46 57 60 62 65 69
c172 42 0 1.67418e-19 $X=3.38 $Y=1.41
c173 41 0 1.12499e-19 $X=3.38 $Y=1.41
c174 38 0 2.638e-20 $X=5.47 $Y=1.41
c175 37 0 1.35287e-19 $X=5.47 $Y=1.41
c176 17 0 1.267e-19 $X=5.395 $Y=2.235
c177 5 0 1.91229e-19 $X=1.86 $Y=1.245
r178 63 65 2.94811 $w=2.13e-07 $l=5.5e-08 $layer=LI1_cond $X=3.545 $Y=2.042
+ $X2=3.6 $Y2=2.042
r179 62 69 0.428816 $w=2.13e-07 $l=8e-09 $layer=LI1_cond $X=4.088 $Y=2.042
+ $X2=4.08 $Y2=2.042
r180 51 53 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.605 $Y=1.41
+ $X2=1.86 $Y2=1.41
r181 46 62 2.14263 $w=2.53e-07 $l=1.12406e-07 $layer=LI1_cond $X=4.126 $Y=1.947
+ $X2=4.088 $Y2=2.042
r182 46 69 2.09048 $w=2.13e-07 $l=3.9e-08 $layer=LI1_cond $X=4.041 $Y=2.042
+ $X2=4.08 $Y2=2.042
r183 45 63 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.042
+ $X2=3.545 $Y2=2.042
r184 45 46 22.8345 $w=2.13e-07 $l=4.26e-07 $layer=LI1_cond $X=3.615 $Y=2.042
+ $X2=4.041 $Y2=2.042
r185 45 65 0.80403 $w=2.13e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=2.042
+ $X2=3.6 $Y2=2.042
r186 42 58 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.575
r187 42 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.245
r188 41 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.575
r189 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.41 $X2=3.38 $Y2=1.41
r190 38 61 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.41
+ $X2=5.47 $Y2=1.575
r191 38 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.41
+ $X2=5.47 $Y2=1.245
r192 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.41 $X2=5.47 $Y2=1.41
r193 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.47 $Y=1.745
+ $X2=5.47 $Y2=1.41
r194 34 46 21.0404 $w=2.53e-07 $l=4.63825e-07 $layer=LI1_cond $X=4.535 $Y=1.83
+ $X2=4.126 $Y2=1.947
r195 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.305 $Y=1.83
+ $X2=5.47 $Y2=1.745
r196 33 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.305 $Y=1.83
+ $X2=4.535 $Y2=1.83
r197 32 45 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.46 $Y=1.935
+ $X2=3.46 $Y2=2.042
r198 32 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.46 $Y=1.935
+ $X2=3.46 $Y2=1.575
r199 29 45 4.65272 $w=1.92e-07 $l=8.84308e-08 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=3.46 $Y2=2.042
r200 29 30 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=3.375 $Y=2.035
+ $X2=2.225 $Y2=2.035
r201 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=1.95
+ $X2=2.225 $Y2=2.035
r202 27 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.14 $Y=1.575
+ $X2=2.14 $Y2=1.95
r203 25 53 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.88 $Y=1.41 $X2=1.86
+ $Y2=1.41
r204 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.41 $X2=1.88 $Y2=1.41
r205 22 27 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=2.055 $Y=1.417
+ $X2=2.14 $Y2=1.575
r206 22 24 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=2.055 $Y=1.417
+ $X2=1.88 $Y2=1.417
r207 21 60 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.52 $Y=0.765
+ $X2=5.52 $Y2=1.245
r208 17 61 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.395 $Y=2.235
+ $X2=5.395 $Y2=1.575
r209 14 57 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.43 $Y=0.765
+ $X2=3.43 $Y2=1.245
r210 10 58 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.34 $Y=2.235
+ $X2=3.34 $Y2=1.575
r211 5 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.245
+ $X2=1.86 $Y2=1.41
r212 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.86 $Y=1.245 $X2=1.86
+ $Y2=0.765
r213 1 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.605 $Y=1.575
+ $X2=1.605 $Y2=1.41
r214 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.605 $Y=1.575
+ $X2=1.605 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%A_339_347# 1 2 9 13 16 20 21 25 27 29 30 32 33
+ 34 36 39 41 45 46 48 51 54 59 61 62 66 70 72 73
c205 46 0 5.68263e-20 $X=4.93 $Y=1.41
c206 45 0 9.88845e-20 $X=4.93 $Y=1.41
c207 25 0 7.90786e-20 $X=7.47 $Y=2.4
r208 72 73 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7 $Y=1.33 $X2=7
+ $Y2=1.255
r209 67 75 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=1.42 $X2=7
+ $Y2=1.585
r210 67 72 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7 $Y=1.42 $X2=7
+ $Y2=1.33
r211 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7 $Y=1.42
+ $X2=7 $Y2=1.42
r212 63 66 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.85 $Y=1.42 $X2=7
+ $Y2=1.42
r213 56 59 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.8 $Y=2.455 $X2=2
+ $Y2=2.455
r214 52 54 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.46 $Y=1.83
+ $X2=1.8 $Y2=1.83
r215 51 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.85 $Y=1.255
+ $X2=6.85 $Y2=1.42
r216 50 51 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.85 $Y=1.09
+ $X2=6.85 $Y2=1.255
r217 49 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=1.005
+ $X2=4.93 $Y2=1.005
r218 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.765 $Y=1.005
+ $X2=6.85 $Y2=1.09
r219 48 49 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=6.765 $Y=1.005
+ $X2=5.095 $Y2=1.005
r220 46 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.93 $Y=1.41
+ $X2=4.93 $Y2=1.575
r221 46 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.93 $Y=1.41
+ $X2=4.93 $Y2=1.245
r222 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.93
+ $Y=1.41 $X2=4.93 $Y2=1.41
r223 43 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.09
+ $X2=4.93 $Y2=1.005
r224 43 45 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.93 $Y=1.09
+ $X2=4.93 $Y2=1.41
r225 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=1.005
+ $X2=2.145 $Y2=1.005
r226 41 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=1.005
+ $X2=4.93 $Y2=1.005
r227 41 42 160.166 $w=1.68e-07 $l=2.455e-06 $layer=LI1_cond $X=4.765 $Y=1.005
+ $X2=2.31 $Y2=1.005
r228 37 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0.92
+ $X2=2.145 $Y2=1.005
r229 37 39 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.145 $Y=0.92
+ $X2=2.145 $Y2=0.54
r230 36 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=2.29 $X2=1.8
+ $Y2=2.455
r231 35 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=1.915
+ $X2=1.8 $Y2=1.83
r232 35 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.8 $Y=1.915
+ $X2=1.8 $Y2=2.29
r233 33 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=1.005
+ $X2=2.145 $Y2=1.005
r234 33 34 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.98 $Y=1.005
+ $X2=1.545 $Y2=1.005
r235 32 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=1.745
+ $X2=1.46 $Y2=1.83
r236 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=1.09
+ $X2=1.545 $Y2=1.005
r237 31 32 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.46 $Y=1.09
+ $X2=1.46 $Y2=1.745
r238 27 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.485 $Y=1.255
+ $X2=7.47 $Y2=1.33
r239 27 29 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.485 $Y=1.255
+ $X2=7.485 $Y2=0.765
r240 23 30 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.47 $Y=1.405
+ $X2=7.47 $Y2=1.33
r241 23 25 386.766 $w=1.8e-07 $l=9.95e-07 $layer=POLY_cond $X=7.47 $Y=1.405
+ $X2=7.47 $Y2=2.4
r242 22 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.33
+ $X2=7 $Y2=1.33
r243 21 30 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.38 $Y=1.33 $X2=7.47
+ $Y2=1.33
r244 21 22 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=7.38 $Y=1.33
+ $X2=7.165 $Y2=1.33
r245 20 73 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.055 $Y=0.765
+ $X2=7.055 $Y2=1.255
r246 16 75 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=6.925 $Y=2.4
+ $X2=6.925 $Y2=1.585
r247 13 70 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.02 $Y=0.765
+ $X2=5.02 $Y2=1.245
r248 9 71 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.885 $Y=2.235
+ $X2=4.885 $Y2=1.575
r249 2 59 600 $w=1.7e-07 $l=8.59069e-07 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=1.735 $X2=2 $Y2=2.455
r250 1 39 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.935
+ $Y=0.395 $X2=2.145 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%B 1 3 4 7 8 9 10 13 16 17 19 22 25 26 28 31 34
+ 35 36 37 38 39 45 48 52
c164 45 0 1.73388e-19 $X=1 $Y=1.41
r165 48 52 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=1.92
r166 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.41
+ $X2=1 $Y2=1.41
r167 42 45 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.75 $Y=1.41 $X2=1
+ $Y2=1.41
r168 40 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.575
+ $X2=0.75 $Y2=1.41
r169 40 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.75 $Y=1.575
+ $X2=0.75 $Y2=1.92
r170 34 39 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.95 $Y=0.765
+ $X2=5.95 $Y2=1.21
r171 29 31 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=5.935 $Y=3.075
+ $X2=5.935 $Y2=2.34
r172 28 39 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.935 $Y=1.3
+ $X2=5.935 $Y2=1.21
r173 28 31 404.258 $w=1.8e-07 $l=1.04e-06 $layer=POLY_cond $X=5.935 $Y=1.3
+ $X2=5.935 $Y2=2.34
r174 27 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.935 $Y=3.15
+ $X2=3.845 $Y2=3.15
r175 26 29 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.845 $Y=3.15
+ $X2=5.935 $Y2=3.075
r176 26 27 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=5.845 $Y=3.15
+ $X2=3.935 $Y2=3.15
r177 25 37 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.86 $Y=0.765
+ $X2=3.86 $Y2=1.21
r178 20 38 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=3.075
+ $X2=3.845 $Y2=3.15
r179 20 22 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=3.845 $Y=3.075
+ $X2=3.845 $Y2=2.39
r180 19 37 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.845 $Y=1.3
+ $X2=3.845 $Y2=1.21
r181 19 22 423.694 $w=1.8e-07 $l=1.09e-06 $layer=POLY_cond $X=3.845 $Y=1.3
+ $X2=3.845 $Y2=2.39
r182 18 36 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.435 $Y=3.15
+ $X2=2.345 $Y2=3.15
r183 17 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.755 $Y=3.15
+ $X2=3.845 $Y2=3.15
r184 17 18 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=3.755 $Y=3.15
+ $X2=2.435 $Y2=3.15
r185 16 35 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.36 $Y=0.765
+ $X2=2.36 $Y2=1.21
r186 11 36 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.345 $Y=3.075
+ $X2=2.345 $Y2=3.15
r187 11 13 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=2.345 $Y=3.075
+ $X2=2.345 $Y2=2.235
r188 10 35 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.345 $Y=1.3
+ $X2=2.345 $Y2=1.21
r189 10 13 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=2.345 $Y=1.3
+ $X2=2.345 $Y2=2.235
r190 8 36 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.255 $Y=3.15
+ $X2=2.345 $Y2=3.15
r191 8 9 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=2.255 $Y=3.15
+ $X2=1.245 $Y2=3.15
r192 5 9 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.155 $Y=3.075
+ $X2=1.245 $Y2=3.15
r193 5 7 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=1.155 $Y=3.075
+ $X2=1.155 $Y2=2.235
r194 4 46 46.8708 $w=3.37e-07 $l=3.07164e-07 $layer=POLY_cond $X=1.155 $Y=1.665
+ $X2=1.04 $Y2=1.41
r195 4 7 221.565 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=1.155 $Y=1.665
+ $X2=1.155 $Y2=2.235
r196 1 46 38.6529 $w=3.37e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.14 $Y=1.245
+ $X2=1.04 $Y2=1.41
r197 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.14 $Y=1.245 $X2=1.14
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%A_995_347# 1 2 9 13 15 19 23 25 26 28 33 35 40
+ 45 47 49
c119 35 0 1.48077e-19 $X=5.17 $Y=2.195
c120 33 0 1.3983e-19 $X=7.965 $Y=2.32
r121 49 50 32.4387 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.087 $Y=1.395
+ $X2=8.087 $Y2=1.32
r122 46 52 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.087 $Y=1.485
+ $X2=8.087 $Y2=1.65
r123 46 49 14.2284 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=8.087 $Y=1.485
+ $X2=8.087 $Y2=1.395
r124 45 48 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.057 $Y=1.485
+ $X2=8.057 $Y2=1.65
r125 45 47 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.057 $Y=1.485
+ $X2=8.057 $Y2=1.32
r126 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.07
+ $Y=1.485 $X2=8.07 $Y2=1.485
r127 40 42 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=5.305 $Y=0.56
+ $X2=5.305 $Y2=0.66
r128 35 37 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.17 $Y=2.195
+ $X2=5.17 $Y2=2.405
r129 33 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.965 $Y=2.32
+ $X2=7.965 $Y2=1.65
r130 30 47 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.965 $Y=0.745
+ $X2=7.965 $Y2=1.32
r131 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=0.66
+ $X2=5.305 $Y2=0.66
r132 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.88 $Y=0.66
+ $X2=7.965 $Y2=0.745
r133 28 29 157.23 $w=1.68e-07 $l=2.41e-06 $layer=LI1_cond $X=7.88 $Y=0.66
+ $X2=5.47 $Y2=0.66
r134 27 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.405
+ $X2=5.17 $Y2=2.405
r135 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.88 $Y=2.405
+ $X2=7.965 $Y2=2.32
r136 26 27 166.037 $w=1.68e-07 $l=2.545e-06 $layer=LI1_cond $X=7.88 $Y=2.405
+ $X2=5.335 $Y2=2.405
r137 21 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.61 $Y2=1.395
r138 21 23 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.625 $Y2=0.765
r139 17 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.61 $Y=1.47
+ $X2=8.61 $Y2=1.395
r140 17 19 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=8.61 $Y=1.47 $X2=8.61
+ $Y2=2.4
r141 16 49 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=8.27 $Y=1.395
+ $X2=8.087 $Y2=1.395
r142 15 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.52 $Y=1.395
+ $X2=8.61 $Y2=1.395
r143 15 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.52 $Y=1.395
+ $X2=8.27 $Y2=1.395
r144 13 50 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.195 $Y=0.765
+ $X2=8.195 $Y2=1.32
r145 9 52 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.16 $Y=2.4 $X2=8.16
+ $Y2=1.65
r146 2 35 300 $w=1.7e-07 $l=5.48908e-07 $layer=licon1_PDIFF $count=2 $X=4.975
+ $Y=1.735 $X2=5.17 $Y2=2.195
r147 1 40 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.095
+ $Y=0.395 $X2=5.305 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%A_27_378# 1 2 9 13 15 17 19
r38 19 21 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.38 $Y=2.25
+ $X2=1.38 $Y2=2.405
r39 16 17 3.9231 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.27 $Y2=2.405
r40 15 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=1.38 $Y2=2.405
r41 15 16 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.215 $Y=2.405
+ $X2=0.445 $Y2=2.405
r42 11 17 2.80976 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.49 $X2=0.27
+ $Y2=2.405
r43 11 13 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.27 $Y=2.49
+ $X2=0.27 $Y2=2.745
r44 7 17 2.80976 $w=3.4e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.26 $Y=2.32
+ $X2=0.27 $Y2=2.405
r45 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.26 $Y=2.32 $X2=0.26
+ $Y2=2.035
r46 2 19 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.245
+ $Y=1.735 $X2=1.38 $Y2=2.25
r47 1 13 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.89 $X2=0.28 $Y2=2.745
r48 1 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.89 $X2=0.26 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%VPWR 1 2 3 4 5 6 21 25 29 33 35 37 42 43 45 46
+ 47 49 61 72 76 82 85 88 96
r111 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r112 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 88 91 11.8458 $w=5.18e-07 $l=5.15e-07 $layer=LI1_cond $X=7.79 $Y=2.815
+ $X2=7.79 $Y2=3.33
r114 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r115 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 80 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 80 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r119 77 91 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=8.05 $Y=3.33
+ $X2=7.79 $Y2=3.33
r120 77 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.05 $Y=3.33
+ $X2=8.4 $Y2=3.33
r121 76 95 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.75 $Y=3.33
+ $X2=8.935 $Y2=3.33
r122 76 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.75 $Y=3.33
+ $X2=8.4 $Y2=3.33
r123 75 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r124 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r125 72 91 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=7.53 $Y=3.33
+ $X2=7.79 $Y2=3.33
r126 72 74 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.53 $Y=3.33 $X2=7.44
+ $Y2=3.33
r127 71 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r128 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r129 67 70 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 65 85 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.097 $Y2=3.33
r131 65 67 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.56 $Y2=3.33
r132 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 61 85 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.097 $Y2=3.33
r135 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r139 57 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r141 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 54 82 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=0.812 $Y2=3.33
r143 54 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 52 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 49 82 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.812 $Y2=3.33
r147 49 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 47 71 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r149 47 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 47 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 45 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.535 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=3.33
+ $X2=6.7 $Y2=3.33
r153 44 74 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.865 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.865 $Y=3.33
+ $X2=6.7 $Y2=3.33
r155 42 59 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.64 $Y2=3.33
r156 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.99 $Y2=3.33
r157 41 63 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.6 $Y2=3.33
r158 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=2.99 $Y2=3.33
r159 37 40 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.875 $Y=1.985
+ $X2=8.875 $Y2=2.815
r160 35 95 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=8.875 $Y=3.245
+ $X2=8.935 $Y2=3.33
r161 35 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.875 $Y=3.245
+ $X2=8.875 $Y2=2.815
r162 31 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.7 $Y=3.245 $X2=6.7
+ $Y2=3.33
r163 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.7 $Y=3.245
+ $X2=6.7 $Y2=2.78
r164 27 85 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.097 $Y=3.245
+ $X2=4.097 $Y2=3.33
r165 27 29 14.9668 $w=3.83e-07 $l=5e-07 $layer=LI1_cond $X=4.097 $Y=3.245
+ $X2=4.097 $Y2=2.745
r166 23 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=3.33
r167 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=2.455
r168 19 82 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.812 $Y=3.245
+ $X2=0.812 $Y2=3.33
r169 19 21 14.5879 $w=3.93e-07 $l=5e-07 $layer=LI1_cond $X=0.812 $Y=3.245
+ $X2=0.812 $Y2=2.745
r170 6 40 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.84 $X2=8.835 $Y2=2.815
r171 6 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.84 $X2=8.835 $Y2=1.985
r172 5 88 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=7.56
+ $Y=1.84 $X2=7.79 $Y2=2.815
r173 4 33 600 $w=1.7e-07 $l=1.05986e-06 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=1.84 $X2=6.7 $Y2=2.78
r174 3 29 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.89 $X2=4.095 $Y2=2.745
r175 2 25 600 $w=1.7e-07 $l=7.84602e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.735 $X2=2.99 $Y2=2.455
r176 1 21 600 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.89 $X2=0.81 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%A_686_347# 1 2 9 15 16
c34 15 0 1.267e-19 $X=4.66 $Y=2.44
c35 9 0 1.67707e-19 $X=3.57 $Y=2.405
r36 15 16 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.515
+ $X2=4.495 $Y2=2.515
r37 9 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=2.405 $X2=3.57
+ $Y2=2.485
r38 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=2.405
+ $X2=3.57 $Y2=2.405
r39 8 16 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.735 $Y=2.405
+ $X2=4.495 $Y2=2.405
r40 2 15 600 $w=1.7e-07 $l=7.69545e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.735 $X2=4.66 $Y2=2.44
r41 1 12 600 $w=1.7e-07 $l=8.17007e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.735 $X2=3.57 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%COUT 1 2 7 12 13 16
c29 7 0 1.1376e-19 $X=7.385 $Y=1
r30 13 16 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.985
+ $X2=7.385 $Y2=1.985
r31 13 16 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.37 $Y=1.985
+ $X2=7.385 $Y2=1.985
r32 13 18 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.37 $Y=1.985
+ $X2=7.195 $Y2=1.985
r33 12 13 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=1.82
+ $X2=7.47 $Y2=1.985
r34 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=7.47 $Y=1.085
+ $X2=7.47 $Y2=1.82
r35 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=1
+ $X2=7.47 $Y2=1.085
r36 7 9 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.385 $Y=1 $X2=7.27
+ $Y2=1
r37 2 18 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=1.84 $X2=7.195 $Y2=1.985
r38 1 9 182 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.395 $X2=7.27 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%SUM 1 2 9 13 14 15 16 23 32
c41 14 0 7.90786e-20 $X=8.315 $Y=1.95
r42 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=8.397 $Y=1.997
+ $X2=8.397 $Y2=2.035
r43 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=8.397 $Y=2.405
+ $X2=8.397 $Y2=2.775
r44 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=8.397 $Y=1.973
+ $X2=8.397 $Y2=1.997
r45 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=8.397 $Y=1.973
+ $X2=8.397 $Y2=1.82
r46 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=8.397 $Y=2.058
+ $X2=8.397 $Y2=2.405
r47 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=8.397 $Y=2.058
+ $X2=8.397 $Y2=2.035
r48 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.49 $Y=1.15
+ $X2=8.49 $Y2=1.82
r49 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.41 $Y=0.985
+ $X2=8.41 $Y2=1.15
r50 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.41 $Y=0.985
+ $X2=8.41 $Y2=0.54
r51 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.25
+ $Y=1.84 $X2=8.385 $Y2=1.985
r52 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.25
+ $Y=1.84 $X2=8.385 $Y2=2.815
r53 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.395 $X2=8.41 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%A_27_79# 1 2 9 11 12 14 15 17
c36 11 0 1.91229e-19 $X=1.035 $Y=0.99
r37 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.205 $Y=0.585
+ $X2=1.5 $Y2=0.585
r38 13 15 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.12 $Y=0.75
+ $X2=1.205 $Y2=0.585
r39 13 14 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.12 $Y=0.75
+ $X2=1.12 $Y2=0.905
r40 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=0.99
+ $X2=1.12 $Y2=0.905
r41 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.035 $Y=0.99
+ $X2=0.445 $Y2=0.99
r42 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.905
+ $X2=0.445 $Y2=0.99
r43 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.28 $Y=0.905
+ $X2=0.28 $Y2=0.54
r44 2 17 182 $w=1.7e-07 $l=3.67933e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.395 $X2=1.5 $Y2=0.585
r45 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.395 $X2=0.28 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%VGND 1 2 3 4 5 6 21 25 27 29 31 33 38 46 51 56
+ 61 67 70 74 88 95
r100 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r101 88 91 8.50545 $w=4.48e-07 $l=3.2e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.84
+ $Y2=0.32
r102 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r103 74 77 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.155 $Y=0
+ $X2=4.155 $Y2=0.325
r104 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r106 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 65 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r108 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r109 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r110 62 88 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.065 $Y=0 $X2=7.84
+ $Y2=0
r111 62 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.065 $Y=0 $X2=8.4
+ $Y2=0
r112 61 94 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.937 $Y2=0
r113 61 64 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=0 $X2=8.4
+ $Y2=0
r114 60 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r115 60 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r116 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r117 57 59 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.925 $Y=0
+ $X2=7.44 $Y2=0
r118 56 88 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.84
+ $Y2=0
r119 56 59 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.615 $Y=0
+ $X2=7.44 $Y2=0
r120 52 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.155
+ $Y2=0
r121 52 54 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.56
+ $Y2=0
r122 51 84 8.41198 $w=4.53e-07 $l=3.2e-07 $layer=LI1_cond $X=6.697 $Y=0
+ $X2=6.697 $Y2=0.32
r123 51 57 6.56868 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=6.697 $Y=0
+ $X2=6.925 $Y2=0
r124 51 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r125 51 54 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=6.47 $Y=0 $X2=4.56
+ $Y2=0
r126 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r127 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r128 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r129 47 70 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.055
+ $Y2=0
r130 47 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.6
+ $Y2=0
r131 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.155
+ $Y2=0
r132 46 49 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.6
+ $Y2=0
r133 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r134 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r135 42 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r136 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r137 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r138 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r139 39 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.74
+ $Y2=0
r140 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r141 38 70 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.055
+ $Y2=0
r142 38 44 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r143 36 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r144 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r145 33 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.74
+ $Y2=0
r146 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r147 31 82 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r148 31 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r149 31 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r150 27 94 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.937 $Y2=0
r151 27 29 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0.54
r152 23 70 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r153 23 25 10.6709 $w=5.08e-07 $l=4.55e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.54
r154 19 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r155 19 21 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.555
r156 6 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.395 $X2=8.84 $Y2=0.54
r157 5 91 182 $w=1.7e-07 $l=3.15278e-07 $layer=licon1_NDIFF $count=1 $X=7.56
+ $Y=0.395 $X2=7.84 $Y2=0.32
r158 4 84 182 $w=1.7e-07 $l=3.15278e-07 $layer=licon1_NDIFF $count=1 $X=6.415
+ $Y=0.395 $X2=6.695 $Y2=0.32
r159 3 77 182 $w=1.7e-07 $l=2.52587e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.395 $X2=4.155 $Y2=0.325
r160 2 25 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.395 $X2=3.055 $Y2=0.54
r161 1 21 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.395 $X2=0.78 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__FA_2%A_701_79# 1 2 10 15 16
r29 15 16 10.9068 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.735 $Y=0.585
+ $X2=4.5 $Y2=0.585
r30 10 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.645 $Y=0.56
+ $X2=3.645 $Y2=0.665
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0.665
+ $X2=3.645 $Y2=0.665
r32 8 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.81 $Y=0.665 $X2=4.5
+ $Y2=0.665
r33 2 15 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.395 $X2=4.735 $Y2=0.585
r34 1 10 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.395 $X2=3.645 $Y2=0.56
.ends


* File: sky130_fd_sc_ms__and4bb_1.pxi.spice
* Created: Fri Aug 28 17:14:25 2020
* 
x_PM_SKY130_FD_SC_MS__AND4BB_1%A_N N_A_N_M1002_g N_A_N_M1013_g A_N N_A_N_c_102_n
+ N_A_N_c_103_n PM_SKY130_FD_SC_MS__AND4BB_1%A_N
x_PM_SKY130_FD_SC_MS__AND4BB_1%A_179_48# N_A_179_48#_M1003_s N_A_179_48#_M1008_d
+ N_A_179_48#_M1005_d N_A_179_48#_M1001_g N_A_179_48#_M1012_g
+ N_A_179_48#_c_132_n N_A_179_48#_c_133_n N_A_179_48#_c_134_n
+ N_A_179_48#_c_135_n N_A_179_48#_c_136_n N_A_179_48#_c_142_n
+ N_A_179_48#_c_143_n N_A_179_48#_c_144_n N_A_179_48#_c_137_n
+ N_A_179_48#_c_138_n N_A_179_48#_c_139_n N_A_179_48#_c_145_n
+ PM_SKY130_FD_SC_MS__AND4BB_1%A_179_48#
x_PM_SKY130_FD_SC_MS__AND4BB_1%A_27_74# N_A_27_74#_M1013_s N_A_27_74#_M1002_s
+ N_A_27_74#_M1008_g N_A_27_74#_M1003_g N_A_27_74#_c_238_n N_A_27_74#_c_239_n
+ N_A_27_74#_c_240_n N_A_27_74#_c_241_n N_A_27_74#_c_246_n N_A_27_74#_c_242_n
+ N_A_27_74#_c_243_n N_A_27_74#_c_249_n PM_SKY130_FD_SC_MS__AND4BB_1%A_27_74#
x_PM_SKY130_FD_SC_MS__AND4BB_1%A_503_48# N_A_503_48#_M1009_d N_A_503_48#_M1010_d
+ N_A_503_48#_M1004_g N_A_503_48#_M1007_g N_A_503_48#_c_323_n
+ N_A_503_48#_c_324_n N_A_503_48#_c_325_n N_A_503_48#_c_326_n
+ N_A_503_48#_c_327_n N_A_503_48#_c_349_n N_A_503_48#_c_328_n
+ N_A_503_48#_c_335_n N_A_503_48#_c_336_n N_A_503_48#_c_329_n
+ N_A_503_48#_c_330_n PM_SKY130_FD_SC_MS__AND4BB_1%A_503_48#
x_PM_SKY130_FD_SC_MS__AND4BB_1%C N_C_M1011_g N_C_M1005_g N_C_c_413_n N_C_c_418_n
+ C N_C_c_414_n N_C_c_415_n PM_SKY130_FD_SC_MS__AND4BB_1%C
x_PM_SKY130_FD_SC_MS__AND4BB_1%D N_D_M1000_g N_D_M1006_g N_D_c_456_n N_D_c_461_n
+ D N_D_c_457_n N_D_c_458_n PM_SKY130_FD_SC_MS__AND4BB_1%D
x_PM_SKY130_FD_SC_MS__AND4BB_1%B_N N_B_N_M1010_g N_B_N_M1009_g B_N N_B_N_c_500_n
+ N_B_N_c_501_n PM_SKY130_FD_SC_MS__AND4BB_1%B_N
x_PM_SKY130_FD_SC_MS__AND4BB_1%VPWR N_VPWR_M1002_d N_VPWR_M1008_s N_VPWR_M1007_d
+ N_VPWR_M1006_d N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n
+ N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_536_n N_VPWR_c_537_n
+ N_VPWR_c_538_n VPWR N_VPWR_c_539_n N_VPWR_c_528_n N_VPWR_c_541_n
+ PM_SKY130_FD_SC_MS__AND4BB_1%VPWR
x_PM_SKY130_FD_SC_MS__AND4BB_1%X N_X_M1001_d N_X_M1012_d N_X_c_593_n N_X_c_594_n
+ N_X_c_595_n N_X_c_599_n X N_X_c_597_n PM_SKY130_FD_SC_MS__AND4BB_1%X
x_PM_SKY130_FD_SC_MS__AND4BB_1%VGND N_VGND_M1013_d N_VGND_M1000_d N_VGND_c_629_n
+ N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n VGND N_VGND_c_633_n
+ N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n PM_SKY130_FD_SC_MS__AND4BB_1%VGND
cc_1 VNB N_A_N_M1002_g 0.00164739f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_2 VNB N_A_N_M1013_g 0.0410018f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_3 VNB N_A_N_c_102_n 0.00427511f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A_N_c_103_n 0.0580678f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_5 VNB N_A_179_48#_M1001_g 0.027508f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_6 VNB N_A_179_48#_M1012_g 0.00188615f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_7 VNB N_A_179_48#_c_132_n 0.0173958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_179_48#_c_133_n 0.00566753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_179_48#_c_134_n 0.0108078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_179_48#_c_135_n 0.00552356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_179_48#_c_136_n 0.00371726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_179_48#_c_137_n 0.0429901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_179_48#_c_138_n 0.00402396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_179_48#_c_139_n 0.0156032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_M1003_g 0.0304942f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_16 VNB N_A_27_74#_c_238_n 0.0252878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_239_n 0.00307298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_240_n 0.00912492f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.665
cc_19 VNB N_A_27_74#_c_241_n 0.00471389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_242_n 0.00288195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_243_n 0.0418726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_503_48#_c_323_n 0.0180921f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_23 VNB N_A_503_48#_c_324_n 0.0233755f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_24 VNB N_A_503_48#_c_325_n 0.0024279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_503_48#_c_326_n 0.00106996f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.665
cc_26 VNB N_A_503_48#_c_327_n 0.0166374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_503_48#_c_328_n 0.00741585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_503_48#_c_329_n 0.0290446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_503_48#_c_330_n 0.0184362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_M1011_g 0.0235303f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_31 VNB N_C_c_413_n 0.0187725f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_32 VNB N_C_c_414_n 0.0152048f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_33 VNB N_C_c_415_n 0.00452729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_M1000_g 0.0243691f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_35 VNB N_D_c_456_n 0.0191427f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_36 VNB N_D_c_457_n 0.0153308f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_37 VNB N_D_c_458_n 0.0035566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_N_M1010_g 0.00151951f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_39 VNB N_B_N_M1009_g 0.0394675f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_40 VNB N_B_N_c_500_n 0.0607038f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_41 VNB N_B_N_c_501_n 0.00477584f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_42 VNB N_VPWR_c_528_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_593_n 0.00354223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_594_n 0.00216891f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_45 VNB N_X_c_595_n 0.00202082f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_46 VNB N_VGND_c_629_n 0.00647573f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_47 VNB N_VGND_c_630_n 0.00961301f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_48 VNB N_VGND_c_631_n 0.0844452f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_49 VNB N_VGND_c_632_n 0.007312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_633_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.252 $Y2=1.665
cc_51 VNB N_VGND_c_634_n 0.0219533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_635_n 0.295025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_636_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VPB N_A_N_M1002_g 0.0285752f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_55 VPB N_A_N_c_102_n 0.00810644f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_56 VPB N_A_179_48#_M1012_g 0.0277691f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_57 VPB N_A_179_48#_c_136_n 0.00312957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_179_48#_c_142_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_179_48#_c_143_n 0.0139431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_179_48#_c_144_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_179_48#_c_145_n 0.00606315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_74#_M1008_g 0.0235767f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_63 VPB N_A_27_74#_c_241_n 0.00110211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_74#_c_246_n 0.0131844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_74#_c_242_n 0.00534047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_74#_c_243_n 0.0397806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_74#_c_249_n 0.0343789f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_503_48#_M1007_g 0.0330815f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_69 VPB N_A_503_48#_c_325_n 0.0132216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_503_48#_c_326_n 0.00115078f $X=-0.19 $Y=1.66 $X2=0.252 $Y2=1.665
cc_71 VPB N_A_503_48#_c_328_n 0.00242007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_503_48#_c_335_n 0.0139052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_503_48#_c_336_n 0.0358457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_C_M1005_g 0.0282876f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_75 VPB N_C_c_413_n 0.00209955f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_76 VPB N_C_c_418_n 0.0145689f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_77 VPB N_C_c_415_n 0.00289358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_D_M1006_g 0.0289646f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_79 VPB N_D_c_456_n 0.00214097f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_80 VPB N_D_c_461_n 0.016036f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_81 VPB N_D_c_458_n 0.00194081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_B_N_M1010_g 0.048426f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_83 VPB N_B_N_c_501_n 0.00929358f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_84 VPB N_VPWR_c_529_n 0.0169261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_530_n 0.0118941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_531_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_532_n 0.00976275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_533_n 0.0257133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_534_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_535_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_536_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_537_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_538_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_539_n 0.0204244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_528_n 0.0746133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_541_n 0.0274712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_X_c_593_n 0.00103109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_X_c_597_n 0.00636858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 N_A_N_M1013_g N_A_179_48#_M1001_g 0.0215682f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_100 N_A_N_M1002_g N_A_179_48#_M1012_g 0.0203866f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_101 N_A_N_c_103_n N_A_179_48#_c_132_n 0.0265647f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_102 N_A_N_M1013_g N_A_27_74#_c_238_n 0.00509125f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_103 N_A_N_M1013_g N_A_27_74#_c_239_n 0.0197241f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_104 N_A_N_c_102_n N_A_27_74#_c_239_n 0.00260541f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_105 N_A_N_c_103_n N_A_27_74#_c_239_n 0.00104609f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_106 N_A_N_c_102_n N_A_27_74#_c_240_n 0.0217424f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_107 N_A_N_c_103_n N_A_27_74#_c_240_n 0.00197868f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_108 N_A_N_M1002_g N_A_27_74#_c_241_n 0.0114233f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_109 N_A_N_M1013_g N_A_27_74#_c_241_n 0.00443834f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_110 N_A_N_c_102_n N_A_27_74#_c_241_n 0.0345406f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_111 N_A_N_c_103_n N_A_27_74#_c_241_n 0.00850438f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_112 N_A_N_M1002_g N_A_27_74#_c_249_n 0.0316039f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_113 N_A_N_c_102_n N_A_27_74#_c_249_n 0.023616f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_114 N_A_N_c_103_n N_A_27_74#_c_249_n 0.0014745f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A_N_M1002_g N_VPWR_c_529_n 0.00339971f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_116 N_A_N_M1002_g N_VPWR_c_528_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_117 N_A_N_M1002_g N_VPWR_c_541_n 0.0046462f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_118 N_A_N_c_103_n N_X_c_593_n 0.00102244f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_119 N_A_N_M1002_g N_X_c_599_n 2.8446e-19 $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_120 N_A_N_M1013_g N_VGND_c_629_n 0.0124836f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_121 N_A_N_M1013_g N_VGND_c_633_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_122 N_A_N_M1013_g N_VGND_c_635_n 0.00761198f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_123 N_A_179_48#_c_136_n N_A_27_74#_M1008_g 0.00143909f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_124 N_A_179_48#_c_142_n N_A_27_74#_M1008_g 0.0010204f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_125 N_A_179_48#_c_145_n N_A_27_74#_M1008_g 0.00653712f $X=2.42 $Y=2.115 $X2=0
+ $Y2=0
cc_126 N_A_179_48#_c_133_n N_A_27_74#_M1003_g 0.00398916f $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_127 N_A_179_48#_c_136_n N_A_27_74#_M1003_g 0.0074719f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_128 N_A_179_48#_c_139_n N_A_27_74#_M1003_g 0.0201006f $X=1.985 $Y=0.515 $X2=0
+ $Y2=0
cc_129 N_A_179_48#_M1001_g N_A_27_74#_c_239_n 0.00122398f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_179_48#_M1001_g N_A_27_74#_c_241_n 0.00215077f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_131 N_A_179_48#_c_132_n N_A_27_74#_c_241_n 0.00151958f $X=0.895 $Y=1.3 $X2=0
+ $Y2=0
cc_132 N_A_179_48#_M1012_g N_A_27_74#_c_246_n 0.0156128f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_133 N_A_179_48#_M1012_g N_A_27_74#_c_242_n 0.00542795f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_134 N_A_179_48#_c_133_n N_A_27_74#_c_242_n 7.3914e-19 $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_135 N_A_179_48#_c_134_n N_A_27_74#_c_242_n 0.00226272f $X=1.82 $Y=0.945 $X2=0
+ $Y2=0
cc_136 N_A_179_48#_c_136_n N_A_27_74#_c_242_n 0.0521373f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_137 N_A_179_48#_c_137_n N_A_27_74#_c_242_n 3.42035e-19 $X=1.38 $Y=1.465 $X2=0
+ $Y2=0
cc_138 N_A_179_48#_c_138_n N_A_27_74#_c_242_n 0.0258568f $X=1.525 $Y=1.465 $X2=0
+ $Y2=0
cc_139 N_A_179_48#_c_139_n N_A_27_74#_c_242_n 0.0144437f $X=1.985 $Y=0.515 $X2=0
+ $Y2=0
cc_140 N_A_179_48#_c_145_n N_A_27_74#_c_242_n 0.010758f $X=2.42 $Y=2.115 $X2=0
+ $Y2=0
cc_141 N_A_179_48#_M1012_g N_A_27_74#_c_243_n 0.00492004f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_179_48#_c_134_n N_A_27_74#_c_243_n 0.00121947f $X=1.82 $Y=0.945 $X2=0
+ $Y2=0
cc_143 N_A_179_48#_c_136_n N_A_27_74#_c_243_n 0.0166905f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_144 N_A_179_48#_c_137_n N_A_27_74#_c_243_n 0.0213513f $X=1.38 $Y=1.465 $X2=0
+ $Y2=0
cc_145 N_A_179_48#_c_138_n N_A_27_74#_c_243_n 0.00207719f $X=1.525 $Y=1.465
+ $X2=0 $Y2=0
cc_146 N_A_179_48#_c_139_n N_A_27_74#_c_243_n 0.00516793f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_147 N_A_179_48#_M1012_g N_A_27_74#_c_249_n 0.00584805f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_148 N_A_179_48#_c_136_n N_A_503_48#_M1007_g 0.00411626f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_149 N_A_179_48#_c_142_n N_A_503_48#_M1007_g 0.012829f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_150 N_A_179_48#_c_143_n N_A_503_48#_M1007_g 0.0138343f $X=3.295 $Y=2.115
+ $X2=0 $Y2=0
cc_151 N_A_179_48#_c_144_n N_A_503_48#_M1007_g 3.9273e-19 $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_152 N_A_179_48#_c_145_n N_A_503_48#_M1007_g 0.00215558f $X=2.42 $Y=2.115
+ $X2=0 $Y2=0
cc_153 N_A_179_48#_c_139_n N_A_503_48#_c_323_n 0.00961636f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_154 N_A_179_48#_c_136_n N_A_503_48#_c_324_n 0.00961636f $X=2.3 $Y=2.03 $X2=0
+ $Y2=0
cc_155 N_A_179_48#_c_143_n N_A_503_48#_c_325_n 4.47545e-19 $X=3.295 $Y=2.115
+ $X2=0 $Y2=0
cc_156 N_A_179_48#_c_145_n N_A_503_48#_c_325_n 0.00213307f $X=2.42 $Y=2.115
+ $X2=0 $Y2=0
cc_157 N_A_179_48#_c_143_n N_A_503_48#_c_326_n 0.012887f $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_158 N_A_179_48#_c_139_n N_A_503_48#_c_326_n 0.0571916f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_159 N_A_179_48#_c_145_n N_A_503_48#_c_326_n 0.00460395f $X=2.42 $Y=2.115
+ $X2=0 $Y2=0
cc_160 N_A_179_48#_c_139_n N_A_503_48#_c_349_n 0.0145967f $X=1.985 $Y=0.515
+ $X2=0 $Y2=0
cc_161 N_A_179_48#_c_143_n N_A_503_48#_c_335_n 0.00386511f $X=3.295 $Y=2.115
+ $X2=0 $Y2=0
cc_162 N_A_179_48#_c_142_n N_C_M1005_g 3.9273e-19 $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_163 N_A_179_48#_c_143_n N_C_M1005_g 0.0153389f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_164 N_A_179_48#_c_144_n N_C_M1005_g 0.0128377f $X=3.46 $Y=2.265 $X2=0 $Y2=0
cc_165 N_A_179_48#_c_143_n N_C_c_418_n 0.00274264f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_166 N_A_179_48#_c_136_n N_C_c_415_n 0.0022031f $X=2.3 $Y=2.03 $X2=0 $Y2=0
cc_167 N_A_179_48#_c_143_n N_C_c_415_n 0.0260806f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_168 N_A_179_48#_c_143_n N_D_M1006_g 0.00482442f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_169 N_A_179_48#_c_144_n N_D_M1006_g 0.0123693f $X=3.46 $Y=2.265 $X2=0 $Y2=0
cc_170 N_A_179_48#_c_143_n N_D_c_458_n 0.00997848f $X=3.295 $Y=2.115 $X2=0 $Y2=0
cc_171 N_A_179_48#_c_143_n N_B_N_M1010_g 4.33296e-19 $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_172 N_A_179_48#_c_143_n N_VPWR_M1007_d 0.00276506f $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_173 N_A_179_48#_M1012_g N_VPWR_c_529_n 0.0224743f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_179_48#_M1012_g N_VPWR_c_530_n 0.00970676f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_179_48#_c_142_n N_VPWR_c_530_n 0.0127976f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_176 N_A_179_48#_c_142_n N_VPWR_c_531_n 0.0236791f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_177 N_A_179_48#_c_143_n N_VPWR_c_531_n 0.0208278f $X=3.295 $Y=2.115 $X2=0
+ $Y2=0
cc_178 N_A_179_48#_c_144_n N_VPWR_c_531_n 0.0236791f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_179 N_A_179_48#_c_144_n N_VPWR_c_532_n 0.0244142f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_180 N_A_179_48#_M1012_g N_VPWR_c_533_n 0.00460063f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_179_48#_c_142_n N_VPWR_c_535_n 0.014549f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_182 N_A_179_48#_c_144_n N_VPWR_c_537_n 0.0144623f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_183 N_A_179_48#_M1012_g N_VPWR_c_528_n 0.00465993f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_179_48#_c_142_n N_VPWR_c_528_n 0.0119743f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_185 N_A_179_48#_c_144_n N_VPWR_c_528_n 0.0118344f $X=3.46 $Y=2.265 $X2=0
+ $Y2=0
cc_186 N_A_179_48#_M1001_g N_X_c_593_n 0.00581287f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_179_48#_M1012_g N_X_c_593_n 0.00679574f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_179_48#_c_132_n N_X_c_593_n 0.0122329f $X=0.895 $Y=1.3 $X2=0 $Y2=0
cc_189 N_A_179_48#_c_133_n N_X_c_593_n 0.00761824f $X=1.525 $Y=1.3 $X2=0 $Y2=0
cc_190 N_A_179_48#_c_138_n N_X_c_593_n 0.023711f $X=1.525 $Y=1.465 $X2=0 $Y2=0
cc_191 N_A_179_48#_M1001_g N_X_c_594_n 0.00163355f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_179_48#_c_135_n N_X_c_594_n 0.00798712f $X=1.61 $Y=0.945 $X2=0 $Y2=0
cc_193 N_A_179_48#_c_139_n N_X_c_594_n 0.0181191f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_194 N_A_179_48#_M1001_g N_X_c_595_n 0.0096135f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_179_48#_c_132_n N_X_c_595_n 0.00721571f $X=0.895 $Y=1.3 $X2=0 $Y2=0
cc_196 N_A_179_48#_c_133_n N_X_c_595_n 0.00777787f $X=1.525 $Y=1.3 $X2=0 $Y2=0
cc_197 N_A_179_48#_c_135_n N_X_c_595_n 0.0057961f $X=1.61 $Y=0.945 $X2=0 $Y2=0
cc_198 N_A_179_48#_c_138_n N_X_c_595_n 0.00150313f $X=1.525 $Y=1.465 $X2=0 $Y2=0
cc_199 N_A_179_48#_M1012_g N_X_c_599_n 0.00784453f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_179_48#_M1012_g N_X_c_597_n 0.0110388f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_179_48#_c_137_n N_X_c_597_n 0.01137f $X=1.38 $Y=1.465 $X2=0 $Y2=0
cc_202 N_A_179_48#_c_138_n N_X_c_597_n 0.0230181f $X=1.525 $Y=1.465 $X2=0 $Y2=0
cc_203 N_A_179_48#_M1001_g N_VGND_c_629_n 0.00364992f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_204 N_A_179_48#_M1001_g N_VGND_c_631_n 0.00461464f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_179_48#_c_139_n N_VGND_c_631_n 0.0246732f $X=1.985 $Y=0.515 $X2=0
+ $Y2=0
cc_206 N_A_179_48#_M1001_g N_VGND_c_635_n 0.00913048f $X=0.97 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_179_48#_c_134_n N_VGND_c_635_n 0.00711624f $X=1.82 $Y=0.945 $X2=0
+ $Y2=0
cc_208 N_A_179_48#_c_135_n N_VGND_c_635_n 0.00631461f $X=1.61 $Y=0.945 $X2=0
+ $Y2=0
cc_209 N_A_179_48#_c_139_n N_VGND_c_635_n 0.02007f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_210 N_A_179_48#_c_139_n A_455_74# 0.00765047f $X=1.985 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_211 N_A_27_74#_c_243_n N_A_503_48#_M1007_g 0.0218313f $X=1.92 $Y=1.455 $X2=0
+ $Y2=0
cc_212 N_A_27_74#_M1003_g N_A_503_48#_c_323_n 0.0397166f $X=2.2 $Y=0.69 $X2=0
+ $Y2=0
cc_213 N_A_27_74#_c_243_n N_A_503_48#_c_324_n 0.0397166f $X=1.92 $Y=1.455 $X2=0
+ $Y2=0
cc_214 N_A_27_74#_M1003_g N_A_503_48#_c_326_n 7.44855e-19 $X=2.2 $Y=0.69 $X2=0
+ $Y2=0
cc_215 N_A_27_74#_c_241_n N_VPWR_M1002_d 9.23293e-19 $X=0.655 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_27_74#_c_246_n N_VPWR_M1002_d 0.00739353f $X=1.78 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_27_74#_c_249_n N_VPWR_M1002_d 0.00508114f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_218 N_A_27_74#_c_246_n N_VPWR_M1008_s 0.0044551f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_219 N_A_27_74#_c_242_n N_VPWR_M1008_s 0.00217969f $X=1.92 $Y=1.455 $X2=0
+ $Y2=0
cc_220 N_A_27_74#_c_246_n N_VPWR_c_529_n 0.0142591f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_221 N_A_27_74#_c_249_n N_VPWR_c_529_n 0.00969384f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_222 N_A_27_74#_M1008_g N_VPWR_c_530_n 0.0105369f $X=2.185 $Y=2.54 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_246_n N_VPWR_c_530_n 0.0213589f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_243_n N_VPWR_c_530_n 6.89412e-19 $X=1.92 $Y=1.455 $X2=0
+ $Y2=0
cc_225 N_A_27_74#_M1008_g N_VPWR_c_535_n 0.00460063f $X=2.185 $Y=2.54 $X2=0
+ $Y2=0
cc_226 N_A_27_74#_M1008_g N_VPWR_c_528_n 0.00909121f $X=2.185 $Y=2.54 $X2=0
+ $Y2=0
cc_227 N_A_27_74#_c_246_n N_VPWR_c_528_n 0.0288733f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_228 N_A_27_74#_c_249_n N_VPWR_c_528_n 0.0177556f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_249_n N_VPWR_c_541_n 0.006683f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_230 N_A_27_74#_c_246_n N_X_M1012_d 0.0129431f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_241_n N_X_c_593_n 0.0506331f $X=0.655 $Y=1.95 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_243_n N_X_c_593_n 0.00109412f $X=1.92 $Y=1.455 $X2=0 $Y2=0
cc_233 N_A_27_74#_c_239_n N_X_c_595_n 0.0139665f $X=0.57 $Y=1.045 $X2=0 $Y2=0
cc_234 N_A_27_74#_c_241_n N_X_c_599_n 0.00561332f $X=0.655 $Y=1.95 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_246_n N_X_c_599_n 0.00986066f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_246_n N_X_c_597_n 0.0324778f $X=1.78 $Y=2.405 $X2=0 $Y2=0
cc_237 N_A_27_74#_c_242_n N_X_c_597_n 0.0235675f $X=1.92 $Y=1.455 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_243_n N_X_c_597_n 0.00166447f $X=1.92 $Y=1.455 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_239_n N_VGND_M1013_d 0.00233685f $X=0.57 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_27_74#_c_238_n N_VGND_c_629_n 0.0164982f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_239_n N_VGND_c_629_n 0.0146425f $X=0.57 $Y=1.045 $X2=0 $Y2=0
cc_242 N_A_27_74#_M1003_g N_VGND_c_631_n 0.00291513f $X=2.2 $Y=0.69 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_238_n N_VGND_c_633_n 0.011066f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_244 N_A_27_74#_M1003_g N_VGND_c_635_n 0.00363725f $X=2.2 $Y=0.69 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_238_n N_VGND_c_635_n 0.00915947f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_246 N_A_503_48#_c_323_n N_C_M1011_g 0.0281202f $X=2.68 $Y=1.12 $X2=0 $Y2=0
cc_247 N_A_503_48#_c_326_n N_C_M1011_g 0.00266937f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_248 N_A_503_48#_c_327_n N_C_M1011_g 0.00388845f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_249 N_A_503_48#_c_330_n N_C_M1011_g 0.0129618f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_250 N_A_503_48#_M1007_g N_C_M1005_g 0.017142f $X=2.685 $Y=2.54 $X2=0 $Y2=0
cc_251 N_A_503_48#_c_324_n N_C_c_413_n 0.012461f $X=2.68 $Y=1.625 $X2=0 $Y2=0
cc_252 N_A_503_48#_M1007_g N_C_c_418_n 0.00291082f $X=2.685 $Y=2.54 $X2=0 $Y2=0
cc_253 N_A_503_48#_c_325_n N_C_c_418_n 0.012461f $X=2.68 $Y=1.79 $X2=0 $Y2=0
cc_254 N_A_503_48#_c_326_n N_C_c_414_n 6.90861e-19 $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_255 N_A_503_48#_c_327_n N_C_c_414_n 0.012461f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_256 N_A_503_48#_c_330_n N_C_c_414_n 0.00265283f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_257 N_A_503_48#_M1007_g N_C_c_415_n 6.97875e-19 $X=2.685 $Y=2.54 $X2=0 $Y2=0
cc_258 N_A_503_48#_c_326_n N_C_c_415_n 0.0469689f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_259 N_A_503_48#_c_327_n N_C_c_415_n 0.00337482f $X=2.68 $Y=1.285 $X2=0 $Y2=0
cc_260 N_A_503_48#_c_330_n N_C_c_415_n 0.0257971f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_261 N_A_503_48#_c_328_n N_D_M1000_g 0.00303034f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_262 N_A_503_48#_c_329_n N_D_M1000_g 0.001133f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_263 N_A_503_48#_c_330_n N_D_M1000_g 0.0129805f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_264 N_A_503_48#_c_328_n N_D_M1006_g 0.00171397f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_265 N_A_503_48#_c_335_n N_D_M1006_g 0.0027246f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_266 N_A_503_48#_c_336_n N_D_M1006_g 9.11033e-19 $X=4.48 $Y=2.265 $X2=0 $Y2=0
cc_267 N_A_503_48#_c_328_n N_D_c_457_n 0.00418923f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_268 N_A_503_48#_c_330_n N_D_c_457_n 0.00521595f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_269 N_A_503_48#_c_328_n N_D_c_458_n 0.050868f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_270 N_A_503_48#_c_330_n N_D_c_458_n 0.0295937f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_271 N_A_503_48#_c_328_n N_B_N_M1010_g 0.0117678f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_272 N_A_503_48#_c_335_n N_B_N_M1010_g 0.0197662f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_273 N_A_503_48#_c_336_n N_B_N_M1010_g 0.0153897f $X=4.48 $Y=2.265 $X2=0 $Y2=0
cc_274 N_A_503_48#_c_328_n N_B_N_M1009_g 0.00739013f $X=4.145 $Y=1.95 $X2=0
+ $Y2=0
cc_275 N_A_503_48#_c_329_n N_B_N_M1009_g 0.0261445f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_276 N_A_503_48#_c_328_n N_B_N_c_500_n 0.00949279f $X=4.145 $Y=1.95 $X2=0
+ $Y2=0
cc_277 N_A_503_48#_c_335_n N_B_N_c_500_n 0.0031002f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_278 N_A_503_48#_c_329_n N_B_N_c_500_n 0.00276952f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_279 N_A_503_48#_c_328_n N_B_N_c_501_n 0.0345409f $X=4.145 $Y=1.95 $X2=0 $Y2=0
cc_280 N_A_503_48#_c_335_n N_B_N_c_501_n 0.0200264f $X=4.48 $Y=2.12 $X2=0 $Y2=0
cc_281 N_A_503_48#_c_329_n N_B_N_c_501_n 0.0156602f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_282 N_A_503_48#_M1007_g N_VPWR_c_530_n 4.24825e-19 $X=2.685 $Y=2.54 $X2=0
+ $Y2=0
cc_283 N_A_503_48#_M1007_g N_VPWR_c_531_n 0.00203999f $X=2.685 $Y=2.54 $X2=0
+ $Y2=0
cc_284 N_A_503_48#_c_335_n N_VPWR_c_532_n 0.00529238f $X=4.48 $Y=2.12 $X2=0
+ $Y2=0
cc_285 N_A_503_48#_c_336_n N_VPWR_c_532_n 0.0266809f $X=4.48 $Y=2.265 $X2=0
+ $Y2=0
cc_286 N_A_503_48#_M1007_g N_VPWR_c_535_n 0.005209f $X=2.685 $Y=2.54 $X2=0 $Y2=0
cc_287 N_A_503_48#_c_336_n N_VPWR_c_539_n 0.014549f $X=4.48 $Y=2.265 $X2=0 $Y2=0
cc_288 N_A_503_48#_M1007_g N_VPWR_c_528_n 0.00983143f $X=2.685 $Y=2.54 $X2=0
+ $Y2=0
cc_289 N_A_503_48#_c_336_n N_VPWR_c_528_n 0.0119743f $X=4.48 $Y=2.265 $X2=0
+ $Y2=0
cc_290 N_A_503_48#_c_329_n N_VGND_M1000_d 0.00182175f $X=4.52 $Y=0.85 $X2=0
+ $Y2=0
cc_291 N_A_503_48#_c_330_n N_VGND_M1000_d 0.00379698f $X=4.06 $Y=0.94 $X2=0
+ $Y2=0
cc_292 N_A_503_48#_c_329_n N_VGND_c_630_n 0.0142603f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_293 N_A_503_48#_c_330_n N_VGND_c_630_n 0.0262201f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_294 N_A_503_48#_c_323_n N_VGND_c_631_n 0.00461464f $X=2.68 $Y=1.12 $X2=0
+ $Y2=0
cc_295 N_A_503_48#_c_329_n N_VGND_c_634_n 0.0102877f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_296 N_A_503_48#_c_323_n N_VGND_c_635_n 0.00585788f $X=2.68 $Y=1.12 $X2=0
+ $Y2=0
cc_297 N_A_503_48#_c_349_n N_VGND_c_635_n 0.0104896f $X=2.845 $Y=0.935 $X2=0
+ $Y2=0
cc_298 N_A_503_48#_c_329_n N_VGND_c_635_n 0.0193098f $X=4.52 $Y=0.85 $X2=0 $Y2=0
cc_299 N_A_503_48#_c_330_n N_VGND_c_635_n 0.029238f $X=4.06 $Y=0.94 $X2=0 $Y2=0
cc_300 N_A_503_48#_c_349_n A_533_74# 0.00294599f $X=2.845 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_301 N_A_503_48#_c_330_n A_533_74# 0.00398078f $X=4.06 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_302 N_A_503_48#_c_330_n A_647_74# 0.00498776f $X=4.06 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_303 N_C_M1011_g N_D_M1000_g 0.034747f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_304 N_C_M1005_g N_D_M1006_g 0.0268601f $X=3.235 $Y=2.54 $X2=0 $Y2=0
cc_305 N_C_c_413_n N_D_c_456_n 0.013848f $X=3.22 $Y=1.695 $X2=0 $Y2=0
cc_306 N_C_c_418_n N_D_c_461_n 0.013848f $X=3.22 $Y=1.86 $X2=0 $Y2=0
cc_307 N_C_c_414_n N_D_c_457_n 0.013848f $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_308 N_C_c_415_n N_D_c_457_n 6.62791e-19 $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_309 N_C_c_414_n N_D_c_458_n 0.00412737f $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_310 N_C_c_415_n N_D_c_458_n 0.0535897f $X=3.22 $Y=1.355 $X2=0 $Y2=0
cc_311 N_C_M1005_g N_VPWR_c_531_n 0.00343717f $X=3.235 $Y=2.54 $X2=0 $Y2=0
cc_312 N_C_M1005_g N_VPWR_c_537_n 0.005209f $X=3.235 $Y=2.54 $X2=0 $Y2=0
cc_313 N_C_M1005_g N_VPWR_c_528_n 0.00982687f $X=3.235 $Y=2.54 $X2=0 $Y2=0
cc_314 N_C_M1011_g N_VGND_c_630_n 0.00207664f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_315 N_C_M1011_g N_VGND_c_631_n 0.00461464f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_316 N_C_M1011_g N_VGND_c_635_n 0.00469123f $X=3.16 $Y=0.69 $X2=0 $Y2=0
cc_317 N_D_M1006_g N_B_N_M1010_g 0.0210205f $X=3.685 $Y=2.54 $X2=0 $Y2=0
cc_318 N_D_c_456_n N_B_N_M1010_g 0.0146356f $X=3.76 $Y=1.695 $X2=0 $Y2=0
cc_319 N_D_M1000_g N_B_N_M1009_g 0.0168987f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_320 N_D_c_457_n N_B_N_M1009_g 0.00363085f $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_321 N_D_c_457_n N_B_N_c_500_n 0.0146356f $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_322 N_D_c_458_n N_B_N_c_500_n 5.47444e-19 $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_323 N_D_M1006_g N_VPWR_c_532_n 0.00741505f $X=3.685 $Y=2.54 $X2=0 $Y2=0
cc_324 N_D_c_461_n N_VPWR_c_532_n 0.0028675f $X=3.76 $Y=1.86 $X2=0 $Y2=0
cc_325 N_D_c_458_n N_VPWR_c_532_n 0.002774f $X=3.76 $Y=1.355 $X2=0 $Y2=0
cc_326 N_D_M1006_g N_VPWR_c_537_n 0.005209f $X=3.685 $Y=2.54 $X2=0 $Y2=0
cc_327 N_D_M1006_g N_VPWR_c_528_n 0.00983291f $X=3.685 $Y=2.54 $X2=0 $Y2=0
cc_328 N_D_M1000_g N_VGND_c_630_n 0.0168272f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_329 N_D_M1000_g N_VGND_c_631_n 0.00383152f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_330 N_D_M1000_g N_VGND_c_635_n 0.00386851f $X=3.67 $Y=0.69 $X2=0 $Y2=0
cc_331 N_B_N_M1010_g N_VPWR_c_532_n 0.00369134f $X=4.255 $Y=2.54 $X2=0 $Y2=0
cc_332 N_B_N_M1010_g N_VPWR_c_539_n 0.005209f $X=4.255 $Y=2.54 $X2=0 $Y2=0
cc_333 N_B_N_M1010_g N_VPWR_c_528_n 0.00986606f $X=4.255 $Y=2.54 $X2=0 $Y2=0
cc_334 N_B_N_M1009_g N_VGND_c_630_n 0.00548248f $X=4.305 $Y=0.735 $X2=0 $Y2=0
cc_335 N_B_N_M1009_g N_VGND_c_634_n 0.00491683f $X=4.305 $Y=0.735 $X2=0 $Y2=0
cc_336 N_B_N_M1009_g N_VGND_c_635_n 0.00517496f $X=4.305 $Y=0.735 $X2=0 $Y2=0
cc_337 N_X_c_594_n N_VGND_c_629_n 0.00133028f $X=1.185 $Y=0.515 $X2=0 $Y2=0
cc_338 N_X_c_594_n N_VGND_c_631_n 0.00832263f $X=1.185 $Y=0.515 $X2=0 $Y2=0
cc_339 N_X_c_594_n N_VGND_c_635_n 0.00691792f $X=1.185 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__nand4_1.pxi.spice
* Created: Fri Aug 28 17:44:19 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4_1%D N_D_M1001_g N_D_M1000_g D N_D_c_49_n N_D_c_50_n
+ PM_SKY130_FD_SC_MS__NAND4_1%D
x_PM_SKY130_FD_SC_MS__NAND4_1%C N_C_M1003_g N_C_M1002_g C N_C_c_78_n N_C_c_79_n
+ N_C_c_80_n PM_SKY130_FD_SC_MS__NAND4_1%C
x_PM_SKY130_FD_SC_MS__NAND4_1%B N_B_M1006_g N_B_M1005_g B N_B_c_113_n
+ N_B_c_114_n PM_SKY130_FD_SC_MS__NAND4_1%B
x_PM_SKY130_FD_SC_MS__NAND4_1%A N_A_c_147_n N_A_M1007_g N_A_M1004_g A
+ N_A_c_150_n PM_SKY130_FD_SC_MS__NAND4_1%A
x_PM_SKY130_FD_SC_MS__NAND4_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_M1004_d
+ N_VPWR_c_171_n N_VPWR_c_172_n N_VPWR_c_173_n N_VPWR_c_174_n N_VPWR_c_175_n
+ N_VPWR_c_176_n N_VPWR_c_177_n N_VPWR_c_178_n VPWR N_VPWR_c_179_n
+ N_VPWR_c_170_n PM_SKY130_FD_SC_MS__NAND4_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND4_1%Y N_Y_M1007_d N_Y_M1001_d N_Y_M1005_d N_Y_c_210_n
+ N_Y_c_211_n N_Y_c_212_n N_Y_c_215_n N_Y_c_216_n N_Y_c_217_n N_Y_c_218_n
+ N_Y_c_219_n N_Y_c_213_n N_Y_c_220_n N_Y_c_221_n Y
+ PM_SKY130_FD_SC_MS__NAND4_1%Y
x_PM_SKY130_FD_SC_MS__NAND4_1%VGND N_VGND_M1000_s VGND N_VGND_c_288_n
+ N_VGND_c_289_n N_VGND_c_290_n PM_SKY130_FD_SC_MS__NAND4_1%VGND
cc_1 VNB N_D_M1001_g 0.00688438f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=2.4
cc_2 VNB D 0.00341988f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_D_c_49_n 0.0347653f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_4 VNB N_D_c_50_n 0.0194922f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.22
cc_5 VNB N_C_M1002_g 0.00681246f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.74
cc_6 VNB N_C_c_78_n 0.0282144f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_7 VNB N_C_c_79_n 0.00766751f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_8 VNB N_C_c_80_n 0.0183508f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.22
cc_9 VNB N_B_M1005_g 0.00701818f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.74
cc_10 VNB B 0.0119609f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_B_c_113_n 0.0283504f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_12 VNB N_B_c_114_n 0.0199072f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.22
cc_13 VNB N_A_c_147_n 0.0243771f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.55
cc_14 VNB N_A_M1004_g 0.00957504f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.74
cc_15 VNB A 0.00941175f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A_c_150_n 0.0590986f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.55
cc_17 VNB N_VPWR_c_170_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_210_n 0.0314733f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_19 VNB N_Y_c_211_n 0.0122962f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_20 VNB N_Y_c_212_n 0.00970183f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.22
cc_21 VNB N_Y_c_213_n 0.021252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_288_n 0.0660892f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB N_VGND_c_289_n 0.186373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_290_n 0.0431564f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.385
cc_25 VPB N_D_M1001_g 0.0247393f $X=-0.19 $Y=1.66 $X2=0.815 $Y2=2.4
cc_26 VPB N_C_M1002_g 0.0243208f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=0.74
cc_27 VPB N_B_M1005_g 0.0254654f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=0.74
cc_28 VPB N_A_M1004_g 0.0301467f $X=-0.19 $Y=1.66 $X2=0.83 $Y2=0.74
cc_29 VPB N_VPWR_c_171_n 0.0476283f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.385
cc_30 VPB N_VPWR_c_172_n 0.00983862f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.385
cc_31 VPB N_VPWR_c_173_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_174_n 0.0555518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_175_n 0.0140765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_176_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_177_n 0.0194903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_178_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_179_n 0.0196506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_170_n 0.0657728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_Y_c_210_n 0.00301672f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.385
cc_40 VPB N_Y_c_215_n 0.00729924f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.55
cc_41 VPB N_Y_c_216_n 0.0138507f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.295
cc_42 VPB N_Y_c_217_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.74 $Y2=1.385
cc_43 VPB N_Y_c_218_n 0.00325836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_Y_c_219_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_220_n 0.00807857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_221_n 0.0104108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 N_D_M1001_g N_C_M1002_g 0.0230875f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_48 N_D_c_49_n N_C_c_78_n 0.0359258f $X=0.74 $Y=1.385 $X2=0 $Y2=0
cc_49 D N_C_c_79_n 0.0283697f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_50 N_D_c_50_n N_C_c_79_n 0.00224093f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_51 D N_C_c_80_n 4.15144e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_D_c_50_n N_C_c_80_n 0.0359258f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_53 N_D_M1001_g N_VPWR_c_171_n 0.00534567f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_54 N_D_M1001_g N_VPWR_c_177_n 0.005209f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_55 N_D_M1001_g N_VPWR_c_170_n 0.00986837f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_56 N_D_M1001_g N_Y_c_210_n 0.00503397f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_57 D N_Y_c_210_n 0.027973f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_D_c_49_n N_Y_c_210_n 0.00739878f $X=0.74 $Y=1.385 $X2=0 $Y2=0
cc_59 N_D_c_50_n N_Y_c_210_n 0.00497484f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_60 D N_Y_c_211_n 0.0228656f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_61 N_D_c_49_n N_Y_c_211_n 0.001011f $X=0.74 $Y=1.385 $X2=0 $Y2=0
cc_62 N_D_c_50_n N_Y_c_211_n 0.0131907f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_63 N_D_M1001_g N_Y_c_215_n 0.0147493f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_64 D N_Y_c_215_n 0.0221856f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_D_c_49_n N_Y_c_215_n 0.00105037f $X=0.74 $Y=1.385 $X2=0 $Y2=0
cc_66 N_D_M1001_g N_Y_c_217_n 0.0108099f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_67 N_D_M1001_g N_Y_c_220_n 0.0114456f $X=0.815 $Y=2.4 $X2=0 $Y2=0
cc_68 D N_Y_c_220_n 0.00234631f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_D_c_50_n N_VGND_c_288_n 0.0036777f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_70 N_D_c_50_n N_VGND_c_289_n 0.00366857f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_71 N_D_c_50_n N_VGND_c_290_n 0.0112037f $X=0.74 $Y=1.22 $X2=0 $Y2=0
cc_72 N_C_M1002_g N_B_M1005_g 0.0360708f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_73 N_C_c_78_n B 4.18645e-19 $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_74 N_C_c_79_n B 0.02242f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_75 N_C_c_78_n N_B_c_113_n 0.0181621f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_76 N_C_c_79_n N_B_c_113_n 4.20537e-19 $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_77 N_C_c_80_n N_B_c_114_n 0.032462f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_78 N_C_M1002_g N_VPWR_c_172_n 0.00755984f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_79 N_C_M1002_g N_VPWR_c_177_n 0.005209f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_80 N_C_M1002_g N_VPWR_c_170_n 0.00983699f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_81 N_C_c_78_n N_Y_c_211_n 0.00101617f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_82 N_C_c_79_n N_Y_c_211_n 0.0255539f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_83 N_C_c_80_n N_Y_c_211_n 0.0122562f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_84 N_C_M1002_g N_Y_c_217_n 0.0126469f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_85 N_C_M1002_g N_Y_c_219_n 9.00138e-19 $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_86 N_C_M1002_g N_Y_c_220_n 0.0050215f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_87 N_C_c_78_n N_Y_c_220_n 8.17195e-19 $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_88 N_C_c_79_n N_Y_c_220_n 0.0103162f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_89 N_C_M1002_g N_Y_c_221_n 0.0196884f $X=1.265 $Y=2.4 $X2=0 $Y2=0
cc_90 N_C_c_78_n N_Y_c_221_n 0.0025662f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_91 N_C_c_79_n N_Y_c_221_n 0.014607f $X=1.31 $Y=1.385 $X2=0 $Y2=0
cc_92 N_C_c_80_n N_VGND_c_288_n 0.00461464f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_93 N_C_c_80_n N_VGND_c_289_n 0.00465551f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_94 N_C_c_80_n N_VGND_c_290_n 0.00180509f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_95 B N_A_c_147_n 0.00346899f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_96 N_B_c_114_n N_A_c_147_n 0.029851f $X=1.88 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_97 N_B_M1005_g N_A_M1004_g 0.0195543f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_98 B A 0.0306948f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B_c_113_n A 2.22676e-19 $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_100 N_B_c_113_n N_A_c_150_n 0.0176224f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_101 N_B_M1005_g N_VPWR_c_172_n 0.00743436f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_102 N_B_M1005_g N_VPWR_c_174_n 8.41409e-19 $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_103 N_B_M1005_g N_VPWR_c_179_n 0.005209f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_104 N_B_M1005_g N_VPWR_c_170_n 0.00984379f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_105 B N_Y_c_211_n 0.0392923f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B_c_113_n N_Y_c_211_n 0.00101286f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_107 N_B_c_114_n N_Y_c_211_n 0.013201f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_108 N_B_M1005_g N_Y_c_217_n 8.93548e-19 $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_109 N_B_M1005_g N_Y_c_218_n 0.00167657f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_110 B N_Y_c_218_n 0.0206854f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B_c_113_n N_Y_c_218_n 0.00176239f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_112 N_B_M1005_g N_Y_c_219_n 0.0128032f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_113 N_B_c_114_n N_Y_c_213_n 0.00223389f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_114 N_B_M1005_g N_Y_c_220_n 4.42656e-19 $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_115 N_B_M1005_g N_Y_c_221_n 0.0196884f $X=1.875 $Y=2.4 $X2=0 $Y2=0
cc_116 B N_Y_c_221_n 0.0117795f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B_c_113_n N_Y_c_221_n 0.00174473f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_118 N_B_c_114_n N_VGND_c_288_n 0.00461464f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_119 N_B_c_114_n N_VGND_c_289_n 0.00467093f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_120 N_A_M1004_g N_VPWR_c_174_n 0.0207018f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_121 A N_VPWR_c_174_n 0.0191168f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A_c_150_n N_VPWR_c_174_n 0.00223706f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_123 N_A_M1004_g N_VPWR_c_179_n 0.00460063f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_M1004_g N_VPWR_c_170_n 0.00909121f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_c_147_n N_Y_c_211_n 0.0145395f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_126 A N_Y_c_211_n 0.0237695f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A_c_150_n N_Y_c_211_n 0.0019436f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A_M1004_g N_Y_c_219_n 4.37331e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_c_147_n N_Y_c_213_n 0.0109821f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_c_147_n N_VGND_c_288_n 0.00434272f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A_c_147_n N_VGND_c_289_n 0.0045104f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_132 N_VPWR_M1001_s N_Y_c_215_n 0.0031621f $X=0.395 $Y=1.84 $X2=0 $Y2=0
cc_133 N_VPWR_c_171_n N_Y_c_215_n 0.0213608f $X=0.54 $Y=2.145 $X2=0 $Y2=0
cc_134 N_VPWR_c_171_n N_Y_c_216_n 0.00268187f $X=0.54 $Y=2.145 $X2=0 $Y2=0
cc_135 N_VPWR_c_171_n N_Y_c_217_n 0.0318965f $X=0.54 $Y=2.145 $X2=0 $Y2=0
cc_136 N_VPWR_c_172_n N_Y_c_217_n 0.0229058f $X=1.565 $Y=2.405 $X2=0 $Y2=0
cc_137 N_VPWR_c_177_n N_Y_c_217_n 0.0144623f $X=1.4 $Y=3.33 $X2=0 $Y2=0
cc_138 N_VPWR_c_170_n N_Y_c_217_n 0.0118344f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_139 N_VPWR_c_174_n N_Y_c_218_n 0.0133269f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_140 N_VPWR_c_172_n N_Y_c_219_n 0.0220125f $X=1.565 $Y=2.405 $X2=0 $Y2=0
cc_141 N_VPWR_c_174_n N_Y_c_219_n 0.031934f $X=2.6 $Y=1.985 $X2=0 $Y2=0
cc_142 N_VPWR_c_179_n N_Y_c_219_n 0.014549f $X=2.435 $Y=3.33 $X2=0 $Y2=0
cc_143 N_VPWR_c_170_n N_Y_c_219_n 0.0119743f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_144 N_VPWR_M1002_d N_Y_c_221_n 0.00462564f $X=1.355 $Y=1.84 $X2=0 $Y2=0
cc_145 N_VPWR_c_172_n N_Y_c_221_n 0.0269118f $X=1.565 $Y=2.405 $X2=0 $Y2=0
cc_146 N_Y_c_211_n N_VGND_M1000_s 0.00674372f $X=2.41 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_147 N_Y_c_213_n N_VGND_c_288_n 0.0145323f $X=2.575 $Y=0.515 $X2=0 $Y2=0
cc_148 N_Y_c_211_n N_VGND_c_289_n 0.0536444f $X=2.41 $Y=0.925 $X2=0 $Y2=0
cc_149 N_Y_c_212_n N_VGND_c_289_n 7.38843e-19 $X=0.405 $Y=0.925 $X2=0 $Y2=0
cc_150 N_Y_c_213_n N_VGND_c_289_n 0.0119861f $X=2.575 $Y=0.515 $X2=0 $Y2=0
cc_151 N_Y_c_211_n N_VGND_c_290_n 0.0192102f $X=2.41 $Y=0.925 $X2=0 $Y2=0
cc_152 N_Y_c_212_n N_VGND_c_290_n 0.0114495f $X=0.405 $Y=0.925 $X2=0 $Y2=0
cc_153 N_Y_c_211_n A_181_74# 0.00722635f $X=2.41 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_154 N_Y_c_211_n A_259_74# 0.0147367f $X=2.41 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_155 N_Y_c_211_n A_373_74# 0.00970428f $X=2.41 $Y=0.925 $X2=-0.19 $Y2=-0.245

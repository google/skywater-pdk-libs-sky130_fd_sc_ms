* File: sky130_fd_sc_ms__dfsbp_2.spice
* Created: Fri Aug 28 17:23:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfsbp_2.pex.spice"
.subckt sky130_fd_sc_ms__dfsbp_2  VNB VPB D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_D_M1033_g N_A_27_74#_M1033_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_CLK_M1035_g N_A_225_74#_M1035_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_398_74#_M1019_d N_A_225_74#_M1019_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_595_97#_M1017_d N_A_225_74#_M1017_g N_A_27_74#_M1017_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1036 A_731_97# N_A_398_74#_M1036_g N_A_595_97#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=0.95 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_757_401#_M1025_g A_731_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 A_1001_74# N_A_595_97#_M1032_g N_A_757_401#_M1032_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_SET_B_M1028_g A_1001_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.15326 AS=0.0441 PD=1.13321 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1012 A_1261_74# N_A_595_97#_M1012_g N_VGND_M1028_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.23354 PD=0.88 PS=1.72679 NRD=12.18 NRS=3.744 M=1 R=4.26667
+ SA=75001.1 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_1339_74#_M1022_d N_A_398_74#_M1022_g A_1261_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.139713 AS=0.0768 PD=1.28 PS=0.88 NRD=13.116 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1037 A_1453_118# N_A_225_74#_M1037_g N_A_1339_74#_M1022_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0916868 PD=0.66 PS=0.84 NRD=18.564 NRS=19.992 M=1 R=2.8
+ SA=75001.8 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1023 A_1531_118# N_A_1501_92#_M1023_g A_1453_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_SET_B_M1002_g A_1531_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.260625 AS=0.0504 PD=1.505 PS=0.66 NRD=161.58 NRS=18.564 M=1 R=2.8
+ SA=75002.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_1501_92#_M1003_d N_A_1339_74#_M1003_g N_VGND_M1002_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1533 AS=0.260625 PD=1.57 PS=1.505 NRD=22.848 NRS=161.58 M=1
+ R=2.8 SA=75003.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 N_Q_N_M1013_d N_A_1339_74#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1024 N_Q_N_M1013_d N_A_1339_74#_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_1339_74#_M1007_g N_A_2221_74#_M1007_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1007_d N_A_2221_74#_M1004_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157545 AS=0.1036 PD=1.24406 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_2221_74#_M1016_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1029 N_VPWR_M1029_d N_D_M1029_g N_A_27_74#_M1029_s VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1018 N_VPWR_M1018_d N_CLK_M1018_g N_A_225_74#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1021 N_A_398_74#_M1021_d N_A_225_74#_M1021_g N_VPWR_M1018_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_595_97#_M1001_d N_A_398_74#_M1001_g N_A_27_74#_M1001_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90004.5 A=0.0756 P=1.2 MULT=1
MM1005 A_709_463# N_A_225_74#_M1005_g N_A_595_97#_M1001_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0567 PD=0.66 PS=0.69 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90004 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_A_757_401#_M1009_g A_709_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.1898 AS=0.0504 PD=1.395 PS=0.66 NRD=186.165 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90003.6 A=0.0756 P=1.2 MULT=1
MM1020 N_A_757_401#_M1020_d N_A_595_97#_M1020_g N_VPWR_M1009_d VPB PSHORT L=0.18
+ W=0.42 AD=0.07035 AS=0.1898 PD=0.755 PS=1.395 NRD=0 NRS=186.165 M=1 R=2.33333
+ SA=90002 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_SET_B_M1000_g N_A_757_401#_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.144131 AS=0.07035 PD=1.09732 PS=0.755 NRD=161.816 NRS=28.1316 M=1
+ R=2.33333 SA=90002.5 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1006 A_1261_341# N_A_595_97#_M1006_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.184812 AS=0.343169 PD=1.58 PS=2.61268 NRD=25.5706 NRS=20.6653 M=1
+ R=5.55556 SA=90001.4 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1027 N_A_1339_74#_M1027_d N_A_225_74#_M1027_g A_1261_341# VPB PSHORT L=0.18
+ W=1 AD=0.300704 AS=0.184812 PD=2.29577 PS=1.58 NRD=0 NRS=25.5706 M=1 R=5.55556
+ SA=90001.8 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1010 A_1524_508# N_A_398_74#_M1010_g N_A_1339_74#_M1027_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.126296 PD=0.66 PS=0.964225 NRD=30.4759 NRS=83.2522 M=1
+ R=2.33333 SA=90002.4 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1031 N_VPWR_M1031_d N_A_1501_92#_M1031_g A_1524_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.0504 PD=0.69 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90002.9
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1034 N_A_1339_74#_M1034_d N_SET_B_M1034_g N_VPWR_M1031_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1155 AS=0.0567 PD=1.39 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90003.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1026 N_VPWR_M1026_d N_A_1339_74#_M1026_g N_A_1501_92#_M1026_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0941182 AS=0.2481 PD=0.804545 PS=2.24 NRD=79.2925
+ NRS=251.274 M=1 R=2.33333 SA=90000.3 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1008 N_Q_N_M1008_d N_A_1339_74#_M1008_g N_VPWR_M1026_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.250982 PD=1.39 PS=2.14545 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.4 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1030 N_Q_N_M1008_d N_A_1339_74#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1015 N_VPWR_M1015_d N_A_1339_74#_M1015_g N_A_2221_74#_M1015_s VPB PSHORT
+ L=0.18 W=1 AD=0.18066 AS=0.28 PD=1.38679 PS=2.56 NRD=14.775 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1011 N_Q_M1011_d N_A_2221_74#_M1011_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.20234 PD=1.39 PS=1.55321 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_Q_M1011_d N_A_2221_74#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX38_noxref VNB VPB NWDIODE A=25.1893 P=30.67
c_142 VNB 0 1.55885e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dfsbp_2.pxi.spice"
*
.ends
*
*

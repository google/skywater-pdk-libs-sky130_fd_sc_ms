* NGSPICE file created from sky130_fd_sc_ms__xor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__xor3_1 A B C VGND VNB VPB VPWR X
M1000 a_84_108# A VGND VNB nlowvt w=640000u l=150000u
+  ad=6.252e+11p pd=4.99e+06u as=1.3258e+12p ps=8.35e+06u
M1001 a_1218_396# a_1157_298# a_416_86# VPB pshort w=840000u l=180000u
+  ad=4.83e+11p pd=2.83e+06u as=5.8575e+11p ps=4.8e+06u
M1002 a_84_108# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.354e+11p pd=5.57e+06u as=1.2444e+12p ps=9e+06u
M1003 a_387_392# C a_1218_396# VPB pshort w=840000u l=180000u
+  ad=5.436e+11p pd=4.69e+06u as=0p ps=0u
M1004 X a_1218_396# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 VPWR a_84_108# a_27_134# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.656e+11p ps=4.42e+06u
M1006 a_27_134# a_452_288# a_416_86# VNB nlowvt w=420000u l=150000u
+  ad=4.987e+11p pd=4.17e+06u as=4.475e+11p ps=4.01e+06u
M1007 a_416_86# C a_1218_396# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.392e+11p ps=2.34e+06u
M1008 a_27_134# a_452_288# a_387_392# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_416_86# B a_27_134# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_84_108# a_452_288# a_416_86# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_452_288# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
M1012 a_387_392# B a_84_108# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR C a_1157_298# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.432e+11p ps=2.04e+06u
M1014 a_387_392# B a_27_134# VNB nlowvt w=640000u l=150000u
+  ad=5.1415e+11p pd=4.38e+06u as=0p ps=0u
M1015 a_416_86# B a_84_108# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1218_396# a_1157_298# a_387_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C a_1157_298# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 X a_1218_396# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 VGND a_84_108# a_27_134# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_84_108# a_452_288# a_387_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B a_452_288# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
.ends


* NGSPICE file created from sky130_fd_sc_ms__o2bb2a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR B1 a_41_392# VPB pshort w=1e+06u l=180000u
+  ad=2.2314e+12p pd=1.735e+07u as=8.3e+11p ps=7.66e+06u
M1001 a_41_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_476_48# A2_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1003 VPWR a_313_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.224e+11p ps=5.77e+06u
M1004 X a_313_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=1.3531e+12p ps=1.093e+07u
M1005 a_27_74# a_476_48# a_313_392# VNB nlowvt w=640000u l=150000u
+  ad=7.648e+11p pd=7.51e+06u as=2.016e+11p ps=1.91e+06u
M1006 a_313_392# B2 a_41_392# VPB pshort w=1e+06u l=180000u
+  ad=5.556e+11p pd=4.9e+06u as=0p ps=0u
M1007 VPWR A1_N a_476_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_313_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_41_392# B2 a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_476_48# a_313_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_313_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_313_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_313_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_313_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B2 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A1_N a_835_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1018 VGND a_313_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_313_392# a_476_48# a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_835_94# A2_N a_476_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.952e+11p ps=1.89e+06u
M1021 a_313_392# a_476_48# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B1 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_74# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* NGSPICE file created from sky130_fd_sc_ms__nand4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.239e+12p ps=8.97e+06u
M1001 VPWR a_27_112# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_443_74# B a_341_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=2.664e+11p ps=2.2e+06u
M1003 Y a_27_112# a_443_74# VNB nlowvt w=740000u l=150000u
+  ad=3.404e+11p pd=2.4e+06u as=0p ps=0u
M1004 VPWR A_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1005 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=2.696e+11p pd=2.26e+06u as=2.695e+11p ps=2.08e+06u
M1007 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_263_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_341_74# C a_263_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__nand4b_2.pex.spice
* Created: Fri Aug 28 17:45:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4B_2%A_N 3 7 9 10 17 18
c32 17 0 1.48501e-19 $X=0.82 $Y=1.345
r33 16 18 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.82 $Y=1.345
+ $X2=0.895 $Y2=1.345
r34 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.82
+ $Y=1.345 $X2=0.82 $Y2=1.345
r35 13 16 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.82 $Y2=1.345
r36 10 17 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.72 $Y=1.345 $X2=0.82
+ $Y2=1.345
r37 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.72 $Y2=1.345
r38 5 18 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.51
+ $X2=0.895 $Y2=1.345
r39 5 7 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=0.895 $Y=1.51
+ $X2=0.895 $Y2=2.34
r40 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=1.345
r41 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%A_27_74# 1 2 9 13 17 21 25 27 28 31 35 36
+ 38 40 48
c85 48 0 1.48501e-19 $X=1.945 $Y=1.515
c86 21 0 9.65687e-20 $X=1.945 $Y=0.74
c87 13 0 4.22696e-20 $X=1.485 $Y=0.74
r88 47 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.885 $Y=1.515
+ $X2=1.945 $Y2=1.515
r89 43 45 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.435 $Y=1.515
+ $X2=1.485 $Y2=1.515
r90 41 47 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.555 $Y=1.515
+ $X2=1.885 $Y2=1.515
r91 41 45 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.555 $Y=1.515
+ $X2=1.485 $Y2=1.515
r92 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.555
+ $Y=1.515 $X2=1.555 $Y2=1.515
r93 38 40 9.29987 $w=4.3e-07 $l=2.67047e-07 $layer=LI1_cond $X=1.24 $Y=1.35
+ $X2=1.437 $Y2=1.515
r94 37 38 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.24 $Y=1.01
+ $X2=1.24 $Y2=1.35
r95 35 40 7.09302 $w=4.3e-07 $l=3.87329e-07 $layer=LI1_cond $X=1.155 $Y=1.765
+ $X2=1.437 $Y2=1.515
r96 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.155 $Y=1.765
+ $X2=0.835 $Y2=1.765
r97 31 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.67 $Y=1.985
+ $X2=0.67 $Y2=2.695
r98 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.67 $Y=1.85
+ $X2=0.835 $Y2=1.765
r99 29 31 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.67 $Y=1.85
+ $X2=0.67 $Y2=1.985
r100 27 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=1.24 $Y2=1.01
r101 27 28 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=0.365 $Y2=0.925
r102 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.365 $Y2=0.925
r103 23 25 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.24 $Y2=0.68
r104 19 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.35
+ $X2=1.945 $Y2=1.515
r105 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.945 $Y=1.35
+ $X2=1.945 $Y2=0.74
r106 15 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.68
+ $X2=1.885 $Y2=1.515
r107 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.885 $Y=1.68
+ $X2=1.885 $Y2=2.4
r108 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.35
+ $X2=1.485 $Y2=1.515
r109 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.485 $Y=1.35
+ $X2=1.485 $Y2=0.74
r110 7 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.68
+ $X2=1.435 $Y2=1.515
r111 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.435 $Y=1.68
+ $X2=1.435 $Y2=2.4
r112 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.84 $X2=0.67 $Y2=2.695
r113 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.84 $X2=0.67 $Y2=1.985
r114 1 25 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%B 3 7 11 15 17 23 26
c60 3 0 3.91537e-20 $X=2.375 $Y=0.74
r61 25 26 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.965 $Y=1.515
+ $X2=3.15 $Y2=1.515
r62 24 25 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.965 $Y2=1.515
r63 22 24 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.425 $Y=1.515
+ $X2=2.7 $Y2=1.515
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.425
+ $Y=1.515 $X2=2.425 $Y2=1.515
r65 19 22 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.375 $Y=1.515
+ $X2=2.425 $Y2=1.515
r66 17 23 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.425 $Y2=1.565
r67 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.68
+ $X2=3.15 $Y2=1.515
r68 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.15 $Y=1.68
+ $X2=3.15 $Y2=2.4
r69 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.35
+ $X2=2.965 $Y2=1.515
r70 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.965 $Y=1.35
+ $X2=2.965 $Y2=0.74
r71 5 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.68 $X2=2.7
+ $Y2=1.515
r72 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.7 $Y=1.68 $X2=2.7
+ $Y2=2.4
r73 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.35
+ $X2=2.375 $Y2=1.515
r74 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.375 $Y=1.35
+ $X2=2.375 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%C 3 7 11 15 17 18 26
c57 3 0 1.0617e-19 $X=3.7 $Y=2.4
r58 24 26 20.1533 $w=2.87e-07 $l=1.2e-07 $layer=POLY_cond $X=4.03 $Y=1.515
+ $X2=4.15 $Y2=1.515
r59 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.03
+ $Y=1.515 $X2=4.03 $Y2=1.515
r60 22 24 12.5958 $w=2.87e-07 $l=7.5e-08 $layer=POLY_cond $X=3.955 $Y=1.515
+ $X2=4.03 $Y2=1.515
r61 21 22 42.8258 $w=2.87e-07 $l=2.55e-07 $layer=POLY_cond $X=3.7 $Y=1.515
+ $X2=3.955 $Y2=1.515
r62 18 25 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.03
+ $Y2=1.565
r63 17 25 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.03 $Y2=1.565
r64 13 26 39.4669 $w=2.87e-07 $l=3.06594e-07 $layer=POLY_cond $X=4.385 $Y=1.35
+ $X2=4.15 $Y2=1.515
r65 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.385 $Y=1.35
+ $X2=4.385 $Y2=0.79
r66 9 26 13.6964 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.15 $Y=1.68
+ $X2=4.15 $Y2=1.515
r67 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.15 $Y=1.68 $X2=4.15
+ $Y2=2.4
r68 5 22 17.9292 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.955 $Y=1.35
+ $X2=3.955 $Y2=1.515
r69 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.955 $Y=1.35
+ $X2=3.955 $Y2=0.79
r70 1 21 13.6964 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.7 $Y=1.68 $X2=3.7
+ $Y2=1.515
r71 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.7 $Y=1.68 $X2=3.7
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%D 1 3 6 8 10 14 16 17 18
r46 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.905
+ $Y=1.515 $X2=4.905 $Y2=1.515
r47 23 25 12.7588 $w=3.4e-07 $l=9e-08 $layer=POLY_cond $X=4.815 $Y=1.56
+ $X2=4.905 $Y2=1.56
r48 22 23 2.12647 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=4.8 $Y=1.56
+ $X2=4.815 $Y2=1.56
r49 17 18 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r50 17 26 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.905 $Y2=1.565
r51 16 26 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.905 $Y2=1.565
r52 12 28 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=1.56
r53 12 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=0.79
r54 8 28 2.12647 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=5.25 $Y=1.56
+ $X2=5.265 $Y2=1.56
r55 8 25 48.9088 $w=3.4e-07 $l=3.45e-07 $layer=POLY_cond $X=5.25 $Y=1.56
+ $X2=4.905 $Y2=1.56
r56 8 10 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.25 $Y=1.68 $X2=5.25
+ $Y2=2.4
r57 4 23 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.815 $Y=1.35
+ $X2=4.815 $Y2=1.56
r58 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.815 $Y=1.35
+ $X2=4.815 $Y2=0.79
r59 1 22 17.6285 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.8 $Y=1.77 $X2=4.8
+ $Y2=1.56
r60 1 3 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=4.8 $Y=1.77 $X2=4.8
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%VPWR 1 2 3 4 5 18 24 28 32 34 36 41 42 43
+ 45 50 59 63 69 72 75 79
r75 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r76 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 67 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 67 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 64 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=4.485 $Y2=3.33
r83 64 66 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 63 78 4.31409 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=5.36 $Y=3.33 $X2=5.56
+ $Y2=3.33
r85 63 66 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=3.33 $X2=5.04
+ $Y2=3.33
r86 62 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 59 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.485 $Y2=3.33
r89 59 61 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 58 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 55 72 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=2.292 $Y2=3.33
r93 55 57 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r96 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r97 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.205 $Y2=3.33
r98 51 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 50 72 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.292 $Y2=3.33
r100 50 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=1.205 $Y2=3.33
r104 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 43 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 43 73 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r107 41 57 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.425 $Y2=3.33
r109 40 61 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=3.425 $Y2=3.33
r111 36 39 28.3056 $w=2.83e-07 $l=7e-07 $layer=LI1_cond $X=5.502 $Y=2.115
+ $X2=5.502 $Y2=2.815
r112 34 78 3.08458 $w=2.85e-07 $l=1.1025e-07 $layer=LI1_cond $X=5.502 $Y=3.245
+ $X2=5.56 $Y2=3.33
r113 34 39 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=5.502 $Y=3.245
+ $X2=5.502 $Y2=2.815
r114 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=3.33
r115 30 32 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=2.41
r116 26 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=3.33
r117 26 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=2.415
r118 22 72 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.292 $Y=3.245
+ $X2=2.292 $Y2=3.33
r119 22 24 15.8807 $w=5.93e-07 $l=7.9e-07 $layer=LI1_cond $X=2.292 $Y=3.245
+ $X2=2.292 $Y2=2.455
r120 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.205 $Y=2.105
+ $X2=1.205 $Y2=2.785
r121 16 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=3.33
r122 16 21 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=2.785
r123 5 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.84 $X2=5.475 $Y2=2.815
r124 5 36 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.84 $X2=5.475 $Y2=2.115
r125 4 32 300 $w=1.7e-07 $l=6.81579e-07 $layer=licon1_PDIFF $count=2 $X=4.24
+ $Y=1.84 $X2=4.485 $Y2=2.41
r126 3 28 300 $w=1.7e-07 $l=6.6106e-07 $layer=licon1_PDIFF $count=2 $X=3.24
+ $Y=1.84 $X2=3.425 $Y2=2.415
r127 2 24 150 $w=1.7e-07 $l=8.28085e-07 $layer=licon1_PDIFF $count=4 $X=1.975
+ $Y=1.84 $X2=2.475 $Y2=2.455
r128 1 21 600 $w=1.7e-07 $l=1.04925e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.84 $X2=1.205 $Y2=2.785
r129 1 18 300 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.84 $X2=1.205 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%Y 1 2 3 4 5 16 18 20 22 26 28 32 34 36 38
+ 41 49 55 58 59
c102 49 0 1.0617e-19 $X=2.925 $Y=1.985
c103 22 0 4.22696e-20 $X=3.005 $Y=1.095
r104 58 59 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.665
r105 53 58 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.18
+ $X2=3.12 $Y2=1.295
r106 50 59 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.12 $Y=1.82
+ $X2=3.12 $Y2=1.665
r107 49 50 7.34574 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.997 $Y=1.985
+ $X2=2.997 $Y2=1.82
r108 41 43 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=1.715 $Y=0.965
+ $X2=1.715 $Y2=1.095
r109 36 57 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=2.12
+ $X2=5.025 $Y2=2.035
r110 36 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.025 $Y=2.12
+ $X2=5.025 $Y2=2.815
r111 35 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=3.925 $Y2=2.035
r112 34 57 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=5.025 $Y2=2.035
r113 34 35 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.09 $Y2=2.035
r114 30 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=2.035
r115 30 32 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=2.815
r116 28 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=2.035
+ $X2=3.925 $Y2=2.035
r117 28 29 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.76 $Y=2.035
+ $X2=3.235 $Y2=2.035
r118 26 52 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.925 $Y=2.815
+ $X2=2.925 $Y2=2.12
r119 23 43 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.895 $Y=1.095
+ $X2=1.715 $Y2=1.095
r120 22 53 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=3.12 $Y2=1.18
r121 22 23 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=1.895 $Y2=1.095
r122 21 46 4.26175 $w=1.7e-07 $l=1.61071e-07 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.687 $Y2=1.985
r123 20 52 3.26684 $w=4.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.997 $Y=2.035
+ $X2=2.997 $Y2=2.12
r124 20 29 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=2.997 $Y=2.035
+ $X2=3.235 $Y2=2.035
r125 20 49 1.25903 $w=4.73e-07 $l=5e-08 $layer=LI1_cond $X=2.997 $Y=2.035
+ $X2=2.997 $Y2=1.985
r126 20 21 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.76 $Y=2.035 $X2=1.825
+ $Y2=2.035
r127 16 46 3.0603 $w=2.75e-07 $l=1.35e-07 $layer=LI1_cond $X=1.687 $Y=2.12
+ $X2=1.687 $Y2=1.985
r128 16 18 29.1254 $w=2.73e-07 $l=6.95e-07 $layer=LI1_cond $X=1.687 $Y=2.12
+ $X2=1.687 $Y2=2.815
r129 5 57 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.025 $Y2=2.035
r130 5 38 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.84 $X2=5.025 $Y2=2.815
r131 4 55 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.79
+ $Y=1.84 $X2=3.925 $Y2=2.035
r132 4 32 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.79
+ $Y=1.84 $X2=3.925 $Y2=2.815
r133 3 49 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.84 $X2=2.925 $Y2=1.985
r134 3 26 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.84 $X2=2.925 $Y2=2.815
r135 2 46 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.66 $Y2=2.015
r136 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.84 $X2=1.66 $Y2=2.815
r137 1 41 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.715 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r56 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r57 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r59 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r60 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.03
+ $Y2=0
r61 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.52
+ $Y2=0
r62 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r63 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r64 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r65 25 28 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r66 25 26 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r67 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r68 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r69 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=0 $X2=5.03
+ $Y2=0
r70 22 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.865 $Y=0 $X2=4.56
+ $Y2=0
r71 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r72 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r74 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r75 15 29 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r76 15 26 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r77 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r78 11 13 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.58
r79 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r80 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.55
r81 2 13 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.42 $X2=5.03 $Y2=0.58
r82 1 9 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.57 $Y=0.37
+ $X2=0.71 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%A_225_74# 1 2 3 10 16 23 24
c37 16 0 9.65687e-20 $X=2.2 $Y=0.49
c38 10 0 3.91537e-20 $X=2.075 $Y=0.49
r39 23 24 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0.717
+ $X2=3.015 $Y2=0.717
r40 19 20 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.2 $Y=0.595 $X2=2.2
+ $Y2=0.755
r41 16 19 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.2 $Y=0.49 $X2=2.2
+ $Y2=0.595
r42 15 20 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=0.755
+ $X2=2.2 $Y2=0.755
r43 15 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.325 $Y=0.755
+ $X2=3.015 $Y2=0.755
r44 10 16 0.0129374 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.49
+ $X2=2.2 $Y2=0.49
r45 10 12 33.1327 $w=2.78e-07 $l=8.05e-07 $layer=LI1_cond $X=2.075 $Y=0.49
+ $X2=1.27 $Y2=0.49
r46 3 23 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.37 $X2=3.18 $Y2=0.715
r47 2 19 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.37 $X2=2.16 $Y2=0.595
r48 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%A_490_74# 1 2 7 11 16
r27 14 16 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0.377
+ $X2=2.835 $Y2=0.377
r28 9 11 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.17 $Y=0.425
+ $X2=4.17 $Y2=0.58
r29 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.005 $Y=0.34
+ $X2=4.17 $Y2=0.425
r30 7 16 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.005 $Y=0.34
+ $X2=2.835 $Y2=0.34
r31 2 11 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.42 $X2=4.17 $Y2=0.58
r32 1 14 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.37 $X2=2.67 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_2%A_719_123# 1 2 3 10 13 14 17 19 21 23 26
r42 21 28 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=0.93
+ $X2=5.52 $Y2=1.055
r43 21 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=5.52 $Y=0.93
+ $X2=5.52 $Y2=0.565
r44 20 26 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.695 $Y=1.055
+ $X2=4.6 $Y2=1.055
r45 19 28 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.395 $Y=1.055
+ $X2=5.52 $Y2=1.055
r46 19 20 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.395 $Y=1.055
+ $X2=4.695 $Y2=1.055
r47 15 26 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.6 $Y=0.93 $X2=4.6
+ $Y2=1.055
r48 15 17 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=4.6 $Y=0.93 $X2=4.6
+ $Y2=0.565
r49 13 26 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.505 $Y=1.055
+ $X2=4.6 $Y2=1.055
r50 13 14 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.505 $Y=1.055
+ $X2=3.825 $Y2=1.055
r51 10 14 6.81649 $w=2.5e-07 $l=1.76777e-07 $layer=LI1_cond $X=3.7 $Y=0.93
+ $X2=3.825 $Y2=1.055
r52 10 12 2.196 $w=2.5e-07 $l=4.5e-08 $layer=LI1_cond $X=3.7 $Y=0.93 $X2=3.7
+ $Y2=0.885
r53 3 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.42 $X2=5.48 $Y2=1.015
r54 3 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.42 $X2=5.48 $Y2=0.565
r55 2 26 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.42 $X2=4.6 $Y2=1.015
r56 2 17 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.42 $X2=4.6 $Y2=0.565
r57 1 12 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.615 $X2=3.74 $Y2=0.885
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o31ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.715000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.835000 1.350000 6.115000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.847200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 7.790000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.702400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.550000 4.665000 1.950000 ;
        RECT 3.965000 1.950000 8.525000 2.120000 ;
        RECT 3.965000 2.120000 4.970000 2.150000 ;
        RECT 4.495000 1.010000 8.095000 1.180000 ;
        RECT 4.495000 1.180000 4.665000 1.550000 ;
        RECT 4.700000 2.150000 4.970000 2.735000 ;
        RECT 5.600000 2.120000 5.930000 2.735000 ;
        RECT 6.550000 2.120000 6.880000 2.980000 ;
        RECT 6.905000 0.920000 8.095000 1.010000 ;
        RECT 8.195000 1.820000 8.525000 1.950000 ;
        RECT 8.195000 2.120000 8.525000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.390000 0.445000 0.920000 ;
      RECT 0.115000  0.920000 2.305000 1.010000 ;
      RECT 0.115000  1.010000 4.325000 1.180000 ;
      RECT 0.120000  1.950000 3.300000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.570000  2.290000 0.900000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.750000 ;
      RECT 1.100000  2.120000 1.270000 2.980000 ;
      RECT 1.470000  2.290000 1.800000 3.245000 ;
      RECT 1.475000  0.085000 1.805000 0.750000 ;
      RECT 1.970000  1.820000 2.300000 1.950000 ;
      RECT 1.970000  2.120000 2.300000 2.980000 ;
      RECT 1.975000  0.390000 2.305000 0.920000 ;
      RECT 2.470000  2.290000 2.800000 2.905000 ;
      RECT 2.470000  2.905000 6.380000 3.075000 ;
      RECT 2.495000  0.085000 2.960000 0.805000 ;
      RECT 2.970000  2.120000 3.300000 2.370000 ;
      RECT 2.970000  2.370000 4.470000 2.540000 ;
      RECT 2.970000  2.540000 3.300000 2.735000 ;
      RECT 3.145000  0.390000 3.475000 1.010000 ;
      RECT 3.640000  2.710000 3.970000 2.905000 ;
      RECT 3.645000  0.085000 3.975000 0.840000 ;
      RECT 4.140000  2.540000 4.470000 2.735000 ;
      RECT 4.155000  0.390000 4.325000 0.670000 ;
      RECT 4.155000  0.670000 6.805000 0.750000 ;
      RECT 4.155000  0.750000 5.775000 0.840000 ;
      RECT 4.155000  0.840000 4.325000 1.010000 ;
      RECT 4.585000  0.085000 5.265000 0.500000 ;
      RECT 5.150000  2.290000 5.400000 2.905000 ;
      RECT 5.445000  0.390000 5.775000 0.580000 ;
      RECT 5.445000  0.580000 6.805000 0.670000 ;
      RECT 5.955000  0.085000 6.295000 0.410000 ;
      RECT 6.130000  2.290000 6.380000 2.905000 ;
      RECT 6.475000  0.390000 8.525000 0.560000 ;
      RECT 6.475000  0.560000 6.805000 0.580000 ;
      RECT 7.050000  2.290000 8.025000 3.245000 ;
      RECT 7.335000  0.560000 7.665000 0.750000 ;
      RECT 8.265000  0.560000 8.525000 1.170000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ms__o31ai_4
END LIBRARY

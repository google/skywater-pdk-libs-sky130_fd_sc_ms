* File: sky130_fd_sc_ms__and2_2.spice
* Created: Fri Aug 28 17:10:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and2_2.pex.spice"
.subckt sky130_fd_sc_ms__and2_2  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 A_118_74# N_A_M1006_g N_A_31_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g A_118_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1332
+ AS=0.0888 PD=1.1 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_A_31_74#_M1005_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1332 PD=1.02 PS=1.1 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1005_d N_A_31_74#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2553 PD=1.02 PS=2.17 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75001.5
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1002 N_A_31_74#_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.275 PD=1.27 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_31_74#_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.167453 AS=0.135 PD=1.36321 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_X_M1001_d N_A_31_74#_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.187547 PD=1.39 PS=1.52679 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1004 N_X_M1001_d N_A_31_74#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__and2_2.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__o31ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.296e+11p ps=8.38e+06u
M1001 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_300_368# A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1003 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=1.2616e+12p pd=7.93e+06u as=1.0582e+12p ps=1.026e+07u
M1004 a_28_368# A2 a_300_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=0p ps=0u
M1008 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_300_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=9.856e+11p ps=8.48e+06u
M1010 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A3 a_300_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* NGSPICE file created from sky130_fd_sc_ms__o41a_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_27_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=6.364e+11p pd=6.16e+06u as=1.2691e+12p ps=9.35e+06u
M1001 X a_431_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1002 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=1.6872e+12p ps=9.9e+06u
M1003 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR B1 a_431_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.236e+11p ps=3.02e+06u
M1005 a_203_368# A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1006 a_431_368# A4 a_317_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=4.368e+11p ps=3.02e+06u
M1007 VGND a_431_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_317_368# A3 a_203_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_431_368# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1010 X a_431_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_431_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


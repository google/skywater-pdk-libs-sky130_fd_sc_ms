* NGSPICE file created from sky130_fd_sc_ms__sdfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1529_74# a_612_74# a_1243_398# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=6.216e+11p ps=3.16e+06u
M1001 a_1723_48# a_1529_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=1.8401e+12p ps=1.538e+07u
M1002 VPWR a_1723_48# a_1694_508# VPB pshort w=420000u l=180000u
+  ad=2.5456e+12p pd=2.012e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_434_74# SCE a_296_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.423e+11p ps=3.31e+06u
M1004 VPWR a_1723_48# a_2216_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1005 Q a_1723_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1006 a_1157_100# a_828_74# a_1021_100# VNB nlowvt w=420000u l=150000u
+  ad=1.932e+11p pd=1.76e+06u as=2.226e+11p ps=1.9e+06u
M1007 a_218_74# a_31_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1008 a_296_74# D a_218_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR SCD a_410_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1010 a_1529_74# a_828_74# a_1243_398# VNB nlowvt w=550000u l=150000u
+  ad=2.887e+11p pd=2.32e+06u as=1.5675e+11p ps=1.67e+06u
M1011 a_1243_398# a_1021_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q a_1723_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 a_612_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1014 a_1723_48# a_1529_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1015 a_828_74# a_612_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1016 VGND a_1243_398# a_1157_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1681_74# a_612_74# a_1529_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1018 a_236_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 a_1243_398# a_1021_100# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1694_508# a_828_74# a_1529_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1723_48# a_1681_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR SCE a_31_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1023 a_612_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 VGND SCE a_31_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1025 a_828_74# a_612_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1026 Q_N a_2216_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1027 VGND SCD a_434_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_296_74# D a_236_464# VPB pshort w=640000u l=180000u
+  ad=2.841e+11p pd=3.19e+06u as=0p ps=0u
M1029 a_1021_100# a_828_74# a_296_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1030 a_1021_100# a_612_74# a_296_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR a_1243_398# a_1183_496# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1032 a_410_464# a_31_74# a_296_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1183_496# a_612_74# a_1021_100# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q_N a_2216_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1035 VGND a_1723_48# a_2216_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__edfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__edfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.316800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.110000 1.845000 1.440000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.502100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.015000 0.350000 12.345000 1.130000 ;
        RECT 12.075000 1.130000 12.345000 1.550000 ;
        RECT 12.075000 1.550000 12.405000 2.980000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.180000 3.780000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.960000 0.085000 ;
        RECT  1.020000  0.085000  1.350000 0.600000 ;
        RECT  2.000000  0.085000  2.330000 0.875000 ;
        RECT  3.440000  0.085000  3.610000 1.010000 ;
        RECT  4.335000  0.085000  4.585000 1.130000 ;
        RECT  7.170000  0.085000  7.420000 0.765000 ;
        RECT  8.610000  0.085000  8.860000 0.765000 ;
        RECT 10.350000  0.085000 11.310000 0.665000 ;
        RECT 12.515000  0.085000 12.845000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.960000 3.415000 ;
        RECT  0.945000 2.520000  1.195000 3.245000 ;
        RECT  2.385000 2.290000  2.635000 3.245000 ;
        RECT  3.670000 2.650000  4.000000 3.245000 ;
        RECT  5.020000 2.650000  5.270000 3.245000 ;
        RECT  7.410000 2.750000  7.740000 3.245000 ;
        RECT  8.505000 2.750000  8.835000 3.245000 ;
        RECT 10.845000 2.525000 11.385000 3.245000 ;
        RECT 12.605000 1.820000 12.855000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.340000  0.530000 0.810000 ;
      RECT  0.085000 0.810000  0.255000 2.180000 ;
      RECT  0.085000 2.180000  1.535000 2.350000 ;
      RECT  0.085000 2.350000  0.435000 2.980000 ;
      RECT  0.975000 0.770000  1.820000 0.940000 ;
      RECT  0.975000 0.940000  1.305000 1.610000 ;
      RECT  0.975000 1.610000  2.385000 1.780000 ;
      RECT  0.975000 1.780000  1.305000 2.010000 ;
      RECT  1.365000 2.350000  1.535000 2.905000 ;
      RECT  1.365000 2.905000  2.215000 3.075000 ;
      RECT  1.570000 0.415000  1.820000 0.770000 ;
      RECT  1.705000 1.780000  1.875000 2.735000 ;
      RECT  2.045000 1.950000  3.270000 2.120000 ;
      RECT  2.045000 2.120000  2.215000 2.905000 ;
      RECT  2.055000 1.385000  2.385000 1.610000 ;
      RECT  2.555000 1.045000  2.930000 1.780000 ;
      RECT  2.790000 0.415000  3.270000 0.875000 ;
      RECT  3.100000 0.875000  3.270000 1.950000 ;
      RECT  3.100000 2.120000  3.475000 2.310000 ;
      RECT  3.100000 2.310000  5.610000 2.480000 ;
      RECT  3.100000 2.480000  3.475000 2.620000 ;
      RECT  3.790000 0.350000  4.120000 1.010000 ;
      RECT  3.950000 1.010000  4.120000 1.470000 ;
      RECT  3.950000 1.470000  4.900000 2.140000 ;
      RECT  4.765000 0.255000  6.960000 0.425000 ;
      RECT  4.765000 0.425000  5.095000 1.130000 ;
      RECT  5.130000 1.480000  5.655000 1.650000 ;
      RECT  5.130000 1.650000  5.300000 2.310000 ;
      RECT  5.325000 0.595000  5.655000 1.480000 ;
      RECT  5.440000 2.480000  5.610000 2.520000 ;
      RECT  5.440000 2.520000  6.245000 2.690000 ;
      RECT  5.470000 1.820000  5.995000 1.970000 ;
      RECT  5.470000 1.970000  6.245000 2.140000 ;
      RECT  5.825000 0.425000  5.995000 1.820000 ;
      RECT  5.825000 2.140000  6.245000 2.300000 ;
      RECT  5.995000 2.690000  6.245000 2.980000 ;
      RECT  6.165000 0.595000  6.620000 0.765000 ;
      RECT  6.165000 0.765000  6.335000 1.630000 ;
      RECT  6.165000 1.630000  8.030000 1.800000 ;
      RECT  6.415000 1.800000  6.585000 2.520000 ;
      RECT  6.415000 2.520000  6.775000 2.980000 ;
      RECT  6.505000 0.935000  7.760000 1.105000 ;
      RECT  6.505000 1.105000  6.960000 1.310000 ;
      RECT  6.755000 2.000000  7.115000 2.330000 ;
      RECT  6.790000 0.425000  6.960000 0.935000 ;
      RECT  6.945000 2.330000  7.115000 2.410000 ;
      RECT  6.945000 2.410000  9.800000 2.580000 ;
      RECT  7.130000 1.275000  8.940000 1.445000 ;
      RECT  7.130000 1.445000  7.460000 1.460000 ;
      RECT  7.590000 0.255000  8.440000 0.425000 ;
      RECT  7.590000 0.425000  7.760000 0.935000 ;
      RECT  7.700000 1.615000  8.030000 1.630000 ;
      RECT  7.700000 1.800000  8.030000 1.830000 ;
      RECT  7.930000 0.595000  8.100000 1.275000 ;
      RECT  7.945000 2.070000  8.440000 2.240000 ;
      RECT  8.270000 0.425000  8.440000 0.935000 ;
      RECT  8.270000 0.935000  9.280000 1.105000 ;
      RECT  8.270000 1.445000  8.940000 1.605000 ;
      RECT  8.270000 1.605000  8.440000 2.070000 ;
      RECT  9.110000 1.105000  9.280000 1.205000 ;
      RECT  9.110000 1.205000 10.605000 1.375000 ;
      RECT  9.110000 1.375000  9.460000 1.550000 ;
      RECT  9.450000 0.350000  9.780000 0.835000 ;
      RECT  9.450000 0.835000 10.945000 1.005000 ;
      RECT  9.630000 1.545000 10.065000 1.725000 ;
      RECT  9.630000 1.725000  9.800000 2.410000 ;
      RECT  9.970000 1.925000 10.405000 2.095000 ;
      RECT  9.970000 2.095000 10.220000 3.000000 ;
      RECT 10.235000 1.755000 10.945000 1.925000 ;
      RECT 10.275000 1.375000 10.605000 1.585000 ;
      RECT 10.665000 2.095000 11.885000 2.320000 ;
      RECT 10.775000 1.005000 11.505000 1.335000 ;
      RECT 10.775000 1.335000 10.945000 1.755000 ;
      RECT 11.490000 0.335000 11.845000 0.810000 ;
      RECT 11.555000 2.320000 11.885000 2.950000 ;
      RECT 11.645000 1.550000 11.885000 2.095000 ;
      RECT 11.675000 0.810000 11.845000 1.550000 ;
    LAYER mcon ;
      RECT  2.555000 1.580000  2.725000 1.750000 ;
      RECT 11.675000 1.580000 11.845000 1.750000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 11.905000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 11.615000 1.550000 11.905000 1.595000 ;
      RECT 11.615000 1.735000 11.905000 1.780000 ;
  END
END sky130_fd_sc_ms__edfxtp_1

* File: sky130_fd_sc_ms__o2bb2a_2.spice
* Created: Fri Aug 28 17:59:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2bb2a_2.pex.spice"
.subckt sky130_fd_sc_ms__o2bb2a_2  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_B1_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_B2_M1010_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1005 N_A_204_392#_M1005_d N_A_270_48#_M1005_g N_A_27_74#_M1010_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 A_500_74# N_A2_N_M1003_g N_A_270_48#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A1_N_M1007_g A_500_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.134771 AS=0.0768 PD=1.0713 PS=0.88 NRD=3.744 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_X_M1001_d N_A_204_392#_M1001_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.155829 PD=1.02 PS=1.2387 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75001 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1001_d N_A_204_392#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 A_120_392# N_B1_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90003.1
+ A=0.18 P=2.36 MULT=1
MM1011 N_A_204_392#_M1011_d N_B2_M1011_g A_120_392# VPB PSHORT L=0.18 W=1
+ AD=0.165 AS=0.12 PD=1.33 PS=1.24 NRD=10.8153 NRS=12.7853 M=1 R=5.55556
+ SA=90000.6 SB=90002.7 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_270_48#_M1004_g N_A_204_392#_M1011_d VPB PSHORT L=0.18
+ W=1 AD=0.260367 AS=0.165 PD=1.68478 PS=1.33 NRD=18.6953 NRS=0 M=1 R=5.55556
+ SA=90001.1 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_270_48#_M1000_d N_A2_N_M1000_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1512 AS=0.218708 PD=1.2 PS=1.41522 NRD=9.3772 NRS=48.1468 M=1
+ R=4.66667 SA=90001.8 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1002 N_VPWR_M1002_d N_A1_N_M1002_g N_A_270_48#_M1000_d VPB PSHORT L=0.18
+ W=0.84 AD=0.262146 AS=0.1512 PD=1.51286 PS=1.2 NRD=60.282 NRS=9.3772 M=1
+ R=4.66667 SA=90002.3 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1008 N_X_M1008_d N_A_204_392#_M1008_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.349529 PD=1.39 PS=2.01714 NRD=0 NRS=25.4918 M=1 R=6.22222
+ SA=90002.4 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1008_d N_A_204_392#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__o2bb2a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand2_1.spice
* Created: Fri Aug 28 17:41:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand2_1.pex.spice"
.subckt sky130_fd_sc_ms__nand2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 A_117_74# N_B_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g A_117_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1001_d VPB PSHORT L=0.18 W=1.12 AD=0.3024
+ AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_ms__nand2_1.pxi.spice"
*
.ends
*
*

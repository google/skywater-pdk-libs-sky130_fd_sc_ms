* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__einvn_8 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR TE_B a_126_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VGND TE_B a_126_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

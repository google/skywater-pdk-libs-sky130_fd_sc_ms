* File: sky130_fd_sc_ms__a2bb2oi_1.pex.spice
* Created: Fri Aug 28 17:04:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%A1_N 3 7 9 13 14
r27 14 15 6.79937 $w=3.19e-07 $l=4.5e-08 $layer=POLY_cond $X=0.51 $Y=1.425
+ $X2=0.555 $Y2=1.425
r28 12 14 36.2633 $w=3.19e-07 $l=2.4e-07 $layer=POLY_cond $X=0.27 $Y=1.425
+ $X2=0.51 $Y2=1.425
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.425 $X2=0.27 $Y2=1.425
r30 9 13 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.425
r31 5 15 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.26
+ $X2=0.555 $Y2=1.425
r32 5 7 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.555 $Y=1.26
+ $X2=0.555 $Y2=0.835
r33 1 14 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.59 $X2=0.51
+ $Y2=1.425
r34 1 3 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=0.51 $Y=1.59 $X2=0.51
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%A2_N 1 3 7 9 13
c42 13 0 8.79615e-20 $X=1.005 $Y=1.615
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.005
+ $Y=1.615 $X2=1.005 $Y2=1.615
r44 9 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=1.005 $Y2=1.615
r45 5 12 38.832 $w=3.54e-07 $l=1.67481e-07 $layer=POLY_cond $X=0.985 $Y=1.45
+ $X2=0.99 $Y2=1.615
r46 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.985 $Y=1.45
+ $X2=0.985 $Y2=0.835
r47 1 12 40.8926 $w=3.54e-07 $l=2.56076e-07 $layer=POLY_cond $X=0.9 $Y=1.83
+ $X2=0.99 $Y2=1.615
r48 1 3 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.9 $Y=1.83 $X2=0.9
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%A_126_112# 1 2 9 11 13 14 15 18 20 21 24
+ 26 29 30
c74 15 0 8.02067e-21 $X=1.92 $Y=1.385
c75 14 0 8.79615e-20 $X=1.83 $Y=1.385
c76 11 0 1.45091e-19 $X=1.935 $Y=1.22
c77 9 0 1.19783e-19 $X=1.92 $Y=2.4
r78 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.545
+ $Y=1.385 $X2=1.545 $Y2=1.385
r79 29 31 1.30231 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=2.115 $X2=1.2
+ $Y2=2.12
r80 29 30 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=2.115
+ $X2=1.2 $Y2=1.95
r81 26 34 8.95599 $w=3.21e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.355 $Y=1.55
+ $X2=1.49 $Y2=1.385
r82 26 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.355 $Y=1.55
+ $X2=1.355 $Y2=1.95
r83 24 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.125 $Y=2.815
+ $X2=1.125 $Y2=2.12
r84 20 34 12.9221 $w=3.21e-07 $l=4.36348e-07 $layer=LI1_cond $X=1.27 $Y=1.045
+ $X2=1.49 $Y2=1.385
r85 20 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.27 $Y=1.045
+ $X2=0.935 $Y2=1.045
r86 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.77 $Y=0.96
+ $X2=0.935 $Y2=1.045
r87 16 18 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.77 $Y=0.96
+ $X2=0.77 $Y2=0.835
r88 14 35 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=1.385
+ $X2=1.545 $Y2=1.385
r89 14 15 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.83 $Y=1.385 $X2=1.92
+ $Y2=1.385
r90 11 15 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.935 $Y=1.22
+ $X2=1.92 $Y2=1.385
r91 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.935 $Y=1.22
+ $X2=1.935 $Y2=0.74
r92 7 15 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.55
+ $X2=1.92 $Y2=1.385
r93 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.92 $Y=1.55 $X2=1.92
+ $Y2=2.4
r94 2 29 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.96 $X2=1.125 $Y2=2.115
r95 2 24 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.96 $X2=1.125 $Y2=2.815
r96 1 18 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.56 $X2=0.77 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%B2 3 7 10 12 15 16 20
c45 15 0 8.02067e-21 $X=2.64 $Y=1.665
r46 15 16 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r47 13 15 6.26328 $w=2.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.54
+ $X2=2.64 $Y2=1.665
r48 12 13 2.67223 $w=2.3e-07 $l=1.6e-07 $layer=LI1_cond $X=2.64 $Y=1.38 $X2=2.64
+ $Y2=1.54
r49 10 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.385
+ $X2=2.385 $Y2=1.55
r50 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.385
+ $X2=2.385 $Y2=1.22
r51 9 12 9.18353 $w=3.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.385 $Y=1.38
+ $X2=2.64 $Y2=1.38
r52 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.385 $X2=2.385 $Y2=1.385
r53 7 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.365 $Y=0.74
+ $X2=2.365 $Y2=1.22
r54 3 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.37 $Y=2.4 $X2=2.37
+ $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%B1 1 3 6 8 14
r29 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r30 12 14 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=2.85 $Y=1.385
+ $X2=3.09 $Y2=1.385
r31 10 12 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.835 $Y=1.385
+ $X2=2.85 $Y2=1.385
r32 8 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r33 4 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.55
+ $X2=2.85 $Y2=1.385
r34 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.85 $Y=1.55 $X2=2.85
+ $Y2=2.4
r35 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.22
+ $X2=2.835 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.835 $Y=1.22 $X2=2.835
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%VPWR 1 2 7 9 14 18 21 22 23 33 34
c43 18 0 1.19783e-19 $X=2.61 $Y=2.815
r44 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 25 37 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r52 25 27 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=0.72
+ $Y2=3.33
r53 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 23 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 21 30 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.43 $Y=3.33 $X2=2.16
+ $Y2=3.33
r56 21 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=3.33
+ $X2=2.515 $Y2=3.33
r57 20 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.6 $Y=3.33 $X2=3.12
+ $Y2=3.33
r58 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=3.33 $X2=2.515
+ $Y2=3.33
r59 15 18 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.515 $Y=2.855
+ $X2=2.61 $Y2=2.855
r60 14 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=3.33
r61 13 15 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=2.98
+ $X2=2.515 $Y2=2.855
r62 13 14 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.515 $Y=2.98
+ $X2=2.515 $Y2=3.245
r63 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.285 $Y=2.115
+ $X2=0.285 $Y2=2.815
r64 7 37 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r65 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.815
r66 2 18 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.84 $X2=2.61 $Y2=2.815
r67 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.96 $X2=0.285 $Y2=2.815
r68 1 9 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.96 $X2=0.285 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%Y 1 2 10 11 13 19 23
c47 13 0 1.45091e-19 $X=2.15 $Y=0.515
r48 23 25 7.73239 $w=4.26e-07 $l=2.7e-07 $layer=LI1_cond $X=1.695 $Y=2.082
+ $X2=1.965 $Y2=2.082
r49 19 25 5.58451 $w=4.26e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=2.082
+ $X2=1.965 $Y2=2.082
r50 11 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.185 $Y=0.965
+ $X2=1.965 $Y2=0.965
r51 11 13 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=2.185 $Y=0.88
+ $X2=2.185 $Y2=0.515
r52 10 25 6.16288 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=1.965 $Y=1.75
+ $X2=1.965 $Y2=2.082
r53 9 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=1.05
+ $X2=1.965 $Y2=0.965
r54 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.965 $Y=1.05 $X2=1.965
+ $Y2=1.75
r55 2 23 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=1.57
+ $Y=1.84 $X2=1.695 $Y2=2.4
r56 2 23 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.84 $X2=1.695 $Y2=1.985
r57 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.37 $X2=2.15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%A_402_368# 1 2 9 11 12 15 19 21
r27 17 21 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.56
+ $X2=3.115 $Y2=2.475
r28 17 19 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.115 $Y=2.56
+ $X2=3.115 $Y2=2.815
r29 13 21 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.39
+ $X2=3.115 $Y2=2.475
r30 13 15 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=3.115 $Y=2.39
+ $X2=3.115 $Y2=1.985
r31 11 21 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=3.115 $Y2=2.475
r32 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=2.23 $Y2=2.475
r33 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.105 $Y=2.56
+ $X2=2.23 $Y2=2.475
r34 7 9 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=2.56
+ $X2=2.105 $Y2=2.685
r35 2 19 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.84 $X2=3.075 $Y2=2.815
r36 2 15 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.84 $X2=3.075 $Y2=1.985
r37 1 9 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=2.01 $Y=1.84
+ $X2=2.145 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_1%VGND 1 2 3 10 12 14 16 18 20 25 39 44
r43 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 39 41 1.27749 $w=7.64e-07 $l=8e-08 $layer=LI1_cond $X=1.495 $Y=0.625
+ $X2=1.495 $Y2=0.705
r45 34 39 9.98037 $w=7.64e-07 $l=6.25e-07 $layer=LI1_cond $X=1.495 $Y=0
+ $X2=1.495 $Y2=0.625
r46 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 29 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r49 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 26 34 9.90117 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.495
+ $Y2=0
r51 26 28 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.64
+ $Y2=0
r52 25 43 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.122
+ $Y2=0
r53 25 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.64
+ $Y2=0
r54 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r55 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r56 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 21 31 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r58 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r59 20 34 9.90117 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.495
+ $Y2=0
r60 20 23 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.72
+ $Y2=0
r61 18 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r62 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 14 43 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.122 $Y2=0
r65 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0.515
r66 10 31 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.212 $Y2=0
r67 10 12 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.815
r68 3 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.91
+ $Y=0.37 $X2=3.05 $Y2=0.515
r69 2 41 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.56 $X2=1.27 $Y2=0.705
r70 2 39 182 $w=1.7e-07 $l=6.91737e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.56 $X2=1.72 $Y2=0.625
r71 1 12 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.56 $X2=0.34 $Y2=0.815
.ends


* File: sky130_fd_sc_ms__and4b_2.pxi.spice
* Created: Wed Sep  2 11:58:42 2020
* 
x_PM_SKY130_FD_SC_MS__AND4B_2%A_N N_A_N_M1005_g N_A_N_M1010_g A_N N_A_N_c_80_n
+ N_A_N_c_81_n PM_SKY130_FD_SC_MS__AND4B_2%A_N
x_PM_SKY130_FD_SC_MS__AND4B_2%A_186_48# N_A_186_48#_M1012_d N_A_186_48#_M1002_d
+ N_A_186_48#_M1003_d N_A_186_48#_M1004_g N_A_186_48#_M1007_g
+ N_A_186_48#_M1013_g N_A_186_48#_M1009_g N_A_186_48#_c_112_n
+ N_A_186_48#_c_113_n N_A_186_48#_c_183_p N_A_186_48#_c_164_p
+ N_A_186_48#_c_126_p N_A_186_48#_c_114_n N_A_186_48#_c_115_n
+ N_A_186_48#_c_116_n N_A_186_48#_c_117_n PM_SKY130_FD_SC_MS__AND4B_2%A_186_48#
x_PM_SKY130_FD_SC_MS__AND4B_2%D N_D_M1002_g N_D_M1000_g D N_D_c_218_n
+ N_D_c_219_n PM_SKY130_FD_SC_MS__AND4B_2%D
x_PM_SKY130_FD_SC_MS__AND4B_2%C N_C_M1006_g N_C_M1001_g C N_C_c_254_n
+ N_C_c_255_n PM_SKY130_FD_SC_MS__AND4B_2%C
x_PM_SKY130_FD_SC_MS__AND4B_2%B N_B_M1008_g N_B_M1003_g B N_B_c_288_n
+ N_B_c_289_n PM_SKY130_FD_SC_MS__AND4B_2%B
x_PM_SKY130_FD_SC_MS__AND4B_2%A_27_112# N_A_27_112#_M1010_s N_A_27_112#_M1005_s
+ N_A_27_112#_M1012_g N_A_27_112#_M1011_g N_A_27_112#_c_323_n
+ N_A_27_112#_c_324_n N_A_27_112#_c_325_n N_A_27_112#_c_326_n
+ N_A_27_112#_c_355_n N_A_27_112#_c_331_n N_A_27_112#_c_332_n
+ N_A_27_112#_c_327_n N_A_27_112#_c_328_n PM_SKY130_FD_SC_MS__AND4B_2%A_27_112#
x_PM_SKY130_FD_SC_MS__AND4B_2%VPWR N_VPWR_M1005_d N_VPWR_M1009_s N_VPWR_M1006_d
+ N_VPWR_M1011_d N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n VPWR
+ N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_408_n
+ PM_SKY130_FD_SC_MS__AND4B_2%VPWR
x_PM_SKY130_FD_SC_MS__AND4B_2%X N_X_M1004_s N_X_M1007_d N_X_c_462_n N_X_c_463_n
+ N_X_c_464_n X PM_SKY130_FD_SC_MS__AND4B_2%X
x_PM_SKY130_FD_SC_MS__AND4B_2%VGND N_VGND_M1010_d N_VGND_M1013_d N_VGND_c_499_n
+ N_VGND_c_500_n VGND N_VGND_c_501_n N_VGND_c_502_n N_VGND_c_503_n
+ N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n PM_SKY130_FD_SC_MS__AND4B_2%VGND
cc_1 VNB N_A_N_M1005_g 0.00201544f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_2 VNB N_A_N_M1010_g 0.0304431f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB N_A_N_c_80_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_A_N_c_81_n 0.0584835f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_5 VNB N_A_186_48#_M1004_g 0.021717f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_6 VNB N_A_186_48#_M1007_g 0.00156209f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_7 VNB N_A_186_48#_M1013_g 0.0244852f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_8 VNB N_A_186_48#_M1009_g 0.00168247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_186_48#_c_112_n 4.01658e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_186_48#_c_113_n 0.0433786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_186_48#_c_114_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_186_48#_c_115_n 0.00565042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_186_48#_c_116_n 0.00320654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_186_48#_c_117_n 0.0553269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_M1000_g 0.0266603f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_16 VNB N_D_c_218_n 0.0267803f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_17 VNB N_D_c_219_n 0.00182951f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_18 VNB N_C_M1001_g 0.0256596f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_19 VNB N_C_c_254_n 0.0266074f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_20 VNB N_C_c_255_n 0.00181929f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_21 VNB N_B_M1008_g 0.0276909f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_22 VNB N_B_c_288_n 0.0246954f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_23 VNB N_B_c_289_n 0.00442487f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_24 VNB N_A_27_112#_M1012_g 0.0358374f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_A_27_112#_c_323_n 0.0195128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_112#_c_324_n 0.00140869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_112#_c_325_n 0.00927871f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_28 VNB N_A_27_112#_c_326_n 0.00959177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_112#_c_327_n 0.027381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_112#_c_328_n 0.0141382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_408_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_462_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_X_c_463_n 0.00156999f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_34 VNB N_X_c_464_n 0.00417716f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_35 VNB N_VGND_c_499_n 0.0157594f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_VGND_c_500_n 0.00951062f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_37 VNB N_VGND_c_501_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_502_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_503_n 0.0679994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_504_n 0.292092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_505_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_506_n 0.0115483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A_N_M1005_g 0.0304908f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_44 VPB N_A_N_c_80_n 0.00716464f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_45 VPB N_A_186_48#_M1007_g 0.0240125f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_46 VPB N_A_186_48#_M1009_g 0.0243322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_186_48#_c_112_n 0.00288026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_D_M1002_g 0.0221449f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_49 VPB N_D_c_218_n 0.00571233f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_50 VPB N_D_c_219_n 0.00273725f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_51 VPB N_C_M1006_g 0.0227334f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_52 VPB N_C_c_254_n 0.00564812f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_53 VPB N_C_c_255_n 0.00203503f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_54 VPB N_B_M1003_g 0.022337f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_55 VPB N_B_c_288_n 0.00550506f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_56 VPB N_B_c_289_n 0.00366259f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_57 VPB N_A_27_112#_M1011_g 0.022679f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_58 VPB N_A_27_112#_c_326_n 0.00315737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_27_112#_c_331_n 0.00692364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_112#_c_332_n 0.0350794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_27_112#_c_327_n 0.00581541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_112#_c_328_n 9.55674e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_409_n 0.0164086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_410_n 0.02094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_411_n 0.013668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_412_n 0.0191428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_413_n 0.0126731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_414_n 0.0288985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_415_n 0.0242802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_416_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_417_n 0.0247575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_418_n 0.0274817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_419_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_408_n 0.0765579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_X_c_463_n 0.00152646f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_76 VPB X 0.00445124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 N_A_N_M1010_g N_A_186_48#_M1004_g 0.0179601f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_78 N_A_N_M1005_g N_A_186_48#_M1007_g 0.0181549f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_79 N_A_N_c_81_n N_A_186_48#_c_117_n 0.0231581f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A_N_M1010_g N_A_27_112#_c_323_n 0.00822581f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_81 N_A_N_M1010_g N_A_27_112#_c_324_n 0.0142232f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_82 N_A_N_c_80_n N_A_27_112#_c_324_n 6.31955e-19 $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_83 N_A_N_c_81_n N_A_27_112#_c_324_n 0.00103766f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_84 N_A_N_M1010_g N_A_27_112#_c_325_n 0.00275868f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_85 N_A_N_c_80_n N_A_27_112#_c_325_n 0.0273182f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_86 N_A_N_c_81_n N_A_27_112#_c_325_n 0.00228689f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_87 N_A_N_M1010_g N_A_27_112#_c_326_n 0.00420609f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_88 N_A_N_c_80_n N_A_27_112#_c_326_n 0.0360322f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_89 N_A_N_c_81_n N_A_27_112#_c_326_n 0.00676086f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_90 N_A_N_M1005_g N_A_27_112#_c_332_n 0.0328168f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_91 N_A_N_c_80_n N_A_27_112#_c_332_n 0.0264887f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_92 N_A_N_c_81_n N_A_27_112#_c_332_n 0.00146577f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_93 N_A_N_M1005_g N_VPWR_c_409_n 0.00284156f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_94 N_A_N_M1005_g N_VPWR_c_418_n 0.0046462f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_95 N_A_N_M1005_g N_VPWR_c_408_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_96 N_A_N_M1010_g N_X_c_462_n 7.4905e-19 $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_97 N_A_N_M1005_g X 2.1398e-19 $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_98 N_A_N_M1010_g N_VGND_c_499_n 0.00430723f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_99 N_A_N_M1010_g N_VGND_c_501_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_100 N_A_N_M1010_g N_VGND_c_504_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_101 N_A_186_48#_M1009_g N_D_M1002_g 0.0311369f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_186_48#_c_112_n N_D_M1002_g 0.00375262f $X=1.695 $Y=1.95 $X2=0 $Y2=0
cc_103 N_A_186_48#_c_126_p N_D_M1002_g 0.0129328f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_104 N_A_186_48#_M1013_g N_D_M1000_g 0.00908327f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_186_48#_c_113_n N_D_M1000_g 0.0156497f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_106 N_A_186_48#_c_116_n N_D_M1000_g 0.00418176f $X=1.587 $Y=1.3 $X2=0 $Y2=0
cc_107 N_A_186_48#_c_117_n N_D_M1000_g 0.00120051f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_108 N_A_186_48#_M1009_g N_D_c_218_n 0.00123737f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_186_48#_c_113_n N_D_c_218_n 0.00118546f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_110 N_A_186_48#_c_126_p N_D_c_218_n 6.00553e-19 $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A_186_48#_c_115_n N_D_c_218_n 0.00208763f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_112 N_A_186_48#_c_117_n N_D_c_218_n 0.0148535f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_113 N_A_186_48#_c_113_n N_D_c_219_n 0.0202397f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_114 N_A_186_48#_c_126_p N_D_c_219_n 0.0212976f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_186_48#_c_115_n N_D_c_219_n 0.032015f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_116 N_A_186_48#_c_117_n N_D_c_219_n 3.17162e-19 $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_117 N_A_186_48#_c_126_p N_C_M1006_g 0.0132054f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_118 N_A_186_48#_c_113_n N_C_M1001_g 0.0155906f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_119 N_A_186_48#_c_113_n N_C_c_254_n 0.00118572f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_120 N_A_186_48#_c_126_p N_C_c_254_n 7.23988e-19 $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_121 N_A_186_48#_c_113_n N_C_c_255_n 0.0202359f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_122 N_A_186_48#_c_126_p N_C_c_255_n 0.0235433f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_123 N_A_186_48#_c_113_n N_B_M1008_g 0.0164071f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_124 N_A_186_48#_c_114_n N_B_M1008_g 0.00282462f $X=3.905 $Y=0.515 $X2=0 $Y2=0
cc_125 N_A_186_48#_c_126_p N_B_M1003_g 0.0132054f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_126 N_A_186_48#_c_113_n N_B_c_288_n 0.00118828f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_127 N_A_186_48#_c_126_p N_B_c_288_n 4.43489e-19 $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_128 N_A_186_48#_c_113_n N_B_c_289_n 0.0249816f $X=3.74 $Y=1.045 $X2=0 $Y2=0
cc_129 N_A_186_48#_c_126_p N_B_c_289_n 0.027051f $X=3.46 $Y=2.035 $X2=0 $Y2=0
cc_130 N_A_186_48#_c_113_n N_A_27_112#_M1012_g 0.0131028f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_131 N_A_186_48#_c_114_n N_A_27_112#_M1012_g 0.0139597f $X=3.905 $Y=0.515
+ $X2=0 $Y2=0
cc_132 N_A_186_48#_c_126_p N_A_27_112#_M1011_g 0.0038447f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_133 N_A_186_48#_M1004_g N_A_27_112#_c_323_n 5.13233e-19 $X=1.005 $Y=0.74
+ $X2=0 $Y2=0
cc_134 N_A_186_48#_M1004_g N_A_27_112#_c_324_n 0.00156766f $X=1.005 $Y=0.74
+ $X2=0 $Y2=0
cc_135 N_A_186_48#_M1004_g N_A_27_112#_c_326_n 0.00275641f $X=1.005 $Y=0.74
+ $X2=0 $Y2=0
cc_136 N_A_186_48#_c_117_n N_A_27_112#_c_326_n 0.00415156f $X=1.5 $Y=1.465 $X2=0
+ $Y2=0
cc_137 N_A_186_48#_M1002_d N_A_27_112#_c_355_n 0.00539181f $X=2.21 $Y=1.84 $X2=0
+ $Y2=0
cc_138 N_A_186_48#_M1003_d N_A_27_112#_c_355_n 0.00582957f $X=3.305 $Y=1.84
+ $X2=0 $Y2=0
cc_139 N_A_186_48#_M1007_g N_A_27_112#_c_355_n 0.0163543f $X=1.05 $Y=2.4 $X2=0
+ $Y2=0
cc_140 N_A_186_48#_M1009_g N_A_27_112#_c_355_n 0.0185309f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_141 N_A_186_48#_c_164_p N_A_27_112#_c_355_n 0.0107758f $X=1.78 $Y=2.075 $X2=0
+ $Y2=0
cc_142 N_A_186_48#_c_126_p N_A_27_112#_c_355_n 0.106612f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_143 N_A_186_48#_M1007_g N_A_27_112#_c_332_n 0.00760665f $X=1.05 $Y=2.4 $X2=0
+ $Y2=0
cc_144 N_A_186_48#_c_113_n N_A_27_112#_c_327_n 0.00419666f $X=3.74 $Y=1.045
+ $X2=0 $Y2=0
cc_145 N_A_186_48#_c_113_n N_A_27_112#_c_328_n 0.0243261f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_146 N_A_186_48#_c_126_p N_A_27_112#_c_328_n 0.00149841f $X=3.46 $Y=2.035
+ $X2=0 $Y2=0
cc_147 N_A_186_48#_c_112_n N_VPWR_M1009_s 0.0021392f $X=1.695 $Y=1.95 $X2=0
+ $Y2=0
cc_148 N_A_186_48#_c_164_p N_VPWR_M1009_s 0.00324346f $X=1.78 $Y=2.075 $X2=0
+ $Y2=0
cc_149 N_A_186_48#_c_126_p N_VPWR_M1009_s 0.0104748f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_150 N_A_186_48#_c_126_p N_VPWR_M1006_d 0.0129639f $X=3.46 $Y=2.035 $X2=0
+ $Y2=0
cc_151 N_A_186_48#_M1007_g N_VPWR_c_409_n 0.0107954f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_186_48#_M1009_g N_VPWR_c_409_n 0.00113074f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_186_48#_M1007_g N_VPWR_c_410_n 0.00490827f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_186_48#_M1009_g N_VPWR_c_410_n 0.00553757f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_186_48#_M1009_g N_VPWR_c_411_n 0.00536428f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_186_48#_M1007_g N_VPWR_c_408_n 0.00478018f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_186_48#_M1009_g N_VPWR_c_408_n 0.00545239f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_186_48#_M1004_g N_X_c_462_n 0.00909182f $X=1.005 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_186_48#_M1013_g N_X_c_462_n 0.0132513f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_186_48#_c_183_p N_X_c_462_n 0.0113177f $X=1.78 $Y=1.045 $X2=0 $Y2=0
cc_161 N_A_186_48#_M1004_g N_X_c_463_n 0.00331189f $X=1.005 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_186_48#_M1007_g N_X_c_463_n 0.00455437f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_186_48#_M1013_g N_X_c_463_n 0.00142748f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_186_48#_M1009_g N_X_c_463_n 0.00145866f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A_186_48#_c_112_n N_X_c_463_n 0.00807612f $X=1.695 $Y=1.95 $X2=0 $Y2=0
cc_166 N_A_186_48#_c_115_n N_X_c_463_n 0.0238617f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_167 N_A_186_48#_c_116_n N_X_c_463_n 0.00718069f $X=1.587 $Y=1.3 $X2=0 $Y2=0
cc_168 N_A_186_48#_c_117_n N_X_c_463_n 0.0143033f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_169 N_A_186_48#_M1004_g N_X_c_464_n 0.00225198f $X=1.005 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_186_48#_M1013_g N_X_c_464_n 0.00346455f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_186_48#_c_117_n N_X_c_464_n 0.00201958f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_172 N_A_186_48#_M1007_g X 0.0081643f $X=1.05 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A_186_48#_M1009_g X 0.0053955f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_186_48#_c_112_n X 0.00566345f $X=1.695 $Y=1.95 $X2=0 $Y2=0
cc_175 N_A_186_48#_c_115_n X 0.00312735f $X=1.56 $Y=1.465 $X2=0 $Y2=0
cc_176 N_A_186_48#_c_117_n X 0.00381194f $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_177 N_A_186_48#_c_113_n N_VGND_M1013_d 0.00478095f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_178 N_A_186_48#_c_183_p N_VGND_M1013_d 0.00472321f $X=1.78 $Y=1.045 $X2=0
+ $Y2=0
cc_179 N_A_186_48#_M1004_g N_VGND_c_499_n 0.00603022f $X=1.005 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_A_186_48#_M1013_g N_VGND_c_500_n 0.00456117f $X=1.435 $Y=0.74 $X2=0
+ $Y2=0
cc_181 N_A_186_48#_c_113_n N_VGND_c_500_n 0.0264272f $X=3.74 $Y=1.045 $X2=0
+ $Y2=0
cc_182 N_A_186_48#_c_183_p N_VGND_c_500_n 0.0153275f $X=1.78 $Y=1.045 $X2=0
+ $Y2=0
cc_183 N_A_186_48#_c_115_n N_VGND_c_500_n 0.00168337f $X=1.56 $Y=1.465 $X2=0
+ $Y2=0
cc_184 N_A_186_48#_c_117_n N_VGND_c_500_n 7.5336e-19 $X=1.5 $Y=1.465 $X2=0 $Y2=0
cc_185 N_A_186_48#_M1004_g N_VGND_c_502_n 0.00434272f $X=1.005 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_186_48#_M1013_g N_VGND_c_502_n 0.00434272f $X=1.435 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_186_48#_c_114_n N_VGND_c_503_n 0.0145639f $X=3.905 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_186_48#_M1004_g N_VGND_c_504_n 0.00825283f $X=1.005 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_186_48#_M1013_g N_VGND_c_504_n 0.00822601f $X=1.435 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_186_48#_c_114_n N_VGND_c_504_n 0.0119984f $X=3.905 $Y=0.515 $X2=0
+ $Y2=0
cc_191 N_A_186_48#_c_113_n A_459_74# 0.0048076f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_186_48#_c_113_n A_537_74# 0.0107783f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_186_48#_c_113_n A_645_74# 0.0107783f $X=3.74 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_194 N_D_M1002_g N_C_M1006_g 0.0401329f $X=2.12 $Y=2.34 $X2=0 $Y2=0
cc_195 N_D_c_219_n N_C_M1006_g 6.21071e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_196 N_D_M1000_g N_C_M1001_g 0.0614519f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_197 N_D_c_218_n N_C_c_254_n 0.0201104f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_198 N_D_c_219_n N_C_c_254_n 0.00114936f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_199 N_D_c_218_n N_C_c_255_n 0.00114936f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_200 N_D_c_219_n N_C_c_255_n 0.0276388f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_201 N_D_M1002_g N_A_27_112#_c_355_n 0.0139734f $X=2.12 $Y=2.34 $X2=0 $Y2=0
cc_202 N_D_M1002_g N_VPWR_c_411_n 0.00463f $X=2.12 $Y=2.34 $X2=0 $Y2=0
cc_203 N_D_M1002_g N_VPWR_c_415_n 0.0059286f $X=2.12 $Y=2.34 $X2=0 $Y2=0
cc_204 N_D_M1002_g N_VPWR_c_408_n 0.00610055f $X=2.12 $Y=2.34 $X2=0 $Y2=0
cc_205 N_D_M1000_g N_VGND_c_500_n 0.0145292f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_206 N_D_M1000_g N_VGND_c_503_n 0.00398535f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_207 N_D_M1000_g N_VGND_c_504_n 0.00787244f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_208 N_C_M1001_g N_B_M1008_g 0.0402276f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_209 N_C_M1006_g N_B_M1003_g 0.0348318f $X=2.595 $Y=2.34 $X2=0 $Y2=0
cc_210 N_C_c_255_n N_B_M1003_g 2.95591e-19 $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_211 N_C_c_254_n N_B_c_288_n 0.0173872f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_212 N_C_c_255_n N_B_c_288_n 3.65288e-19 $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_213 N_C_M1006_g N_B_c_289_n 2.85078e-19 $X=2.595 $Y=2.34 $X2=0 $Y2=0
cc_214 N_C_c_254_n N_B_c_289_n 0.00202953f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_215 N_C_c_255_n N_B_c_289_n 0.0349699f $X=2.67 $Y=1.515 $X2=0 $Y2=0
cc_216 N_C_M1006_g N_A_27_112#_c_355_n 0.0139383f $X=2.595 $Y=2.34 $X2=0 $Y2=0
cc_217 N_C_M1006_g N_VPWR_c_412_n 0.00463f $X=2.595 $Y=2.34 $X2=0 $Y2=0
cc_218 N_C_M1006_g N_VPWR_c_415_n 0.0059286f $X=2.595 $Y=2.34 $X2=0 $Y2=0
cc_219 N_C_M1006_g N_VPWR_c_408_n 0.00610055f $X=2.595 $Y=2.34 $X2=0 $Y2=0
cc_220 N_C_M1001_g N_VGND_c_500_n 0.00269307f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_221 N_C_M1001_g N_VGND_c_503_n 0.00461464f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_222 N_C_M1001_g N_VGND_c_504_n 0.00910057f $X=2.61 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B_M1008_g N_A_27_112#_M1012_g 0.0370849f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_224 N_B_M1003_g N_A_27_112#_M1011_g 0.0370952f $X=3.215 $Y=2.34 $X2=0 $Y2=0
cc_225 N_B_c_289_n N_A_27_112#_M1011_g 8.91029e-19 $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_226 N_B_M1003_g N_A_27_112#_c_355_n 0.0140575f $X=3.215 $Y=2.34 $X2=0 $Y2=0
cc_227 N_B_c_289_n N_A_27_112#_c_331_n 0.00436141f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_228 N_B_c_288_n N_A_27_112#_c_327_n 0.0207808f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_229 N_B_c_289_n N_A_27_112#_c_327_n 4.1329e-19 $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_230 N_B_c_288_n N_A_27_112#_c_328_n 0.00114347f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_231 N_B_c_289_n N_A_27_112#_c_328_n 0.0213706f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B_M1003_g N_VPWR_c_412_n 0.00463f $X=3.215 $Y=2.34 $X2=0 $Y2=0
cc_233 N_B_M1003_g N_VPWR_c_417_n 0.0059286f $X=3.215 $Y=2.34 $X2=0 $Y2=0
cc_234 N_B_M1003_g N_VPWR_c_408_n 0.00610055f $X=3.215 $Y=2.34 $X2=0 $Y2=0
cc_235 N_B_M1008_g N_VGND_c_503_n 0.00461464f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B_M1008_g N_VGND_c_504_n 0.00911376f $X=3.15 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_27_112#_c_326_n N_VPWR_M1005_d 0.00119203f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_238 N_A_27_112#_c_355_n N_VPWR_M1005_d 0.00519989f $X=3.815 $Y=2.455
+ $X2=-0.19 $Y2=-0.245
cc_239 N_A_27_112#_c_332_n N_VPWR_M1005_d 0.00680924f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_27_112#_c_355_n N_VPWR_M1009_s 0.0076027f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_241 N_A_27_112#_c_355_n N_VPWR_M1006_d 0.00755633f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_242 N_A_27_112#_c_355_n N_VPWR_M1011_d 0.00919766f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_243 N_A_27_112#_c_331_n N_VPWR_M1011_d 0.0226986f $X=3.9 $Y=2.37 $X2=0 $Y2=0
cc_244 N_A_27_112#_c_355_n N_VPWR_c_409_n 0.00991706f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_245 N_A_27_112#_c_332_n N_VPWR_c_409_n 0.0125888f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_246 N_A_27_112#_c_355_n N_VPWR_c_411_n 0.0258995f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_247 N_A_27_112#_c_355_n N_VPWR_c_412_n 0.0258995f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_248 N_A_27_112#_M1011_g N_VPWR_c_414_n 0.00819554f $X=3.705 $Y=2.34 $X2=0
+ $Y2=0
cc_249 N_A_27_112#_c_355_n N_VPWR_c_414_n 0.0116318f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_250 N_A_27_112#_M1011_g N_VPWR_c_417_n 0.0059286f $X=3.705 $Y=2.34 $X2=0
+ $Y2=0
cc_251 N_A_27_112#_c_332_n N_VPWR_c_418_n 0.006683f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_252 N_A_27_112#_M1011_g N_VPWR_c_408_n 0.00610055f $X=3.705 $Y=2.34 $X2=0
+ $Y2=0
cc_253 N_A_27_112#_c_355_n N_VPWR_c_408_n 0.0786444f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_254 N_A_27_112#_c_332_n N_VPWR_c_408_n 0.0183785f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_255 N_A_27_112#_c_355_n N_X_M1007_d 0.00466364f $X=3.815 $Y=2.455 $X2=0 $Y2=0
cc_256 N_A_27_112#_c_323_n N_X_c_462_n 0.00441257f $X=0.28 $Y=0.835 $X2=0 $Y2=0
cc_257 N_A_27_112#_c_324_n N_X_c_462_n 0.0101363f $X=0.625 $Y=1.045 $X2=0 $Y2=0
cc_258 N_A_27_112#_c_326_n N_X_c_463_n 0.0358559f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_259 N_A_27_112#_c_326_n X 0.00697846f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_260 N_A_27_112#_c_355_n X 0.0202465f $X=3.815 $Y=2.455 $X2=0 $Y2=0
cc_261 N_A_27_112#_c_332_n X 0.0150412f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_262 N_A_27_112#_c_324_n N_VGND_M1010_d 0.00376661f $X=0.625 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_263 N_A_27_112#_c_323_n N_VGND_c_499_n 0.0096883f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_264 N_A_27_112#_c_324_n N_VGND_c_499_n 0.0151472f $X=0.625 $Y=1.045 $X2=0
+ $Y2=0
cc_265 N_A_27_112#_c_323_n N_VGND_c_501_n 0.00806442f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_266 N_A_27_112#_M1012_g N_VGND_c_503_n 0.00434272f $X=3.69 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_27_112#_M1012_g N_VGND_c_504_n 0.00826337f $X=3.69 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_27_112#_c_323_n N_VGND_c_504_n 0.0105742f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_269 N_X_c_462_n N_VGND_c_499_n 0.0164982f $X=1.22 $Y=0.515 $X2=0 $Y2=0
cc_270 N_X_c_462_n N_VGND_c_500_n 0.0173772f $X=1.22 $Y=0.515 $X2=0 $Y2=0
cc_271 N_X_c_462_n N_VGND_c_502_n 0.0144922f $X=1.22 $Y=0.515 $X2=0 $Y2=0
cc_272 N_X_c_462_n N_VGND_c_504_n 0.0118826f $X=1.22 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o32a_1.pex.spice
* Created: Wed Sep  2 12:26:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O32A_1%A_83_264# 1 2 9 13 16 17 18 21 23 25 26 29 31
+ 34
c93 25 0 1.9056e-19 $X=3.15 $Y=1.18
r94 29 39 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.485
+ $X2=0.58 $Y2=1.65
r95 29 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.485
+ $X2=0.58 $Y2=1.32
r96 28 31 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.58 $Y=1.485 $X2=0.7
+ $Y2=1.485
r97 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.485 $X2=0.58 $Y2=1.485
r98 25 36 13.3697 $w=4.98e-07 $l=3.90058e-07 $layer=LI1_cond $X=3.15 $Y=1.18
+ $X2=2.982 $Y2=0.865
r99 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.15 $Y=1.18
+ $X2=3.15 $Y2=1.95
r100 24 34 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.595 $Y=2.035
+ $X2=2.4 $Y2=2.035
r101 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.15 $Y2=1.95
r102 23 24 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=2.595 $Y2=2.035
r103 19 34 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.12 $X2=2.4
+ $Y2=2.035
r104 19 21 17.5821 $w=3.88e-07 $l=5.95e-07 $layer=LI1_cond $X=2.4 $Y=2.12
+ $X2=2.4 $Y2=2.715
r105 17 34 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.205 $Y=2.035
+ $X2=2.4 $Y2=2.035
r106 17 18 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=2.205 $Y=2.035
+ $X2=0.785 $Y2=2.035
r107 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.95
+ $X2=0.785 $Y2=2.035
r108 15 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=1.65 $X2=0.7
+ $Y2=1.485
r109 15 16 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.7 $Y=1.65 $X2=0.7
+ $Y2=1.95
r110 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.61 $Y=0.74
+ $X2=0.61 $Y2=1.32
r111 9 39 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.65
r112 2 34 400 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_PDIFF $count=1 $X=2.215
+ $Y=1.84 $X2=2.395 $Y2=2.035
r113 2 21 400 $w=1.7e-07 $l=9.60794e-07 $layer=licon1_PDIFF $count=1 $X=2.215
+ $Y=1.84 $X2=2.395 $Y2=2.715
r114 1 36 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.37 $X2=2.975 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%A1 3 7 9 12 13
c41 3 0 2.36033e-19 $X=1.165 $Y=2.34
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.515
+ $X2=1.12 $Y2=1.68
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.515
+ $X2=1.12 $Y2=1.35
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.515 $X2=1.12 $Y2=1.515
r45 9 13 4.80185 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.135 $Y=1.665
+ $X2=1.135 $Y2=1.515
r46 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.18 $Y=0.69 $X2=1.18
+ $Y2=1.35
r47 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.165 $Y=2.34
+ $X2=1.165 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%A2 3 7 9 12 13
c36 13 0 1.13074e-19 $X=1.66 $Y=1.515
c37 3 0 1.02106e-19 $X=1.585 $Y=2.34
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.515
+ $X2=1.66 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.515
+ $X2=1.66 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.515 $X2=1.66 $Y2=1.515
r41 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=1.515
r42 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.61 $Y=0.69 $X2=1.61
+ $Y2=1.35
r43 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.585 $Y=2.34
+ $X2=1.585 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%A3 3 7 9 12 13
c38 13 0 1.02106e-19 $X=2.2 $Y=1.515
c39 7 0 1.9056e-19 $X=2.18 $Y=0.69
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.515
+ $X2=2.2 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.515
+ $X2=2.2 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.2
+ $Y=1.515 $X2=2.2 $Y2=1.515
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=1.515
r44 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.18 $Y=0.69 $X2=2.18
+ $Y2=1.35
r45 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.125 $Y=2.34
+ $X2=2.125 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%B2 3 7 9 12 13
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.515
+ $X2=2.74 $Y2=1.68
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.515
+ $X2=2.74 $Y2=1.35
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.515 $X2=2.74 $Y2=1.515
r44 9 13 4.80185 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=2.715 $Y=1.665
+ $X2=2.715 $Y2=1.515
r45 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.68 $Y=0.69 $X2=2.68
+ $Y2=1.35
r46 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.665 $Y=2.34
+ $X2=2.665 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%B1 3 7 9 10 17
r30 15 17 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.275 $Y=1.345
+ $X2=3.57 $Y2=1.345
r31 13 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.26 $Y=1.345
+ $X2=3.275 $Y2=1.345
r32 9 10 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=3.572 $Y=1.295
+ $X2=3.572 $Y2=1.665
r33 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.345 $X2=3.57 $Y2=1.345
r34 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.18
+ $X2=3.275 $Y2=1.345
r35 5 7 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.275 $Y=1.18
+ $X2=3.275 $Y2=0.69
r36 1 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.51
+ $X2=3.26 $Y2=1.345
r37 1 3 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=3.26 $Y=1.51 $X2=3.26
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%X 1 2 11 14 15 16 17 23 29
c27 14 0 1.22959e-19 $X=0.28 $Y=1.985
r28 21 29 0.805779 $w=4.73e-07 $l=3.2e-08 $layer=LI1_cond $X=0.322 $Y=0.893
+ $X2=0.322 $Y2=0.925
r29 17 31 9.71933 $w=4.73e-07 $l=1.79e-07 $layer=LI1_cond $X=0.322 $Y=0.951
+ $X2=0.322 $Y2=1.13
r30 17 29 0.654696 $w=4.73e-07 $l=2.6e-08 $layer=LI1_cond $X=0.322 $Y=0.951
+ $X2=0.322 $Y2=0.925
r31 17 21 0.679876 $w=4.73e-07 $l=2.7e-08 $layer=LI1_cond $X=0.322 $Y=0.866
+ $X2=0.322 $Y2=0.893
r32 16 17 7.83117 $w=4.73e-07 $l=3.11e-07 $layer=LI1_cond $X=0.322 $Y=0.555
+ $X2=0.322 $Y2=0.866
r33 16 23 1.00722 $w=4.73e-07 $l=4e-08 $layer=LI1_cond $X=0.322 $Y=0.555
+ $X2=0.322 $Y2=0.515
r34 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.82 $X2=0.17
+ $Y2=1.13
r35 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=1.82
r36 9 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=1.985
r37 9 11 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=2.815
r38 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r39 2 11 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r40 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.25
+ $Y=0.37 $X2=0.395 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%VPWR 1 2 9 13 14 16 19 22 24 29 38 42
r41 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 36 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r49 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 29 41 4.5891 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.32 $Y=3.33 $X2=3.58
+ $Y2=3.33
r51 29 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.32 $Y=3.33 $X2=3.12
+ $Y2=3.33
r52 27 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r55 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 22 36 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 22 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 19 21 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.53 $Y=2.135
+ $X2=3.53 $Y2=2.29
r59 14 41 3.17707 $w=3.3e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.485 $Y=3.245
+ $X2=3.58 $Y2=3.33
r60 14 16 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.485 $Y=3.245
+ $X2=3.485 $Y2=2.695
r61 13 21 6.63994 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=2.455
+ $X2=3.485 $Y2=2.29
r62 13 16 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.485 $Y=2.455
+ $X2=3.485 $Y2=2.695
r63 9 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.78 $Y=2.455
+ $X2=0.78 $Y2=2.815
r64 7 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r65 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.815
r66 2 19 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=1.84 $X2=3.495 $Y2=2.135
r67 2 16 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=1.84 $X2=3.485 $Y2=2.695
r68 1 12 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.815
r69 1 9 600 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 32 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r46 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r47 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r50 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 21 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r52 21 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r53 19 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.68
+ $Y2=0
r54 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.895
+ $Y2=0
r55 18 31 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=2.16
+ $Y2=0
r56 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=0 $X2=1.895
+ $Y2=0
r57 16 24 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.73 $Y=0 $X2=0.72
+ $Y2=0
r58 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0 $X2=0.895
+ $Y2=0
r59 15 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=1.68
+ $Y2=0
r60 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.895
+ $Y2=0
r61 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.085
+ $X2=1.895 $Y2=0
r62 11 13 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=1.895 $Y=0.085
+ $X2=1.895 $Y2=0.655
r63 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0
r64 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0.515
r65 2 13 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.37 $X2=1.895 $Y2=0.655
r66 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.685
+ $Y=0.37 $X2=0.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_1%A_251_74# 1 2 3 12 14 15 16 17 18 25
r48 19 23 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0.43
+ $X2=2.395 $Y2=0.43
r49 18 25 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.405 $Y=0.43
+ $X2=3.53 $Y2=0.43
r50 18 19 52.0657 $w=1.78e-07 $l=8.45e-07 $layer=LI1_cond $X=3.405 $Y=0.43
+ $X2=2.56 $Y2=0.43
r51 16 23 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.395 $Y=0.52 $X2=2.395
+ $Y2=0.43
r52 16 17 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.395 $Y=0.52
+ $X2=2.395 $Y2=1.01
r53 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.23 $Y=1.095
+ $X2=2.395 $Y2=1.01
r54 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.23 $Y=1.095
+ $X2=1.56 $Y2=1.095
r55 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.395 $Y=1.01
+ $X2=1.56 $Y2=1.095
r56 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.395 $Y=1.01
+ $X2=1.395 $Y2=0.515
r57 3 25 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.35
+ $Y=0.37 $X2=3.49 $Y2=0.505
r58 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.255
+ $Y=0.37 $X2=2.395 $Y2=0.515
r59 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.255
+ $Y=0.37 $X2=1.395 $Y2=0.515
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor3_4 A B C VGND VNB VPB VPWR X
M1000 VPWR C a_1155_284# VPB pshort w=640000u l=180000u
+  ad=2.1152e+12p pd=1.487e+07u as=1.792e+11p ps=1.84e+06u
M1001 VGND C a_1155_284# VNB nlowvt w=420000u l=150000u
+  ad=1.6131e+12p pd=1.223e+07u as=2.121e+11p ps=1.85e+06u
M1002 VPWR a_74_294# a_27_118# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6055e+11p ps=4.93e+06u
M1003 a_1221_388# a_1155_284# a_416_118# VPB pshort w=840000u l=180000u
+  ad=4.2e+11p pd=2.68e+06u as=6.5265e+11p ps=4.95e+06u
M1004 VGND a_1221_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1005 VGND a_74_294# a_27_118# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.264e+11p ps=4.03e+06u
M1006 a_326_392# B a_27_118# VNB nlowvt w=640000u l=150000u
+  ad=4.6775e+11p pd=4.06e+06u as=0p ps=0u
M1007 a_326_392# C a_1221_388# VPB pshort w=840000u l=180000u
+  ad=5.184e+11p pd=4.63e+06u as=0p ps=0u
M1008 a_1221_388# a_1155_284# a_326_392# VNB nlowvt w=640000u l=150000u
+  ad=3.392e+11p pd=2.34e+06u as=0p ps=0u
M1009 a_326_392# B a_74_294# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=8.764e+11p ps=5.66e+06u
M1010 X a_1221_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_1221_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_1221_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1013 a_416_118# B a_74_294# VNB nlowvt w=640000u l=150000u
+  ad=3.899e+11p pd=3.83e+06u as=7.264e+11p ps=4.83e+06u
M1014 a_74_294# a_397_320# a_416_118# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR B a_397_320# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1016 a_416_118# C a_1221_388# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_1221_388# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_118# a_397_320# a_416_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_118# a_397_320# a_326_392# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1221_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_416_118# B a_27_118# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1221_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_74_294# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B a_397_320# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1025 a_74_294# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1221_388# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_74_294# a_397_320# a_326_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__inv_8.spice
* Created: Fri Aug 28 17:38:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__inv_8.pex.spice"
.subckt sky130_fd_sc_ms__inv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75003.4
+ A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75003
+ A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1001_d N_A_M1010_g N_Y_M1010_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1 SB=75002.6
+ A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1010_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1011_d N_A_M1012_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.4 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1013_d N_A_M1014_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.2146
+ AS=0.1036 PD=2.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90003.5
+ A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6 SB=90003
+ A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.1 SB=90002.5
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6 SB=90002.1
+ A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002 SB=90001.6
+ A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5 SB=90001.2
+ A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1008_d N_A_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.4 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__inv_8.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__a311o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_261_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=8.9e+11p ps=5.96e+06u
M1001 VGND B1 a_89_270# VNB nlowvt w=640000u l=150000u
+  ad=5.289e+11p pd=4.33e+06u as=3.488e+11p ps=3.65e+06u
M1002 VPWR A2 a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_89_270# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_264_120# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=2.10625e+11p pd=1.96e+06u as=0p ps=0u
M1005 a_89_270# C1 a_549_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1006 VGND a_89_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1007 a_89_270# A1 a_359_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1008 a_261_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_549_392# B1 a_261_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_89_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1011 a_359_123# A2 a_264_120# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


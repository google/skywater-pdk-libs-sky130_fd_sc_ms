* File: sky130_fd_sc_ms__and2_1.pex.spice
* Created: Fri Aug 28 17:10:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND2_1%A 3 6 9 12 13 14 18
c33 12 0 9.98687e-20 $X=0.7 $Y=1.545
r34 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=0.405 $X2=0.61 $Y2=0.405
r35 14 19 3.05467 $w=4.13e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=0.462
+ $X2=0.61 $Y2=0.462
r36 13 19 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.462
+ $X2=0.61 $Y2=0.462
r37 11 12 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.7 $Y=1.395 $X2=0.7
+ $Y2=1.545
r38 9 12 386.766 $w=1.8e-07 $l=9.95e-07 $layer=POLY_cond $X=0.745 $Y=2.54
+ $X2=0.745 $Y2=1.545
r39 6 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.64 $Y=1 $X2=0.64
+ $Y2=1.395
r40 3 18 20.9154 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.64 $Y=0.57
+ $X2=0.67 $Y2=0.405
r41 3 6 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.64 $Y=0.57 $X2=0.64
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_1%B 3 6 8 11 13
r44 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.24 $Y=1.515
+ $X2=1.24 $Y2=1.68
r45 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.24 $Y=1.515
+ $X2=1.24 $Y2=1.35
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.515 $X2=1.24 $Y2=1.515
r47 8 12 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.24 $Y=1.295
+ $X2=1.24 $Y2=1.515
r48 6 14 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=1.245 $Y=2.54
+ $X2=1.245 $Y2=1.68
r49 3 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.21 $Y=0.92 $X2=1.21
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_1%A_56_136# 1 2 9 13 16 18 19 22 24 27 28 32 33
+ 36
c67 27 0 1.10419e-19 $X=1.665 $Y=1.85
r68 33 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.515
+ $X2=1.81 $Y2=1.68
r69 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.515
+ $X2=1.81 $Y2=1.35
r70 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.515 $X2=1.81 $Y2=1.515
r71 29 32 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.665 $Y=1.515
+ $X2=1.81 $Y2=1.515
r72 26 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=1.68
+ $X2=1.665 $Y2=1.515
r73 26 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.665 $Y=1.68
+ $X2=1.665 $Y2=1.85
r74 25 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=1.935
+ $X2=1.02 $Y2=1.935
r75 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=1.935
+ $X2=1.665 $Y2=1.85
r76 24 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.58 $Y=1.935
+ $X2=1.185 $Y2=1.935
r77 20 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=2.02 $X2=1.02
+ $Y2=1.935
r78 20 22 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.02 $Y=2.02
+ $X2=1.02 $Y2=2.265
r79 18 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=1.935
+ $X2=1.02 $Y2=1.935
r80 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.855 $Y=1.935
+ $X2=0.59 $Y2=1.935
r81 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.425 $Y=1.85
+ $X2=0.59 $Y2=1.935
r82 14 16 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=0.425 $Y=1.85
+ $X2=0.425 $Y2=1.03
r83 13 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.79 $Y=0.87 $X2=1.79
+ $Y2=1.35
r84 9 37 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.78 $Y=2.4 $X2=1.78
+ $Y2=1.68
r85 2 22 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.835
+ $Y=2.12 $X2=1.02 $Y2=2.265
r86 1 16 182 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_NDIFF $count=1 $X=0.28
+ $Y=0.68 $X2=0.425 $Y2=1.03
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_1%VPWR 1 2 9 13 16 17 19 20 21 31 32
c30 9 0 9.98687e-20 $X=0.515 $Y=2.295
c31 2 0 1.10419e-19 $X=1.335 $Y=2.12
r32 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 21 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r37 19 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.555 $Y2=3.33
r39 18 31 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.555 $Y2=3.33
r41 16 24 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.35 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 16 17 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.35 $Y=3.33
+ $X2=0.517 $Y2=3.33
r43 15 28 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=0.685 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 15 17 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.685 $Y=3.33
+ $X2=0.517 $Y2=3.33
r45 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=3.245
+ $X2=1.555 $Y2=3.33
r46 11 13 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=1.555 $Y=3.245
+ $X2=1.555 $Y2=2.355
r47 7 17 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.517 $Y=3.245
+ $X2=0.517 $Y2=3.33
r48 7 9 32.6812 $w=3.33e-07 $l=9.5e-07 $layer=LI1_cond $X=0.517 $Y=3.245
+ $X2=0.517 $Y2=2.295
r49 2 13 300 $w=1.7e-07 $l=3.26994e-07 $layer=licon1_PDIFF $count=2 $X=1.335
+ $Y=2.12 $X2=1.555 $Y2=2.355
r50 1 9 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.37
+ $Y=2.12 $X2=0.515 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_1%X 1 2 10 13 14 15 30 34
r22 32 34 0.583515 $w=3.93e-07 $l=2e-08 $layer=LI1_cond $X=2.117 $Y=2.015
+ $X2=2.117 $Y2=2.035
r23 20 34 0.350109 $w=3.93e-07 $l=1.2e-08 $layer=LI1_cond $X=2.117 $Y=2.047
+ $X2=2.117 $Y2=2.035
r24 15 27 1.16703 $w=3.93e-07 $l=4e-08 $layer=LI1_cond $X=2.117 $Y=2.775
+ $X2=2.117 $Y2=2.815
r25 14 15 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.117 $Y=2.405
+ $X2=2.117 $Y2=2.775
r26 13 32 0.495988 $w=3.93e-07 $l=1.7e-08 $layer=LI1_cond $X=2.117 $Y=1.998
+ $X2=2.117 $Y2=2.015
r27 13 30 8.13121 $w=3.93e-07 $l=1.48e-07 $layer=LI1_cond $X=2.117 $Y=1.998
+ $X2=2.117 $Y2=1.85
r28 13 14 9.3946 $w=3.93e-07 $l=3.22e-07 $layer=LI1_cond $X=2.117 $Y=2.083
+ $X2=2.117 $Y2=2.405
r29 13 20 1.05033 $w=3.93e-07 $l=3.6e-08 $layer=LI1_cond $X=2.117 $Y=2.083
+ $X2=2.117 $Y2=2.047
r30 12 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.23 $Y=1.18
+ $X2=2.23 $Y2=1.85
r31 10 12 18.6836 $w=4.73e-07 $l=5.35e-07 $layer=LI1_cond $X=2.077 $Y=0.645
+ $X2=2.077 $Y2=1.18
r32 2 32 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.84 $X2=2.005 $Y2=2.015
r33 2 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.84 $X2=2.005 $Y2=2.815
r34 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.5 $X2=2.005 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_1%VGND 1 6 9 10 11 21 22
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 14 18 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r28 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r30 11 15 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r31 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 9 18 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.34 $Y=0 $X2=1.2
+ $Y2=0
r33 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=0 $X2=1.505
+ $Y2=0
r34 8 21 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=2.16
+ $Y2=0
r35 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.505
+ $Y2=0
r36 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=0.085
+ $X2=1.505 $Y2=0
r37 4 6 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.505 $Y=0.085
+ $X2=1.505 $Y2=0.845
r38 1 6 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=1.285
+ $Y=0.6 $X2=1.505 $Y2=0.845
.ends


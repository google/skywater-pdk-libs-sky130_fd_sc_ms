# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a32oi_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__a32oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.805000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.735000 1.350000 8.515000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.350000 10.435000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 4.195000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.252600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.950000 6.350000 2.120000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.515000 2.120000 1.845000 2.735000 ;
        RECT 2.400000 0.595000 2.730000 0.880000 ;
        RECT 2.400000 0.880000 3.660000 1.010000 ;
        RECT 2.400000 1.010000 6.350000 1.130000 ;
        RECT 2.400000 1.130000 5.150000 1.180000 ;
        RECT 2.515000 2.120000 2.845000 2.735000 ;
        RECT 3.515000 2.120000 3.845000 2.735000 ;
        RECT 4.820000 0.770000 6.350000 1.010000 ;
        RECT 6.180000 1.130000 6.350000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 10.560000 0.085000 ;
        RECT  0.615000  0.085000  0.945000 0.840000 ;
        RECT  1.475000  0.085000  1.805000 0.840000 ;
        RECT  8.395000  0.085000  8.725000 0.840000 ;
        RECT  9.255000  0.085000  9.585000 0.840000 ;
        RECT 10.115000  0.085000 10.445000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.560000 3.415000 ;
        RECT 4.605000 2.630000  4.935000 3.245000 ;
        RECT 5.605000 2.630000  5.935000 3.245000 ;
        RECT 6.605000 2.630000  6.935000 3.245000 ;
        RECT 7.605000 2.290000  7.935000 3.245000 ;
        RECT 8.605000 2.290000  8.935000 3.245000 ;
        RECT 9.605000 2.290000  9.935000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.350000  0.445000 1.010000 ;
      RECT  0.115000 1.010000  2.220000 1.180000 ;
      RECT  0.115000 1.950000  0.445000 2.905000 ;
      RECT  0.115000 2.905000  4.345000 3.075000 ;
      RECT  1.125000 0.350000  1.295000 1.010000 ;
      RECT  1.145000 2.290000  1.315000 2.905000 ;
      RECT  2.015000 2.290000  2.345000 2.905000 ;
      RECT  2.050000 0.255000  4.090000 0.425000 ;
      RECT  2.050000 0.425000  2.220000 1.010000 ;
      RECT  2.900000 0.425000  3.230000 0.710000 ;
      RECT  3.015000 2.290000  3.345000 2.905000 ;
      RECT  3.760000 0.425000  4.090000 0.710000 ;
      RECT  4.015000 2.290000  7.435000 2.460000 ;
      RECT  4.015000 2.460000  4.345000 2.905000 ;
      RECT  4.320000 0.350000  8.165000 0.600000 ;
      RECT  4.320000 0.600000  4.650000 0.840000 ;
      RECT  5.105000 2.460000  5.435000 2.980000 ;
      RECT  6.105000 2.460000  6.435000 2.980000 ;
      RECT  6.540000 0.770000  6.870000 0.850000 ;
      RECT  6.540000 0.850000  7.735000 1.010000 ;
      RECT  6.540000 1.010000  9.935000 1.180000 ;
      RECT  7.105000 1.950000 10.440000 2.120000 ;
      RECT  7.105000 2.120000  7.435000 2.290000 ;
      RECT  7.105000 2.460000  7.435000 2.980000 ;
      RECT  7.835000 0.600000  8.165000 0.680000 ;
      RECT  8.105000 2.120000  8.435000 2.980000 ;
      RECT  8.905000 0.350000  9.075000 1.010000 ;
      RECT  9.105000 2.120000  9.435000 2.980000 ;
      RECT  9.765000 0.350000  9.935000 1.010000 ;
      RECT 10.110000 2.120000 10.440000 2.980000 ;
  END
END sky130_fd_sc_ms__a32oi_4

* File: sky130_fd_sc_ms__o21ba_2.pex.spice
* Created: Fri Aug 28 17:55:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21BA_2%B1_N 3 7 9 13 16
c28 7 0 1.06953e-19 $X=0.505 $Y=2.26
c29 3 0 5.63373e-20 $X=0.485 $Y=0.645
r30 15 16 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.485 $Y=1.465
+ $X2=0.505 $Y2=1.465
r31 12 15 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.485 $Y2=1.465
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r33 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r34 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r35 5 7 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.26
r36 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.3
+ $X2=0.485 $Y2=1.465
r37 1 3 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.485 $Y=1.3
+ $X2=0.485 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%A_177_48# 1 2 9 13 17 21 23 27 33 35 40 43
+ 44 49
c102 40 0 1.9148e-19 $X=2.465 $Y=1.095
r103 48 49 18.4097 $w=2.88e-07 $l=1.1e-07 $layer=POLY_cond $X=1.39 $Y=1.465
+ $X2=1.5 $Y2=1.465
r104 43 45 12.7457 $w=3.93e-07 $l=4.25e-07 $layer=LI1_cond $X=2.577 $Y=1.985
+ $X2=2.577 $Y2=2.41
r105 43 44 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.577 $Y=1.985
+ $X2=2.577 $Y2=1.82
r106 38 49 2.51042 $w=2.88e-07 $l=1.5e-08 $layer=POLY_cond $X=1.515 $Y=1.465
+ $X2=1.5 $Y2=1.465
r107 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=1.465 $X2=1.515 $Y2=1.465
r108 35 37 17.702 $w=2.55e-07 $l=3.7e-07 $layer=LI1_cond $X=1.515 $Y=1.095
+ $X2=1.515 $Y2=1.465
r109 33 45 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.61 $Y=2.695
+ $X2=2.61 $Y2=2.41
r110 29 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.18
+ $X2=2.465 $Y2=1.095
r111 29 44 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.465 $Y=1.18
+ $X2=2.465 $Y2=1.82
r112 25 40 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.105 $Y=1.095
+ $X2=2.465 $Y2=1.095
r113 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.105 $Y=1.01
+ $X2=2.105 $Y2=0.515
r114 24 35 3.11056 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.095
+ $X2=1.515 $Y2=1.095
r115 23 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.98 $Y=1.095
+ $X2=2.105 $Y2=1.095
r116 23 24 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=1.095
+ $X2=1.68 $Y2=1.095
r117 19 49 13.7767 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.63
+ $X2=1.5 $Y2=1.465
r118 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.5 $Y=1.63 $X2=1.5
+ $Y2=2.4
r119 15 48 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=1.465
r120 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=0.74
r121 11 48 56.9028 $w=2.88e-07 $l=3.4e-07 $layer=POLY_cond $X=1.05 $Y=1.465
+ $X2=1.39 $Y2=1.465
r122 11 13 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=1.05 $Y=1.6 $X2=1.05
+ $Y2=2.4
r123 7 11 15.0625 $w=2.88e-07 $l=9e-08 $layer=POLY_cond $X=0.96 $Y=1.465
+ $X2=1.05 $Y2=1.465
r124 7 9 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.96 $Y=1.345
+ $X2=0.96 $Y2=0.74
r125 2 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.84 $X2=2.61 $Y2=1.985
r126 2 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.84 $X2=2.61 $Y2=2.695
r127 1 27 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.37 $X2=2.145 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%A_27_74# 1 2 9 13 15 16 19 21 22 24 25 29 33
c88 16 0 1.9148e-19 $X=2.38 $Y=1.515
c89 9 0 2.05372e-19 $X=2.36 $Y=0.74
r90 33 34 4.70956 $w=5.44e-07 $l=2.1e-07 $layer=LI1_cond $X=0.455 $Y=2.115
+ $X2=0.455 $Y2=2.325
r91 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.515 $X2=2.055 $Y2=1.515
r92 27 29 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=2.05 $Y=2.24 $X2=2.05
+ $Y2=1.515
r93 26 34 7.68949 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=0.795 $Y=2.325
+ $X2=0.455 $Y2=2.325
r94 25 27 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.89 $Y=2.325
+ $X2=2.05 $Y2=2.24
r95 25 26 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=1.89 $Y=2.325
+ $X2=0.795 $Y2=2.325
r96 24 33 9.98939 $w=5.44e-07 $l=3.27261e-07 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.455 $Y2=2.115
r97 23 24 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r98 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.71 $Y2=1.13
r99 21 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.355 $Y2=1.045
r100 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=0.96
+ $X2=0.355 $Y2=1.045
r101 17 19 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.23 $Y=0.96
+ $X2=0.23 $Y2=0.645
r102 15 30 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.055 $Y2=1.515
r103 15 16 3.90195 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.38 $Y2=1.515
r104 11 16 34.7346 $w=1.65e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.385 $Y=1.68
+ $X2=2.38 $Y2=1.515
r105 11 13 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.385 $Y=1.68
+ $X2=2.385 $Y2=2.34
r106 7 16 34.7346 $w=1.65e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.36 $Y=1.35
+ $X2=2.38 $Y2=1.515
r107 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.36 $Y=1.35 $X2=2.36
+ $Y2=0.74
r108 2 33 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r109 1 19 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.27 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%A2 3 6 8 11 13
c35 13 0 2.53695e-20 $X=2.88 $Y=1.22
c36 8 0 1.75261e-19 $X=3.12 $Y=1.295
r37 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.385
+ $X2=2.88 $Y2=1.55
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.385
+ $X2=2.88 $Y2=1.22
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.385 $X2=2.88 $Y2=1.385
r40 8 12 7.47531 $w=3.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.88 $Y2=1.365
r41 6 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.835 $Y=2.34
+ $X2=2.835 $Y2=1.55
r42 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.79 $Y=0.74 $X2=2.79
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%A1 1 3 5 7 8
c25 8 0 2.53695e-20 $X=3.6 $Y=1.295
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.385 $X2=3.57 $Y2=1.385
r27 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.57 $Y=1.295 $X2=3.57
+ $Y2=1.385
r28 5 11 39.4323 $w=3.92e-07 $l=2.22486e-07 $layer=POLY_cond $X=3.36 $Y=1.22
+ $X2=3.495 $Y2=1.385
r29 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.36 $Y=1.22 $X2=3.36
+ $Y2=0.74
r30 1 11 45.5886 $w=3.92e-07 $l=3.21364e-07 $layer=POLY_cond $X=3.345 $Y=1.64
+ $X2=3.495 $Y2=1.385
r31 1 3 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=3.345 $Y=1.64 $X2=3.345
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%VPWR 1 2 3 14 16 18 22 24 29 35 38 48
r45 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 41 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 38 41 10.9789 $w=6.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.9 $Y=2.715
+ $X2=1.9 $Y2=3.33
r49 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 33 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 33 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 30 41 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=1.9 $Y2=3.33
r54 30 32 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 29 47 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.622 $Y2=3.33
r56 29 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r61 25 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 24 41 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.9 $Y2=3.33
r63 24 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 22 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.57 $Y=1.985
+ $X2=3.57 $Y2=2.695
r67 16 47 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.622 $Y2=3.33
r68 16 21 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.695
r69 12 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r70 12 14 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.745
r71 3 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.84 $X2=3.57 $Y2=2.695
r72 3 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.84 $X2=3.57 $Y2=1.985
r73 2 38 300 $w=1.7e-07 $l=1.08886e-06 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.84 $X2=2.07 $Y2=2.715
r74 1 14 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%X 1 2 8 12 14 15 26
c35 15 0 5.63373e-20 $X=1.115 $Y=0.84
c36 12 0 1.06953e-19 $X=1.275 $Y=1.985
r37 19 26 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.175 $Y=0.965
+ $X2=1.175 $Y2=0.925
r38 15 28 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=1.175 $Y=0.987
+ $X2=1.175 $Y2=1.13
r39 15 19 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=1.175 $Y=0.987
+ $X2=1.175 $Y2=0.965
r40 15 26 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=1.175 $Y=0.902
+ $X2=1.175 $Y2=0.925
r41 14 15 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=1.175 $Y=0.515
+ $X2=1.175 $Y2=0.902
r42 9 12 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.095 $Y=1.945
+ $X2=1.275 $Y2=1.945
r43 8 9 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.82
+ $X2=1.095 $Y2=1.945
r44 8 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.82
+ $X2=1.095 $Y2=1.13
r45 2 12 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.84 $X2=1.275 $Y2=1.985
r46 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%VGND 1 2 3 12 16 20 23 24 25 31 35 42 43 46
+ 49
r56 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 43 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r59 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.075
+ $Y2=0
r61 40 42 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.6
+ $Y2=0
r62 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r63 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 36 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.645
+ $Y2=0
r65 36 38 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.64
+ $Y2=0
r66 35 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.075
+ $Y2=0
r67 35 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.64
+ $Y2=0
r68 34 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r69 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r70 31 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.645
+ $Y2=0
r71 31 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.2
+ $Y2=0
r72 29 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r73 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 25 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r75 25 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r76 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r77 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.66
+ $Y2=0
r78 22 33 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=1.2
+ $Y2=0
r79 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.66
+ $Y2=0
r80 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0
r81 18 20 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0.335
r82 14 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r83 14 16 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.64
r84 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=0.085
+ $X2=0.66 $Y2=0
r85 10 12 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=0.66 $Y=0.085
+ $X2=0.66 $Y2=0.61
r86 3 20 182 $w=1.7e-07 $l=2.26826e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.37 $X2=3.075 $Y2=0.335
r87 2 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.64
r88 1 12 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.37 $X2=0.7 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_2%A_487_74# 1 2 7 10 15
c28 7 0 3.01108e-20 $X=3.41 $Y=0.755
r29 15 17 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.575 $Y=0.515
+ $X2=3.575 $Y2=0.755
r30 10 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.575 $Y=0.595
+ $X2=2.575 $Y2=0.755
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=0.755
+ $X2=2.575 $Y2=0.755
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=0.755
+ $X2=3.575 $Y2=0.755
r33 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.41 $Y=0.755 $X2=2.74
+ $Y2=0.755
r34 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.37 $X2=3.575 $Y2=0.515
r35 1 10 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.37 $X2=2.575 $Y2=0.595
.ends


* File: sky130_fd_sc_ms__o21ai_4.pxi.spice
* Created: Fri Aug 28 17:55:09 2020
* 
x_PM_SKY130_FD_SC_MS__O21AI_4%A1 N_A1_M1004_g N_A1_M1009_g N_A1_M1018_g
+ N_A1_M1005_g N_A1_M1019_g N_A1_M1006_g N_A1_M1021_g N_A1_M1007_g A1 A1
+ N_A1_c_105_n N_A1_c_134_p PM_SKY130_FD_SC_MS__O21AI_4%A1
x_PM_SKY130_FD_SC_MS__O21AI_4%B1 N_B1_c_185_n N_B1_M1002_g N_B1_M1011_g
+ N_B1_c_187_n N_B1_M1003_g N_B1_M1012_g N_B1_c_189_n N_B1_M1010_g N_B1_c_190_n
+ N_B1_c_191_n N_B1_M1017_g B1 B1 N_B1_c_192_n N_B1_c_193_n
+ PM_SKY130_FD_SC_MS__O21AI_4%B1
x_PM_SKY130_FD_SC_MS__O21AI_4%A2 N_A2_c_263_n N_A2_M1013_g N_A2_M1000_g
+ N_A2_c_264_n N_A2_M1014_g N_A2_M1001_g N_A2_c_265_n N_A2_M1015_g N_A2_M1008_g
+ N_A2_c_266_n N_A2_M1020_g N_A2_M1016_g A2 A2 A2 A2 N_A2_c_262_n
+ PM_SKY130_FD_SC_MS__O21AI_4%A2
x_PM_SKY130_FD_SC_MS__O21AI_4%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1007_s
+ N_VPWR_M1012_s N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n VPWR N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_335_n N_VPWR_c_347_n N_VPWR_c_348_n
+ PM_SKY130_FD_SC_MS__O21AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O21AI_4%A_119_368# N_A_119_368#_M1004_d
+ N_A_119_368#_M1006_d N_A_119_368#_M1013_d N_A_119_368#_M1014_d
+ N_A_119_368#_M1020_d N_A_119_368#_c_404_n N_A_119_368#_c_405_n
+ N_A_119_368#_c_423_n N_A_119_368#_c_428_n N_A_119_368#_c_432_n
+ N_A_119_368#_c_406_n N_A_119_368#_c_407_n N_A_119_368#_c_408_n
+ N_A_119_368#_c_409_n N_A_119_368#_c_410_n N_A_119_368#_c_411_n
+ N_A_119_368#_c_487_p N_A_119_368#_c_412_n N_A_119_368#_c_413_n
+ N_A_119_368#_c_438_n N_A_119_368#_c_414_n
+ PM_SKY130_FD_SC_MS__O21AI_4%A_119_368#
x_PM_SKY130_FD_SC_MS__O21AI_4%Y N_Y_M1002_d N_Y_M1010_d N_Y_M1011_d N_Y_M1013_s
+ N_Y_M1015_s N_Y_c_495_n N_Y_c_503_n N_Y_c_519_n N_Y_c_520_n N_Y_c_507_n
+ N_Y_c_510_n N_Y_c_524_n N_Y_c_528_n Y N_Y_c_494_n
+ PM_SKY130_FD_SC_MS__O21AI_4%Y
x_PM_SKY130_FD_SC_MS__O21AI_4%A_27_74# N_A_27_74#_M1009_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1021_s N_A_27_74#_M1003_s N_A_27_74#_M1017_s N_A_27_74#_M1001_s
+ N_A_27_74#_M1016_s N_A_27_74#_c_563_n N_A_27_74#_c_564_n N_A_27_74#_c_565_n
+ N_A_27_74#_c_566_n N_A_27_74#_c_585_n N_A_27_74#_c_567_n N_A_27_74#_c_568_n
+ N_A_27_74#_c_569_n N_A_27_74#_c_598_n N_A_27_74#_c_570_n N_A_27_74#_c_571_n
+ N_A_27_74#_c_572_n N_A_27_74#_c_573_n N_A_27_74#_c_574_n N_A_27_74#_c_575_n
+ N_A_27_74#_c_576_n N_A_27_74#_c_577_n PM_SKY130_FD_SC_MS__O21AI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O21AI_4%VGND N_VGND_M1009_d N_VGND_M1019_d N_VGND_M1000_d
+ N_VGND_M1008_d N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ N_VGND_c_668_n VGND N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n
+ N_VGND_c_672_n N_VGND_c_673_n N_VGND_c_674_n N_VGND_c_675_n N_VGND_c_676_n
+ N_VGND_c_677_n PM_SKY130_FD_SC_MS__O21AI_4%VGND
cc_1 VNB N_A1_M1004_g 7.56802e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A1_M1009_g 0.0301354f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_A1_M1018_g 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_A1_M1005_g 4.76178e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_5 VNB N_A1_M1019_g 0.0217592f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_6 VNB N_A1_M1006_g 4.03451e-19 $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_7 VNB N_A1_M1021_g 0.0222874f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_8 VNB N_A1_M1007_g 4.57629e-19 $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_9 VNB N_A1_c_105_n 0.095325f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.485
cc_10 VNB N_B1_c_185_n 0.0144853f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_11 VNB N_B1_M1011_g 0.00599169f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_12 VNB N_B1_c_187_n 0.0143176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1012_g 0.00705436f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.65
cc_14 VNB N_B1_c_189_n 0.0142846f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_15 VNB N_B1_c_190_n 0.0246434f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_16 VNB N_B1_c_191_n 0.0143551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_192_n 0.0170818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_193_n 0.0696617f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_19 VNB N_A2_M1000_g 0.0233837f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_A2_M1001_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.65
cc_21 VNB N_A2_M1008_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_M1016_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_23 VNB A2 0.0166485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_262_n 0.0782675f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.485
cc_25 VNB N_VPWR_c_335_n 0.243291f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.485
cc_26 VNB Y 0.00850576f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.485
cc_27 VNB N_Y_c_494_n 0.00427957f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.485
cc_28 VNB N_A_27_74#_c_563_n 0.0255089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_564_n 0.00456647f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_30 VNB N_A_27_74#_c_565_n 0.0115038f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_31 VNB N_A_27_74#_c_566_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_32 VNB N_A_27_74#_c_567_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_33 VNB N_A_27_74#_c_568_n 0.00213254f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_34 VNB N_A_27_74#_c_569_n 0.00477762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_570_n 0.00337922f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.485
cc_36 VNB N_A_27_74#_c_571_n 0.00405692f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.485
cc_37 VNB N_A_27_74#_c_572_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.485
cc_38 VNB N_A_27_74#_c_573_n 0.0132288f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.485
cc_39 VNB N_A_27_74#_c_574_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.485
cc_40 VNB N_A_27_74#_c_575_n 0.00167779f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.55
cc_41 VNB N_A_27_74#_c_576_n 0.00202117f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.55
cc_42 VNB N_A_27_74#_c_577_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_664_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_44 VNB N_VGND_c_665_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_45 VNB N_VGND_c_666_n 0.0539351f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.65
cc_46 VNB N_VGND_c_667_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.32
cc_47 VNB N_VGND_c_668_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.65
cc_48 VNB N_VGND_c_669_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.485
cc_49 VNB N_VGND_c_670_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_50 VNB N_VGND_c_671_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_672_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.485
cc_52 VNB N_VGND_c_673_n 0.31955f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.485
cc_53 VNB N_VGND_c_674_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.485
cc_54 VNB N_VGND_c_675_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.485
cc_55 VNB N_VGND_c_676_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.55
cc_56 VNB N_VGND_c_677_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.55
cc_57 VPB N_A1_M1004_g 0.0280872f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_58 VPB N_A1_M1005_g 0.0223011f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_59 VPB N_A1_M1006_g 0.0214382f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_60 VPB N_A1_M1007_g 0.022493f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_61 VPB A1 0.00595134f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_62 VPB N_B1_M1011_g 0.0220746f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_63 VPB N_B1_M1012_g 0.0251845f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.65
cc_64 VPB N_A2_c_263_n 0.0210764f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_65 VPB N_A2_c_264_n 0.0181093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A2_c_265_n 0.0176212f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_67 VPB N_A2_c_266_n 0.0225686f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_68 VPB A2 0.0177343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A2_c_262_n 0.0235132f $X=-0.19 $Y=1.66 $X2=1.29 $Y2=1.485
cc_70 VPB N_VPWR_c_336_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.65
cc_71 VPB N_VPWR_c_337_n 0.0587237f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_72 VPB N_VPWR_c_338_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.65
cc_73 VPB N_VPWR_c_339_n 0.00498113f $X=-0.19 $Y=1.66 $X2=1.8 $Y2=1.32
cc_74 VPB N_VPWR_c_340_n 0.012174f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.65
cc_75 VPB N_VPWR_c_341_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_342_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.485
cc_77 VPB N_VPWR_c_343_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_344_n 0.0206218f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.485
cc_79 VPB N_VPWR_c_345_n 0.061582f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.485
cc_80 VPB N_VPWR_c_335_n 0.0910135f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.485
cc_81 VPB N_VPWR_c_347_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_348_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.55
cc_83 VPB N_A_119_368#_c_404_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_119_368#_c_405_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_85 VPB N_A_119_368#_c_406_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.8 $Y2=0.74
cc_86 VPB N_A_119_368#_c_407_n 0.0118988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_119_368#_c_408_n 3.13193e-19 $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_88 VPB N_A_119_368#_c_409_n 0.00522274f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_89 VPB N_A_119_368#_c_410_n 0.00262732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_119_368#_c_411_n 0.00418606f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.485
cc_91 VPB N_A_119_368#_c_412_n 0.0119149f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_92 VPB N_A_119_368#_c_413_n 0.0351758f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.485
cc_93 VPB N_A_119_368#_c_414_n 0.00123754f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.485
cc_94 VPB N_Y_c_495_n 0.0106719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB Y 0.00932227f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.485
cc_96 N_A1_M1021_g N_B1_c_185_n 0.0181168f $X=1.8 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_97 A1 N_B1_M1011_g 0.00107565f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A1_c_105_n N_B1_M1011_g 0.0570771f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_99 N_A1_M1021_g N_B1_c_192_n 0.00382458f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_100 A1 N_B1_c_192_n 0.0151989f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A1_c_105_n N_B1_c_192_n 0.00213182f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_102 N_A1_c_105_n N_B1_c_193_n 0.0151767f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_103 N_A1_M1004_g N_VPWR_c_337_n 0.00649184f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A1_M1005_g N_VPWR_c_338_n 0.0027763f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A1_M1006_g N_VPWR_c_338_n 0.0027763f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A1_M1007_g N_VPWR_c_339_n 0.002979f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A1_M1004_g N_VPWR_c_341_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A1_M1005_g N_VPWR_c_341_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A1_M1006_g N_VPWR_c_343_n 0.005209f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A1_M1007_g N_VPWR_c_343_n 0.005209f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A1_M1004_g N_VPWR_c_335_n 0.00986008f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A1_M1005_g N_VPWR_c_335_n 0.00982266f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A1_M1006_g N_VPWR_c_335_n 0.00982266f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A1_M1007_g N_VPWR_c_335_n 0.00982376f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A1_M1004_g N_A_119_368#_c_404_n 0.00442661f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A1_M1005_g N_A_119_368#_c_404_n 0.00361305f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A1_M1006_g N_A_119_368#_c_404_n 6.1989e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A1_c_105_n N_A_119_368#_c_404_n 0.00215577f $X=1.855 $Y=1.485 $X2=0
+ $Y2=0
cc_119 N_A1_c_134_p N_A_119_368#_c_404_n 0.0275631f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_120 N_A1_M1004_g N_A_119_368#_c_405_n 0.0118478f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A1_M1005_g N_A_119_368#_c_405_n 0.0125215f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A1_M1006_g N_A_119_368#_c_405_n 6.50516e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A1_M1005_g N_A_119_368#_c_423_n 0.0136654f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A1_M1006_g N_A_119_368#_c_423_n 0.012931f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_125 A1 N_A_119_368#_c_423_n 0.0267057f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A1_c_105_n N_A_119_368#_c_423_n 4.56682e-19 $X=1.855 $Y=1.485 $X2=0
+ $Y2=0
cc_127 N_A1_c_134_p N_A_119_368#_c_423_n 0.00770917f $X=1.085 $Y=1.55 $X2=0
+ $Y2=0
cc_128 N_A1_M1006_g N_A_119_368#_c_428_n 8.84614e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A1_M1007_g N_A_119_368#_c_428_n 0.00366667f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_130 A1 N_A_119_368#_c_428_n 0.0236942f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A1_c_105_n N_A_119_368#_c_428_n 5.1677e-19 $X=1.855 $Y=1.485 $X2=0
+ $Y2=0
cc_132 N_A1_M1005_g N_A_119_368#_c_432_n 4.31538e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A1_M1006_g N_A_119_368#_c_432_n 0.00321805f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A1_M1007_g N_A_119_368#_c_432_n 0.00320621f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A1_M1006_g N_A_119_368#_c_406_n 0.00667044f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A1_M1007_g N_A_119_368#_c_406_n 0.00788893f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A1_M1007_g N_A_119_368#_c_407_n 0.0172079f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A1_M1006_g N_A_119_368#_c_438_n 0.0020266f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A1_M1007_g N_A_119_368#_c_438_n 4.64231e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A1_M1007_g N_Y_c_495_n 0.00110035f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A1_M1009_g N_A_27_74#_c_563_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A1_M1009_g N_A_27_74#_c_564_n 0.0137615f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1018_g N_A_27_74#_c_564_n 0.0124568f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_c_105_n N_A_27_74#_c_564_n 0.00254808f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_145 N_A1_c_134_p N_A_27_74#_c_564_n 0.0448197f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_146 N_A1_M1018_g N_A_27_74#_c_566_n 3.92313e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A1_M1019_g N_A_27_74#_c_566_n 3.92313e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A1_M1019_g N_A_27_74#_c_585_n 0.0104439f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A1_M1021_g N_A_27_74#_c_585_n 0.0125823f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_150 A1 N_A_27_74#_c_585_n 0.0227309f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A1_c_105_n N_A_27_74#_c_585_n 0.00314046f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_152 N_A1_M1021_g N_A_27_74#_c_568_n 9.83948e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1019_g N_A_27_74#_c_575_n 9.34957e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_c_105_n N_A_27_74#_c_575_n 0.00250705f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_155 N_A1_c_134_p N_A_27_74#_c_575_n 0.0144048f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_156 N_A1_M1009_g N_VGND_c_664_n 0.0127296f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_M1018_g N_VGND_c_664_n 0.00970341f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A1_M1019_g N_VGND_c_664_n 4.62684e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A1_M1018_g N_VGND_c_665_n 4.20905e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_M1019_g N_VGND_c_665_n 0.00765209f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A1_M1021_g N_VGND_c_665_n 0.00617842f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A1_M1021_g N_VGND_c_666_n 0.00429299f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A1_M1009_g N_VGND_c_669_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_M1018_g N_VGND_c_670_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1019_g N_VGND_c_670_n 0.00383152f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1009_g N_VGND_c_673_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_M1018_g N_VGND_c_673_n 0.0075754f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_M1019_g N_VGND_c_673_n 0.00383967f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A1_M1021_g N_VGND_c_673_n 0.00429576f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B1_c_191_n N_A2_M1000_g 0.0164408f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_171 N_B1_M1011_g N_VPWR_c_339_n 0.0114971f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_172 N_B1_M1012_g N_VPWR_c_339_n 0.0013933f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B1_M1012_g N_VPWR_c_340_n 0.010463f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B1_M1011_g N_VPWR_c_344_n 0.00460063f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B1_M1012_g N_VPWR_c_344_n 0.00553757f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_176 N_B1_M1011_g N_VPWR_c_335_n 0.00908554f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_177 N_B1_M1012_g N_VPWR_c_335_n 0.010939f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B1_M1011_g N_A_119_368#_c_428_n 4.9654e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B1_M1011_g N_A_119_368#_c_432_n 8.03925e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_180 N_B1_M1011_g N_A_119_368#_c_406_n 8.83197e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_181 N_B1_M1011_g N_A_119_368#_c_407_n 0.0205784f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_182 N_B1_M1012_g N_A_119_368#_c_407_n 0.0190001f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_183 N_B1_M1012_g N_A_119_368#_c_409_n 0.00445711f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_184 N_B1_M1011_g N_Y_c_495_n 0.00705962f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_185 N_B1_M1012_g N_Y_c_495_n 0.0176688f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_186 N_B1_c_190_n N_Y_c_495_n 0.00492945f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_187 N_B1_c_192_n N_Y_c_495_n 0.04402f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_188 N_B1_c_193_n N_Y_c_495_n 0.00991009f $X=3.165 $Y=1.367 $X2=0 $Y2=0
cc_189 N_B1_c_187_n N_Y_c_503_n 0.00950771f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_190 N_B1_c_189_n N_Y_c_503_n 0.00950771f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_191 N_B1_c_192_n N_Y_c_503_n 0.0418422f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_192 N_B1_c_193_n N_Y_c_503_n 6.92962e-19 $X=3.165 $Y=1.367 $X2=0 $Y2=0
cc_193 N_B1_c_185_n N_Y_c_507_n 0.00516423f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_194 N_B1_c_192_n N_Y_c_507_n 0.0183113f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_195 N_B1_c_193_n N_Y_c_507_n 7.37755e-19 $X=3.165 $Y=1.367 $X2=0 $Y2=0
cc_196 N_B1_c_190_n N_Y_c_510_n 0.00304357f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_197 N_B1_c_191_n N_Y_c_510_n 0.00625443f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_198 N_B1_M1012_g Y 0.00814452f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_199 N_B1_c_190_n Y 0.0040411f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_200 N_B1_c_189_n N_Y_c_494_n 0.00351883f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_201 N_B1_c_190_n N_Y_c_494_n 0.0112144f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_202 N_B1_c_191_n N_Y_c_494_n 0.00324088f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B1_c_192_n N_Y_c_494_n 0.0288059f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_204 N_B1_c_193_n N_Y_c_494_n 0.00148844f $X=3.165 $Y=1.367 $X2=0 $Y2=0
cc_205 N_B1_c_192_n N_A_27_74#_c_585_n 0.00471836f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_206 N_B1_c_185_n N_A_27_74#_c_567_n 0.0120041f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_207 N_B1_c_187_n N_A_27_74#_c_567_n 0.00785166f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_208 N_B1_c_189_n N_A_27_74#_c_569_n 0.00785166f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_209 N_B1_c_191_n N_A_27_74#_c_569_n 0.0110523f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_210 N_B1_c_191_n N_A_27_74#_c_598_n 0.00271595f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_211 N_B1_c_191_n N_A_27_74#_c_571_n 9.24829e-19 $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_212 N_B1_c_185_n N_A_27_74#_c_576_n 6.25215e-19 $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_213 N_B1_c_187_n N_A_27_74#_c_576_n 0.00663416f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_214 N_B1_c_189_n N_A_27_74#_c_576_n 0.00669566f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_215 N_B1_c_191_n N_A_27_74#_c_576_n 6.30166e-19 $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B1_c_185_n N_VGND_c_666_n 0.00278271f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_217 N_B1_c_187_n N_VGND_c_666_n 0.00279469f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_218 N_B1_c_189_n N_VGND_c_666_n 0.00279469f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_219 N_B1_c_191_n N_VGND_c_666_n 0.00278271f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_220 N_B1_c_185_n N_VGND_c_673_n 0.00353526f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_221 N_B1_c_187_n N_VGND_c_673_n 0.00352518f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_222 N_B1_c_189_n N_VGND_c_673_n 0.00352518f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_223 N_B1_c_191_n N_VGND_c_673_n 0.00353754f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_224 N_A2_c_263_n N_VPWR_c_340_n 0.00136573f $X=3.85 $Y=1.725 $X2=0 $Y2=0
cc_225 N_A2_c_263_n N_VPWR_c_345_n 0.00333896f $X=3.85 $Y=1.725 $X2=0 $Y2=0
cc_226 N_A2_c_264_n N_VPWR_c_345_n 0.00333926f $X=4.35 $Y=1.725 $X2=0 $Y2=0
cc_227 N_A2_c_265_n N_VPWR_c_345_n 0.00333926f $X=4.8 $Y=1.725 $X2=0 $Y2=0
cc_228 N_A2_c_266_n N_VPWR_c_345_n 0.00333926f $X=5.25 $Y=1.725 $X2=0 $Y2=0
cc_229 N_A2_c_263_n N_VPWR_c_335_n 0.00428307f $X=3.85 $Y=1.725 $X2=0 $Y2=0
cc_230 N_A2_c_264_n N_VPWR_c_335_n 0.00423176f $X=4.35 $Y=1.725 $X2=0 $Y2=0
cc_231 N_A2_c_265_n N_VPWR_c_335_n 0.00422687f $X=4.8 $Y=1.725 $X2=0 $Y2=0
cc_232 N_A2_c_266_n N_VPWR_c_335_n 0.00426447f $X=5.25 $Y=1.725 $X2=0 $Y2=0
cc_233 N_A2_c_263_n N_A_119_368#_c_408_n 0.00234398f $X=3.85 $Y=1.725 $X2=0
+ $Y2=0
cc_234 N_A2_c_263_n N_A_119_368#_c_409_n 0.00643885f $X=3.85 $Y=1.725 $X2=0
+ $Y2=0
cc_235 N_A2_c_264_n N_A_119_368#_c_409_n 7.24402e-19 $X=4.35 $Y=1.725 $X2=0
+ $Y2=0
cc_236 N_A2_c_263_n N_A_119_368#_c_410_n 0.0119307f $X=3.85 $Y=1.725 $X2=0 $Y2=0
cc_237 N_A2_c_264_n N_A_119_368#_c_410_n 0.0143183f $X=4.35 $Y=1.725 $X2=0 $Y2=0
cc_238 N_A2_c_263_n N_A_119_368#_c_411_n 0.00291744f $X=3.85 $Y=1.725 $X2=0
+ $Y2=0
cc_239 N_A2_c_265_n N_A_119_368#_c_412_n 0.0140221f $X=4.8 $Y=1.725 $X2=0 $Y2=0
cc_240 N_A2_c_266_n N_A_119_368#_c_412_n 0.0149887f $X=5.25 $Y=1.725 $X2=0 $Y2=0
cc_241 A2 N_A_119_368#_c_413_n 0.0213263f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A2_c_263_n N_Y_c_519_n 0.0197647f $X=3.85 $Y=1.725 $X2=0 $Y2=0
cc_243 N_A2_c_264_n N_Y_c_520_n 0.012931f $X=4.35 $Y=1.725 $X2=0 $Y2=0
cc_244 N_A2_c_265_n N_Y_c_520_n 0.012931f $X=4.8 $Y=1.725 $X2=0 $Y2=0
cc_245 A2 N_Y_c_520_n 0.0391868f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_262_n N_Y_c_520_n 5.42978e-19 $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_247 N_A2_c_264_n N_Y_c_524_n 0.0105459f $X=4.35 $Y=1.725 $X2=0 $Y2=0
cc_248 N_A2_c_265_n N_Y_c_524_n 5.73047e-19 $X=4.8 $Y=1.725 $X2=0 $Y2=0
cc_249 A2 N_Y_c_524_n 0.024482f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_250 N_A2_c_262_n N_Y_c_524_n 9.5024e-19 $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_251 N_A2_c_264_n N_Y_c_528_n 5.73047e-19 $X=4.35 $Y=1.725 $X2=0 $Y2=0
cc_252 N_A2_c_265_n N_Y_c_528_n 0.010564f $X=4.8 $Y=1.725 $X2=0 $Y2=0
cc_253 N_A2_c_266_n N_Y_c_528_n 0.0114036f $X=5.25 $Y=1.725 $X2=0 $Y2=0
cc_254 A2 N_Y_c_528_n 0.0235494f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_255 N_A2_c_262_n N_Y_c_528_n 6.14241e-19 $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_256 A2 Y 0.0147816f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A2_c_262_n Y 0.0118f $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_258 N_A2_M1000_g N_Y_c_494_n 0.00579798f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_259 A2 N_Y_c_494_n 0.00747454f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_260 N_A2_M1000_g N_A_27_74#_c_569_n 9.86481e-19 $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_M1000_g N_A_27_74#_c_570_n 0.0149208f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1001_g N_A_27_74#_c_570_n 0.0130453f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_263 A2 N_A_27_74#_c_570_n 0.0428095f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A2_c_262_n N_A_27_74#_c_570_n 0.00432092f $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_265 N_A2_c_262_n N_A_27_74#_c_571_n 0.00324053f $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_266 N_A2_M1001_g N_A_27_74#_c_572_n 3.92313e-19 $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A2_M1008_g N_A_27_74#_c_572_n 3.92313e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A2_M1008_g N_A_27_74#_c_573_n 0.0130918f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A2_M1016_g N_A_27_74#_c_573_n 0.0136535f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_270 A2 N_A_27_74#_c_573_n 0.073609f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_271 N_A2_c_262_n N_A_27_74#_c_573_n 0.00240215f $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_272 N_A2_M1016_g N_A_27_74#_c_574_n 0.00159319f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_273 A2 N_A_27_74#_c_577_n 0.0146029f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_274 N_A2_c_262_n N_A_27_74#_c_577_n 0.00255673f $X=5.25 $Y=1.537 $X2=0 $Y2=0
cc_275 N_A2_M1000_g N_VGND_c_666_n 0.00383152f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A2_M1000_g N_VGND_c_667_n 0.00971294f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A2_M1001_g N_VGND_c_667_n 0.0103289f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A2_M1008_g N_VGND_c_667_n 4.71636e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A2_M1001_g N_VGND_c_668_n 4.71636e-19 $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A2_M1008_g N_VGND_c_668_n 0.0103289f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A2_M1016_g N_VGND_c_668_n 0.0133724f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A2_M1001_g N_VGND_c_671_n 0.00383152f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A2_M1008_g N_VGND_c_671_n 0.00383152f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A2_M1016_g N_VGND_c_672_n 0.00383152f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A2_M1000_g N_VGND_c_673_n 0.00757866f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A2_M1001_g N_VGND_c_673_n 0.0075754f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A2_M1008_g N_VGND_c_673_n 0.0075754f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A2_M1016_g N_VGND_c_673_n 0.00761198f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_289 N_VPWR_c_337_n N_A_119_368#_c_404_n 0.0112654f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_337_n N_A_119_368#_c_405_n 0.0289761f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_338_n N_A_119_368#_c_405_n 0.0233699f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_341_n N_A_119_368#_c_405_n 0.0144623f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_335_n N_A_119_368#_c_405_n 0.0118344f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_M1005_s N_A_119_368#_c_423_n 0.00315327f $X=1.045 $Y=1.84 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_338_n N_A_119_368#_c_423_n 0.0126919f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_338_n N_A_119_368#_c_406_n 0.0177362f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_339_n N_A_119_368#_c_406_n 0.0122069f $X=2.08 $Y=2.805 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_343_n N_A_119_368#_c_406_n 0.0144623f $X=1.995 $Y=3.33 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_335_n N_A_119_368#_c_406_n 0.0118344f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_M1007_s N_A_119_368#_c_407_n 0.00761058f $X=1.945 $Y=1.84 $X2=0
+ $Y2=0
cc_301 N_VPWR_M1012_s N_A_119_368#_c_407_n 0.00827647f $X=2.845 $Y=1.84 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_339_n N_A_119_368#_c_407_n 0.0148589f $X=2.08 $Y=2.805 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_340_n N_A_119_368#_c_407_n 0.0266632f $X=3.065 $Y=2.805 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_340_n N_A_119_368#_c_409_n 0.0185065f $X=3.065 $Y=2.805 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_345_n N_A_119_368#_c_410_n 0.0440768f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_335_n N_A_119_368#_c_410_n 0.0248093f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_340_n N_A_119_368#_c_411_n 0.0121618f $X=3.065 $Y=2.805 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_345_n N_A_119_368#_c_411_n 0.0235512f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_335_n N_A_119_368#_c_411_n 0.0126924f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_345_n N_A_119_368#_c_412_n 0.0638408f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_335_n N_A_119_368#_c_412_n 0.0355196f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_345_n N_A_119_368#_c_414_n 0.0121867f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_335_n N_A_119_368#_c_414_n 0.00660921f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_M1012_s N_Y_c_495_n 0.0061969f $X=2.845 $Y=1.84 $X2=0 $Y2=0
cc_315 N_VPWR_c_337_n N_A_27_74#_c_565_n 0.00886035f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_119_368#_c_407_n N_Y_M1011_d 0.00761462f $X=3.46 $Y=2.375 $X2=0 $Y2=0
cc_317 N_A_119_368#_c_410_n N_Y_M1013_s 0.00218982f $X=4.49 $Y=2.99 $X2=0 $Y2=0
cc_318 N_A_119_368#_c_412_n N_Y_M1015_s 0.00165831f $X=5.39 $Y=2.99 $X2=0 $Y2=0
cc_319 N_A_119_368#_c_428_n N_Y_c_495_n 0.00524697f $X=1.63 $Y=2.12 $X2=0 $Y2=0
cc_320 N_A_119_368#_c_407_n N_Y_c_495_n 0.0598415f $X=3.46 $Y=2.375 $X2=0 $Y2=0
cc_321 N_A_119_368#_c_408_n N_Y_c_519_n 0.00224313f $X=3.625 $Y=2.46 $X2=0 $Y2=0
cc_322 N_A_119_368#_M1014_d N_Y_c_520_n 0.00313001f $X=4.44 $Y=1.84 $X2=0 $Y2=0
cc_323 N_A_119_368#_c_487_p N_Y_c_520_n 0.0126919f $X=4.575 $Y=2.455 $X2=0 $Y2=0
cc_324 N_A_119_368#_c_410_n N_Y_c_524_n 0.0177084f $X=4.49 $Y=2.99 $X2=0 $Y2=0
cc_325 N_A_119_368#_c_412_n N_Y_c_528_n 0.0159318f $X=5.39 $Y=2.99 $X2=0 $Y2=0
cc_326 N_A_119_368#_M1013_d Y 0.00400582f $X=3.48 $Y=1.84 $X2=0 $Y2=0
cc_327 N_A_119_368#_c_407_n Y 0.0104353f $X=3.46 $Y=2.375 $X2=0 $Y2=0
cc_328 N_A_119_368#_c_408_n Y 0.0217495f $X=3.625 $Y=2.46 $X2=0 $Y2=0
cc_329 N_Y_c_503_n N_A_27_74#_M1003_s 0.00328233f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_330 N_Y_M1002_d N_A_27_74#_c_567_n 0.00176461f $X=2.305 $Y=0.37 $X2=0 $Y2=0
cc_331 N_Y_c_503_n N_A_27_74#_c_567_n 0.0035136f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_332 N_Y_c_507_n N_A_27_74#_c_567_n 0.0138155f $X=2.445 $Y=0.8 $X2=0 $Y2=0
cc_333 N_Y_M1010_d N_A_27_74#_c_569_n 0.00176461f $X=3.165 $Y=0.37 $X2=0 $Y2=0
cc_334 N_Y_c_503_n N_A_27_74#_c_569_n 0.0035136f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_335 N_Y_c_510_n N_A_27_74#_c_569_n 0.0165223f $X=3.305 $Y=0.8 $X2=0 $Y2=0
cc_336 N_Y_c_510_n N_A_27_74#_c_598_n 0.03026f $X=3.305 $Y=0.8 $X2=0 $Y2=0
cc_337 Y N_A_27_74#_c_571_n 0.0020972f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_338 N_Y_c_494_n N_A_27_74#_c_571_n 0.0135061f $X=3.525 $Y=1.55 $X2=0 $Y2=0
cc_339 N_Y_c_503_n N_A_27_74#_c_576_n 0.0160355f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_340 N_Y_c_503_n N_VGND_c_673_n 0.00146755f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_564_n N_VGND_M1009_d 0.00176461f $X=1.055 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_342 N_A_27_74#_c_585_n N_VGND_M1019_d 0.00412925f $X=1.93 $Y=0.925 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_570_n N_VGND_M1000_d 0.00176461f $X=4.535 $Y=1.095 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_573_n N_VGND_M1008_d 0.00176461f $X=5.395 $Y=1.095 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_563_n N_VGND_c_664_n 0.017215f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_346 N_A_27_74#_c_564_n N_VGND_c_664_n 0.0170777f $X=1.055 $Y=1.065 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_566_n N_VGND_c_664_n 0.0171736f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_348 N_A_27_74#_c_566_n N_VGND_c_665_n 0.0121558f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_349 N_A_27_74#_c_585_n N_VGND_c_665_n 0.0167779f $X=1.93 $Y=0.925 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_568_n N_VGND_c_665_n 0.010561f $X=2.1 $Y=0.34 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_567_n N_VGND_c_666_n 0.0384655f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_568_n N_VGND_c_666_n 0.0121867f $X=2.1 $Y=0.34 $X2=0 $Y2=0
cc_353 N_A_27_74#_c_569_n N_VGND_c_666_n 0.0522627f $X=3.675 $Y=0.34 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_576_n N_VGND_c_666_n 0.0225055f $X=2.875 $Y=0.34 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_569_n N_VGND_c_667_n 0.0112234f $X=3.675 $Y=0.34 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_570_n N_VGND_c_667_n 0.0171619f $X=4.535 $Y=1.095 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_572_n N_VGND_c_667_n 0.0182488f $X=4.62 $Y=0.515 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_572_n N_VGND_c_668_n 0.0182488f $X=4.62 $Y=0.515 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_573_n N_VGND_c_668_n 0.0171619f $X=5.395 $Y=1.095 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_574_n N_VGND_c_668_n 0.0182902f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_563_n N_VGND_c_669_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_566_n N_VGND_c_670_n 0.00749631f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_572_n N_VGND_c_671_n 0.00749631f $X=4.62 $Y=0.515 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_574_n N_VGND_c_672_n 0.011066f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_563_n N_VGND_c_673_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_566_n N_VGND_c_673_n 0.0062048f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_585_n N_VGND_c_673_n 0.0120697f $X=1.93 $Y=0.925 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_567_n N_VGND_c_673_n 0.0216792f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_568_n N_VGND_c_673_n 0.00660921f $X=2.1 $Y=0.34 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_569_n N_VGND_c_673_n 0.0292284f $X=3.675 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_572_n N_VGND_c_673_n 0.0062048f $X=4.62 $Y=0.515 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_574_n N_VGND_c_673_n 0.00915947f $X=5.48 $Y=0.515 $X2=0
+ $Y2=0
cc_373 N_A_27_74#_c_576_n N_VGND_c_673_n 0.0123739f $X=2.875 $Y=0.34 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o311a_4.spice
* Created: Wed Sep  2 12:25:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o311a_4.pex.spice"
.subckt sky130_fd_sc_ms__o311a_4  VNB VPB B1 C1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_83_244#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=5.664 M=1 R=4.93333 SA=75000.3
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1001_d N_A_83_244#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.20165 PD=1.02 PS=1.285 NRD=0 NRS=21.072 M=1 R=4.93333
+ SA=75000.7 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1014 N_X_M1014_d N_A_83_244#_M1014_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.20165 PD=1.09 PS=1.285 NRD=0 NRS=21.888 M=1 R=4.93333
+ SA=75001.4 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_X_M1014_d N_A_83_244#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_651_78#_M1007_d N_B1_M1007_g N_A_564_78#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2544 AS=0.178025 PD=1.435 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_83_244#_M1017_d N_C1_M1017_g N_A_651_78#_M1007_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.171975 AS=0.2544 PD=1.295 PS=1.435 NRD=40.068 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75004.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_83_244#_M1017_d N_C1_M1023_g N_A_651_78#_M1023_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.171975 AS=0.0896 PD=1.295 PS=0.92 NRD=40.068 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75003.6 A=0.096 P=1.58 MULT=1
MM1026 N_A_651_78#_M1023_s N_B1_M1026_g N_A_564_78#_M1026_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1216 PD=0.92 PS=1.02 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.2 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1021 N_A_564_78#_M1026_s N_A3_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.1232 PD=1.02 PS=1.025 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75002.7 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1024 N_A_564_78#_M1024_d N_A3_M1024_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0912 AS=0.1232 PD=0.925 PS=1.025 NRD=0.936 NRS=12.18 M=1 R=4.26667
+ SA=75003.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1015 N_A_564_78#_M1024_d N_A2_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0912 AS=0.12 PD=0.925 PS=1.015 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75003.7
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 N_A_564_78#_M1006_d N_A1_M1006_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.12 PD=1.02 PS=1.015 NRD=8.436 NRS=4.68 M=1 R=4.26667 SA=75004.2
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1027 N_A_564_78#_M1006_d N_A1_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.0944 PD=1.02 PS=0.935 NRD=10.308 NRS=2.808 M=1 R=4.26667
+ SA=75004.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1022 N_A_564_78#_M1022_d N_A2_M1022_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0944 PD=1.85 PS=0.935 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_X_M1009_d N_A_83_244#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004 A=0.2016 P=2.6 MULT=1
MM1010 N_X_M1009_d N_A_83_244#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1011_d N_A_83_244#_M1011_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2548 AS=0.1792 PD=1.575 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1018 N_X_M1011_d N_A_83_244#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2548 AS=0.187547 PD=1.575 PS=1.52679 NRD=22.852 NRS=0 M=1 R=6.22222
+ SA=90001.8 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1003 N_A_83_244#_M1003_d N_B1_M1003_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.167453 PD=1.39 PS=1.36321 NRD=0 NRS=9.8303 M=1 R=5.55556
+ SA=90002.3 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_A_83_244#_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.3425 AS=0.195 PD=1.685 PS=1.39 NRD=0 NRS=22.6353 M=1 R=5.55556 SA=90002.8
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1000_d N_C1_M1019_g N_A_83_244#_M1019_s VPB PSHORT L=0.18 W=1
+ AD=0.3425 AS=0.16 PD=1.685 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90003.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1020 N_A_83_244#_M1019_s N_B1_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90004.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_83_244#_M1008_d N_A3_M1008_g N_A_1034_392#_M1008_s VPB PSHORT L=0.18
+ W=1 AD=0.145 AS=0.43 PD=1.29 PS=2.86 NRD=0.9653 NRS=13.7703 M=1 R=5.55556
+ SA=90000.3 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1012 N_A_83_244#_M1008_d N_A3_M1012_g N_A_1034_392#_M1012_s VPB PSHORT L=0.18
+ W=1 AD=0.145 AS=0.1375 PD=1.29 PS=1.275 NRD=0.9653 NRS=0 M=1 R=5.55556
+ SA=90000.8 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_1341_392#_M1004_d N_A2_M1004_g N_A_1034_392#_M1012_s VPB PSHORT
+ L=0.18 W=1 AD=0.195 AS=0.1375 PD=1.39 PS=1.275 NRD=14.7553 NRS=0 M=1 R=5.55556
+ SA=90001.3 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_1341_392#_M1004_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.195 PD=1.27 PS=1.39 NRD=0 NRS=6.8753 M=1 R=5.55556 SA=90001.8
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1002_d N_A1_M1005_g N_A_1341_392#_M1005_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.3
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1016 N_A_1341_392#_M1005_s N_A2_M1016_g N_A_1034_392#_M1016_s VPB PSHORT
+ L=0.18 W=1 AD=0.145 AS=0.31 PD=1.29 PS=2.62 NRD=2.9353 NRS=4.9053 M=1
+ R=5.55556 SA=90002.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__o311a_4.pxi.spice"
*
.ends
*
*

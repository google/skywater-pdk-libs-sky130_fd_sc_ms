* File: sky130_fd_sc_ms__and4b_1.pex.spice
* Created: Fri Aug 28 17:13:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4B_1%A_N 3 7 11 12 13 16 17
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.43
+ $Y=1.355 $X2=0.43 $Y2=1.355
r40 13 17 3.39186 $w=6.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.525
+ $X2=0.43 $Y2=1.525
r41 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.43 $Y=1.695
+ $X2=0.43 $Y2=1.355
r42 11 12 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.695
+ $X2=0.43 $Y2=1.86
r43 10 16 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.19
+ $X2=0.43 $Y2=1.355
r44 7 10 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.495 $Y=0.645
+ $X2=0.495 $Y2=1.19
r45 3 12 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.505 $Y=2.54
+ $X2=0.505 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%A_27_74# 1 2 9 13 14 15 17 20 24 26 27 28 29
+ 31 33 37 38 41
r84 38 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.715
+ $X2=1.09 $Y2=1.88
r85 38 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.715
+ $X2=1.09 $Y2=1.55
r86 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.715 $X2=1.09 $Y2=1.715
r87 34 37 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.86 $Y=1.715
+ $X2=1.09 $Y2=1.715
r88 32 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.88
+ $X2=0.86 $Y2=1.715
r89 32 33 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.86 $Y=1.88 $X2=0.86
+ $Y2=2.03
r90 31 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.55
+ $X2=0.86 $Y2=1.715
r91 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.86 $Y=1.02
+ $X2=0.86 $Y2=1.55
r92 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.775 $Y=2.115
+ $X2=0.86 $Y2=2.03
r93 28 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.775 $Y=2.115
+ $X2=0.445 $Y2=2.115
r94 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.775 $Y=0.935
+ $X2=0.86 $Y2=1.02
r95 26 27 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.775 $Y=0.935
+ $X2=0.405 $Y2=0.935
r96 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.2
+ $X2=0.445 $Y2=2.115
r97 22 24 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=0.28 $Y=2.2 $X2=0.28
+ $Y2=2.265
r98 18 27 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.26 $Y=0.85
+ $X2=0.405 $Y2=0.935
r99 18 20 8.14658 $w=2.88e-07 $l=2.05e-07 $layer=LI1_cond $X=0.26 $Y=0.85
+ $X2=0.26 $Y2=0.645
r100 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.69 $Y=0.545
+ $X2=1.69 $Y2=0.94
r101 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.615 $Y=0.47
+ $X2=1.69 $Y2=0.545
r102 13 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.615 $Y=0.47
+ $X2=1.255 $Y2=0.47
r103 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.18 $Y=0.545
+ $X2=1.255 $Y2=0.47
r104 11 41 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.18 $Y=0.545
+ $X2=1.18 $Y2=1.55
r105 9 42 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.055 $Y=2.54
+ $X2=1.055 $Y2=1.88
r106 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r107 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%B 3 7 9 10 11 12
c37 12 0 7.31803e-20 $X=2.16 $Y=1.665
c38 9 0 1.33077e-19 $X=1.675 $Y=1.795
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.075
+ $Y=1.795 $X2=2.075 $Y2=1.795
r40 12 17 2.38921 $w=4.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.755
+ $X2=2.075 $Y2=1.755
r41 11 17 11.1028 $w=4.08e-07 $l=3.95e-07 $layer=LI1_cond $X=1.68 $Y=1.755
+ $X2=2.075 $Y2=1.755
r42 10 16 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.09 $Y=1.795
+ $X2=2.075 $Y2=1.795
r43 9 16 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=1.675 $Y=1.795
+ $X2=2.075 $Y2=1.795
r44 5 10 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.165 $Y=1.63
+ $X2=2.09 $Y2=1.795
r45 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.165 $Y=1.63
+ $X2=2.165 $Y2=1.015
r46 1 9 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.585 $Y=1.96
+ $X2=1.675 $Y2=1.795
r47 1 3 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.585 $Y=1.96
+ $X2=1.585 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%C 4 7 10 11 12 16 17
c43 10 0 7.31803e-20 $X=2.612 $Y=1.56
r44 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=0.42
+ $X2=2.645 $Y2=0.585
r45 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=0.42 $X2=2.645 $Y2=0.42
r46 12 17 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=2.64 $Y=0.462
+ $X2=2.645 $Y2=0.462
r47 11 12 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=2.64 $Y2=0.462
r48 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.612 $Y=1.41
+ $X2=2.612 $Y2=1.56
r49 7 10 380.935 $w=1.8e-07 $l=9.8e-07 $layer=POLY_cond $X=2.655 $Y=2.54
+ $X2=2.655 $Y2=1.56
r50 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.555 $Y=1.015
+ $X2=2.555 $Y2=1.41
r51 4 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.555 $Y=1.015
+ $X2=2.555 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%D 3 7 9 12
c40 12 0 1.01275e-19 $X=3.15 $Y=1.715
c41 9 0 1.57025e-19 $X=3.12 $Y=1.665
r42 12 15 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.152 $Y=1.715
+ $X2=3.152 $Y2=1.88
r43 12 14 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.152 $Y=1.715
+ $X2=3.152 $Y2=1.55
r44 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.715 $X2=3.15 $Y2=1.715
r45 7 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.245 $Y=0.92
+ $X2=3.245 $Y2=1.55
r46 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.155 $Y=2.54
+ $X2=3.155 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%A_229_424# 1 2 3 12 16 19 23 24 26 27 31 36
+ 37 39 41 46 48
c103 46 0 1.57025e-19 $X=3.725 $Y=1.515
c104 23 0 1.33077e-19 $X=2.595 $Y=1.295
r105 46 49 40.7387 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.732 $Y=1.515
+ $X2=3.732 $Y2=1.68
r106 46 48 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.732 $Y=1.515
+ $X2=3.732 $Y2=1.35
r107 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.725
+ $Y=1.515 $X2=3.725 $Y2=1.515
r108 38 41 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.68 $Y=2.225
+ $X2=2.93 $Y2=2.225
r109 38 39 4.11343 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=2.225
+ $X2=2.595 $Y2=2.225
r110 36 39 59.4556 $w=2.18e-07 $l=1.135e-06 $layer=LI1_cond $X=1.46 $Y=2.24
+ $X2=2.595 $Y2=2.24
r111 34 36 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=2.295
+ $X2=1.46 $Y2=2.295
r112 31 41 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.93 $Y=2.815
+ $X2=2.93 $Y2=2.35
r113 28 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=1.295
+ $X2=2.68 $Y2=1.295
r114 27 45 8.97659 $w=2.99e-07 $l=2.95533e-07 $layer=LI1_cond $X=3.535 $Y=1.295
+ $X2=3.712 $Y2=1.515
r115 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.535 $Y=1.295
+ $X2=2.765 $Y2=1.295
r116 26 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.68 $Y=2.1
+ $X2=2.68 $Y2=2.225
r117 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.38
+ $X2=2.68 $Y2=1.295
r118 25 26 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.68 $Y=1.38
+ $X2=2.68 $Y2=2.1
r119 23 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.295
+ $X2=2.68 $Y2=1.295
r120 23 24 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.595 $Y=1.295
+ $X2=1.64 $Y2=1.295
r121 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=1.21
+ $X2=1.64 $Y2=1.295
r122 17 19 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.475 $Y=1.21
+ $X2=1.475 $Y2=0.765
r123 16 48 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.825 $Y=0.87
+ $X2=3.825 $Y2=1.35
r124 12 49 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.815 $Y=2.4
+ $X2=3.815 $Y2=1.68
r125 3 41 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.12 $X2=2.93 $Y2=2.265
r126 3 31 600 $w=1.7e-07 $l=7.82049e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.12 $X2=2.93 $Y2=2.815
r127 2 34 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=2.12 $X2=1.295 $Y2=2.295
r128 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.62 $X2=1.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%VPWR 1 2 3 12 18 21 22 23 25 35 36 39 44 50
r48 49 50 12.1537 $w=8.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=2.975
+ $X2=2.595 $Y2=2.975
r49 46 49 3.74318 $w=8.78e-07 $l=2.7e-07 $layer=LI1_cond $X=2.16 $Y=2.975
+ $X2=2.43 $Y2=2.975
r50 42 46 6.65455 $w=8.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.975
+ $X2=2.16 $Y2=2.975
r51 42 44 10.3515 $w=8.78e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=2.975
+ $X2=1.645 $Y2=2.975
r52 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 32 50 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.595 $Y2=3.33
r58 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 28 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r62 25 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 23 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 23 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 23 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 21 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r68 20 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r69 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r70 16 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r71 16 18 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=2.265
r72 15 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r73 15 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.645 $Y2=3.33
r74 10 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r75 10 12 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.455
r76 3 18 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=3.245
+ $Y=2.12 $X2=3.5 $Y2=2.265
r77 2 49 300 $w=1.7e-07 $l=9.98299e-07 $layer=licon1_PDIFF $count=2 $X=1.675
+ $Y=2.12 $X2=2.43 $Y2=2.685
r78 1 12 300 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.12 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%X 1 2 9 13 14 15 16 23 32
c24 14 0 1.01275e-19 $X=3.995 $Y=1.95
r25 21 23 0.259705 $w=3.53e-07 $l=8e-09 $layer=LI1_cond $X=4.052 $Y=2.027
+ $X2=4.052 $Y2=2.035
r26 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=4.052 $Y=2.405
+ $X2=4.052 $Y2=2.775
r27 14 21 1.26606 $w=3.53e-07 $l=3.9e-08 $layer=LI1_cond $X=4.052 $Y=1.988
+ $X2=4.052 $Y2=2.027
r28 14 32 7.62255 $w=3.53e-07 $l=1.38e-07 $layer=LI1_cond $X=4.052 $Y=1.988
+ $X2=4.052 $Y2=1.85
r29 14 15 10.7778 $w=3.53e-07 $l=3.32e-07 $layer=LI1_cond $X=4.052 $Y=2.073
+ $X2=4.052 $Y2=2.405
r30 14 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=4.052 $Y=2.073
+ $X2=4.052 $Y2=2.035
r31 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.145 $Y=1.18
+ $X2=4.145 $Y2=1.85
r32 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=4.052 $Y=1.003
+ $X2=4.052 $Y2=1.18
r33 7 9 11.6218 $w=3.53e-07 $l=3.58e-07 $layer=LI1_cond $X=4.052 $Y=1.003
+ $X2=4.052 $Y2=0.645
r34 2 14 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=2.015
r35 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9 $Y=0.5
+ $X2=4.04 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r45 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r46 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.54
+ $Y2=0
r47 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=4.08
+ $Y2=0
r48 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r49 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 25 28 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r52 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 23 36 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.725
+ $Y2=0
r54 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r55 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.54
+ $Y2=0
r56 22 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.12
+ $Y2=0
r57 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 17 36 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.725
+ $Y2=0
r60 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r61 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r62 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r63 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=0.085
+ $X2=3.54 $Y2=0
r64 11 13 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.54 $Y=0.085
+ $X2=3.54 $Y2=0.875
r65 7 36 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r66 7 9 16.5184 $w=2.98e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.515
r67 2 13 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.6 $X2=3.54 $Y2=0.875
r68 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends


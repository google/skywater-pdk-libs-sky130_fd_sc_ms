* File: sky130_fd_sc_ms__o2bb2ai_2.pex.spice
* Created: Wed Sep  2 12:24:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%A1_N 3 7 9 11 12 14 16 17 19 20 23 25 26
+ 31 33 38 43
c96 23 0 1.08648e-19 $X=2.25 $Y=2.45
c97 17 0 7.66098e-20 $X=0.5 $Y=1.3
c98 12 0 1.89231e-19 $X=2.205 $Y=1.68
r99 41 43 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.63
+ $X2=0.24 $Y2=1.665
r100 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.465 $X2=0.315 $Y2=1.465
r101 33 38 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=0.24 $Y=1.465
+ $X2=0.315 $Y2=1.465
r102 33 41 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.465
+ $X2=0.24 $Y2=1.63
r103 33 43 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=1.69
+ $X2=0.24 $Y2=1.665
r104 28 31 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.13 $Y=1.515
+ $X2=2.25 $Y2=1.515
r105 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r106 25 26 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=0.65 $Y=2.517
+ $X2=0.82 $Y2=2.517
r107 24 33 36.327 $w=2.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.24 $Y=2.415
+ $X2=0.24 $Y2=1.69
r108 22 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=1.68
+ $X2=2.25 $Y2=1.515
r109 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.25 $Y=1.68
+ $X2=2.25 $Y2=2.45
r110 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=2.535
+ $X2=2.25 $Y2=2.45
r111 20 26 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.165 $Y=2.535
+ $X2=0.82 $Y2=2.535
r112 19 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.5
+ $X2=0.24 $Y2=2.415
r113 19 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.355 $Y=2.5
+ $X2=0.65 $Y2=2.5
r114 16 37 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.5 $Y=1.465
+ $X2=0.315 $Y2=1.465
r115 16 17 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.465
+ $X2=0.5 $Y2=1.3
r116 12 29 34.8237 $w=2.7e-07 $l=2.14942e-07 $layer=POLY_cond $X=2.205 $Y=1.68
+ $X2=2.09 $Y2=1.515
r117 12 14 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.205 $Y=1.68
+ $X2=2.205 $Y2=2.26
r118 9 29 86.21 $w=2.7e-07 $l=4.90714e-07 $layer=POLY_cond $X=1.96 $Y=1.085
+ $X2=2.09 $Y2=1.515
r119 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.96 $Y=1.085
+ $X2=1.96 $Y2=0.69
r120 5 17 34.7346 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=0.595 $Y=1.3
+ $X2=0.5 $Y2=1.3
r121 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.595 $Y=1.3
+ $X2=0.595 $Y2=0.69
r122 1 17 34.7346 $w=1.65e-07 $l=4.62817e-07 $layer=POLY_cond $X=0.59 $Y=1.72
+ $X2=0.5 $Y2=1.3
r123 1 3 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=0.59 $Y=1.72
+ $X2=0.59 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%A2_N 3 7 11 15 17 26
c63 26 0 1.08648e-19 $X=1.66 $Y=1.61
c64 17 0 7.66098e-20 $X=1.68 $Y=1.665
c65 7 0 1.51381e-19 $X=1.04 $Y=2.355
r66 24 26 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.54 $Y=1.61
+ $X2=1.66 $Y2=1.61
r67 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.61 $X2=1.54 $Y2=1.61
r68 22 24 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.53 $Y=1.61 $X2=1.54
+ $Y2=1.61
r69 21 22 85.682 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=1.04 $Y=1.61 $X2=1.53
+ $Y2=1.61
r70 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.025 $Y=1.61
+ $X2=1.04 $Y2=1.61
r71 17 25 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.612
+ $X2=1.54 $Y2=1.612
r72 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.775
+ $X2=1.66 $Y2=1.61
r73 13 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.66 $Y=1.775
+ $X2=1.66 $Y2=2.355
r74 9 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=1.445
+ $X2=1.53 $Y2=1.61
r75 9 11 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.53 $Y=1.445
+ $X2=1.53 $Y2=0.69
r76 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.775
+ $X2=1.04 $Y2=1.61
r77 5 7 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.04 $Y=1.775 $X2=1.04
+ $Y2=2.355
r78 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.445
+ $X2=1.025 $Y2=1.61
r79 1 3 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.025 $Y=1.445
+ $X2=1.025 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%A_136_387# 1 2 3 12 16 18 20 24 27 28 29
+ 34 36 40 42 43 45
c102 42 0 1.51381e-19 $X=1.895 $Y=2.115
c103 24 0 1.70695e-19 $X=3.38 $Y=0.74
r104 50 51 7.60252 $w=3.17e-07 $l=5e-08 $layer=POLY_cond $X=2.9 $Y=1.465
+ $X2=2.95 $Y2=1.465
r105 48 50 34.9716 $w=3.17e-07 $l=2.3e-07 $layer=POLY_cond $X=2.67 $Y=1.465
+ $X2=2.9 $Y2=1.465
r106 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.465 $X2=2.67 $Y2=1.465
r107 45 47 17.702 $w=2.55e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.095
+ $X2=2.67 $Y2=1.465
r108 42 43 6.26754 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.895 $Y=2.115
+ $X2=1.72 $Y2=2.115
r109 37 40 7.02821 $w=1.7e-07 $l=1.46629e-07 $layer=LI1_cond $X=1.405 $Y=1.095
+ $X2=1.28 $Y2=1.142
r110 36 45 3.11056 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.095
+ $X2=2.67 $Y2=1.095
r111 36 37 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.505 $Y=1.095
+ $X2=1.405 $Y2=1.095
r112 32 40 0.00168595 $w=2.5e-07 $l=1.32e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=1.142
r113 32 34 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.78
r114 31 39 3.6196 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=2.097
+ $X2=0.815 $Y2=2.097
r115 31 43 28.9087 $w=2.93e-07 $l=7.4e-07 $layer=LI1_cond $X=0.98 $Y=2.097
+ $X2=1.72 $Y2=2.097
r116 28 40 7.02821 $w=1.7e-07 $l=1.47054e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=1.28 $Y2=1.142
r117 28 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=0.98 $Y2=1.19
r118 27 39 3.22473 $w=3.3e-07 $l=1.47e-07 $layer=LI1_cond $X=0.815 $Y=1.95
+ $X2=0.815 $Y2=2.097
r119 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.815 $Y=1.275
+ $X2=0.98 $Y2=1.19
r120 26 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.815 $Y=1.275
+ $X2=0.815 $Y2=1.95
r121 22 53 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.3
+ $X2=3.38 $Y2=1.465
r122 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.38 $Y=1.3
+ $X2=3.38 $Y2=0.74
r123 18 53 2.28076 $w=3.17e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.465
+ $X2=3.38 $Y2=1.465
r124 18 51 63.1009 $w=3.17e-07 $l=4.15e-07 $layer=POLY_cond $X=3.365 $Y=1.465
+ $X2=2.95 $Y2=1.465
r125 18 20 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=3.365 $Y=1.605
+ $X2=3.365 $Y2=2.4
r126 14 51 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.3
+ $X2=2.95 $Y2=1.465
r127 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.95 $Y=1.3
+ $X2=2.95 $Y2=0.74
r128 10 50 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.9 $Y=1.63
+ $X2=2.9 $Y2=1.465
r129 10 12 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.9 $Y=1.63 $X2=2.9
+ $Y2=2.4
r130 3 42 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=1.935 $X2=1.895 $Y2=2.115
r131 2 39 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.935 $X2=0.815 $Y2=2.08
r132 1 34 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.37 $X2=1.24 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%B1 3 7 11 15 19 20 22 23 24 30
c87 30 0 1.34056e-19 $X=5.33 $Y=1.515
r88 30 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.33 $Y=1.515
+ $X2=5.33 $Y2=1.68
r89 30 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.33 $Y=1.515
+ $X2=5.33 $Y2=1.35
r90 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.515 $X2=5.33 $Y2=1.515
r91 24 31 3.75 $w=4.88e-07 $l=1.5e-07 $layer=LI1_cond $X=5.21 $Y=1.665 $X2=5.21
+ $Y2=1.515
r92 22 24 3.5 $w=4.88e-07 $l=3.4803e-07 $layer=LI1_cond $X=4.925 $Y=1.805
+ $X2=5.21 $Y2=1.665
r93 22 23 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.925 $Y=1.805
+ $X2=4.025 $Y2=1.805
r94 20 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.86 $Y=1.515
+ $X2=3.86 $Y2=1.68
r95 20 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.86 $Y=1.515
+ $X2=3.86 $Y2=1.35
r96 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.86
+ $Y=1.515 $X2=3.86 $Y2=1.515
r97 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.86 $Y=1.72
+ $X2=4.025 $Y2=1.805
r98 17 19 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.86 $Y=1.72
+ $X2=3.86 $Y2=1.515
r99 15 32 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.265 $Y=0.74
+ $X2=5.265 $Y2=1.35
r100 11 33 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.255 $Y=2.4
+ $X2=5.255 $Y2=1.68
r101 7 28 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.905 $Y=2.4
+ $X2=3.905 $Y2=1.68
r102 3 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.84 $Y=0.74
+ $X2=3.84 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%B2 1 3 6 10 12 14 15 24
c56 15 0 1.34056e-19 $X=4.56 $Y=1.295
c57 1 0 9.27061e-20 $X=4.34 $Y=1.22
r58 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.805 $Y=1.385
+ $X2=4.82 $Y2=1.385
r59 21 23 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=4.51 $Y=1.385
+ $X2=4.805 $Y2=1.385
r60 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.385 $X2=4.51 $Y2=1.385
r61 19 21 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=4.355 $Y=1.385
+ $X2=4.51 $Y2=1.385
r62 17 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.34 $Y=1.385
+ $X2=4.355 $Y2=1.385
r63 15 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.51 $Y=1.295 $X2=4.51
+ $Y2=1.385
r64 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.82 $Y=1.22
+ $X2=4.82 $Y2=1.385
r65 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.82 $Y=1.22 $X2=4.82
+ $Y2=0.74
r66 8 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.55
+ $X2=4.805 $Y2=1.385
r67 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.805 $Y=1.55
+ $X2=4.805 $Y2=2.4
r68 4 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.55
+ $X2=4.355 $Y2=1.385
r69 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.355 $Y=1.55
+ $X2=4.355 $Y2=2.4
r70 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.34 $Y=1.22
+ $X2=4.34 $Y2=1.385
r71 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.34 $Y=1.22 $X2=4.34
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%VPWR 1 2 3 4 5 16 18 20 24 28 34 36 38 42
+ 44 49 54 66 69 72 76
r79 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r84 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 61 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r86 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 58 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=5.04
+ $Y2=3.33
r90 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 55 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=3.625 $Y2=3.33
r92 55 57 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 54 75 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.577 $Y2=3.33
r94 54 60 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 53 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r96 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 50 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=3.33
r98 50 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.625 $Y2=3.33
r100 49 52 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 48 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 45 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.35 $Y2=3.33
r105 45 47 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 44 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.67 $Y2=3.33
r107 44 47 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 42 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 42 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 38 41 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.52 $Y=2.115
+ $X2=5.52 $Y2=2.815
r111 36 75 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.577 $Y2=3.33
r112 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=2.815
r113 32 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=3.245
+ $X2=3.625 $Y2=3.33
r114 32 34 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=3.625 $Y=3.245
+ $X2=3.625 $Y2=2.485
r115 28 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.67 $Y=1.985
+ $X2=2.67 $Y2=2.815
r116 26 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r117 26 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.815
r118 22 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=3.245
+ $X2=1.35 $Y2=3.33
r119 22 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.35 $Y=3.245
+ $X2=1.35 $Y2=2.875
r120 21 63 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r121 20 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=1.35 $Y2=3.33
r122 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=0.445 $Y2=3.33
r123 16 63 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r124 16 18 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.84
r125 5 41 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.84 $X2=5.48 $Y2=2.815
r126 5 38 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.84 $X2=5.48 $Y2=2.115
r127 4 34 300 $w=1.7e-07 $l=7.25034e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.84 $X2=3.625 $Y2=2.485
r128 3 31 600 $w=1.7e-07 $l=1.14728e-06 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.84 $X2=2.67 $Y2=2.815
r129 3 28 300 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=2 $X=2.295
+ $Y=1.84 $X2=2.67 $Y2=1.985
r130 2 24 600 $w=1.7e-07 $l=1.04422e-06 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.935 $X2=1.35 $Y2=2.875
r131 1 18 600 $w=1.7e-07 $l=9.74808e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.935 $X2=0.28 $Y2=2.84
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%Y 1 2 3 12 14 19 20 21 22 23 35 45
c44 20 0 1.39855e-19 $X=3.035 $Y=0.84
r45 37 45 1.01091 $w=2.83e-07 $l=2.5e-08 $layer=LI1_cond $X=3.147 $Y=2.06
+ $X2=3.147 $Y2=2.035
r46 30 35 2.38436 $w=2.88e-07 $l=6e-08 $layer=LI1_cond $X=3.145 $Y=0.985
+ $X2=3.145 $Y2=0.925
r47 23 37 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.147 $Y=2.145
+ $X2=3.147 $Y2=2.06
r48 23 45 2.02183 $w=2.83e-07 $l=5e-08 $layer=LI1_cond $X=3.147 $Y=1.985
+ $X2=3.147 $Y2=2.035
r49 22 23 12.9397 $w=2.83e-07 $l=3.2e-07 $layer=LI1_cond $X=3.147 $Y=1.665
+ $X2=3.147 $Y2=1.985
r50 21 22 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.147 $Y=1.295
+ $X2=3.147 $Y2=1.665
r51 21 47 6.67204 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.147 $Y=1.295
+ $X2=3.147 $Y2=1.13
r52 20 47 5.28534 $w=2.88e-07 $l=1.33e-07 $layer=LI1_cond $X=3.145 $Y=0.997
+ $X2=3.145 $Y2=1.13
r53 20 30 0.476873 $w=2.88e-07 $l=1.2e-08 $layer=LI1_cond $X=3.145 $Y=0.997
+ $X2=3.145 $Y2=0.985
r54 20 35 2.58306 $w=2.88e-07 $l=6.5e-08 $layer=LI1_cond $X=3.145 $Y=0.86
+ $X2=3.145 $Y2=0.925
r55 15 23 3.25423 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.29 $Y=2.145
+ $X2=3.147 $Y2=2.145
r56 14 19 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.465 $Y=2.145
+ $X2=4.58 $Y2=2.145
r57 14 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=4.465 $Y=2.145
+ $X2=3.29 $Y2=2.145
r58 10 23 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.147 $Y=2.23
+ $X2=3.147 $Y2=2.145
r59 10 12 23.6554 $w=2.83e-07 $l=5.85e-07 $layer=LI1_cond $X=3.147 $Y=2.23
+ $X2=3.147 $Y2=2.815
r60 3 19 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=4.445
+ $Y=1.84 $X2=4.58 $Y2=2.225
r61 2 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.125 $Y2=1.985
r62 2 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.125 $Y2=2.815
r63 1 20 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%A_799_368# 1 2 9 11 12 15
r28 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.03 $Y=2.145
+ $X2=5.03 $Y2=2.825
r29 13 18 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.03 $Y=2.905 $X2=5.03
+ $Y2=2.825
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.865 $Y=2.99
+ $X2=5.03 $Y2=2.905
r31 11 12 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.865 $Y=2.99
+ $X2=4.295 $Y2=2.99
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.13 $Y=2.905
+ $X2=4.295 $Y2=2.99
r33 7 9 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.13 $Y=2.905 $X2=4.13
+ $Y2=2.485
r34 2 18 400 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.84 $X2=5.03 $Y2=2.825
r35 2 15 400 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.84 $X2=5.03 $Y2=2.145
r36 1 9 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=3.995
+ $Y=1.84 $X2=4.13 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%VGND 1 2 3 4 13 15 19 23 27 29 31 36 44 51
+ 52 58 61 64
c72 19 0 1.89231e-19 $X=2.175 $Y=0.66
r73 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r74 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r75 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r76 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r78 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r79 49 64 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.042
+ $Y2=0
r80 49 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.52
+ $Y2=0
r81 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r82 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r83 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.125
+ $Y2=0
r85 45 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.56
+ $Y2=0
r86 44 64 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.87 $Y=0 $X2=5.042
+ $Y2=0
r87 44 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.87 $Y=0 $X2=4.56
+ $Y2=0
r88 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r89 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r90 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r91 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r92 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r93 37 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.21
+ $Y2=0
r94 37 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.64
+ $Y2=0
r95 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=4.125
+ $Y2=0
r96 36 42 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.6
+ $Y2=0
r97 35 59 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r98 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r99 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r100 32 55 4.66755 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=0
+ $X2=0.237 $Y2=0
r101 32 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=0 $X2=0.72
+ $Y2=0
r102 31 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.08 $Y=0 $X2=2.21
+ $Y2=0
r103 31 34 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.08 $Y=0 $X2=0.72
+ $Y2=0
r104 29 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r105 29 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r106 25 64 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.042 $Y=0.085
+ $X2=5.042 $Y2=0
r107 25 27 14.3638 $w=3.43e-07 $l=4.3e-07 $layer=LI1_cond $X=5.042 $Y=0.085
+ $X2=5.042 $Y2=0.515
r108 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0.085
+ $X2=4.125 $Y2=0
r109 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.125 $Y=0.085
+ $X2=4.125 $Y2=0.55
r110 17 58 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r111 17 19 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.66
r112 13 55 3.09863 $w=3.3e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.237 $Y2=0
r113 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.31 $Y2=0.515
r114 4 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.895
+ $Y=0.37 $X2=5.04 $Y2=0.515
r115 3 23 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.37 $X2=4.125 $Y2=0.55
r116 2 19 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.37 $X2=2.175 $Y2=0.66
r117 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%A_134_74# 1 2 9 11 12 15
r24 13 15 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.745 $Y=0.425
+ $X2=1.745 $Y2=0.66
r25 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.58 $Y=0.34
+ $X2=1.745 $Y2=0.425
r26 11 12 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.58 $Y=0.34
+ $X2=0.975 $Y2=0.34
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.81 $Y=0.425
+ $X2=0.975 $Y2=0.34
r28 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=0.81 $Y=0.425 $X2=0.81
+ $Y2=0.495
r29 2 15 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.37 $X2=1.745 $Y2=0.66
r30 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.67
+ $Y=0.37 $X2=0.81 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2AI_2%A_518_74# 1 2 3 4 15 17 18 22 23 24 27 29
+ 31 33 36
c60 24 0 1.70695e-19 $X=3.79 $Y=0.925
c61 17 0 9.27061e-20 $X=3.46 $Y=0.34
r62 31 38 3.37178 $w=2.5e-07 $l=1.98997e-07 $layer=LI1_cond $X=5.52 $Y=0.77
+ $X2=5.48 $Y2=0.95
r63 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.52 $Y=0.77
+ $X2=5.52 $Y2=0.515
r64 30 36 5.47651 $w=2.05e-07 $l=1.1e-07 $layer=LI1_cond $X=4.69 $Y=0.89
+ $X2=4.58 $Y2=0.89
r65 29 38 3.44841 $w=2.4e-07 $l=1.92678e-07 $layer=LI1_cond $X=5.315 $Y=0.89
+ $X2=5.48 $Y2=0.95
r66 29 30 30.0115 $w=2.38e-07 $l=6.25e-07 $layer=LI1_cond $X=5.315 $Y=0.89
+ $X2=4.69 $Y2=0.89
r67 25 36 1.08954 $w=2.2e-07 $l=1.2e-07 $layer=LI1_cond $X=4.58 $Y=0.77 $X2=4.58
+ $Y2=0.89
r68 25 27 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=4.58 $Y=0.77
+ $X2=4.58 $Y2=0.515
r69 23 36 5.47651 $w=2.05e-07 $l=1.26293e-07 $layer=LI1_cond $X=4.47 $Y=0.925
+ $X2=4.58 $Y2=0.89
r70 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.47 $Y=0.925
+ $X2=3.79 $Y2=0.925
r71 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.625 $Y=0.84
+ $X2=3.79 $Y2=0.925
r72 20 22 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.625 $Y=0.84
+ $X2=3.625 $Y2=0.515
r73 19 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.625 $Y=0.425
+ $X2=3.625 $Y2=0.515
r74 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.46 $Y=0.34
+ $X2=3.625 $Y2=0.425
r75 17 18 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.46 $Y=0.34 $X2=2.82
+ $Y2=0.34
r76 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.695 $Y=0.425
+ $X2=2.82 $Y2=0.34
r77 13 15 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=2.695 $Y=0.425
+ $X2=2.695 $Y2=0.66
r78 4 38 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.95
r79 4 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.515
r80 3 36 182 $w=1.7e-07 $l=6.32139e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.37 $X2=4.58 $Y2=0.925
r81 3 27 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.415
+ $Y=0.37 $X2=4.58 $Y2=0.515
r82 2 22 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.37 $X2=3.625 $Y2=0.515
r83 1 15 182 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.37 $X2=2.735 $Y2=0.66
.ends


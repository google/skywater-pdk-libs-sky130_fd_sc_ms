# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.310000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.502100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.470000 0.350000 13.835000 1.130000 ;
        RECT 13.555000 1.820000 13.835000 2.980000 ;
        RECT 13.665000 1.130000 13.835000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.520800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.015000 0.350000 12.345000 2.980000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.455400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.785000 1.820000  4.165000 2.150000 ;
        RECT  7.745000 1.820000  8.035000 2.150000 ;
        RECT 10.695000 1.685000 11.065000 2.150000 ;
      LAYER mcon ;
        RECT  3.995000 1.950000  4.165000 2.120000 ;
        RECT  7.835000 1.950000  8.005000 2.120000 ;
        RECT 10.715000 1.950000 10.885000 2.120000 ;
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.935000 1.440000 3.265000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.490000 2.725000 1.660000 ;
        RECT 0.605000 1.660000 1.795000 1.880000 ;
        RECT 2.395000 1.260000 2.725000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.785000 1.180000 4.645000 1.650000 ;
        RECT 4.395000 1.650000 4.645000 1.775000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.920000 0.085000 ;
        RECT  0.545000  0.085000  0.875000 0.810000 ;
        RECT  3.560000  0.085000  3.865000 0.750000 ;
        RECT  4.660000  0.085000  4.990000 0.670000 ;
        RECT  7.440000  0.085000  7.770000 0.425000 ;
        RECT 10.165000  0.085000 10.495000 0.760000 ;
        RECT 11.510000  0.085000 11.840000 0.410000 ;
        RECT 13.120000  0.085000 13.290000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.920000 3.415000 ;
        RECT  1.225000 2.390000  1.555000 3.245000 ;
        RECT  3.085000 2.730000  3.445000 3.245000 ;
        RECT  4.705000 2.795000  5.035000 3.245000 ;
        RECT  7.090000 2.660000  7.420000 3.245000 ;
        RECT  8.235000 1.715000  8.485000 3.245000 ;
        RECT 10.305000 2.660000 10.650000 3.245000 ;
        RECT 11.370000 2.695000 11.815000 3.245000 ;
        RECT 11.585000 1.970000 11.815000 2.695000 ;
        RECT 13.045000 1.820000 13.325000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.350000  0.365000 0.980000 ;
      RECT  0.115000 0.980000  1.395000 1.310000 ;
      RECT  0.115000 1.310000  0.285000 2.050000 ;
      RECT  0.115000 2.050000  2.695000 2.220000 ;
      RECT  0.115000 2.220000  1.055000 2.975000 ;
      RECT  1.105000 0.255000  3.390000 0.425000 ;
      RECT  1.105000 0.425000  1.355000 0.810000 ;
      RECT  2.095000 2.390000  3.985000 2.445000 ;
      RECT  2.095000 2.445000  5.975000 2.560000 ;
      RECT  2.095000 2.560000  2.425000 3.000000 ;
      RECT  2.270000 0.595000  2.600000 0.920000 ;
      RECT  2.270000 0.920000  3.615000 1.090000 ;
      RECT  2.365000 1.830000  2.695000 2.050000 ;
      RECT  3.060000 0.425000  3.390000 0.750000 ;
      RECT  3.445000 1.090000  3.615000 2.320000 ;
      RECT  3.445000 2.320000  3.985000 2.390000 ;
      RECT  3.615000 2.560000  5.975000 2.625000 ;
      RECT  3.615000 2.625000  3.985000 3.000000 ;
      RECT  4.225000 0.595000  4.490000 0.840000 ;
      RECT  4.225000 0.840000  4.985000 1.010000 ;
      RECT  4.335000 1.945000  4.985000 2.115000 ;
      RECT  4.335000 2.115000  4.585000 2.275000 ;
      RECT  4.815000 1.010000  4.985000 1.445000 ;
      RECT  4.815000 1.445000  5.215000 1.775000 ;
      RECT  4.815000 1.775000  4.985000 1.945000 ;
      RECT  5.155000 1.945000  5.620000 2.275000 ;
      RECT  5.170000 0.255000  7.185000 0.425000 ;
      RECT  5.170000 0.425000  5.420000 1.105000 ;
      RECT  5.170000 1.105000  5.620000 1.275000 ;
      RECT  5.385000 1.275000  5.620000 1.575000 ;
      RECT  5.385000 1.575000  6.165000 1.905000 ;
      RECT  5.385000 1.905000  5.620000 1.945000 ;
      RECT  5.725000 2.625000  5.975000 2.755000 ;
      RECT  5.790000 2.075000  6.505000 2.245000 ;
      RECT  5.790000 2.245000  5.975000 2.445000 ;
      RECT  5.800000 0.595000  5.980000 1.095000 ;
      RECT  5.800000 1.095000  6.505000 1.265000 ;
      RECT  6.150000 0.595000  6.845000 0.925000 ;
      RECT  6.175000 2.415000  7.945000 2.490000 ;
      RECT  6.175000 2.490000  6.845000 2.755000 ;
      RECT  6.335000 1.265000  6.505000 2.075000 ;
      RECT  6.675000 0.925000  6.845000 2.320000 ;
      RECT  6.675000 2.320000  7.945000 2.415000 ;
      RECT  7.015000 0.425000  7.185000 0.595000 ;
      RECT  7.015000 0.595000  8.110000 0.765000 ;
      RECT  7.015000 0.935000  8.610000 1.105000 ;
      RECT  7.015000 1.105000  7.235000 1.780000 ;
      RECT  7.405000 1.275000  8.270000 1.545000 ;
      RECT  7.405000 1.545000  7.575000 2.320000 ;
      RECT  7.615000 2.490000  7.945000 2.755000 ;
      RECT  7.940000 0.255000  8.950000 0.425000 ;
      RECT  7.940000 0.425000  8.110000 0.595000 ;
      RECT  8.280000 0.595000  8.610000 0.935000 ;
      RECT  8.440000 1.105000  8.610000 1.245000 ;
      RECT  8.440000 1.245000  8.935000 1.415000 ;
      RECT  8.685000 1.415000  8.935000 2.755000 ;
      RECT  8.780000 0.425000  8.950000 0.905000 ;
      RECT  8.780000 0.905000  9.435000 1.075000 ;
      RECT  9.105000 1.075000  9.435000 1.345000 ;
      RECT  9.105000 1.345000  9.755000 1.575000 ;
      RECT  9.105000 1.755000  9.325000 2.425000 ;
      RECT  9.105000 2.425000 10.095000 2.755000 ;
      RECT  9.135000 0.405000  9.775000 0.735000 ;
      RECT  9.505000 1.575000  9.755000 2.230000 ;
      RECT  9.605000 0.735000  9.775000 1.005000 ;
      RECT  9.605000 1.005000 11.425000 1.175000 ;
      RECT  9.925000 1.175000 11.425000 1.435000 ;
      RECT  9.925000 1.435000 10.095000 2.425000 ;
      RECT 10.265000 1.650000 10.525000 2.320000 ;
      RECT 10.265000 2.320000 11.405000 2.490000 ;
      RECT 10.855000 2.490000 11.185000 2.885000 ;
      RECT 10.955000 0.350000 11.285000 0.580000 ;
      RECT 10.955000 0.580000 11.845000 0.750000 ;
      RECT 11.235000 1.630000 11.845000 1.800000 ;
      RECT 11.235000 1.800000 11.405000 2.320000 ;
      RECT 11.675000 0.750000 11.845000 1.630000 ;
      RECT 12.570000 0.455000 12.855000 1.300000 ;
      RECT 12.570000 1.300000 13.485000 1.630000 ;
      RECT 12.570000 1.630000 12.855000 2.980000 ;
  END
END sky130_fd_sc_ms__sdfrbp_1

* File: sky130_fd_sc_ms__o32a_4.pxi.spice
* Created: Fri Aug 28 18:03:57 2020
* 
x_PM_SKY130_FD_SC_MS__O32A_4%A_83_256# N_A_83_256#_M1010_d N_A_83_256#_M1021_s
+ N_A_83_256#_M1016_d N_A_83_256#_M1000_s N_A_83_256#_M1003_g
+ N_A_83_256#_M1015_g N_A_83_256#_c_160_n N_A_83_256#_M1006_g
+ N_A_83_256#_M1020_g N_A_83_256#_M1008_g N_A_83_256#_M1024_g
+ N_A_83_256#_M1009_g N_A_83_256#_M1027_g N_A_83_256#_c_167_n
+ N_A_83_256#_c_168_n N_A_83_256#_c_169_n N_A_83_256#_c_170_n
+ N_A_83_256#_c_171_n N_A_83_256#_c_172_n N_A_83_256#_c_192_p
+ N_A_83_256#_c_173_n N_A_83_256#_c_180_n N_A_83_256#_c_229_p
+ N_A_83_256#_c_174_n PM_SKY130_FD_SC_MS__O32A_4%A_83_256#
x_PM_SKY130_FD_SC_MS__O32A_4%B1 N_B1_M1018_g N_B1_c_328_n N_B1_c_329_n
+ N_B1_c_330_n N_B1_c_331_n N_B1_M1010_g N_B1_c_332_n N_B1_c_333_n N_B1_M1025_g
+ N_B1_c_340_n N_B1_M1023_g N_B1_c_341_n N_B1_c_342_n N_B1_c_343_n N_B1_c_334_n
+ N_B1_c_344_n N_B1_c_345_n N_B1_c_430_p N_B1_c_346_n N_B1_c_347_n N_B1_c_335_n
+ N_B1_c_336_n B1 N_B1_c_337_n N_B1_c_338_n PM_SKY130_FD_SC_MS__O32A_4%B1
x_PM_SKY130_FD_SC_MS__O32A_4%B2 N_B2_c_480_n N_B2_M1016_g N_B2_c_481_n
+ N_B2_c_482_n N_B2_c_472_n N_B2_M1019_g N_B2_c_473_n N_B2_c_474_n N_B2_M1021_g
+ N_B2_c_475_n N_B2_c_476_n N_B2_M1022_g N_B2_c_477_n B2 N_B2_c_478_n
+ N_B2_c_479_n PM_SKY130_FD_SC_MS__O32A_4%B2
x_PM_SKY130_FD_SC_MS__O32A_4%A3 N_A3_M1002_g N_A3_M1000_g N_A3_c_556_n
+ N_A3_M1017_g N_A3_M1012_g N_A3_c_552_n A3 N_A3_c_554_n
+ PM_SKY130_FD_SC_MS__O32A_4%A3
x_PM_SKY130_FD_SC_MS__O32A_4%A2 N_A2_M1001_g N_A2_c_612_n N_A2_M1004_g
+ N_A2_c_613_n N_A2_M1007_g N_A2_M1013_g N_A2_c_614_n N_A2_c_615_n A2 A2 A2 A2
+ N_A2_c_617_n N_A2_c_638_n N_A2_c_618_n A2 N_A2_c_619_n
+ PM_SKY130_FD_SC_MS__O32A_4%A2
x_PM_SKY130_FD_SC_MS__O32A_4%A1 N_A1_c_710_n N_A1_M1011_g N_A1_c_704_n
+ N_A1_M1005_g N_A1_c_711_n N_A1_M1026_g N_A1_c_705_n N_A1_c_706_n N_A1_M1014_g
+ N_A1_c_707_n A1 N_A1_c_708_n N_A1_c_709_n PM_SKY130_FD_SC_MS__O32A_4%A1
x_PM_SKY130_FD_SC_MS__O32A_4%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1009_d
+ N_VPWR_M1023_s N_VPWR_M1011_s N_VPWR_c_767_n N_VPWR_c_768_n N_VPWR_c_769_n
+ N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n N_VPWR_c_774_n
+ N_VPWR_c_775_n VPWR N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n
+ N_VPWR_c_766_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n
+ PM_SKY130_FD_SC_MS__O32A_4%VPWR
x_PM_SKY130_FD_SC_MS__O32A_4%X N_X_M1015_d N_X_M1024_d N_X_M1003_s N_X_M1008_s
+ N_X_c_865_n N_X_c_866_n N_X_c_867_n N_X_c_874_n N_X_c_868_n N_X_c_875_n
+ N_X_c_869_n N_X_c_876_n N_X_c_870_n N_X_c_871_n N_X_c_906_n X N_X_c_873_n
+ PM_SKY130_FD_SC_MS__O32A_4%X
x_PM_SKY130_FD_SC_MS__O32A_4%A_537_388# N_A_537_388#_M1018_d
+ N_A_537_388#_M1019_s N_A_537_388#_c_938_n
+ PM_SKY130_FD_SC_MS__O32A_4%A_537_388#
x_PM_SKY130_FD_SC_MS__O32A_4%A_961_392# N_A_961_392#_M1000_d
+ N_A_961_392#_M1017_d N_A_961_392#_M1013_s N_A_961_392#_c_955_n
+ N_A_961_392#_c_969_n N_A_961_392#_c_973_n N_A_961_392#_c_966_n
+ N_A_961_392#_c_956_n N_A_961_392#_c_957_n N_A_961_392#_c_958_n
+ PM_SKY130_FD_SC_MS__O32A_4%A_961_392#
x_PM_SKY130_FD_SC_MS__O32A_4%A_1237_392# N_A_1237_392#_M1001_d
+ N_A_1237_392#_M1026_d N_A_1237_392#_c_1007_n N_A_1237_392#_c_1014_n
+ N_A_1237_392#_c_1006_n N_A_1237_392#_c_1016_n
+ PM_SKY130_FD_SC_MS__O32A_4%A_1237_392#
x_PM_SKY130_FD_SC_MS__O32A_4%VGND N_VGND_M1015_s N_VGND_M1020_s N_VGND_M1027_s
+ N_VGND_M1002_s N_VGND_M1004_s N_VGND_M1005_d N_VGND_c_1027_n N_VGND_c_1028_n
+ N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n N_VGND_c_1032_n
+ N_VGND_c_1033_n N_VGND_c_1034_n N_VGND_c_1035_n N_VGND_c_1036_n
+ N_VGND_c_1037_n N_VGND_c_1038_n N_VGND_c_1039_n N_VGND_c_1040_n VGND
+ N_VGND_c_1041_n N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n
+ N_VGND_c_1045_n PM_SKY130_FD_SC_MS__O32A_4%VGND
x_PM_SKY130_FD_SC_MS__O32A_4%A_564_74# N_A_564_74#_M1010_s N_A_564_74#_M1025_s
+ N_A_564_74#_M1022_d N_A_564_74#_M1012_d N_A_564_74#_M1007_d
+ N_A_564_74#_M1014_s N_A_564_74#_c_1134_n N_A_564_74#_c_1135_n
+ N_A_564_74#_c_1136_n N_A_564_74#_c_1150_n N_A_564_74#_c_1137_n
+ N_A_564_74#_c_1138_n N_A_564_74#_c_1172_n N_A_564_74#_c_1139_n
+ N_A_564_74#_c_1182_n N_A_564_74#_c_1140_n N_A_564_74#_c_1141_n
+ N_A_564_74#_c_1142_n N_A_564_74#_c_1143_n N_A_564_74#_c_1178_n
+ N_A_564_74#_c_1191_n PM_SKY130_FD_SC_MS__O32A_4%A_564_74#
cc_1 VNB N_A_83_256#_M1003_g 0.0139124f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_256#_M1015_g 0.0224732f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_3 VNB N_A_83_256#_c_160_n 0.00585843f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.355
cc_4 VNB N_A_83_256#_M1006_g 0.0110137f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_5 VNB N_A_83_256#_M1020_g 0.0208918f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_6 VNB N_A_83_256#_M1008_g 0.00293103f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_7 VNB N_A_83_256#_M1024_g 0.0229607f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=0.74
cc_8 VNB N_A_83_256#_M1009_g 0.0031281f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.4
cc_9 VNB N_A_83_256#_M1027_g 0.0231429f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=0.74
cc_10 VNB N_A_83_256#_c_167_n 0.0132856f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.355
cc_11 VNB N_A_83_256#_c_168_n 0.00163584f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.445
cc_12 VNB N_A_83_256#_c_169_n 0.0799573f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_13 VNB N_A_83_256#_c_170_n 0.0226784f $X=-0.19 $Y=-0.245 $X2=3.23 $Y2=1.195
cc_14 VNB N_A_83_256#_c_171_n 0.0013403f $X=-0.19 $Y=-0.245 $X2=3.395 $Y2=1.28
cc_15 VNB N_A_83_256#_c_172_n 0.00846832f $X=-0.19 $Y=-0.245 $X2=3.395 $Y2=1.92
cc_16 VNB N_A_83_256#_c_173_n 0.00267952f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.015
cc_17 VNB N_A_83_256#_c_174_n 0.00527666f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.195
cc_18 VNB N_B1_c_328_n 0.013557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_329_n 0.016436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_330_n 0.0119858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_331_n 0.0189724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_332_n 0.020595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_333_n 0.0145703f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_24 VNB N_B1_c_334_n 0.00530224f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_25 VNB N_B1_c_335_n 0.00489941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_336_n 0.0213149f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.28
cc_27 VNB N_B1_c_337_n 0.0220325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B1_c_338_n 0.00267016f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_29 VNB N_B2_c_472_n 0.0142058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B2_c_473_n 0.0274709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B2_c_474_n 0.0151192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B2_c_475_n 0.0302534f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_33 VNB N_B2_c_476_n 0.0158157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B2_c_477_n 0.0110645f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.355
cc_35 VNB N_B2_c_478_n 0.0236629f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_36 VNB N_B2_c_479_n 9.04634e-19 $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_37 VNB N_A3_M1002_g 0.022736f $X=-0.19 $Y=-0.245 $X2=3.275 $Y2=1.94
cc_38 VNB N_A3_M1000_g 0.0084209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A3_M1012_g 0.0217763f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_40 VNB N_A3_c_552_n 0.00799726f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_41 VNB A3 0.0124579f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_42 VNB N_A3_c_554_n 0.044114f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_43 VNB N_A2_c_612_n 0.0162939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A2_c_613_n 0.0156098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A2_c_614_n 0.029645f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.28
cc_46 VNB N_A2_c_615_n 0.00499367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB A2 0.0116853f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_48 VNB N_A2_c_617_n 0.0326934f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_49 VNB N_A2_c_618_n 0.0235028f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.28
cc_50 VNB N_A2_c_619_n 0.00960991f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_51 VNB N_A1_c_704_n 0.0172606f $X=-0.19 $Y=-0.245 $X2=5.265 $Y2=1.96
cc_52 VNB N_A1_c_705_n 0.0298031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A1_c_706_n 0.0223976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A1_c_707_n 0.00981662f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.355
cc_55 VNB N_A1_c_708_n 0.0352436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A1_c_709_n 0.0111425f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_57 VNB N_VPWR_c_766_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_X_c_865_n 0.00341655f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.43
cc_59 VNB N_X_c_866_n 0.00221303f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_60 VNB N_X_c_867_n 0.00932569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_X_c_868_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_62 VNB N_X_c_869_n 0.00162994f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_63 VNB N_X_c_870_n 0.00282884f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.61
cc_64 VNB N_X_c_871_n 0.00154309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB X 0.00825292f $X=-0.19 $Y=-0.245 $X2=2.185 $Y2=1.445
cc_66 VNB N_X_c_873_n 0.011349f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_67 VNB N_VGND_c_1027_n 0.0144497f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.74
cc_68 VNB N_VGND_c_1028_n 0.0355428f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.355
cc_69 VNB N_VGND_c_1029_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.43
cc_70 VNB N_VGND_c_1030_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.28
cc_71 VNB N_VGND_c_1031_n 0.011586f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.61
cc_72 VNB N_VGND_c_1032_n 0.00867401f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.28
cc_73 VNB N_VGND_c_1033_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.61
cc_74 VNB N_VGND_c_1034_n 0.00947287f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=1.28
cc_75 VNB N_VGND_c_1035_n 0.020287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1036_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.355
cc_77 VNB N_VGND_c_1037_n 0.0627424f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_78 VNB N_VGND_c_1038_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_79 VNB N_VGND_c_1039_n 0.0186748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1040_n 0.00613276f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_81 VNB N_VGND_c_1041_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1042_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1043_n 0.436015f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=1.445
cc_84 VNB N_VGND_c_1044_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.43
cc_85 VNB N_VGND_c_1045_n 0.00737978f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.445
cc_86 VNB N_A_564_74#_c_1134_n 0.00465679f $X=-0.19 $Y=-0.245 $X2=0.865
+ $Y2=1.355
cc_87 VNB N_A_564_74#_c_1135_n 0.00230691f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.43
cc_88 VNB N_A_564_74#_c_1136_n 0.00418558f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_89 VNB N_A_564_74#_c_1137_n 0.00670648f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.74
cc_90 VNB N_A_564_74#_c_1138_n 0.00400232f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_91 VNB N_A_564_74#_c_1139_n 0.00256835f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.61
cc_92 VNB N_A_564_74#_c_1140_n 0.00206225f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=0.74
cc_93 VNB N_A_564_74#_c_1141_n 0.0139705f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.355
cc_94 VNB N_A_564_74#_c_1142_n 0.0189752f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.445
cc_95 VNB N_A_564_74#_c_1143_n 0.00220179f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.445
cc_96 VPB N_A_83_256#_M1003_g 0.0274205f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_97 VPB N_A_83_256#_M1006_g 0.0219998f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_98 VPB N_A_83_256#_M1008_g 0.0233198f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_99 VPB N_A_83_256#_M1009_g 0.0250827f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=2.4
cc_100 VPB N_A_83_256#_c_172_n 9.11378e-19 $X=-0.19 $Y=1.66 $X2=3.395 $Y2=1.92
cc_101 VPB N_A_83_256#_c_180_n 0.00230942f $X=-0.19 $Y=1.66 $X2=5.4 $Y2=2.105
cc_102 VPB N_B1_M1018_g 0.0234822f $X=-0.19 $Y=1.66 $X2=3.275 $Y2=1.94
cc_103 VPB N_B1_c_340_n 0.0151012f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.28
cc_104 VPB N_B1_c_341_n 0.0364563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_B1_c_342_n 0.0136199f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.355
cc_106 VPB N_B1_c_343_n 0.0698096f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.43
cc_107 VPB N_B1_c_344_n 0.00274485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_B1_c_345_n 0.00329833f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.28
cc_109 VPB N_B1_c_346_n 0.0201001f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_110 VPB N_B1_c_347_n 0.00197943f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_111 VPB N_B1_c_335_n 0.00338539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_B1_c_336_n 0.013955f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.28
cc_113 VPB N_B1_c_337_n 0.0141581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_B1_c_338_n 0.00123343f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.445
cc_115 VPB N_B2_c_480_n 0.0163479f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=0.37
cc_116 VPB N_B2_c_481_n 0.0120921f $X=-0.19 $Y=1.66 $X2=5.265 $Y2=1.96
cc_117 VPB N_B2_c_482_n 0.010564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B2_c_472_n 0.0270867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_B2_c_479_n 0.0045594f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_120 VPB N_A3_M1000_g 0.0291583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A3_c_556_n 0.0245654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A3_c_552_n 0.00408276f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_123 VPB N_A2_M1001_g 0.0240552f $X=-0.19 $Y=1.66 $X2=3.275 $Y2=1.94
cc_124 VPB N_A2_M1013_g 0.0318255f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.43
cc_125 VPB N_A2_c_615_n 0.0172522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB A2 0.00227558f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.355
cc_127 VPB A2 0.00614495f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_128 VPB N_A2_c_618_n 0.0129154f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.28
cc_129 VPB N_A2_c_619_n 0.00476546f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.445
cc_130 VPB N_A1_c_710_n 0.0181274f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=0.37
cc_131 VPB N_A1_c_711_n 0.044222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A1_c_708_n 0.00513583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_767_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_768_n 0.0570215f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_135 VPB N_VPWR_c_769_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_136 VPB N_VPWR_c_770_n 0.0190152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_771_n 0.00708345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_772_n 0.00517516f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=0.74
cc_139 VPB N_VPWR_c_773_n 0.00396467f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=2.4
cc_140 VPB N_VPWR_c_774_n 0.0456572f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=1.28
cc_141 VPB N_VPWR_c_775_n 0.00510271f $X=-0.19 $Y=1.66 $X2=2.19 $Y2=0.74
cc_142 VPB N_VPWR_c_776_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.355
cc_143 VPB N_VPWR_c_777_n 0.0602951f $X=-0.19 $Y=1.66 $X2=3.395 $Y2=1.92
cc_144 VPB N_VPWR_c_778_n 0.0320405f $X=-0.19 $Y=1.66 $X2=5.4 $Y2=2.105
cc_145 VPB N_VPWR_c_766_n 0.0916216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_780_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_781_n 0.0061274f $X=-0.19 $Y=1.66 $X2=3.395 $Y2=1.015
cc_148 VPB N_VPWR_c_782_n 0.00601668f $X=-0.19 $Y=1.66 $X2=3.41 $Y2=2.095
cc_149 VPB N_X_c_874_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.74
cc_150 VPB N_X_c_875_n 0.00630005f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.28
cc_151 VPB N_X_c_876_n 0.00327433f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_152 VPB N_A_537_388#_c_938_n 0.00832858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_961_392#_c_955_n 0.0103475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_961_392#_c_956_n 0.0185484f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.355
cc_155 VPB N_A_961_392#_c_957_n 0.0188649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_961_392#_c_958_n 0.00704942f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.74
cc_157 VPB N_A_1237_392#_c_1006_n 0.00249696f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_158 N_A_83_256#_c_169_n N_B1_c_328_n 0.00426339f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_159 N_A_83_256#_c_170_n N_B1_c_328_n 0.00402633f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_160 N_A_83_256#_c_172_n N_B1_c_328_n 0.005066f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_161 N_A_83_256#_c_174_n N_B1_c_328_n 0.00305315f $X=2.27 $Y=1.195 $X2=0 $Y2=0
cc_162 N_A_83_256#_c_170_n N_B1_c_329_n 0.00795139f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_163 N_A_83_256#_M1027_g N_B1_c_330_n 0.00426339f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_83_256#_c_170_n N_B1_c_330_n 0.00748939f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_165 N_A_83_256#_c_171_n N_B1_c_331_n 0.00255236f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_166 N_A_83_256#_c_171_n N_B1_c_332_n 0.0172734f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_167 N_A_83_256#_c_173_n N_B1_c_332_n 0.00201739f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_168 N_A_83_256#_c_171_n N_B1_c_333_n 0.00114575f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_169 N_A_83_256#_c_192_p N_B1_c_333_n 0.00559119f $X=3.395 $Y=0.81 $X2=0 $Y2=0
cc_170 N_A_83_256#_c_173_n N_B1_c_333_n 0.00713217f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_171 N_A_83_256#_c_172_n N_B1_c_340_n 9.80842e-19 $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_172 N_A_83_256#_c_180_n N_B1_c_340_n 0.0119257f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_173 N_A_83_256#_c_180_n N_B1_c_343_n 0.0114978f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_174 N_A_83_256#_c_170_n N_B1_c_334_n 0.00724703f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_175 N_A_83_256#_c_171_n N_B1_c_334_n 0.0020413f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_176 N_A_83_256#_c_172_n N_B1_c_344_n 0.0170906f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_177 N_A_83_256#_M1016_d N_B1_c_345_n 0.00318494f $X=3.275 $Y=1.94 $X2=0 $Y2=0
cc_178 N_A_83_256#_M1000_s N_B1_c_345_n 0.0037193f $X=5.265 $Y=1.96 $X2=0 $Y2=0
cc_179 N_A_83_256#_c_172_n N_B1_c_345_n 0.0181197f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_180 N_A_83_256#_c_180_n N_B1_c_345_n 0.116747f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_181 N_A_83_256#_c_180_n N_B1_c_346_n 0.0472823f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_182 N_A_83_256#_c_173_n N_B1_c_335_n 0.00281519f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_183 N_A_83_256#_c_180_n N_B1_c_335_n 0.0252946f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_184 N_A_83_256#_c_180_n N_B1_c_336_n 0.00104009f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_185 N_A_83_256#_M1009_g N_B1_c_337_n 0.0243597f $X=2.025 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A_83_256#_c_169_n N_B1_c_337_n 0.00847396f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_187 N_A_83_256#_c_170_n N_B1_c_337_n 0.00549621f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_188 N_A_83_256#_c_172_n N_B1_c_337_n 0.00128966f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_189 N_A_83_256#_c_174_n N_B1_c_337_n 9.65797e-19 $X=2.27 $Y=1.195 $X2=0 $Y2=0
cc_190 N_A_83_256#_M1009_g N_B1_c_338_n 9.61267e-19 $X=2.025 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_83_256#_c_170_n N_B1_c_338_n 0.0242401f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_192 N_A_83_256#_c_172_n N_B1_c_338_n 0.0141794f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_193 N_A_83_256#_c_174_n N_B1_c_338_n 0.0120085f $X=2.27 $Y=1.195 $X2=0 $Y2=0
cc_194 N_A_83_256#_c_172_n N_B2_c_480_n 0.00702087f $X=3.395 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_83_256#_c_172_n N_B2_c_481_n 0.0102798f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_196 N_A_83_256#_c_170_n N_B2_c_482_n 0.00239007f $X=3.23 $Y=1.195 $X2=0 $Y2=0
cc_197 N_A_83_256#_c_172_n N_B2_c_482_n 0.00330886f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_198 N_A_83_256#_c_172_n N_B2_c_472_n 0.0134504f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_199 N_A_83_256#_c_173_n N_B2_c_472_n 0.00770389f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_200 N_A_83_256#_c_180_n N_B2_c_472_n 0.0125999f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_201 N_A_83_256#_c_180_n N_B2_c_473_n 0.00507783f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_202 N_A_83_256#_c_192_p N_B2_c_474_n 4.63525e-19 $X=3.395 $Y=0.81 $X2=0 $Y2=0
cc_203 N_A_83_256#_c_173_n N_B2_c_474_n 0.0101141f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_204 N_A_83_256#_c_173_n N_B2_c_475_n 0.0154786f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_205 N_A_83_256#_c_173_n N_B2_c_476_n 0.00371982f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_206 N_A_83_256#_c_229_p N_B2_c_476_n 0.00399613f $X=4.395 $Y=0.81 $X2=0 $Y2=0
cc_207 N_A_83_256#_c_171_n N_B2_c_477_n 8.09549e-19 $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_208 N_A_83_256#_c_173_n N_B2_c_477_n 0.00676917f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_209 N_A_83_256#_c_171_n N_B2_c_478_n 0.00127419f $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_210 N_A_83_256#_c_172_n N_B2_c_478_n 0.00337625f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_211 N_A_83_256#_c_171_n N_B2_c_479_n 4.77843e-19 $X=3.395 $Y=1.28 $X2=0 $Y2=0
cc_212 N_A_83_256#_c_172_n N_B2_c_479_n 0.0228292f $X=3.395 $Y=1.92 $X2=0 $Y2=0
cc_213 N_A_83_256#_c_173_n N_B2_c_479_n 0.0245197f $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_214 N_A_83_256#_c_180_n N_B2_c_479_n 0.0171032f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_215 N_A_83_256#_c_173_n N_A3_M1002_g 4.24543e-19 $X=4.23 $Y=1.015 $X2=0 $Y2=0
cc_216 N_A_83_256#_c_180_n N_A3_M1000_g 0.0101026f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_217 N_A_83_256#_c_180_n N_A3_c_556_n 0.00189694f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_218 N_A_83_256#_c_180_n N_VPWR_M1023_s 0.0128712f $X=5.4 $Y=2.105 $X2=0 $Y2=0
cc_219 N_A_83_256#_M1003_g N_VPWR_c_768_n 0.00649215f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_220 N_A_83_256#_M1006_g N_VPWR_c_769_n 0.00408927f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_221 N_A_83_256#_M1008_g N_VPWR_c_769_n 0.0161497f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_83_256#_M1009_g N_VPWR_c_769_n 6.81855e-19 $X=2.025 $Y=2.4 $X2=0
+ $Y2=0
cc_223 N_A_83_256#_M1008_g N_VPWR_c_770_n 0.00460063f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_83_256#_M1009_g N_VPWR_c_770_n 0.00460063f $X=2.025 $Y=2.4 $X2=0
+ $Y2=0
cc_225 N_A_83_256#_M1008_g N_VPWR_c_771_n 7.38863e-19 $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_226 N_A_83_256#_M1009_g N_VPWR_c_771_n 0.0174992f $X=2.025 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_83_256#_c_168_n N_VPWR_c_771_n 0.00316131f $X=2.185 $Y=1.445 $X2=0
+ $Y2=0
cc_228 N_A_83_256#_c_169_n N_VPWR_c_771_n 0.00207532f $X=2.1 $Y=1.445 $X2=0
+ $Y2=0
cc_229 N_A_83_256#_c_170_n N_VPWR_c_771_n 0.00179271f $X=3.23 $Y=1.195 $X2=0
+ $Y2=0
cc_230 N_A_83_256#_c_174_n N_VPWR_c_771_n 0.00880609f $X=2.27 $Y=1.195 $X2=0
+ $Y2=0
cc_231 N_A_83_256#_M1003_g N_VPWR_c_776_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_83_256#_M1006_g N_VPWR_c_776_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_83_256#_M1003_g N_VPWR_c_766_n 0.00986008f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_234 N_A_83_256#_M1006_g N_VPWR_c_766_n 0.00982082f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_235 N_A_83_256#_M1008_g N_VPWR_c_766_n 0.00909652f $X=1.455 $Y=2.4 $X2=0
+ $Y2=0
cc_236 N_A_83_256#_M1009_g N_VPWR_c_766_n 0.00909652f $X=2.025 $Y=2.4 $X2=0
+ $Y2=0
cc_237 N_A_83_256#_M1015_g N_X_c_865_n 0.0109683f $X=0.635 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_83_256#_c_167_n N_X_c_865_n 0.00706368f $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_239 N_A_83_256#_M1003_g N_X_c_866_n 0.0150931f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A_83_256#_M1003_g N_X_c_874_n 0.0139766f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_83_256#_M1006_g N_X_c_874_n 0.0143169f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A_83_256#_M1008_g N_X_c_874_n 2.74397e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_83_256#_M1015_g N_X_c_868_n 0.00746201f $X=0.635 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_83_256#_M1020_g N_X_c_868_n 0.00896067f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_83_256#_M1024_g N_X_c_868_n 6.1951e-19 $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_83_256#_M1006_g N_X_c_875_n 0.0158148f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_83_256#_M1008_g N_X_c_875_n 0.0153525f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_83_256#_M1009_g N_X_c_875_n 0.0026697f $X=2.025 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_83_256#_c_168_n N_X_c_875_n 0.0504197f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_250 N_A_83_256#_c_169_n N_X_c_875_n 0.0131384f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_251 N_A_83_256#_M1020_g N_X_c_869_n 0.014323f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_83_256#_M1024_g N_X_c_869_n 0.0126012f $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_83_256#_M1027_g N_X_c_869_n 0.00533726f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_83_256#_c_168_n N_X_c_869_n 0.0539257f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_255 N_A_83_256#_c_169_n N_X_c_869_n 0.0115136f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_256 N_A_83_256#_M1008_g N_X_c_876_n 5.04913e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A_83_256#_M1009_g N_X_c_876_n 0.0062654f $X=2.025 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A_83_256#_M1020_g N_X_c_870_n 6.14947e-19 $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_83_256#_M1024_g N_X_c_870_n 0.00878544f $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_83_256#_M1027_g N_X_c_870_n 0.00535397f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_83_256#_M1003_g N_X_c_871_n 0.014668f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_83_256#_M1006_g N_X_c_871_n 0.0108224f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A_83_256#_M1008_g N_X_c_871_n 0.00132923f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_83_256#_c_167_n N_X_c_871_n 0.0028273f $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_265 N_A_83_256#_c_168_n N_X_c_871_n 0.00562369f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_266 N_A_83_256#_M1015_g N_X_c_906_n 0.0104872f $X=0.635 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_83_256#_c_160_n N_X_c_906_n 0.00361547f $X=0.865 $Y=1.355 $X2=0 $Y2=0
cc_268 N_A_83_256#_M1020_g N_X_c_906_n 0.00636589f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_83_256#_M1024_g N_X_c_906_n 8.53592e-19 $X=1.635 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_83_256#_c_167_n N_X_c_906_n 3.57967e-19 $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_271 N_A_83_256#_c_168_n N_X_c_906_n 0.00175494f $X=2.185 $Y=1.445 $X2=0 $Y2=0
cc_272 N_A_83_256#_c_169_n N_X_c_906_n 0.00487067f $X=2.1 $Y=1.445 $X2=0 $Y2=0
cc_273 N_A_83_256#_c_167_n X 0.00776373f $X=0.562 $Y=1.355 $X2=0 $Y2=0
cc_274 N_A_83_256#_c_180_n N_A_537_388#_M1019_s 0.00385416f $X=5.4 $Y=2.105
+ $X2=0 $Y2=0
cc_275 N_A_83_256#_M1016_d N_A_537_388#_c_938_n 0.00168426f $X=3.275 $Y=1.94
+ $X2=0 $Y2=0
cc_276 N_A_83_256#_c_180_n N_A_961_392#_M1000_d 0.0047023f $X=5.4 $Y=2.105
+ $X2=-0.19 $Y2=-0.245
cc_277 N_A_83_256#_M1000_s N_A_961_392#_c_955_n 0.00190453f $X=5.265 $Y=1.96
+ $X2=0 $Y2=0
cc_278 N_A_83_256#_c_174_n N_VGND_M1027_s 9.75702e-19 $X=2.27 $Y=1.195 $X2=0
+ $Y2=0
cc_279 N_A_83_256#_M1015_g N_VGND_c_1028_n 0.0153292f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_83_256#_c_167_n N_VGND_c_1028_n 5.27357e-19 $X=0.562 $Y=1.355 $X2=0
+ $Y2=0
cc_281 N_A_83_256#_M1015_g N_VGND_c_1029_n 0.00434272f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_83_256#_M1020_g N_VGND_c_1029_n 0.00434272f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_83_256#_M1020_g N_VGND_c_1030_n 0.00441895f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_83_256#_M1024_g N_VGND_c_1030_n 0.00580088f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_83_256#_M1024_g N_VGND_c_1031_n 7.01214e-19 $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_83_256#_M1027_g N_VGND_c_1031_n 0.0125112f $X=2.19 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_83_256#_c_170_n N_VGND_c_1031_n 0.0177292f $X=3.23 $Y=1.195 $X2=0
+ $Y2=0
cc_288 N_A_83_256#_c_174_n N_VGND_c_1031_n 0.00721878f $X=2.27 $Y=1.195 $X2=0
+ $Y2=0
cc_289 N_A_83_256#_M1024_g N_VGND_c_1035_n 0.00434272f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_290 N_A_83_256#_M1027_g N_VGND_c_1035_n 0.00383152f $X=2.19 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_83_256#_M1015_g N_VGND_c_1043_n 0.00824109f $X=0.635 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_83_256#_M1020_g N_VGND_c_1043_n 0.00821294f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_83_256#_M1024_g N_VGND_c_1043_n 0.0082241f $X=1.635 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_83_256#_M1027_g N_VGND_c_1043_n 0.00758657f $X=2.19 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_83_256#_c_173_n N_A_564_74#_M1025_s 0.00250873f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_296 N_A_83_256#_c_170_n N_A_564_74#_c_1134_n 0.0232013f $X=3.23 $Y=1.195
+ $X2=0 $Y2=0
cc_297 N_A_83_256#_M1010_d N_A_564_74#_c_1135_n 0.00168861f $X=3.255 $Y=0.37
+ $X2=0 $Y2=0
cc_298 N_A_83_256#_c_192_p N_A_564_74#_c_1135_n 0.0143448f $X=3.395 $Y=0.81
+ $X2=0 $Y2=0
cc_299 N_A_83_256#_c_173_n N_A_564_74#_c_1135_n 0.00347117f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_300 N_A_83_256#_M1027_g N_A_564_74#_c_1136_n 6.04331e-19 $X=2.19 $Y=0.74
+ $X2=0 $Y2=0
cc_301 N_A_83_256#_c_173_n N_A_564_74#_c_1150_n 0.0204865f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_302 N_A_83_256#_M1021_s N_A_564_74#_c_1137_n 0.00237953f $X=4.185 $Y=0.37
+ $X2=0 $Y2=0
cc_303 N_A_83_256#_c_173_n N_A_564_74#_c_1137_n 0.00347117f $X=4.23 $Y=1.015
+ $X2=0 $Y2=0
cc_304 N_A_83_256#_c_229_p N_A_564_74#_c_1137_n 0.0192294f $X=4.395 $Y=0.81
+ $X2=0 $Y2=0
cc_305 N_B1_c_345_n N_B2_c_480_n 0.0162379f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_306 N_B1_c_334_n N_B2_c_481_n 0.00350641f $X=3.18 $Y=1.165 $X2=0 $Y2=0
cc_307 N_B1_c_345_n N_B2_c_481_n 3.18712e-19 $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_308 N_B1_M1018_g N_B2_c_482_n 0.0330641f $X=2.595 $Y=2.44 $X2=0 $Y2=0
cc_309 N_B1_c_329_n N_B2_c_482_n 0.00350641f $X=3.105 $Y=1.165 $X2=0 $Y2=0
cc_310 N_B1_c_344_n N_B2_c_482_n 0.00689805f $X=2.77 $Y=2.36 $X2=0 $Y2=0
cc_311 N_B1_c_337_n N_B2_c_482_n 0.00365659f $X=2.78 $Y=1.615 $X2=0 $Y2=0
cc_312 N_B1_c_338_n N_B2_c_482_n 2.86983e-19 $X=2.77 $Y=1.615 $X2=0 $Y2=0
cc_313 N_B1_c_332_n N_B2_c_472_n 0.0120737f $X=3.535 $Y=1.165 $X2=0 $Y2=0
cc_314 N_B1_c_340_n N_B2_c_472_n 0.0460345f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_315 N_B1_c_345_n N_B2_c_472_n 0.011587f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_316 N_B1_c_337_n N_B2_c_472_n 0.00236341f $X=2.78 $Y=1.615 $X2=0 $Y2=0
cc_317 N_B1_c_340_n N_B2_c_473_n 0.0118f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_318 N_B1_c_335_n N_B2_c_473_n 6.33942e-19 $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_319 N_B1_c_336_n N_B2_c_473_n 0.00821351f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_320 N_B1_c_333_n N_B2_c_474_n 0.0203621f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_321 N_B1_c_335_n N_B2_c_475_n 0.00123953f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_322 N_B1_c_336_n N_B2_c_475_n 0.0126816f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_323 N_B1_c_332_n N_B2_c_477_n 0.0100546f $X=3.535 $Y=1.165 $X2=0 $Y2=0
cc_324 N_B1_c_340_n N_B2_c_479_n 0.00181036f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_325 N_B1_c_335_n N_B2_c_479_n 0.0195613f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_326 N_B1_c_336_n N_B2_c_479_n 0.00447962f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_327 N_B1_c_343_n N_A3_M1000_g 0.0409389f $X=4.655 $Y=3.015 $X2=0 $Y2=0
cc_328 N_B1_c_345_n N_A3_M1000_g 0.0121608f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_329 N_B1_c_346_n N_A3_M1000_g 0.0117387f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_330 N_B1_c_335_n N_A3_M1000_g 0.0012304f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_331 N_B1_c_336_n N_A3_M1000_g 0.0137874f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_332 N_B1_c_345_n N_A3_c_556_n 0.0128614f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_333 N_B1_c_346_n N_A3_c_556_n 0.00830783f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_334 N_B1_c_347_n N_A3_c_556_n 0.00468894f $X=5.82 $Y=2.36 $X2=0 $Y2=0
cc_335 N_B1_c_346_n N_A3_c_552_n 0.00442139f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_336 N_B1_c_346_n A3 0.0490884f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_337 N_B1_c_335_n A3 0.0035661f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_338 N_B1_c_336_n A3 2.16867e-19 $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_339 N_B1_c_346_n N_A3_c_554_n 0.00366609f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_340 N_B1_c_336_n N_A3_c_554_n 0.00323048f $X=4.66 $Y=1.615 $X2=0 $Y2=0
cc_341 N_B1_c_345_n N_A2_M1001_g 0.0019322f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_342 N_B1_c_347_n N_A2_M1001_g 0.00772651f $X=5.82 $Y=2.36 $X2=0 $Y2=0
cc_343 N_B1_c_346_n N_A2_c_615_n 0.00247363f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_344 N_B1_c_346_n A2 0.0106093f $X=5.735 $Y=1.765 $X2=0 $Y2=0
cc_345 N_B1_c_345_n N_VPWR_M1023_s 0.00590078f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_346 N_B1_M1018_g N_VPWR_c_771_n 0.0160063f $X=2.595 $Y=2.44 $X2=0 $Y2=0
cc_347 N_B1_c_430_p N_VPWR_c_771_n 0.00980088f $X=2.855 $Y=2.445 $X2=0 $Y2=0
cc_348 N_B1_c_340_n N_VPWR_c_772_n 0.00187364f $X=4.085 $Y=3.015 $X2=0 $Y2=0
cc_349 N_B1_c_341_n N_VPWR_c_772_n 0.0217307f $X=4.58 $Y=3.09 $X2=0 $Y2=0
cc_350 N_B1_c_343_n N_VPWR_c_772_n 0.00397506f $X=4.655 $Y=3.015 $X2=0 $Y2=0
cc_351 N_B1_c_345_n N_VPWR_c_772_n 0.0233068f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_352 N_B1_M1018_g N_VPWR_c_774_n 0.00643693f $X=2.595 $Y=2.44 $X2=0 $Y2=0
cc_353 N_B1_c_342_n N_VPWR_c_774_n 0.00661248f $X=4.175 $Y=3.09 $X2=0 $Y2=0
cc_354 N_B1_c_341_n N_VPWR_c_777_n 0.00716255f $X=4.58 $Y=3.09 $X2=0 $Y2=0
cc_355 N_B1_M1018_g N_VPWR_c_766_n 0.00647345f $X=2.595 $Y=2.44 $X2=0 $Y2=0
cc_356 N_B1_c_341_n N_VPWR_c_766_n 0.00812355f $X=4.58 $Y=3.09 $X2=0 $Y2=0
cc_357 N_B1_c_342_n N_VPWR_c_766_n 0.00668088f $X=4.175 $Y=3.09 $X2=0 $Y2=0
cc_358 N_B1_c_345_n N_VPWR_c_766_n 0.0170232f $X=5.735 $Y=2.445 $X2=0 $Y2=0
cc_359 N_B1_c_344_n N_A_537_388#_M1018_d 0.00752828f $X=2.77 $Y=2.36 $X2=-0.19
+ $Y2=-0.245
cc_360 N_B1_c_345_n N_A_537_388#_M1018_d 0.00939564f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_361 N_B1_c_430_p N_A_537_388#_M1018_d 0.00222845f $X=2.855 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_362 N_B1_c_345_n N_A_537_388#_M1019_s 0.00329665f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_363 N_B1_M1018_g N_A_537_388#_c_938_n 0.00913144f $X=2.595 $Y=2.44 $X2=0
+ $Y2=0
cc_364 N_B1_c_340_n N_A_537_388#_c_938_n 0.00393571f $X=4.085 $Y=3.015 $X2=0
+ $Y2=0
cc_365 N_B1_c_345_n N_A_537_388#_c_938_n 0.0624821f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_366 N_B1_c_430_p N_A_537_388#_c_938_n 0.0091325f $X=2.855 $Y=2.445 $X2=0
+ $Y2=0
cc_367 N_B1_c_345_n N_A_961_392#_M1000_d 0.00468357f $X=5.735 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_368 N_B1_c_345_n N_A_961_392#_M1017_d 0.00280996f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_369 N_B1_c_347_n N_A_961_392#_M1017_d 0.00499256f $X=5.82 $Y=2.36 $X2=0 $Y2=0
cc_370 N_B1_c_343_n N_A_961_392#_c_955_n 0.00301582f $X=4.655 $Y=3.015 $X2=0
+ $Y2=0
cc_371 N_B1_c_345_n N_A_961_392#_c_955_n 0.0645321f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_372 N_B1_c_345_n N_A_961_392#_c_966_n 0.0122365f $X=5.735 $Y=2.445 $X2=0
+ $Y2=0
cc_373 N_B1_c_347_n N_A_1237_392#_c_1007_n 0.0144374f $X=5.82 $Y=2.36 $X2=0
+ $Y2=0
cc_374 N_B1_c_331_n N_VGND_c_1031_n 0.00176715f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_375 N_B1_c_331_n N_VGND_c_1037_n 0.00278247f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_376 N_B1_c_333_n N_VGND_c_1037_n 0.00278271f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_377 N_B1_c_331_n N_VGND_c_1043_n 0.00358425f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_378 N_B1_c_333_n N_VGND_c_1043_n 0.0035414f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_379 N_B1_c_330_n N_A_564_74#_c_1134_n 0.00638349f $X=2.855 $Y=1.165 $X2=0
+ $Y2=0
cc_380 N_B1_c_331_n N_A_564_74#_c_1134_n 0.00694622f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_381 N_B1_c_333_n N_A_564_74#_c_1134_n 6.20636e-19 $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_382 N_B1_c_331_n N_A_564_74#_c_1135_n 0.0100711f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_383 N_B1_c_332_n N_A_564_74#_c_1135_n 2.67777e-19 $X=3.535 $Y=1.165 $X2=0
+ $Y2=0
cc_384 N_B1_c_333_n N_A_564_74#_c_1135_n 0.0109066f $X=3.61 $Y=1.09 $X2=0 $Y2=0
cc_385 N_B1_c_331_n N_A_564_74#_c_1136_n 0.00281658f $X=3.18 $Y=1.09 $X2=0 $Y2=0
cc_386 N_B1_c_346_n N_A_564_74#_c_1138_n 0.0063124f $X=5.735 $Y=1.765 $X2=0
+ $Y2=0
cc_387 N_B1_c_335_n N_A_564_74#_c_1138_n 0.00351334f $X=4.66 $Y=1.615 $X2=0
+ $Y2=0
cc_388 N_B1_c_336_n N_A_564_74#_c_1138_n 5.96818e-19 $X=4.66 $Y=1.615 $X2=0
+ $Y2=0
cc_389 N_B2_c_476_n N_A3_M1002_g 0.00961692f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_390 N_B2_c_475_n A3 4.16793e-19 $X=4.535 $Y=1.165 $X2=0 $Y2=0
cc_391 N_B2_c_475_n N_A3_c_554_n 0.00961692f $X=4.535 $Y=1.165 $X2=0 $Y2=0
cc_392 N_B2_c_472_n N_VPWR_c_772_n 2.39237e-19 $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_393 N_B2_c_480_n N_VPWR_c_774_n 0.00481634f $X=3.185 $Y=1.865 $X2=0 $Y2=0
cc_394 N_B2_c_472_n N_VPWR_c_774_n 0.00481634f $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_395 N_B2_c_480_n N_VPWR_c_766_n 0.00647345f $X=3.185 $Y=1.865 $X2=0 $Y2=0
cc_396 N_B2_c_472_n N_VPWR_c_766_n 0.00647345f $X=3.635 $Y=1.865 $X2=0 $Y2=0
cc_397 N_B2_c_480_n N_A_537_388#_c_938_n 0.0157486f $X=3.185 $Y=1.865 $X2=0
+ $Y2=0
cc_398 N_B2_c_472_n N_A_537_388#_c_938_n 0.0118809f $X=3.635 $Y=1.865 $X2=0
+ $Y2=0
cc_399 N_B2_c_474_n N_VGND_c_1037_n 0.00278247f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_400 N_B2_c_476_n N_VGND_c_1037_n 0.00278271f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_401 N_B2_c_474_n N_VGND_c_1043_n 0.00354796f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_402 N_B2_c_476_n N_VGND_c_1043_n 0.00355038f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_403 N_B2_c_474_n N_A_564_74#_c_1150_n 0.00539089f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_404 N_B2_c_476_n N_A_564_74#_c_1150_n 5.81199e-19 $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_405 N_B2_c_477_n N_A_564_74#_c_1150_n 4.55305e-19 $X=4.09 $Y=1.165 $X2=0
+ $Y2=0
cc_406 N_B2_c_474_n N_A_564_74#_c_1137_n 0.00806723f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_407 N_B2_c_475_n N_A_564_74#_c_1137_n 4.55221e-19 $X=4.535 $Y=1.165 $X2=0
+ $Y2=0
cc_408 N_B2_c_476_n N_A_564_74#_c_1137_n 0.0137079f $X=4.61 $Y=1.09 $X2=0 $Y2=0
cc_409 N_B2_c_474_n N_A_564_74#_c_1143_n 0.00253515f $X=4.11 $Y=1.09 $X2=0 $Y2=0
cc_410 N_A3_c_556_n N_A2_M1001_g 0.0178657f $X=5.645 $Y=1.84 $X2=0 $Y2=0
cc_411 N_A3_M1012_g N_A2_c_612_n 0.0110549f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_412 N_A3_M1012_g N_A2_c_614_n 0.0178657f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_413 A3 N_A2_c_614_n 0.00137288f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_414 N_A3_c_552_n N_A2_c_615_n 0.0178657f $X=5.645 $Y=1.75 $X2=0 $Y2=0
cc_415 N_A3_c_552_n A2 6.38672e-19 $X=5.645 $Y=1.75 $X2=0 $Y2=0
cc_416 N_A3_c_554_n N_A2_c_617_n 0.0178657f $X=5.66 $Y=1.345 $X2=0 $Y2=0
cc_417 N_A3_M1012_g N_A2_c_638_n 2.7656e-19 $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_418 A3 N_A2_c_638_n 0.0149466f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_419 N_A3_c_554_n N_A2_c_638_n 7.57327e-19 $X=5.66 $Y=1.345 $X2=0 $Y2=0
cc_420 N_A3_M1000_g N_VPWR_c_772_n 3.24475e-19 $X=5.175 $Y=2.46 $X2=0 $Y2=0
cc_421 N_A3_M1000_g N_VPWR_c_777_n 0.00349978f $X=5.175 $Y=2.46 $X2=0 $Y2=0
cc_422 N_A3_c_556_n N_VPWR_c_777_n 0.00349978f $X=5.645 $Y=1.84 $X2=0 $Y2=0
cc_423 N_A3_M1000_g N_VPWR_c_766_n 0.00430581f $X=5.175 $Y=2.46 $X2=0 $Y2=0
cc_424 N_A3_c_556_n N_VPWR_c_766_n 0.0042983f $X=5.645 $Y=1.84 $X2=0 $Y2=0
cc_425 N_A3_M1000_g N_A_961_392#_c_955_n 0.0126119f $X=5.175 $Y=2.46 $X2=0 $Y2=0
cc_426 N_A3_c_556_n N_A_961_392#_c_955_n 0.0125993f $X=5.645 $Y=1.84 $X2=0 $Y2=0
cc_427 N_A3_c_556_n N_A_961_392#_c_969_n 5.45521e-19 $X=5.645 $Y=1.84 $X2=0
+ $Y2=0
cc_428 N_A3_c_556_n N_A_961_392#_c_966_n 2.84049e-19 $X=5.645 $Y=1.84 $X2=0
+ $Y2=0
cc_429 N_A3_M1002_g N_VGND_c_1032_n 0.00148871f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_430 N_A3_M1012_g N_VGND_c_1032_n 0.00198878f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_431 N_A3_M1002_g N_VGND_c_1037_n 0.00461464f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_432 N_A3_M1012_g N_VGND_c_1039_n 0.00456932f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_433 N_A3_M1002_g N_VGND_c_1043_n 0.00451999f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_434 N_A3_M1012_g N_VGND_c_1043_n 0.00443718f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_435 N_A3_M1002_g N_A_564_74#_c_1137_n 0.00118927f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_436 N_A3_M1002_g N_A_564_74#_c_1172_n 0.0104635f $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_437 N_A3_M1012_g N_A_564_74#_c_1172_n 0.0101963f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_438 A3 N_A_564_74#_c_1172_n 0.036068f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_439 N_A3_c_554_n N_A_564_74#_c_1172_n 0.00430721f $X=5.66 $Y=1.345 $X2=0
+ $Y2=0
cc_440 N_A3_M1002_g N_A_564_74#_c_1139_n 3.11133e-19 $X=5.14 $Y=0.69 $X2=0 $Y2=0
cc_441 N_A3_M1012_g N_A_564_74#_c_1139_n 0.00560871f $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_442 N_A3_M1012_g N_A_564_74#_c_1178_n 2.51849e-19 $X=5.66 $Y=0.69 $X2=0 $Y2=0
cc_443 A3 N_A_564_74#_c_1178_n 2.88494e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_444 N_A2_c_613_n N_A1_c_704_n 0.00828772f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_445 N_A2_M1001_g N_A1_c_711_n 0.0330586f $X=6.095 $Y=2.46 $X2=0 $Y2=0
cc_446 N_A2_M1013_g N_A1_c_711_n 0.0312188f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_447 N_A2_c_614_n N_A1_c_711_n 8.18936e-19 $X=6.205 $Y=1.235 $X2=0 $Y2=0
cc_448 N_A2_c_615_n N_A1_c_711_n 0.00361947f $X=6.205 $Y=1.8 $X2=0 $Y2=0
cc_449 N_A2_c_619_n N_A1_c_711_n 0.0178069f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_450 A2 N_A1_c_705_n 8.24499e-19 $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_451 N_A2_c_618_n N_A1_c_705_n 0.012571f $X=7.73 $Y=1.615 $X2=0 $Y2=0
cc_452 N_A2_c_619_n N_A1_c_705_n 0.00558949f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_453 N_A2_c_614_n N_A1_c_707_n 0.00828772f $X=6.205 $Y=1.235 $X2=0 $Y2=0
cc_454 N_A2_c_617_n N_A1_c_707_n 0.00478184f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_455 N_A2_c_638_n N_A1_c_707_n 2.55438e-19 $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_456 N_A2_c_615_n N_A1_c_708_n 0.00478184f $X=6.205 $Y=1.8 $X2=0 $Y2=0
cc_457 A2 N_A1_c_708_n 8.80533e-19 $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_458 N_A2_c_638_n N_A1_c_708_n 9.78829e-19 $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_459 N_A2_c_618_n N_A1_c_708_n 0.0312188f $X=7.73 $Y=1.615 $X2=0 $Y2=0
cc_460 N_A2_c_619_n N_A1_c_708_n 0.0139494f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_461 N_A2_c_614_n N_A1_c_709_n 0.00142867f $X=6.205 $Y=1.235 $X2=0 $Y2=0
cc_462 N_A2_c_617_n N_A1_c_709_n 0.00149364f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_463 N_A2_c_638_n N_A1_c_709_n 0.0111493f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_464 N_A2_c_619_n N_A1_c_709_n 0.0331366f $X=7.565 $Y=1.615 $X2=0 $Y2=0
cc_465 N_A2_M1001_g N_VPWR_c_773_n 7.10865e-19 $X=6.095 $Y=2.46 $X2=0 $Y2=0
cc_466 N_A2_M1013_g N_VPWR_c_773_n 0.00124657f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_467 N_A2_M1001_g N_VPWR_c_777_n 0.00349879f $X=6.095 $Y=2.46 $X2=0 $Y2=0
cc_468 N_A2_M1013_g N_VPWR_c_778_n 0.005209f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_469 N_A2_M1001_g N_VPWR_c_766_n 0.00431195f $X=6.095 $Y=2.46 $X2=0 $Y2=0
cc_470 N_A2_M1013_g N_VPWR_c_766_n 0.00520375f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_471 N_A2_M1001_g N_A_961_392#_c_955_n 0.0121899f $X=6.095 $Y=2.46 $X2=0 $Y2=0
cc_472 N_A2_M1001_g N_A_961_392#_c_969_n 0.00447932f $X=6.095 $Y=2.46 $X2=0
+ $Y2=0
cc_473 N_A2_M1013_g N_A_961_392#_c_973_n 0.0111746f $X=7.655 $Y=2.46 $X2=0 $Y2=0
cc_474 A2 N_A_961_392#_c_973_n 0.00296232f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_475 N_A2_M1001_g N_A_961_392#_c_966_n 0.00870602f $X=6.095 $Y=2.46 $X2=0
+ $Y2=0
cc_476 A2 N_A_961_392#_c_966_n 0.00237965f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_477 N_A2_M1013_g N_A_961_392#_c_956_n 0.00872239f $X=7.655 $Y=2.46 $X2=0
+ $Y2=0
cc_478 N_A2_M1013_g N_A_961_392#_c_957_n 2.57198e-19 $X=7.655 $Y=2.46 $X2=0
+ $Y2=0
cc_479 A2 N_A_961_392#_c_957_n 0.0232636f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_480 N_A2_c_618_n N_A_961_392#_c_957_n 0.00300514f $X=7.73 $Y=1.615 $X2=0
+ $Y2=0
cc_481 N_A2_M1013_g N_A_961_392#_c_958_n 0.00128025f $X=7.655 $Y=2.46 $X2=0
+ $Y2=0
cc_482 A2 N_A_961_392#_c_958_n 0.00106598f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_483 N_A2_M1001_g N_A_1237_392#_c_1007_n 0.00825781f $X=6.095 $Y=2.46 $X2=0
+ $Y2=0
cc_484 N_A2_c_615_n N_A_1237_392#_c_1007_n 0.00143895f $X=6.205 $Y=1.8 $X2=0
+ $Y2=0
cc_485 A2 N_A_1237_392#_c_1007_n 0.0178903f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_486 N_A2_c_619_n N_A_1237_392#_c_1007_n 0.0515068f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_487 N_A2_M1013_g N_A_1237_392#_c_1006_n 0.00386013f $X=7.655 $Y=2.46 $X2=0
+ $Y2=0
cc_488 N_A2_c_619_n N_A_1237_392#_c_1006_n 0.0254857f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_489 N_A2_c_612_n N_VGND_c_1033_n 0.00312943f $X=6.11 $Y=1.085 $X2=0 $Y2=0
cc_490 N_A2_c_613_n N_VGND_c_1033_n 0.0070913f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_491 N_A2_c_612_n N_VGND_c_1039_n 0.00434272f $X=6.11 $Y=1.085 $X2=0 $Y2=0
cc_492 N_A2_c_613_n N_VGND_c_1041_n 0.00383152f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_493 N_A2_c_612_n N_VGND_c_1043_n 0.00433282f $X=6.11 $Y=1.085 $X2=0 $Y2=0
cc_494 N_A2_c_613_n N_VGND_c_1043_n 0.0037147f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_495 N_A2_c_612_n N_A_564_74#_c_1139_n 0.00639171f $X=6.11 $Y=1.085 $X2=0
+ $Y2=0
cc_496 N_A2_c_613_n N_A_564_74#_c_1139_n 6.25537e-19 $X=6.61 $Y=1.085 $X2=0
+ $Y2=0
cc_497 N_A2_c_612_n N_A_564_74#_c_1182_n 0.00925007f $X=6.11 $Y=1.085 $X2=0
+ $Y2=0
cc_498 N_A2_c_613_n N_A_564_74#_c_1182_n 0.0111557f $X=6.61 $Y=1.085 $X2=0 $Y2=0
cc_499 N_A2_c_614_n N_A_564_74#_c_1182_n 0.00458615f $X=6.205 $Y=1.235 $X2=0
+ $Y2=0
cc_500 N_A2_c_638_n N_A_564_74#_c_1182_n 0.0223703f $X=6.24 $Y=1.295 $X2=0 $Y2=0
cc_501 N_A2_c_619_n N_A_564_74#_c_1182_n 0.00783756f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_502 A2 N_A_564_74#_c_1141_n 0.0183141f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_503 N_A2_c_618_n N_A_564_74#_c_1141_n 0.00348736f $X=7.73 $Y=1.615 $X2=0
+ $Y2=0
cc_504 N_A2_c_619_n N_A_564_74#_c_1141_n 0.00735461f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_505 N_A2_c_612_n N_A_564_74#_c_1178_n 0.00177241f $X=6.11 $Y=1.085 $X2=0
+ $Y2=0
cc_506 N_A2_c_619_n N_A_564_74#_c_1191_n 0.00332297f $X=7.565 $Y=1.615 $X2=0
+ $Y2=0
cc_507 N_A1_c_710_n N_VPWR_c_773_n 0.00937862f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_508 N_A1_c_711_n N_VPWR_c_773_n 0.00893884f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_509 N_A1_c_710_n N_VPWR_c_777_n 0.00490827f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_510 N_A1_c_711_n N_VPWR_c_778_n 0.00490827f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_511 N_A1_c_710_n N_VPWR_c_766_n 0.00474288f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_512 N_A1_c_711_n N_VPWR_c_766_n 0.00472755f $X=7.205 $Y=1.885 $X2=0 $Y2=0
cc_513 N_A1_c_710_n N_A_961_392#_c_955_n 0.00299444f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_514 N_A1_c_710_n N_A_961_392#_c_969_n 0.00237013f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_515 N_A1_c_710_n N_A_961_392#_c_973_n 0.0140372f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_516 N_A1_c_711_n N_A_961_392#_c_973_n 0.0131476f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_517 N_A1_c_711_n N_A_961_392#_c_956_n 0.00154004f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_518 N_A1_c_710_n N_A_1237_392#_c_1014_n 0.00605775f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_519 N_A1_c_711_n N_A_1237_392#_c_1006_n 0.00193207f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_520 N_A1_c_710_n N_A_1237_392#_c_1016_n 0.0103835f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_521 N_A1_c_711_n N_A_1237_392#_c_1016_n 0.0132413f $X=7.205 $Y=1.885 $X2=0
+ $Y2=0
cc_522 N_A1_c_704_n N_VGND_c_1033_n 4.2194e-19 $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_523 N_A1_c_704_n N_VGND_c_1034_n 0.00356619f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_524 N_A1_c_706_n N_VGND_c_1034_n 0.00508961f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_525 N_A1_c_704_n N_VGND_c_1041_n 0.00434272f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_526 N_A1_c_706_n N_VGND_c_1042_n 0.00434272f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_527 N_A1_c_704_n N_VGND_c_1043_n 0.00434075f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_528 N_A1_c_706_n N_VGND_c_1043_n 0.00437635f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_529 N_A1_c_704_n N_A_564_74#_c_1140_n 0.00668866f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_530 N_A1_c_706_n N_A_564_74#_c_1140_n 8.41862e-19 $X=7.665 $Y=1.09 $X2=0
+ $Y2=0
cc_531 N_A1_c_704_n N_A_564_74#_c_1141_n 0.0096489f $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_532 N_A1_c_706_n N_A_564_74#_c_1141_n 0.0126914f $X=7.665 $Y=1.09 $X2=0 $Y2=0
cc_533 N_A1_c_707_n N_A_564_74#_c_1141_n 0.00748895f $X=7.13 $Y=1.165 $X2=0
+ $Y2=0
cc_534 N_A1_c_709_n N_A_564_74#_c_1141_n 0.0198892f $X=7.13 $Y=1.285 $X2=0 $Y2=0
cc_535 N_A1_c_704_n N_A_564_74#_c_1142_n 8.3913e-19 $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_536 N_A1_c_706_n N_A_564_74#_c_1142_n 0.00700896f $X=7.665 $Y=1.09 $X2=0
+ $Y2=0
cc_537 N_A1_c_704_n N_A_564_74#_c_1191_n 7.15802e-19 $X=7.04 $Y=1.09 $X2=0 $Y2=0
cc_538 N_A1_c_709_n N_A_564_74#_c_1191_n 0.00961222f $X=7.13 $Y=1.285 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_768_n N_X_c_866_n 7.22336e-19 $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_540 N_VPWR_c_768_n N_X_c_867_n 0.0210943f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_541 N_VPWR_c_769_n N_X_c_874_n 0.0330597f $X=1.23 $Y=2.285 $X2=0 $Y2=0
cc_542 N_VPWR_c_776_n N_X_c_874_n 0.0144623f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_c_766_n N_X_c_874_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_M1006_d N_X_c_875_n 0.00218982f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_545 N_VPWR_c_769_n N_X_c_875_n 0.0189268f $X=1.23 $Y=2.285 $X2=0 $Y2=0
cc_546 N_VPWR_c_769_n N_X_c_876_n 0.0330597f $X=1.23 $Y=2.285 $X2=0 $Y2=0
cc_547 N_VPWR_c_770_n N_X_c_876_n 0.0146357f $X=2.085 $Y=3.33 $X2=0 $Y2=0
cc_548 N_VPWR_c_771_n N_X_c_876_n 0.0360842f $X=2.25 $Y=2.115 $X2=0 $Y2=0
cc_549 N_VPWR_c_766_n N_X_c_876_n 0.0121141f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_550 N_VPWR_c_768_n N_X_c_871_n 0.0395357f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_551 N_VPWR_c_771_n N_A_537_388#_c_938_n 0.0163152f $X=2.25 $Y=2.115 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_772_n N_A_537_388#_c_938_n 0.01162f $X=4.36 $Y=2.79 $X2=0 $Y2=0
cc_553 N_VPWR_c_774_n N_A_537_388#_c_938_n 0.0515981f $X=4.195 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_766_n N_A_537_388#_c_938_n 0.0479151f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_772_n N_A_961_392#_c_955_n 0.0182355f $X=4.36 $Y=2.79 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_773_n N_A_961_392#_c_955_n 0.0081628f $X=6.97 $Y=2.815 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_777_n N_A_961_392#_c_955_n 0.0598406f $X=6.805 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_766_n N_A_961_392#_c_955_n 0.0499222f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_M1011_s N_A_961_392#_c_973_n 0.00366155f $X=6.825 $Y=1.96 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_773_n N_A_961_392#_c_973_n 0.0166493f $X=6.97 $Y=2.815 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_766_n N_A_961_392#_c_973_n 0.0396753f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_773_n N_A_961_392#_c_956_n 0.00681581f $X=6.97 $Y=2.815 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_778_n N_A_961_392#_c_956_n 0.0145282f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_766_n N_A_961_392#_c_956_n 0.0119657f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_M1011_s N_A_1237_392#_c_1016_n 0.00367556f $X=6.825 $Y=1.96 $X2=0
+ $Y2=0
cc_566 N_X_c_869_n N_VGND_M1020_s 0.00694709f $X=1.685 $Y=1.025 $X2=0 $Y2=0
cc_567 N_X_c_865_n N_VGND_c_1028_n 0.0126161f $X=0.685 $Y=1.225 $X2=0 $Y2=0
cc_568 N_X_c_868_n N_VGND_c_1028_n 0.0240168f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_569 N_X_c_873_n N_VGND_c_1028_n 0.0152345f $X=0.24 $Y=1.31 $X2=0 $Y2=0
cc_570 N_X_c_868_n N_VGND_c_1029_n 0.0144922f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_571 N_X_c_868_n N_VGND_c_1030_n 0.0165499f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_572 N_X_c_869_n N_VGND_c_1030_n 0.0248957f $X=1.685 $Y=1.025 $X2=0 $Y2=0
cc_573 N_X_c_870_n N_VGND_c_1030_n 0.0165499f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_574 N_X_c_870_n N_VGND_c_1031_n 0.0369264f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_575 N_X_c_870_n N_VGND_c_1035_n 0.0145639f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_576 N_X_c_868_n N_VGND_c_1043_n 0.0118826f $X=0.85 $Y=0.515 $X2=0 $Y2=0
cc_577 N_X_c_870_n N_VGND_c_1043_n 0.0119984f $X=1.85 $Y=0.515 $X2=0 $Y2=0
cc_578 N_A_961_392#_c_955_n N_A_1237_392#_M1001_d 0.00419731f $X=6.075 $Y=2.84
+ $X2=-0.19 $Y2=1.66
cc_579 N_A_961_392#_c_969_n N_A_1237_392#_M1001_d 0.00194297f $X=6.16 $Y=2.7
+ $X2=-0.19 $Y2=1.66
cc_580 N_A_961_392#_c_973_n N_A_1237_392#_M1001_d 0.0108847f $X=7.715 $Y=2.475
+ $X2=-0.19 $Y2=1.66
cc_581 N_A_961_392#_c_973_n N_A_1237_392#_M1026_d 0.00468888f $X=7.715 $Y=2.475
+ $X2=0 $Y2=0
cc_582 N_A_961_392#_c_973_n N_A_1237_392#_c_1007_n 0.0276746f $X=7.715 $Y=2.475
+ $X2=0 $Y2=0
cc_583 N_A_961_392#_c_966_n N_A_1237_392#_c_1007_n 0.0025684f $X=6.245 $Y=2.475
+ $X2=0 $Y2=0
cc_584 N_A_961_392#_c_957_n N_A_1237_392#_c_1006_n 0.0106894f $X=7.88 $Y=2.115
+ $X2=0 $Y2=0
cc_585 N_A_961_392#_c_973_n N_A_1237_392#_c_1016_n 0.0455325f $X=7.715 $Y=2.475
+ $X2=0 $Y2=0
cc_586 N_VGND_c_1031_n N_A_564_74#_c_1134_n 0.0346868f $X=2.405 $Y=0.515 $X2=0
+ $Y2=0
cc_587 N_VGND_c_1037_n N_A_564_74#_c_1135_n 0.0377951f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_1043_n N_A_564_74#_c_1135_n 0.0212998f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_1031_n N_A_564_74#_c_1136_n 0.0121616f $X=2.405 $Y=0.515 $X2=0
+ $Y2=0
cc_590 N_VGND_c_1037_n N_A_564_74#_c_1136_n 0.0235818f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_1043_n N_A_564_74#_c_1136_n 0.0127177f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_1032_n N_A_564_74#_c_1137_n 0.0100772f $X=5.395 $Y=0.525 $X2=0
+ $Y2=0
cc_593 N_VGND_c_1037_n N_A_564_74#_c_1137_n 0.065961f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_1043_n N_A_564_74#_c_1137_n 0.0367613f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_M1002_s N_A_564_74#_c_1172_n 0.00534428f $X=5.215 $Y=0.37 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1032_n N_A_564_74#_c_1172_n 0.0203382f $X=5.395 $Y=0.525 $X2=0
+ $Y2=0
cc_597 N_VGND_c_1043_n N_A_564_74#_c_1172_n 0.0112873f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_1032_n N_A_564_74#_c_1139_n 0.0109215f $X=5.395 $Y=0.525 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1033_n N_A_564_74#_c_1139_n 0.0105463f $X=6.395 $Y=0.52 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1039_n N_A_564_74#_c_1139_n 0.0144379f $X=6.23 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1043_n N_A_564_74#_c_1139_n 0.0119346f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_M1004_s N_A_564_74#_c_1182_n 0.0051536f $X=6.185 $Y=0.37 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1033_n N_A_564_74#_c_1182_n 0.0204467f $X=6.395 $Y=0.52 $X2=0
+ $Y2=0
cc_604 N_VGND_c_1043_n N_A_564_74#_c_1182_n 0.0120866f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_1033_n N_A_564_74#_c_1140_n 0.0100467f $X=6.395 $Y=0.52 $X2=0
+ $Y2=0
cc_606 N_VGND_c_1034_n N_A_564_74#_c_1140_n 0.009799f $X=7.35 $Y=0.515 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1041_n N_A_564_74#_c_1140_n 0.0108951f $X=7.16 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1043_n N_A_564_74#_c_1140_n 0.00900503f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_M1005_d N_A_564_74#_c_1141_n 0.00956917f $X=7.115 $Y=0.37 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1034_n N_A_564_74#_c_1141_n 0.027256f $X=7.35 $Y=0.515 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1043_n N_A_564_74#_c_1141_n 0.0119957f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_c_1034_n N_A_564_74#_c_1142_n 0.0101897f $X=7.35 $Y=0.515 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1042_n N_A_564_74#_c_1142_n 0.0145639f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_c_1043_n N_A_564_74#_c_1142_n 0.0119984f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_c_1037_n N_A_564_74#_c_1143_n 0.0230525f $X=5.23 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_1043_n N_A_564_74#_c_1143_n 0.0126179f $X=7.92 $Y=0 $X2=0 $Y2=0

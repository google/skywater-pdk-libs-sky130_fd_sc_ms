* File: sky130_fd_sc_ms__maj3_4.pex.spice
* Created: Fri Aug 28 17:39:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MAJ3_4%B 3 5 7 8 10 12 14 17 19 21 22 24 27 31 35 36
+ 37 50 53
c120 19 0 1.44963e-19 $X=2.935 $Y=1.375
r121 50 51 2.23839 $w=3.23e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.54
+ $X2=3.38 $Y2=1.54
r122 48 50 61.1827 $w=3.23e-07 $l=4.1e-07 $layer=POLY_cond $X=2.955 $Y=1.54
+ $X2=3.365 $Y2=1.54
r123 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.54 $X2=2.955 $Y2=1.54
r124 46 48 2.98452 $w=3.23e-07 $l=2e-08 $layer=POLY_cond $X=2.935 $Y=1.54
+ $X2=2.955 $Y2=1.54
r125 45 46 8.20743 $w=3.23e-07 $l=5.5e-08 $layer=POLY_cond $X=2.88 $Y=1.54
+ $X2=2.935 $Y2=1.54
r126 40 41 9.24189 $w=3.39e-07 $l=6.5e-08 $layer=POLY_cond $X=1.02 $Y=1.585
+ $X2=1.085 $Y2=1.585
r127 37 49 3.43222 $w=5.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.417
+ $X2=2.955 $Y2=1.417
r128 36 49 6.55243 $w=5.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=1.417
+ $X2=2.955 $Y2=1.417
r129 36 53 8.95336 $w=5.73e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.417
+ $X2=2.525 $Y2=1.417
r130 35 53 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.465 $Y=1.215
+ $X2=2.525 $Y2=1.215
r131 32 41 30.5693 $w=3.39e-07 $l=2.15e-07 $layer=POLY_cond $X=1.3 $Y=1.585
+ $X2=1.085 $Y2=1.585
r132 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.3
+ $Y=1.54 $X2=1.3 $Y2=1.54
r133 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.3 $Y=1.3
+ $X2=1.465 $Y2=1.215
r134 29 31 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.3 $Y=1.3 $X2=1.3
+ $Y2=1.54
r135 25 51 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.705
+ $X2=3.38 $Y2=1.54
r136 25 27 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=3.38 $Y=1.705
+ $X2=3.38 $Y2=2.46
r137 22 50 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.375
+ $X2=3.365 $Y2=1.54
r138 22 24 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.365 $Y=1.375
+ $X2=3.365 $Y2=0.945
r139 19 46 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.935 $Y=1.375
+ $X2=2.935 $Y2=1.54
r140 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.935 $Y=1.375
+ $X2=2.935 $Y2=0.945
r141 15 45 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.705
+ $X2=2.88 $Y2=1.54
r142 15 17 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=2.88 $Y=1.705
+ $X2=2.88 $Y2=2.46
r143 12 44 21.8644 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.515 $Y=1.375
+ $X2=1.515 $Y2=1.585
r144 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.515 $Y=1.375
+ $X2=1.515 $Y2=0.945
r145 8 44 6.39823 $w=3.39e-07 $l=4.5e-08 $layer=POLY_cond $X=1.47 $Y=1.585
+ $X2=1.515 $Y2=1.585
r146 8 32 24.1711 $w=3.39e-07 $l=1.7e-07 $layer=POLY_cond $X=1.47 $Y=1.585
+ $X2=1.3 $Y2=1.585
r147 8 10 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=1.47 $Y=1.705
+ $X2=1.47 $Y2=2.46
r148 5 41 21.8644 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.085 $Y=1.375
+ $X2=1.085 $Y2=1.585
r149 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.085 $Y=1.375
+ $X2=1.085 $Y2=0.945
r150 1 40 17.5597 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.02 $Y=1.795
+ $X2=1.02 $Y2=1.585
r151 1 3 258.492 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=1.02 $Y=1.795
+ $X2=1.02 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A 4 7 9 10 13 18 21 26 27 28 31 36 38 40 41
+ 45 46 48 51
c163 41 0 7.45928e-20 $X=4.24 $Y=1.96
c164 31 0 1.41402e-19 $X=5.8 $Y=2.46
c165 18 0 9.20449e-20 $X=2.015 $Y=0.945
c166 7 0 1.06155e-19 $X=0.52 $Y=2.46
r167 51 54 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.635
+ $X2=1.965 $Y2=1.8
r168 51 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.965 $Y=1.635
+ $X2=1.965 $Y2=1.47
r169 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.965
+ $Y=1.635 $X2=1.965 $Y2=1.635
r170 48 52 1.06087 $w=3.45e-07 $l=3e-08 $layer=LI1_cond $X=2.037 $Y=1.665
+ $X2=2.037 $Y2=1.635
r171 46 57 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.635
+ $X2=4.405 $Y2=1.8
r172 46 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.635
+ $X2=4.405 $Y2=1.47
r173 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.635 $X2=4.405 $Y2=1.635
r174 43 45 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.405 $Y=1.875
+ $X2=4.405 $Y2=1.635
r175 42 48 10.4319 $w=3.45e-07 $l=3.96529e-07 $layer=LI1_cond $X=2.275 $Y=1.96
+ $X2=2.037 $Y2=1.665
r176 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.24 $Y=1.96
+ $X2=4.405 $Y2=1.875
r177 41 42 128.198 $w=1.68e-07 $l=1.965e-06 $layer=LI1_cond $X=4.24 $Y=1.96
+ $X2=2.275 $Y2=1.96
r178 39 40 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.805 $Y=1.31
+ $X2=5.805 $Y2=1.46
r179 37 38 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.515 $Y=1.34
+ $X2=0.515 $Y2=1.49
r180 36 39 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.825 $Y=0.915
+ $X2=5.825 $Y2=1.31
r181 33 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.825 $Y=0.255
+ $X2=5.825 $Y2=0.915
r182 31 40 388.71 $w=1.8e-07 $l=1e-06 $layer=POLY_cond $X=5.8 $Y=2.46 $X2=5.8
+ $Y2=1.46
r183 27 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.75 $Y=0.18
+ $X2=5.825 $Y2=0.255
r184 27 28 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=5.75 $Y=0.18
+ $X2=4.53 $Y2=0.18
r185 26 56 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.455 $Y=0.71
+ $X2=4.455 $Y2=1.47
r186 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=0.255
+ $X2=4.53 $Y2=0.18
r187 23 26 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.455 $Y=0.255
+ $X2=4.455 $Y2=0.71
r188 21 57 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.45 $Y=2.46
+ $X2=4.45 $Y2=1.8
r189 18 53 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.015 $Y=0.945
+ $X2=2.015 $Y2=1.47
r190 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.015 $Y=0.255
+ $X2=2.015 $Y2=0.945
r191 13 54 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.92 $Y=2.46
+ $X2=1.92 $Y2=1.8
r192 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.94 $Y=0.18
+ $X2=2.015 $Y2=0.255
r193 9 10 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=1.94 $Y=0.18
+ $X2=0.57 $Y2=0.18
r194 7 38 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=0.52 $Y=2.46
+ $X2=0.52 $Y2=1.49
r195 4 37 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=0.945
+ $X2=0.495 $Y2=1.34
r196 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.57 $Y2=0.18
r197 1 4 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.495 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%C 1 3 8 9 10 13 18 21 25 29 33 36 39 43 46 49
+ 56 58
c142 43 0 1.41402e-19 $X=5.055 $Y=1.635
c143 18 0 1.46446e-19 $X=3.955 $Y=0.71
r144 56 57 6.75701 $w=3.21e-07 $l=4.5e-08 $layer=POLY_cond $X=5.35 $Y=1.635
+ $X2=5.395 $Y2=1.635
r145 53 54 9.76012 $w=3.21e-07 $l=6.5e-08 $layer=POLY_cond $X=4.9 $Y=1.635
+ $X2=4.965 $Y2=1.635
r146 49 52 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.54
+ $X2=3.855 $Y2=1.705
r147 49 51 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.54
+ $X2=3.855 $Y2=1.375
r148 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.54 $X2=3.845 $Y2=1.54
r149 46 50 5.5817 $w=5.23e-07 $l=2.45e-07 $layer=LI1_cond $X=3.747 $Y=1.295
+ $X2=3.747 $Y2=1.54
r150 46 58 1.8226 $w=5.23e-07 $l=8e-08 $layer=LI1_cond $X=3.747 $Y=1.295
+ $X2=3.747 $Y2=1.215
r151 44 56 44.296 $w=3.21e-07 $l=2.95e-07 $layer=POLY_cond $X=5.055 $Y=1.635
+ $X2=5.35 $Y2=1.635
r152 44 54 13.514 $w=3.21e-07 $l=9e-08 $layer=POLY_cond $X=5.055 $Y=1.635
+ $X2=4.965 $Y2=1.635
r153 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.635 $X2=5.055 $Y2=1.635
r154 40 43 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.84 $Y=1.635
+ $X2=5.055 $Y2=1.635
r155 39 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=1.47
+ $X2=4.84 $Y2=1.635
r156 38 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.84 $Y=1.3
+ $X2=4.84 $Y2=1.47
r157 37 58 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=4.01 $Y=1.215
+ $X2=3.747 $Y2=1.215
r158 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.755 $Y=1.215
+ $X2=4.84 $Y2=1.3
r159 36 37 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.755 $Y=1.215
+ $X2=4.01 $Y2=1.215
r160 31 57 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.47
+ $X2=5.395 $Y2=1.635
r161 31 33 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.395 $Y=1.47
+ $X2=5.395 $Y2=0.915
r162 27 56 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.35 $Y=1.8
+ $X2=5.35 $Y2=1.635
r163 27 29 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.35 $Y=1.8
+ $X2=5.35 $Y2=2.46
r164 23 54 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.47
+ $X2=4.965 $Y2=1.635
r165 23 25 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.965 $Y=1.47
+ $X2=4.965 $Y2=0.915
r166 19 53 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.8 $X2=4.9
+ $Y2=1.635
r167 19 21 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.9 $Y=1.8 $X2=4.9
+ $Y2=2.46
r168 18 51 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.955 $Y=0.71
+ $X2=3.955 $Y2=1.375
r169 15 18 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.955 $Y=0.255
+ $X2=3.955 $Y2=0.71
r170 13 52 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=3.88 $Y=2.46
+ $X2=3.88 $Y2=1.705
r171 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.88 $Y=0.18
+ $X2=3.955 $Y2=0.255
r172 9 10 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=3.88 $Y=0.18
+ $X2=2.52 $Y2=0.18
r173 8 35 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.445 $Y=0.945
+ $X2=2.445 $Y2=1.34
r174 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.52 $Y2=0.18
r175 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.445 $Y2=0.945
r176 1 35 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.43 $Y=1.43 $X2=2.43
+ $Y2=1.34
r177 1 3 400.371 $w=1.8e-07 $l=1.03e-06 $layer=POLY_cond $X=2.43 $Y=1.43
+ $X2=2.43 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_222_392# 1 2 3 4 5 6 21 23 25 28 30 32 35
+ 37 39 42 44 46 47 48 49 52 55 57 61 63 65 71 72 78 88 90 92 97 100 111
c224 92 0 1.44963e-19 $X=3.15 $Y=0.78
c225 72 0 1.04369e-19 $X=5.475 $Y=1.97
c226 55 0 1.06155e-19 $X=1.245 $Y=2.57
c227 47 0 9.20449e-20 $X=0.88 $Y=0.96
c228 30 0 1.55372e-19 $X=6.805 $Y=1.345
c229 23 0 1.82103e-19 $X=6.335 $Y=1.345
r230 111 112 1.46505 $w=3.29e-07 $l=1e-08 $layer=POLY_cond $X=7.655 $Y=1.51
+ $X2=7.665 $Y2=1.51
r231 110 111 61.5319 $w=3.29e-07 $l=4.2e-07 $layer=POLY_cond $X=7.235 $Y=1.51
+ $X2=7.655 $Y2=1.51
r232 109 110 4.39514 $w=3.29e-07 $l=3e-08 $layer=POLY_cond $X=7.205 $Y=1.51
+ $X2=7.235 $Y2=1.51
r233 106 107 7.32523 $w=3.29e-07 $l=5e-08 $layer=POLY_cond $X=6.755 $Y=1.51
+ $X2=6.805 $Y2=1.51
r234 105 106 61.5319 $w=3.29e-07 $l=4.2e-07 $layer=POLY_cond $X=6.335 $Y=1.51
+ $X2=6.755 $Y2=1.51
r235 100 102 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.18 $Y=0.76
+ $X2=5.18 $Y2=0.875
r236 92 94 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=3.19 $Y=0.78
+ $X2=3.19 $Y2=0.875
r237 79 109 32.231 $w=3.29e-07 $l=2.2e-07 $layer=POLY_cond $X=6.985 $Y=1.51
+ $X2=7.205 $Y2=1.51
r238 79 107 26.3708 $w=3.29e-07 $l=1.8e-07 $layer=POLY_cond $X=6.985 $Y=1.51
+ $X2=6.805 $Y2=1.51
r239 78 79 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.985
+ $Y=1.51 $X2=6.985 $Y2=1.51
r240 76 105 4.39514 $w=3.29e-07 $l=3e-08 $layer=POLY_cond $X=6.305 $Y=1.51
+ $X2=6.335 $Y2=1.51
r241 75 78 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.305 $Y=1.51
+ $X2=6.985 $Y2=1.51
r242 75 76 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.305
+ $Y=1.51 $X2=6.305 $Y2=1.51
r243 73 75 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=5.56 $Y=1.51
+ $X2=6.305 $Y2=1.51
r244 72 97 14.0461 $w=3.04e-07 $l=4.41531e-07 $layer=LI1_cond $X=5.475 $Y=1.97
+ $X2=5.125 $Y2=2.177
r245 71 73 9.18505 $w=2.62e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.475 $Y=1.675
+ $X2=5.39 $Y2=1.51
r246 71 72 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.475 $Y=1.675
+ $X2=5.475 $Y2=1.97
r247 68 73 19.1965 $w=2.62e-07 $l=4.73498e-07 $layer=LI1_cond $X=5.18 $Y=1.13
+ $X2=5.39 $Y2=1.51
r248 68 70 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.18 $Y=1.13 $X2=5.18
+ $Y2=1.1
r249 67 102 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=0.96
+ $X2=5.18 $Y2=0.875
r250 67 70 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=0.96
+ $X2=5.18 $Y2=1.1
r251 66 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=2.3
+ $X2=3.155 $Y2=2.3
r252 65 97 8.97325 $w=3.04e-07 $l=2.17991e-07 $layer=LI1_cond $X=4.96 $Y=2.3
+ $X2=5.125 $Y2=2.177
r253 65 66 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=4.96 $Y=2.3
+ $X2=3.32 $Y2=2.3
r254 64 94 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.315 $Y=0.875
+ $X2=3.19 $Y2=0.875
r255 63 102 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.875
+ $X2=5.18 $Y2=0.875
r256 63 64 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=5.095 $Y=0.875
+ $X2=3.315 $Y2=0.875
r257 59 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.385
+ $X2=3.155 $Y2=2.3
r258 59 61 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.155 $Y=2.385
+ $X2=3.155 $Y2=2.65
r259 58 88 3.25423 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.41 $Y=2.3
+ $X2=1.252 $Y2=2.3
r260 57 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=2.3
+ $X2=3.155 $Y2=2.3
r261 57 58 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=2.99 $Y=2.3
+ $X2=1.41 $Y2=2.3
r262 53 88 3.29812 $w=2.85e-07 $l=9.88686e-08 $layer=LI1_cond $X=1.222 $Y=2.385
+ $X2=1.252 $Y2=2.3
r263 53 55 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=1.222 $Y=2.385
+ $X2=1.222 $Y2=2.57
r264 50 88 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.252 $Y=2.215
+ $X2=1.252 $Y2=2.3
r265 50 52 2.0122 $w=3.13e-07 $l=5.5e-08 $layer=LI1_cond $X=1.252 $Y=2.215
+ $X2=1.252 $Y2=2.16
r266 49 84 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=1.252 $Y=1.96
+ $X2=0.88 $Y2=1.96
r267 49 52 4.20733 $w=3.13e-07 $l=1.15e-07 $layer=LI1_cond $X=1.252 $Y=2.045
+ $X2=1.252 $Y2=2.16
r268 48 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.875
+ $X2=0.88 $Y2=1.96
r269 47 83 19.6322 $w=2.61e-07 $l=5.35593e-07 $layer=LI1_cond $X=0.88 $Y=0.96
+ $X2=1.3 $Y2=0.697
r270 47 48 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.88 $Y=0.96
+ $X2=0.88 $Y2=1.875
r271 44 112 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.345
+ $X2=7.665 $Y2=1.51
r272 44 46 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.665 $Y=1.345
+ $X2=7.665 $Y2=0.865
r273 40 111 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.675
+ $X2=7.655 $Y2=1.51
r274 40 42 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=7.655 $Y=1.675
+ $X2=7.655 $Y2=2.4
r275 37 110 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.235 $Y=1.345
+ $X2=7.235 $Y2=1.51
r276 37 39 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.235 $Y=1.345
+ $X2=7.235 $Y2=0.865
r277 33 109 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=1.675
+ $X2=7.205 $Y2=1.51
r278 33 35 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=7.205 $Y=1.675
+ $X2=7.205 $Y2=2.4
r279 30 107 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.805 $Y=1.345
+ $X2=6.805 $Y2=1.51
r280 30 32 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.805 $Y=1.345
+ $X2=6.805 $Y2=0.865
r281 26 106 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.755 $Y=1.675
+ $X2=6.755 $Y2=1.51
r282 26 28 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=6.755 $Y=1.675
+ $X2=6.755 $Y2=2.4
r283 23 105 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=1.51
r284 23 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=0.865
r285 19 76 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.675
+ $X2=6.305 $Y2=1.51
r286 19 21 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=6.305 $Y=1.675
+ $X2=6.305 $Y2=2.4
r287 6 97 600 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_PDIFF $count=1 $X=4.99
+ $Y=1.96 $X2=5.125 $Y2=2.215
r288 5 90 600 $w=1.7e-07 $l=4.22493e-07 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.96 $X2=3.155 $Y2=2.3
r289 5 61 600 $w=1.7e-07 $l=7.77013e-07 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.96 $X2=3.155 $Y2=2.65
r290 4 55 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.96 $X2=1.245 $Y2=2.57
r291 4 52 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.96 $X2=1.245 $Y2=2.16
r292 3 100 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.595 $X2=5.18 $Y2=0.76
r293 3 70 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.595 $X2=5.18 $Y2=1.1
r294 2 92 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.625 $X2=3.15 $Y2=0.78
r295 1 83 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.625 $X2=1.3 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 43 45 47
+ 51 53 61 69 74 83 86 89 92 96
c106 2 0 7.45928e-20 $X=2.01 $Y=1.96
r107 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r110 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r111 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 78 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 75 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.145 $Y=3.33
+ $X2=7.02 $Y2=3.33
r117 75 77 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.145 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 74 95 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.937 $Y2=3.33
r119 74 77 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 73 90 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r121 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r122 70 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.155 $Y2=3.33
r123 70 72 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 69 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=6.065 $Y2=3.33
r125 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r127 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r130 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r131 62 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.19 $Y2=3.33
r132 62 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 61 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.155 $Y2=3.33
r134 61 67 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.6 $Y2=3.33
r135 60 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r137 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r138 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 54 80 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.19 $Y2=3.33
r142 54 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 53 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=2.19 $Y2=3.33
r144 53 59 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=1.68 $Y2=3.33
r145 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 51 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r148 47 50 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.88 $Y=1.985
+ $X2=7.88 $Y2=2.815
r149 45 95 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.937 $Y2=3.33
r150 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.815
r151 41 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.02 $Y=3.245
+ $X2=7.02 $Y2=3.33
r152 41 43 41.2575 $w=2.48e-07 $l=8.95e-07 $layer=LI1_cond $X=7.02 $Y=3.245
+ $X2=7.02 $Y2=2.35
r153 40 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.065 $Y2=3.33
r154 39 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.895 $Y=3.33
+ $X2=7.02 $Y2=3.33
r155 39 40 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.895 $Y=3.33
+ $X2=6.19 $Y2=3.33
r156 35 38 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.065 $Y=2.105
+ $X2=6.065 $Y2=2.815
r157 33 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.065 $Y=3.245
+ $X2=6.065 $Y2=3.33
r158 33 38 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.065 $Y=3.245
+ $X2=6.065 $Y2=2.815
r159 29 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=3.33
r160 29 31 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=2.72
r161 25 83 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r162 25 27 23.2705 $w=2.58e-07 $l=5.25e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.72
r163 21 24 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.255 $Y=2.105
+ $X2=0.255 $Y2=2.815
r164 19 80 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.19 $Y2=3.33
r165 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r166 6 50 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=2.815
r167 6 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=1.985
r168 5 43 300 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=2 $X=6.845
+ $Y=1.84 $X2=6.98 $Y2=2.35
r169 4 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.96 $X2=6.025 $Y2=2.815
r170 4 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.96 $X2=6.025 $Y2=2.105
r171 3 31 600 $w=1.7e-07 $l=8.47467e-07 $layer=licon1_PDIFF $count=1 $X=3.97
+ $Y=1.96 $X2=4.155 $Y2=2.72
r172 2 27 600 $w=1.7e-07 $l=8.27043e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.96 $X2=2.15 $Y2=2.72
r173 1 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.96 $X2=0.295 $Y2=2.815
r174 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.96 $X2=0.295 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_122_392# 1 2 9 11 12 15
r24 13 15 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.695 $Y=2.905
+ $X2=1.695 $Y2=2.765
r25 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.53 $Y=2.99
+ $X2=1.695 $Y2=2.905
r26 11 12 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.53 $Y=2.99
+ $X2=0.91 $Y2=2.99
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.745 $Y=2.905
+ $X2=0.91 $Y2=2.99
r28 7 9 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.745 $Y=2.905
+ $X2=0.745 $Y2=2.38
r29 2 15 600 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.96 $X2=1.695 $Y2=2.765
r30 1 9 300 $w=1.7e-07 $l=4.82804e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.96 $X2=0.745 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_504_392# 1 2 9 11 12 15
r27 13 15 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.655 $Y=2.905
+ $X2=3.655 $Y2=2.72
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.49 $Y=2.99
+ $X2=3.655 $Y2=2.905
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.49 $Y=2.99
+ $X2=2.82 $Y2=2.99
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.655 $Y=2.905
+ $X2=2.82 $Y2=2.99
r31 7 9 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.655 $Y=2.905
+ $X2=2.655 $Y2=2.72
r32 2 15 600 $w=1.7e-07 $l=8.47467e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.96 $X2=3.655 $Y2=2.72
r33 1 9 600 $w=1.7e-07 $l=8.24742e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.96 $X2=2.655 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_908_392# 1 2 7 9 14
c25 2 0 1.04369e-19 $X=5.44 $Y=1.96
r26 14 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.575 $Y=2.64 $X2=5.575
+ $Y2=2.72
r27 9 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.675 $Y=2.64 $X2=4.675
+ $Y2=2.72
r28 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=2.64 $X2=4.675
+ $Y2=2.64
r29 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=2.64
+ $X2=5.575 $Y2=2.64
r30 7 8 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.41 $Y=2.64 $X2=4.84
+ $Y2=2.64
r31 2 17 600 $w=1.7e-07 $l=8.24742e-07 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=1.96 $X2=5.575 $Y2=2.72
r32 1 12 600 $w=1.7e-07 $l=8.24742e-07 $layer=licon1_PDIFF $count=1 $X=4.54
+ $Y=1.96 $X2=4.675 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%X 1 2 3 4 13 15 19 21 22 25 28 31 33 34 41
c58 19 0 3.37475e-19 $X=6.59 $Y=0.64
r59 40 41 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.92 $Y=1.48
+ $X2=7.92 $Y2=1.295
r60 39 41 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.92 $Y=1.175
+ $X2=7.92 $Y2=1.295
r61 33 40 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.565
+ $X2=7.92 $Y2=1.48
r62 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.805 $Y=1.565
+ $X2=7.515 $Y2=1.565
r63 29 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=2.015
+ $X2=7.43 $Y2=1.93
r64 29 31 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.43 $Y=2.015 $X2=7.43
+ $Y2=2.815
r65 28 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=1.845
+ $X2=7.43 $Y2=1.93
r66 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.43 $Y=1.65
+ $X2=7.515 $Y2=1.565
r67 27 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.43 $Y=1.65
+ $X2=7.43 $Y2=1.845
r68 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=1.93
+ $X2=6.53 $Y2=1.93
r69 25 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=1.93
+ $X2=7.43 $Y2=1.93
r70 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.345 $Y=1.93
+ $X2=6.695 $Y2=1.93
r71 22 24 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.675 $Y=1.09
+ $X2=7.45 $Y2=1.09
r72 21 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.09
+ $X2=7.92 $Y2=1.175
r73 21 24 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.805 $Y=1.09
+ $X2=7.45 $Y2=1.09
r74 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.55 $Y=1.005
+ $X2=6.675 $Y2=1.09
r75 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=6.55 $Y=1.005
+ $X2=6.55 $Y2=0.64
r76 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=2.015 $X2=6.53
+ $Y2=1.93
r77 13 15 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=6.53 $Y=2.015 $X2=6.53
+ $Y2=2.815
r78 4 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.43 $Y2=1.985
r79 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.43 $Y2=2.815
r80 3 36 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=6.395
+ $Y=1.84 $X2=6.53 $Y2=2.01
r81 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.395
+ $Y=1.84 $X2=6.53 $Y2=2.815
r82 2 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.31
+ $Y=0.495 $X2=7.45 $Y2=1.09
r83 1 19 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=6.41
+ $Y=0.495 $X2=6.59 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 39 41 43
+ 45 50 55 60 65 74 77 80 83 87
r94 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r95 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r96 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r97 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r98 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r99 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r100 69 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r101 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r102 66 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.185 $Y=0 $X2=7.02
+ $Y2=0
r103 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.185 $Y=0
+ $X2=7.44 $Y2=0
r104 65 86 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.937 $Y2=0
r105 65 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.44 $Y2=0
r106 64 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r107 64 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r108 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r109 61 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.08
+ $Y2=0
r110 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=6.48 $Y2=0
r111 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=0 $X2=7.02
+ $Y2=0
r112 60 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.855 $Y=0
+ $X2=6.48 $Y2=0
r113 59 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r114 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r115 56 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.17
+ $Y2=0
r116 56 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.56 $Y2=0
r117 55 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.955 $Y=0 $X2=6.08
+ $Y2=0
r118 55 58 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.955 $Y=0
+ $X2=4.56 $Y2=0
r119 54 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r120 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r121 51 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.23
+ $Y2=0
r122 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.64 $Y2=0
r123 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.17
+ $Y2=0
r124 50 53 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.005 $Y=0
+ $X2=2.64 $Y2=0
r125 49 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r126 49 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r127 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 46 71 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r129 46 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r130 45 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.23
+ $Y2=0
r131 45 48 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.145 $Y=0
+ $X2=0.72 $Y2=0
r132 43 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r133 43 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r134 43 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r135 39 86 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.937 $Y2=0
r136 39 41 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.67
r137 35 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.02 $Y=0.085
+ $X2=7.02 $Y2=0
r138 35 37 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=7.02 $Y=0.085
+ $X2=7.02 $Y2=0.67
r139 31 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.08 $Y=0.085
+ $X2=6.08 $Y2=0
r140 31 33 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=6.08 $Y=0.085
+ $X2=6.08 $Y2=0.64
r141 27 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0
r142 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0.535
r143 23 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=0.085
+ $X2=2.23 $Y2=0
r144 23 25 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.23 $Y=0.085
+ $X2=2.23 $Y2=0.78
r145 19 71 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r146 19 21 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.77
r147 6 41 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=7.74
+ $Y=0.495 $X2=7.88 $Y2=0.67
r148 5 37 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=6.88
+ $Y=0.495 $X2=7.02 $Y2=0.67
r149 4 33 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=5.9
+ $Y=0.595 $X2=6.12 $Y2=0.64
r150 3 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.39 $X2=4.17 $Y2=0.535
r151 2 25 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.625 $X2=2.23 $Y2=0.78
r152 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_114_125# 1 2 7 11 13
r26 13 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.79 $Y=0.35
+ $X2=0.79 $Y2=0.535
r27 9 11 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.8 $Y=0.435 $X2=1.8
+ $Y2=0.78
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0.35
+ $X2=0.79 $Y2=0.35
r29 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.635 $Y=0.35
+ $X2=1.8 $Y2=0.435
r30 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.635 $Y=0.35
+ $X2=0.955 $Y2=0.35
r31 2 11 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.625 $X2=1.8 $Y2=0.78
r32 1 16 182 $w=1.7e-07 $l=2.61151e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.625 $X2=0.79 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_504_125# 1 2 9 11 12 13
r34 13 16 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.66 $Y=0.35
+ $X2=3.66 $Y2=0.53
r35 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=3.66 $Y2=0.35
r36 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=2.885 $Y2=0.35
r37 7 12 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=2.69 $Y=0.435
+ $X2=2.885 $Y2=0.35
r38 7 9 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.69 $Y=0.435
+ $X2=2.69 $Y2=0.77
r39 2 16 182 $w=1.7e-07 $l=2.63249e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.625 $X2=3.66 $Y2=0.53
r40 1 9 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=2.52
+ $Y=0.625 $X2=2.69 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_4%A_906_78# 1 2 7 11 13
c30 13 0 1.46446e-19 $X=4.67 $Y=0.34
r31 13 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.67 $Y=0.34
+ $X2=4.67 $Y2=0.535
r32 9 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.61 $Y2=0.795
r33 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.34
+ $X2=4.67 $Y2=0.34
r34 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=5.61 $Y2=0.425
r35 7 8 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=4.835 $Y2=0.34
r36 2 11 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.595 $X2=5.61 $Y2=0.795
r37 1 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.39 $X2=4.67 $Y2=0.535
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dfbbn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 1.180000 2.755000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.502200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.005000 0.350000 13.340000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.496600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.555000 0.405000 11.925000 1.150000 ;
        RECT 11.575000 1.820000 11.925000 2.980000 ;
        RECT 11.755000 1.150000 11.925000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.350000 11.015000 1.780000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.524700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.675000 5.850000 1.960000 ;
        RECT 5.435000 1.960000 5.635000 2.150000 ;
        RECT 8.730000 1.275000 9.060000 2.120000 ;
      LAYER mcon ;
        RECT 5.435000 1.950000 5.605000 2.120000 ;
        RECT 8.795000 1.950000 8.965000 2.120000 ;
      LAYER met1 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 1.965000 9.025000 2.105000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.495000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.440000 0.085000 ;
        RECT  0.545000  0.085000  0.875000 0.790000 ;
        RECT  2.045000  0.085000  2.410000 0.670000 ;
        RECT  5.815000  0.085000  6.145000 1.035000 ;
        RECT  8.715000  0.085000  8.885000 0.765000 ;
        RECT 11.055000  0.085000 11.385000 0.425000 ;
        RECT 12.580000  0.085000 12.830000 0.810000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.440000 3.415000 ;
        RECT  0.635000 2.290000  0.805000 3.245000 ;
        RECT  2.295000 2.525000  2.465000 3.245000 ;
        RECT  5.040000 2.660000  5.370000 3.245000 ;
        RECT  6.020000 2.660000  6.350000 3.245000 ;
        RECT  7.905000 2.970000  8.270000 3.245000 ;
        RECT  9.035000 2.970000  9.365000 3.245000 ;
        RECT 11.045000 2.630000 11.375000 3.245000 ;
        RECT 12.555000 1.820000 12.805000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.105000 1.950000  0.835000 2.120000 ;
      RECT  0.105000 2.120000  0.435000 2.980000 ;
      RECT  0.115000 0.350000  0.365000 0.960000 ;
      RECT  0.115000 0.960000  0.835000 1.130000 ;
      RECT  0.665000 1.130000  0.835000 1.300000 ;
      RECT  0.665000 1.300000  1.075000 1.630000 ;
      RECT  0.665000 1.630000  0.835000 1.950000 ;
      RECT  1.005000 1.820000  1.415000 2.905000 ;
      RECT  1.005000 2.905000  2.125000 3.075000 ;
      RECT  1.055000 0.350000  1.415000 1.130000 ;
      RECT  1.245000 1.130000  1.415000 1.820000 ;
      RECT  1.585000 0.575000  1.865000 0.840000 ;
      RECT  1.585000 0.840000  2.750000 1.010000 ;
      RECT  1.585000 1.010000  1.755000 2.405000 ;
      RECT  1.585000 2.405000  1.785000 2.735000 ;
      RECT  1.955000 1.685000  3.240000 1.855000 ;
      RECT  1.955000 1.855000  2.125000 2.905000 ;
      RECT  2.370000 2.025000  2.805000 2.355000 ;
      RECT  2.580000 0.255000  4.145000 0.425000 ;
      RECT  2.580000 0.425000  2.750000 0.840000 ;
      RECT  2.635000 2.355000  2.805000 2.905000 ;
      RECT  2.635000 2.905000  4.530000 3.075000 ;
      RECT  2.950000 0.595000  3.280000 0.785000 ;
      RECT  2.950000 0.785000  3.805000 0.955000 ;
      RECT  2.975000 1.125000  3.465000 1.455000 ;
      RECT  2.975000 1.455000  3.240000 1.685000 ;
      RECT  2.975000 1.855000  3.240000 2.355000 ;
      RECT  3.090000 2.565000  3.580000 2.735000 ;
      RECT  3.410000 1.625000  4.135000 1.795000 ;
      RECT  3.410000 1.795000  3.580000 2.565000 ;
      RECT  3.460000 0.425000  4.145000 0.615000 ;
      RECT  3.635000 0.955000  3.805000 1.395000 ;
      RECT  3.635000 1.395000  4.135000 1.625000 ;
      RECT  3.750000 1.965000  4.475000 2.135000 ;
      RECT  3.750000 2.135000  4.000000 2.735000 ;
      RECT  3.975000 0.615000  4.145000 0.995000 ;
      RECT  3.975000 0.995000  4.475000 1.165000 ;
      RECT  4.200000 2.305000  4.815000 2.320000 ;
      RECT  4.200000 2.320000  6.450000 2.490000 ;
      RECT  4.200000 2.490000  4.530000 2.905000 ;
      RECT  4.305000 1.165000  4.475000 1.965000 ;
      RECT  4.315000 0.255000  5.645000 0.425000 ;
      RECT  4.315000 0.425000  4.645000 0.825000 ;
      RECT  4.645000 0.995000  5.145000 1.165000 ;
      RECT  4.645000 1.165000  4.815000 2.305000 ;
      RECT  4.815000 0.715000  5.145000 0.995000 ;
      RECT  4.985000 1.335000  6.485000 1.505000 ;
      RECT  4.985000 1.505000  5.265000 1.665000 ;
      RECT  5.315000 0.425000  5.645000 1.035000 ;
      RECT  5.570000 2.490000  5.820000 2.980000 ;
      RECT  6.120000 1.675000  6.450000 2.320000 ;
      RECT  6.315000 0.340000  8.545000 0.510000 ;
      RECT  6.315000 0.510000  6.485000 1.335000 ;
      RECT  6.710000 1.180000  7.865000 1.560000 ;
      RECT  6.710000 1.560000  7.075000 1.930000 ;
      RECT  6.720000 0.680000  8.205000 1.010000 ;
      RECT  6.860000 2.100000  7.415000 2.980000 ;
      RECT  7.245000 1.730000  8.560000 1.900000 ;
      RECT  7.245000 1.900000  7.415000 2.100000 ;
      RECT  7.890000 2.070000  8.220000 2.630000 ;
      RECT  7.890000 2.630000 10.320000 2.800000 ;
      RECT  8.035000 1.010000  8.205000 1.730000 ;
      RECT  8.375000 0.510000  8.545000 0.935000 ;
      RECT  8.375000 0.935000 10.890000 1.105000 ;
      RECT  8.390000 1.900000  8.560000 2.290000 ;
      RECT  8.390000 2.290000  9.400000 2.460000 ;
      RECT  8.500000 2.800000  8.830000 2.980000 ;
      RECT  9.065000 0.255000 10.360000 0.425000 ;
      RECT  9.065000 0.425000  9.315000 0.765000 ;
      RECT  9.230000 1.950000 10.170000 2.120000 ;
      RECT  9.230000 2.120000  9.400000 2.290000 ;
      RECT  9.300000 1.105000  9.630000 1.560000 ;
      RECT  9.495000 0.595000 11.385000 0.765000 ;
      RECT  9.840000 1.420000 10.170000 1.950000 ;
      RECT  9.990000 2.290000 11.385000 2.460000 ;
      RECT  9.990000 2.460000 10.320000 2.630000 ;
      RECT  9.990000 2.800000 10.320000 2.980000 ;
      RECT 10.345000 1.105000 10.515000 1.950000 ;
      RECT 10.345000 1.950000 10.850000 2.120000 ;
      RECT 11.215000 0.765000 11.385000 1.320000 ;
      RECT 11.215000 1.320000 11.585000 1.650000 ;
      RECT 11.215000 1.650000 11.385000 2.290000 ;
      RECT 12.110000 0.350000 12.360000 1.255000 ;
      RECT 12.110000 1.255000 12.835000 1.585000 ;
      RECT 12.110000 1.585000 12.360000 2.910000 ;
    LAYER mcon ;
      RECT 3.035000 1.210000 3.205000 1.380000 ;
      RECT 6.875000 1.210000 7.045000 1.380000 ;
    LAYER met1 ;
      RECT 2.975000 1.180000 3.265000 1.225000 ;
      RECT 2.975000 1.225000 7.105000 1.365000 ;
      RECT 2.975000 1.365000 3.265000 1.410000 ;
      RECT 6.815000 1.180000 7.105000 1.225000 ;
      RECT 6.815000 1.365000 7.105000 1.410000 ;
  END
END sky130_fd_sc_ms__dfbbn_1

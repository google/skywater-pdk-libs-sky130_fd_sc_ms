* File: sky130_fd_sc_ms__o211a_2.spice
* Created: Wed Sep  2 12:20:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o211a_2.pex.spice"
.subckt sky130_fd_sc_ms__o211a_2  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1011 A_117_74# N_C1_M1011_g N_A_27_368#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1004 N_A_195_74#_M1004_d N_B1_M1004_g A_117_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.0888 PD=1.1 PS=0.98 NRD=12.156 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_195_74#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1751 AS=0.1332 PD=1.33 PS=1.1 NRD=29.448 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_A_195_74#_M1000_d N_A1_M1000_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.1751 PD=2.02 PS=1.33 NRD=0 NRS=29.448 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_X_M1003_d N_A_27_368#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1003_d N_A_27_368#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_C1_M1007_g N_A_27_368#_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1006 N_A_27_368#_M1006_d N_B1_M1006_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1
+ AD=0.14 AS=0.18 PD=1.28 PS=1.36 NRD=0.9653 NRS=6.8753 M=1 R=5.55556 SA=90000.7
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1005 A_317_368# N_A2_M1005_g N_A_27_368#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.145 AS=0.14 PD=1.29 PS=1.28 NRD=17.7103 NRS=0 M=1 R=5.55556 SA=90001.2
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_317_368# VPB PSHORT L=0.18 W=1 AD=0.339623
+ AS=0.145 PD=1.70755 PS=1.29 NRD=0 NRS=17.7103 M=1 R=5.55556 SA=90001.6
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1001 N_X_M1001_d N_A_27_368#_M1001_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.380377 PD=1.39 PS=1.91245 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.3 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1002 N_X_M1001_d N_A_27_368#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
c_37 VNB 0 1.11614e-19 $X=0 $Y=0
c_407 A_117_74# 0 7.65495e-20 $X=0.585 $Y=0.37
*
.include "sky130_fd_sc_ms__o211a_2.pxi.spice"
*
.ends
*
*

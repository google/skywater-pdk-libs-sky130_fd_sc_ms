* File: sky130_fd_sc_ms__clkinv_8.pxi.spice
* Created: Fri Aug 28 17:20:34 2020
* 
x_PM_SKY130_FD_SC_MS__CLKINV_8%A N_A_M1000_g N_A_M1002_g N_A_M1003_g N_A_M1004_g
+ N_A_M1005_g N_A_M1006_g N_A_M1001_g N_A_M1007_g N_A_M1012_g N_A_M1008_g
+ N_A_M1015_g N_A_M1009_g N_A_M1016_g N_A_M1010_g N_A_M1017_g N_A_M1011_g
+ N_A_M1018_g N_A_M1013_g N_A_M1014_g N_A_M1019_g A A A A A A A N_A_c_104_n
+ N_A_c_91_n PM_SKY130_FD_SC_MS__CLKINV_8%A
x_PM_SKY130_FD_SC_MS__CLKINV_8%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1005_s
+ N_VPWR_M1007_s N_VPWR_M1009_s N_VPWR_M1011_s N_VPWR_M1014_s N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n VPWR
+ N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n
+ N_VPWR_c_283_n PM_SKY130_FD_SC_MS__CLKINV_8%VPWR
x_PM_SKY130_FD_SC_MS__CLKINV_8%Y N_Y_M1000_d N_Y_M1012_d N_Y_M1016_d N_Y_M1018_d
+ N_Y_M1002_d N_Y_M1004_d N_Y_M1006_d N_Y_M1008_d N_Y_M1010_d N_Y_M1013_d
+ N_Y_c_381_n N_Y_c_395_n N_Y_c_411_n N_Y_c_414_n N_Y_c_382_n N_Y_c_383_n
+ N_Y_c_396_n N_Y_c_427_n N_Y_c_397_n N_Y_c_384_n N_Y_c_438_n N_Y_c_442_n
+ N_Y_c_398_n N_Y_c_385_n N_Y_c_454_n N_Y_c_458_n N_Y_c_399_n N_Y_c_386_n
+ N_Y_c_470_n N_Y_c_387_n N_Y_c_400_n N_Y_c_388_n N_Y_c_401_n N_Y_c_484_n
+ N_Y_c_389_n N_Y_c_490_n N_Y_c_390_n N_Y_c_498_n N_Y_c_391_n N_Y_c_506_n
+ N_Y_c_392_n N_Y_c_513_n Y PM_SKY130_FD_SC_MS__CLKINV_8%Y
x_PM_SKY130_FD_SC_MS__CLKINV_8%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1015_s
+ N_VGND_M1017_s N_VGND_M1019_s N_VGND_c_574_n N_VGND_c_575_n N_VGND_c_576_n
+ N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n
+ N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n VGND N_VGND_c_585_n
+ N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n PM_SKY130_FD_SC_MS__CLKINV_8%VGND
cc_1 VNB N_A_M1000_g 0.0596095f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.61
cc_2 VNB N_A_M1001_g 0.0529153f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.61
cc_3 VNB N_A_M1012_g 0.0385104f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.61
cc_4 VNB N_A_M1015_g 0.0385105f $X=-0.19 $Y=-0.245 $X2=3.675 $Y2=0.61
cc_5 VNB N_A_M1016_g 0.0385105f $X=-0.19 $Y=-0.245 $X2=4.245 $Y2=0.61
cc_6 VNB N_A_M1017_g 0.0385105f $X=-0.19 $Y=-0.245 $X2=4.675 $Y2=0.61
cc_7 VNB N_A_M1018_g 0.0402814f $X=-0.19 $Y=-0.245 $X2=5.245 $Y2=0.61
cc_8 VNB N_A_M1019_g 0.0480697f $X=-0.19 $Y=-0.245 $X2=5.745 $Y2=0.61
cc_9 VNB N_A_c_91_n 0.268498f $X=-0.19 $Y=-0.245 $X2=5.745 $Y2=1.515
cc_10 VNB N_VPWR_c_283_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.515
cc_11 VNB N_Y_c_381_n 0.0164554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_Y_c_382_n 0.0246541f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=2.4
cc_13 VNB N_Y_c_383_n 0.0177577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_384_n 0.00999295f $X=-0.19 $Y=-0.245 $X2=4.245 $Y2=0.61
cc_15 VNB N_Y_c_385_n 0.00999295f $X=-0.19 $Y=-0.245 $X2=4.78 $Y2=2.4
cc_16 VNB N_Y_c_386_n 0.00999295f $X=-0.19 $Y=-0.245 $X2=5.73 $Y2=2.4
cc_17 VNB N_Y_c_387_n 0.00189504f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_18 VNB N_Y_c_388_n 0.0148487f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=1.58
cc_19 VNB N_Y_c_389_n 0.00436883f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.515
cc_20 VNB N_Y_c_390_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.515
cc_21 VNB N_Y_c_391_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=1.515
cc_22 VNB N_Y_c_392_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=4.245 $Y2=1.515
cc_23 VNB Y 0.0236628f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=1.515
cc_24 VNB N_VGND_c_574_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_575_n 0.0275144f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=2.4
cc_26 VNB N_VGND_c_576_n 0.0109417f $X=-0.19 $Y=-0.245 $X2=2.43 $Y2=2.4
cc_27 VNB N_VGND_c_577_n 0.00966068f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.61
cc_28 VNB N_VGND_c_578_n 0.00966068f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=2.4
cc_29 VNB N_VGND_c_579_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_580_n 0.025863f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=0.61
cc_31 VNB N_VGND_c_581_n 0.0620883f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=1.68
cc_32 VNB N_VGND_c_582_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.38 $Y2=2.4
cc_33 VNB N_VGND_c_583_n 0.0191309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_584_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.675 $Y2=1.35
cc_35 VNB N_VGND_c_585_n 0.0191309f $X=-0.19 $Y=-0.245 $X2=4.33 $Y2=2.4
cc_36 VNB N_VGND_c_586_n 0.0191309f $X=-0.19 $Y=-0.245 $X2=4.675 $Y2=0.61
cc_37 VNB N_VGND_c_587_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=5.245 $Y2=0.61
cc_38 VNB N_VGND_c_588_n 0.368436f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=2.4
cc_39 VPB N_A_M1002_g 0.0238156f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=2.4
cc_40 VPB N_A_M1003_g 0.0210642f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=2.4
cc_41 VPB N_A_M1004_g 0.0210664f $X=-0.19 $Y=1.66 $X2=1.48 $Y2=2.4
cc_42 VPB N_A_M1005_g 0.0210667f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=2.4
cc_43 VPB N_A_M1006_g 0.0210664f $X=-0.19 $Y=1.66 $X2=2.43 $Y2=2.4
cc_44 VPB N_A_M1007_g 0.0210667f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=2.4
cc_45 VPB N_A_M1008_g 0.0210664f $X=-0.19 $Y=1.66 $X2=3.38 $Y2=2.4
cc_46 VPB N_A_M1009_g 0.0210667f $X=-0.19 $Y=1.66 $X2=3.83 $Y2=2.4
cc_47 VPB N_A_M1010_g 0.0210664f $X=-0.19 $Y=1.66 $X2=4.33 $Y2=2.4
cc_48 VPB N_A_M1011_g 0.0210667f $X=-0.19 $Y=1.66 $X2=4.78 $Y2=2.4
cc_49 VPB N_A_M1013_g 0.0210645f $X=-0.19 $Y=1.66 $X2=5.28 $Y2=2.4
cc_50 VPB N_A_M1014_g 0.0223668f $X=-0.19 $Y=1.66 $X2=5.73 $Y2=2.4
cc_51 VPB N_A_c_104_n 0.0305696f $X=-0.19 $Y=1.66 $X2=5.55 $Y2=1.515
cc_52 VPB N_A_c_91_n 0.0479171f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=1.515
cc_53 VPB N_VPWR_c_284_n 0.011133f $X=-0.19 $Y=1.66 $X2=2.43 $Y2=2.4
cc_54 VPB N_VPWR_c_285_n 0.0383003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_286_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.675 $Y2=0.61
cc_56 VPB N_VPWR_c_287_n 0.00884785f $X=-0.19 $Y=1.66 $X2=2.88 $Y2=2.4
cc_57 VPB N_VPWR_c_288_n 0.00884785f $X=-0.19 $Y=1.66 $X2=3.245 $Y2=0.61
cc_58 VPB N_VPWR_c_289_n 0.00884785f $X=-0.19 $Y=1.66 $X2=3.38 $Y2=2.4
cc_59 VPB N_VPWR_c_290_n 0.00884785f $X=-0.19 $Y=1.66 $X2=3.675 $Y2=0.61
cc_60 VPB N_VPWR_c_291_n 0.00884785f $X=-0.19 $Y=1.66 $X2=3.83 $Y2=2.4
cc_61 VPB N_VPWR_c_292_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_293_n 0.0370432f $X=-0.19 $Y=1.66 $X2=4.245 $Y2=0.61
cc_63 VPB N_VPWR_c_294_n 0.0196495f $X=-0.19 $Y=1.66 $X2=4.33 $Y2=2.4
cc_64 VPB N_VPWR_c_295_n 0.0196495f $X=-0.19 $Y=1.66 $X2=4.675 $Y2=0.61
cc_65 VPB N_VPWR_c_296_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_297_n 0.0196495f $X=-0.19 $Y=1.66 $X2=5.28 $Y2=1.68
cc_67 VPB N_VPWR_c_298_n 0.0196495f $X=-0.19 $Y=1.66 $X2=5.73 $Y2=2.4
cc_68 VPB N_VPWR_c_299_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_69 VPB N_VPWR_c_300_n 0.0047828f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=1.58
cc_70 VPB N_VPWR_c_301_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_302_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_303_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.515
cc_73 VPB N_VPWR_c_283_n 0.076034f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=1.515
cc_74 VPB N_Y_c_381_n 0.00618364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_Y_c_395_n 0.00231613f $X=-0.19 $Y=1.66 $X2=3.245 $Y2=0.61
cc_76 VPB N_Y_c_396_n 0.00231613f $X=-0.19 $Y=1.66 $X2=3.675 $Y2=0.61
cc_77 VPB N_Y_c_397_n 0.00231613f $X=-0.19 $Y=1.66 $X2=4.245 $Y2=1.35
cc_78 VPB N_Y_c_398_n 0.00231613f $X=-0.19 $Y=1.66 $X2=4.78 $Y2=1.68
cc_79 VPB N_Y_c_399_n 0.00231613f $X=-0.19 $Y=1.66 $X2=5.73 $Y2=1.68
cc_80 VPB N_Y_c_400_n 0.00231613f $X=-0.19 $Y=1.66 $X2=3.035 $Y2=1.58
cc_81 VPB N_Y_c_401_n 0.00714919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB Y 0.0128198f $X=-0.19 $Y=1.66 $X2=5.28 $Y2=1.515
cc_83 N_A_M1002_g N_VPWR_c_285_n 0.00507182f $X=0.53 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_M1002_g N_VPWR_c_286_n 0.005209f $X=0.53 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_VPWR_c_286_n 0.005209f $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_VPWR_c_287_n 0.00306788f $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_VPWR_c_287_n 0.00318542f $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_M1005_g N_VPWR_c_288_n 0.00306788f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_VPWR_c_288_n 0.00318542f $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_M1007_g N_VPWR_c_289_n 0.00306788f $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_M1008_g N_VPWR_c_289_n 0.00318542f $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_M1009_g N_VPWR_c_290_n 0.00306788f $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A_M1010_g N_VPWR_c_290_n 0.00318542f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A_M1011_g N_VPWR_c_291_n 0.00306788f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A_M1013_g N_VPWR_c_291_n 0.00318542f $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A_M1014_g N_VPWR_c_293_n 0.00501904f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_M1004_g N_VPWR_c_294_n 0.005209f $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_M1005_g N_VPWR_c_294_n 0.005209f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_M1006_g N_VPWR_c_295_n 0.005209f $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_M1007_g N_VPWR_c_295_n 0.005209f $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_M1008_g N_VPWR_c_296_n 0.005209f $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_M1009_g N_VPWR_c_296_n 0.005209f $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_M1010_g N_VPWR_c_297_n 0.005209f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_M1011_g N_VPWR_c_297_n 0.005209f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_M1013_g N_VPWR_c_298_n 0.005209f $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_M1014_g N_VPWR_c_298_n 0.005209f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_M1002_g N_VPWR_c_283_n 0.00986091f $X=0.53 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_M1003_g N_VPWR_c_283_n 0.00982754f $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_M1004_g N_VPWR_c_283_n 0.00982082f $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_M1005_g N_VPWR_c_283_n 0.00982754f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_M1006_g N_VPWR_c_283_n 0.00982082f $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_M1007_g N_VPWR_c_283_n 0.00982754f $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_M1008_g N_VPWR_c_283_n 0.00982082f $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_M1009_g N_VPWR_c_283_n 0.00982754f $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A_M1010_g N_VPWR_c_283_n 0.00982082f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A_M1011_g N_VPWR_c_283_n 0.00982754f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_M1013_g N_VPWR_c_283_n 0.00982082f $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_M1014_g N_VPWR_c_283_n 0.00986025f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_M1000_g N_Y_c_381_n 0.00957473f $X=0.515 $Y=0.61 $X2=0 $Y2=0
cc_120 N_A_M1002_g N_Y_c_381_n 0.00861357f $X=0.53 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_M1003_g N_Y_c_381_n 6.3743e-19 $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_c_104_n N_Y_c_381_n 0.0330139f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_c_91_n N_Y_c_381_n 0.0106828f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_M1002_g N_Y_c_395_n 0.0169136f $X=0.53 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_Y_c_395_n 0.0124648f $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_M1004_g N_Y_c_395_n 6.38607e-19 $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_M1003_g N_Y_c_411_n 0.0132272f $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_M1004_g N_Y_c_411_n 0.0132272f $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_c_91_n N_Y_c_411_n 7.63416e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_M1002_g N_Y_c_414_n 0.0198755f $X=0.53 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A_M1003_g N_Y_c_414_n 9.43996e-19 $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_c_104_n N_Y_c_414_n 0.0624734f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_91_n N_Y_c_414_n 4.90767e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_c_104_n N_Y_c_382_n 0.191911f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A_c_91_n N_Y_c_382_n 0.0403224f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_M1000_g N_Y_c_383_n 0.0311196f $X=0.515 $Y=0.61 $X2=0 $Y2=0
cc_137 N_A_c_104_n N_Y_c_383_n 0.0302039f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_91_n N_Y_c_383_n 0.00768078f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A_M1003_g N_Y_c_396_n 6.10838e-19 $X=0.98 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_M1004_g N_Y_c_396_n 0.0118711f $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_M1005_g N_Y_c_396_n 0.0123563f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1006_g N_Y_c_396_n 6.3785e-19 $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_M1005_g N_Y_c_427_n 0.0132272f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_M1006_g N_Y_c_427_n 0.0132272f $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_c_104_n N_Y_c_427_n 0.0431694f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A_c_91_n N_Y_c_427_n 7.63416e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A_M1005_g N_Y_c_397_n 6.10838e-19 $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_M1006_g N_Y_c_397_n 0.0118711f $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_M1007_g N_Y_c_397_n 0.0123563f $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1008_g N_Y_c_397_n 6.3785e-19 $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_M1001_g N_Y_c_384_n 0.0118691f $X=2.675 $Y=0.61 $X2=0 $Y2=0
cc_152 N_A_M1012_g N_Y_c_384_n 0.0118691f $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_153 N_A_c_91_n N_Y_c_384_n 0.00624771f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_M1007_g N_Y_c_438_n 0.0132272f $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_M1008_g N_Y_c_438_n 0.0132272f $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_c_104_n N_Y_c_438_n 0.0431694f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_157 N_A_c_91_n N_Y_c_438_n 7.54951e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A_M1001_g N_Y_c_442_n 8.00299e-19 $X=2.675 $Y=0.61 $X2=0 $Y2=0
cc_159 N_A_M1012_g N_Y_c_442_n 0.0109339f $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_160 N_A_M1015_g N_Y_c_442_n 0.0109374f $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_161 N_A_M1016_g N_Y_c_442_n 8.00492e-19 $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_162 N_A_M1007_g N_Y_c_398_n 6.10838e-19 $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_M1008_g N_Y_c_398_n 0.0118711f $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_M1009_g N_Y_c_398_n 0.0123563f $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A_M1010_g N_Y_c_398_n 6.3785e-19 $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_M1015_g N_Y_c_385_n 0.0118691f $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_167 N_A_M1016_g N_Y_c_385_n 0.0118691f $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_168 N_A_c_104_n N_Y_c_385_n 0.050393f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A_c_91_n N_Y_c_385_n 0.00605072f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A_M1009_g N_Y_c_454_n 0.0132272f $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_M1010_g N_Y_c_454_n 0.0132272f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_c_104_n N_Y_c_454_n 0.0431694f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A_c_91_n N_Y_c_454_n 7.58478e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A_M1015_g N_Y_c_458_n 8.00492e-19 $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_175 N_A_M1016_g N_Y_c_458_n 0.0109374f $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_176 N_A_M1017_g N_Y_c_458_n 0.0109374f $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_177 N_A_M1018_g N_Y_c_458_n 8.00492e-19 $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_178 N_A_M1009_g N_Y_c_399_n 6.10838e-19 $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_M1010_g N_Y_c_399_n 0.0118711f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_M1011_g N_Y_c_399_n 0.0123563f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_M1013_g N_Y_c_399_n 6.3785e-19 $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_M1017_g N_Y_c_386_n 0.0118691f $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_183 N_A_M1018_g N_Y_c_386_n 0.0118691f $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_184 N_A_c_104_n N_Y_c_386_n 0.050393f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A_c_91_n N_Y_c_386_n 0.00585372f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A_M1011_g N_Y_c_470_n 0.0132272f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_M1013_g N_Y_c_470_n 0.0132272f $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_c_104_n N_Y_c_470_n 0.0431694f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A_c_91_n N_Y_c_470_n 7.62005e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A_M1017_g N_Y_c_387_n 8.00492e-19 $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_191 N_A_M1018_g N_Y_c_387_n 0.0109496f $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_192 N_A_M1019_g N_Y_c_387_n 0.00729782f $X=5.745 $Y=0.61 $X2=0 $Y2=0
cc_193 N_A_M1011_g N_Y_c_400_n 6.10838e-19 $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_M1013_g N_Y_c_400_n 0.0118711f $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_M1014_g N_Y_c_400_n 0.0167812f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_M1019_g N_Y_c_388_n 0.0193631f $X=5.745 $Y=0.61 $X2=0 $Y2=0
cc_197 N_A_c_104_n N_Y_c_388_n 0.00669825f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A_M1014_g N_Y_c_401_n 0.0175619f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_c_104_n N_Y_c_401_n 0.00324945f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A_M1004_g N_Y_c_484_n 8.84614e-19 $X=1.48 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_M1005_g N_Y_c_484_n 8.84614e-19 $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_c_104_n N_Y_c_484_n 0.0235495f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A_c_91_n N_Y_c_484_n 5.54777e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_204 N_A_M1001_g N_Y_c_389_n 0.0177984f $X=2.675 $Y=0.61 $X2=0 $Y2=0
cc_205 N_A_M1012_g N_Y_c_389_n 7.94581e-19 $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_206 N_A_M1006_g N_Y_c_490_n 8.84614e-19 $X=2.43 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_M1007_g N_Y_c_490_n 8.84614e-19 $X=2.88 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_c_104_n N_Y_c_490_n 0.0235495f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_209 N_A_c_91_n N_Y_c_490_n 5.48413e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A_M1012_g N_Y_c_390_n 0.00279308f $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_211 N_A_M1015_g N_Y_c_390_n 0.00279308f $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_212 N_A_c_104_n N_Y_c_390_n 0.0281223f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A_c_91_n N_Y_c_390_n 0.00272398f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_214 N_A_M1008_g N_Y_c_498_n 8.84614e-19 $X=3.38 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_M1009_g N_Y_c_498_n 8.84614e-19 $X=3.83 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A_c_104_n N_Y_c_498_n 0.0235495f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_c_91_n N_Y_c_498_n 5.48413e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_218 N_A_M1016_g N_Y_c_391_n 0.00279308f $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_219 N_A_M1017_g N_Y_c_391_n 0.00279308f $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_220 N_A_c_104_n N_Y_c_391_n 0.0281223f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_221 N_A_c_91_n N_Y_c_391_n 0.00272398f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_222 N_A_M1010_g N_Y_c_506_n 8.84614e-19 $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_M1011_g N_Y_c_506_n 8.84614e-19 $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A_c_104_n N_Y_c_506_n 0.0235495f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_225 N_A_c_91_n N_Y_c_506_n 5.48413e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_226 N_A_M1018_g N_Y_c_392_n 0.00319101f $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_227 N_A_c_104_n N_Y_c_392_n 0.0282341f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A_c_91_n N_Y_c_392_n 0.0042758f $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A_M1013_g N_Y_c_513_n 8.84614e-19 $X=5.28 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A_M1014_g N_Y_c_513_n 8.84614e-19 $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A_c_104_n N_Y_c_513_n 0.0235495f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_232 N_A_c_91_n N_Y_c_513_n 5.54777e-19 $X=5.745 $Y=1.515 $X2=0 $Y2=0
cc_233 N_A_M1019_g Y 0.0257851f $X=5.745 $Y=0.61 $X2=0 $Y2=0
cc_234 N_A_c_104_n Y 0.0349176f $X=5.55 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A_M1000_g N_VGND_c_575_n 0.0138212f $X=0.515 $Y=0.61 $X2=0 $Y2=0
cc_236 N_A_M1001_g N_VGND_c_576_n 0.00605361f $X=2.675 $Y=0.61 $X2=0 $Y2=0
cc_237 N_A_M1012_g N_VGND_c_576_n 0.00441793f $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_238 N_A_M1015_g N_VGND_c_577_n 0.00441793f $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_239 N_A_M1016_g N_VGND_c_577_n 0.00441793f $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_240 N_A_M1017_g N_VGND_c_578_n 0.00441793f $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_241 N_A_M1018_g N_VGND_c_578_n 0.00441793f $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_242 N_A_M1018_g N_VGND_c_580_n 4.79211e-19 $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_243 N_A_M1019_g N_VGND_c_580_n 0.0107071f $X=5.745 $Y=0.61 $X2=0 $Y2=0
cc_244 N_A_M1000_g N_VGND_c_581_n 0.00536147f $X=0.515 $Y=0.61 $X2=0 $Y2=0
cc_245 N_A_M1001_g N_VGND_c_581_n 0.00531206f $X=2.675 $Y=0.61 $X2=0 $Y2=0
cc_246 N_A_M1012_g N_VGND_c_583_n 0.00531901f $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_247 N_A_M1015_g N_VGND_c_583_n 0.00531901f $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_248 N_A_M1016_g N_VGND_c_585_n 0.00531901f $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_249 N_A_M1017_g N_VGND_c_585_n 0.00531901f $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_250 N_A_M1018_g N_VGND_c_586_n 0.00531901f $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_251 N_A_M1019_g N_VGND_c_586_n 0.00462012f $X=5.745 $Y=0.61 $X2=0 $Y2=0
cc_252 N_A_M1000_g N_VGND_c_588_n 0.00521957f $X=0.515 $Y=0.61 $X2=0 $Y2=0
cc_253 N_A_M1001_g N_VGND_c_588_n 0.00536257f $X=2.675 $Y=0.61 $X2=0 $Y2=0
cc_254 N_A_M1012_g N_VGND_c_588_n 0.00536257f $X=3.245 $Y=0.61 $X2=0 $Y2=0
cc_255 N_A_M1015_g N_VGND_c_588_n 0.00536257f $X=3.675 $Y=0.61 $X2=0 $Y2=0
cc_256 N_A_M1016_g N_VGND_c_588_n 0.00536257f $X=4.245 $Y=0.61 $X2=0 $Y2=0
cc_257 N_A_M1017_g N_VGND_c_588_n 0.00536257f $X=4.675 $Y=0.61 $X2=0 $Y2=0
cc_258 N_A_M1018_g N_VGND_c_588_n 0.00536257f $X=5.245 $Y=0.61 $X2=0 $Y2=0
cc_259 N_A_M1019_g N_VGND_c_588_n 0.00450456f $X=5.745 $Y=0.61 $X2=0 $Y2=0
cc_260 N_VPWR_M1002_s N_Y_c_381_n 0.00448393f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_261 N_VPWR_c_285_n N_Y_c_395_n 0.0234181f $X=0.29 $Y=2.455 $X2=0 $Y2=0
cc_262 N_VPWR_c_286_n N_Y_c_395_n 0.0144623f $X=1.12 $Y=3.33 $X2=0 $Y2=0
cc_263 N_VPWR_c_287_n N_Y_c_395_n 0.0234083f $X=1.205 $Y=2.455 $X2=0 $Y2=0
cc_264 N_VPWR_c_283_n N_Y_c_395_n 0.0118344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_M1003_s N_Y_c_411_n 0.00410979f $X=1.07 $Y=1.84 $X2=0 $Y2=0
cc_266 N_VPWR_c_287_n N_Y_c_411_n 0.0167599f $X=1.205 $Y=2.455 $X2=0 $Y2=0
cc_267 N_VPWR_M1002_s N_Y_c_414_n 0.00889652f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_268 N_VPWR_c_285_n N_Y_c_414_n 0.00793666f $X=0.29 $Y=2.455 $X2=0 $Y2=0
cc_269 N_VPWR_c_287_n N_Y_c_396_n 0.0266484f $X=1.205 $Y=2.455 $X2=0 $Y2=0
cc_270 N_VPWR_c_288_n N_Y_c_396_n 0.0234083f $X=2.155 $Y=2.455 $X2=0 $Y2=0
cc_271 N_VPWR_c_294_n N_Y_c_396_n 0.0144623f $X=2.07 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_283_n N_Y_c_396_n 0.0118344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_M1005_s N_Y_c_427_n 0.00410979f $X=2.02 $Y=1.84 $X2=0 $Y2=0
cc_274 N_VPWR_c_288_n N_Y_c_427_n 0.0167599f $X=2.155 $Y=2.455 $X2=0 $Y2=0
cc_275 N_VPWR_c_288_n N_Y_c_397_n 0.0266484f $X=2.155 $Y=2.455 $X2=0 $Y2=0
cc_276 N_VPWR_c_289_n N_Y_c_397_n 0.0234083f $X=3.105 $Y=2.455 $X2=0 $Y2=0
cc_277 N_VPWR_c_295_n N_Y_c_397_n 0.0144623f $X=3.02 $Y=3.33 $X2=0 $Y2=0
cc_278 N_VPWR_c_283_n N_Y_c_397_n 0.0118344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_M1007_s N_Y_c_438_n 0.00410979f $X=2.97 $Y=1.84 $X2=0 $Y2=0
cc_280 N_VPWR_c_289_n N_Y_c_438_n 0.0167599f $X=3.105 $Y=2.455 $X2=0 $Y2=0
cc_281 N_VPWR_c_289_n N_Y_c_398_n 0.0266484f $X=3.105 $Y=2.455 $X2=0 $Y2=0
cc_282 N_VPWR_c_290_n N_Y_c_398_n 0.0234083f $X=4.055 $Y=2.455 $X2=0 $Y2=0
cc_283 N_VPWR_c_296_n N_Y_c_398_n 0.0144623f $X=3.97 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VPWR_c_283_n N_Y_c_398_n 0.0118344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_M1009_s N_Y_c_454_n 0.00410979f $X=3.92 $Y=1.84 $X2=0 $Y2=0
cc_286 N_VPWR_c_290_n N_Y_c_454_n 0.0167599f $X=4.055 $Y=2.455 $X2=0 $Y2=0
cc_287 N_VPWR_c_290_n N_Y_c_399_n 0.0266484f $X=4.055 $Y=2.455 $X2=0 $Y2=0
cc_288 N_VPWR_c_291_n N_Y_c_399_n 0.0234083f $X=5.005 $Y=2.455 $X2=0 $Y2=0
cc_289 N_VPWR_c_297_n N_Y_c_399_n 0.0144623f $X=4.92 $Y=3.33 $X2=0 $Y2=0
cc_290 N_VPWR_c_283_n N_Y_c_399_n 0.0118344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_M1011_s N_Y_c_470_n 0.00410979f $X=4.87 $Y=1.84 $X2=0 $Y2=0
cc_292 N_VPWR_c_291_n N_Y_c_470_n 0.0167599f $X=5.005 $Y=2.455 $X2=0 $Y2=0
cc_293 N_VPWR_c_291_n N_Y_c_400_n 0.0266484f $X=5.005 $Y=2.455 $X2=0 $Y2=0
cc_294 N_VPWR_c_293_n N_Y_c_400_n 0.0234083f $X=5.955 $Y=2.455 $X2=0 $Y2=0
cc_295 N_VPWR_c_298_n N_Y_c_400_n 0.0144623f $X=5.87 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_c_283_n N_Y_c_400_n 0.0118344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_297 N_VPWR_M1014_s N_Y_c_401_n 0.00365063f $X=5.82 $Y=1.84 $X2=0 $Y2=0
cc_298 N_VPWR_c_293_n N_Y_c_401_n 0.0213127f $X=5.955 $Y=2.455 $X2=0 $Y2=0
cc_299 N_VPWR_M1014_s Y 0.00184872f $X=5.82 $Y=1.84 $X2=0 $Y2=0
cc_300 N_Y_c_383_n N_VGND_c_575_n 0.00947664f $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_301 N_Y_c_384_n N_VGND_c_576_n 0.0206815f $X=3.295 $Y=1.095 $X2=0 $Y2=0
cc_302 N_Y_c_385_n N_VGND_c_577_n 0.0206815f $X=4.295 $Y=1.095 $X2=0 $Y2=0
cc_303 N_Y_c_386_n N_VGND_c_578_n 0.0206815f $X=5.295 $Y=1.095 $X2=0 $Y2=0
cc_304 N_Y_c_388_n N_VGND_c_580_n 0.0203245f $X=5.885 $Y=1.095 $X2=0 $Y2=0
cc_305 N_Y_c_382_n N_VGND_c_581_n 0.0483046f $X=2.265 $Y=0.82 $X2=0 $Y2=0
cc_306 N_Y_c_383_n N_VGND_c_581_n 0.0103163f $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_307 N_Y_c_442_n N_VGND_c_583_n 0.00846545f $X=3.46 $Y=0.61 $X2=0 $Y2=0
cc_308 N_Y_c_458_n N_VGND_c_585_n 0.00846545f $X=4.46 $Y=0.61 $X2=0 $Y2=0
cc_309 N_Y_c_387_n N_VGND_c_586_n 0.00918079f $X=5.46 $Y=0.61 $X2=0 $Y2=0
cc_310 N_Y_c_382_n N_VGND_c_588_n 0.0567884f $X=2.265 $Y=0.82 $X2=0 $Y2=0
cc_311 N_Y_c_383_n N_VGND_c_588_n 0.0124117f $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_312 N_Y_c_442_n N_VGND_c_588_n 0.0113241f $X=3.46 $Y=0.61 $X2=0 $Y2=0
cc_313 N_Y_c_458_n N_VGND_c_588_n 0.0113241f $X=4.46 $Y=0.61 $X2=0 $Y2=0
cc_314 N_Y_c_387_n N_VGND_c_588_n 0.0113609f $X=5.46 $Y=0.61 $X2=0 $Y2=0

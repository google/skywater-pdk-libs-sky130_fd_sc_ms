* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_293_74# a_141_385# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_112_119# B a_141_385# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VGND B a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR A a_141_385# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X4 a_141_385# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 VGND A a_112_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 Y a_141_385# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VPWR A a_379_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_293_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_379_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

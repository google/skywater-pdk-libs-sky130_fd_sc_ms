* File: sky130_fd_sc_ms__or3_1.spice
* Created: Fri Aug 28 18:07:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or3_1.pex.spice"
.subckt sky130_fd_sc_ms__or3_1  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_C_M1007_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.15675 PD=0.9 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1003 N_A_27_74#_M1003_d N_B_M1003_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.182875 AS=0.09625 PD=1.215 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_27_74#_M1003_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.11874 AS=0.182875 PD=0.989147 PS=1.215 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1005 N_X_M1005_d N_A_27_74#_M1005_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.15976 PD=2.05 PS=1.33085 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 A_119_368# N_C_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90002.1
+ A=0.18 P=2.36 MULT=1
MM1002 A_203_368# N_B_M1002_g A_119_368# VPB PSHORT L=0.18 W=1 AD=0.195 AS=0.12
+ PD=1.39 PS=1.24 NRD=27.5603 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90001.6
+ A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_203_368# VPB PSHORT L=0.18 W=1 AD=0.34434
+ AS=0.195 PD=1.71698 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90001.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1004_d N_A_27_74#_M1004_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.38566 PD=2.8 PS=1.92302 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__or3_1.pxi.spice"
*
.ends
*
*

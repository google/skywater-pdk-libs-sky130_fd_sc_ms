* File: sky130_fd_sc_ms__nor3_4.pex.spice
* Created: Fri Aug 28 17:48:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR3_4%A 3 7 11 15 17 19 20 22 23 25 28 30 34 35 39
+ 40 44 45 46 57 60
c132 46 0 9.21872e-20 $X=1.68 $Y=2.035
c133 30 0 1.39786e-19 $X=5.805 $Y=2.105
c134 25 0 1.07767e-19 $X=0.77 $Y=1.515
c135 15 0 1.53462e-19 $X=0.95 $Y=2.4
c136 11 0 7.79871e-20 $X=0.935 $Y=0.74
r137 60 71 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.71 $Y=2.045
+ $X2=1.71 $Y2=2.255
r138 57 58 2.21101 $w=3.27e-07 $l=1.5e-08 $layer=POLY_cond $X=0.935 $Y=1.515
+ $X2=0.95 $Y2=1.515
r139 54 55 0.737003 $w=3.27e-07 $l=5e-09 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.5 $Y2=1.515
r140 46 60 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=2.045
r141 46 60 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.61 $Y=2.045
+ $X2=1.625 $Y2=2.045
r142 45 46 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=2.045
+ $X2=1.61 $Y2=2.045
r143 45 61 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=2.045
+ $X2=0.935 $Y2=2.045
r144 44 61 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=2.045
+ $X2=0.935 $Y2=2.045
r145 40 42 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.935 $Y=2.105
+ $X2=3.935 $Y2=2.255
r146 39 51 10.6277 $w=5.7e-07 $l=1.2e-07 $layer=POLY_cond $X=6 $Y=1.515 $X2=6
+ $Y2=1.395
r147 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=1.515 $X2=5.97 $Y2=1.515
r148 35 51 84.4783 $w=5.7e-07 $l=9e-07 $layer=POLY_cond $X=6 $Y=0.495 $X2=6
+ $Y2=1.395
r149 34 38 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=5.97 $Y=0.495
+ $X2=5.97 $Y2=1.515
r150 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=0.495 $X2=5.97 $Y2=0.495
r151 32 38 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=5.97 $Y=2.02
+ $X2=5.97 $Y2=1.515
r152 31 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.105
+ $X2=3.935 $Y2=2.105
r153 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.805 $Y=2.105
+ $X2=5.97 $Y2=2.02
r154 30 31 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=5.805 $Y=2.105
+ $X2=4.02 $Y2=2.105
r155 29 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.255
+ $X2=1.71 $Y2=2.255
r156 28 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.255
+ $X2=3.935 $Y2=2.255
r157 28 29 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=3.85 $Y=2.255
+ $X2=1.795 $Y2=2.255
r158 26 57 24.3211 $w=3.27e-07 $l=1.65e-07 $layer=POLY_cond $X=0.77 $Y=1.515
+ $X2=0.935 $Y2=1.515
r159 26 55 39.7982 $w=3.27e-07 $l=2.7e-07 $layer=POLY_cond $X=0.77 $Y=1.515
+ $X2=0.5 $Y2=1.515
r160 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.515 $X2=0.77 $Y2=1.515
r161 23 44 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.77 $Y=1.92
+ $X2=0.77 $Y2=2.045
r162 23 25 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.77 $Y=1.92
+ $X2=0.77 $Y2=1.515
r163 20 39 48.3446 $w=2.59e-07 $l=3.49857e-07 $layer=POLY_cond $X=6.225 $Y=1.77
+ $X2=6 $Y2=1.515
r164 20 22 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=6.225 $Y=1.77
+ $X2=6.225 $Y2=2.4
r165 17 39 48.3446 $w=2.59e-07 $l=3.49857e-07 $layer=POLY_cond $X=5.775 $Y=1.77
+ $X2=6 $Y2=1.515
r166 17 19 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=5.775 $Y=1.77
+ $X2=5.775 $Y2=2.4
r167 13 58 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.68
+ $X2=0.95 $Y2=1.515
r168 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.95 $Y=1.68
+ $X2=0.95 $Y2=2.4
r169 9 57 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.35
+ $X2=0.935 $Y2=1.515
r170 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.935 $Y=1.35
+ $X2=0.935 $Y2=0.74
r171 5 54 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r172 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
r173 1 55 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.68 $X2=0.5
+ $Y2=1.515
r174 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.5 $Y=1.68 $X2=0.5
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%B 5 7 9 10 12 14 17 21 25 27 32 35 39 41 42
+ 48 53 55 56 60 62 64 66
c118 53 0 1.39786e-19 $X=5.325 $Y=1.345
c119 48 0 9.21872e-20 $X=1.475 $Y=1.68
c120 32 0 1.58468e-19 $X=4.8 $Y=1.345
c121 25 0 6.80408e-20 $X=5.325 $Y=2.4
c122 12 0 4.22428e-20 $X=1.925 $Y=1.185
r123 56 62 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=1.35
+ $X2=2.16 $Y2=1.35
r124 55 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=1.35
+ $X2=2.64 $Y2=1.35
r125 52 53 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=4.875 $Y=1.345
+ $X2=5.325 $Y2=1.345
r126 42 66 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=2.655 $Y=1.35
+ $X2=2.755 $Y2=1.35
r127 42 64 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.655 $Y=1.35
+ $X2=2.64 $Y2=1.35
r128 42 55 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.57 $Y=1.35
+ $X2=2.585 $Y2=1.35
r129 41 62 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=1.35
+ $X2=2.16 $Y2=1.35
r130 41 60 6.26872 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=2.145 $Y=1.35
+ $X2=2.045 $Y2=1.35
r131 41 42 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.23 $Y=1.35
+ $X2=2.57 $Y2=1.35
r132 41 56 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.23 $Y=1.35
+ $X2=2.215 $Y2=1.35
r133 39 48 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.515
+ $X2=1.475 $Y2=1.68
r134 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.475
+ $Y=1.515 $X2=1.475 $Y2=1.515
r135 35 38 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.475 $Y=1.435
+ $X2=1.475 $Y2=1.515
r136 33 52 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.8 $Y=1.345
+ $X2=4.875 $Y2=1.345
r137 33 49 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.8 $Y=1.345
+ $X2=4.425 $Y2=1.345
r138 32 66 71.4165 $w=3.28e-07 $l=2.045e-06 $layer=LI1_cond $X=4.8 $Y=1.345
+ $X2=2.755 $Y2=1.345
r139 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.8
+ $Y=1.345 $X2=4.8 $Y2=1.345
r140 29 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=1.435
+ $X2=1.475 $Y2=1.435
r141 29 60 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.64 $Y=1.435
+ $X2=2.045 $Y2=1.435
r142 23 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.51
+ $X2=5.325 $Y2=1.345
r143 23 25 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=5.325 $Y=1.51
+ $X2=5.325 $Y2=2.4
r144 19 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.51
+ $X2=4.875 $Y2=1.345
r145 19 21 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=4.875 $Y=1.51
+ $X2=4.875 $Y2=2.4
r146 15 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.51
+ $X2=4.425 $Y2=1.345
r147 15 17 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=4.425 $Y=1.51
+ $X2=4.425 $Y2=2.4
r148 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.925 $Y=1.185
+ $X2=1.925 $Y2=0.74
r149 11 27 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.26
+ $X2=1.475 $Y2=1.26
r150 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.85 $Y=1.26
+ $X2=1.925 $Y2=1.185
r151 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.85 $Y=1.26
+ $X2=1.64 $Y2=1.26
r152 7 27 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=1.495 $Y=1.185
+ $X2=1.475 $Y2=1.26
r153 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.495 $Y=1.185
+ $X2=1.495 $Y2=0.74
r154 5 48 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.4 $Y=2.4 $X2=1.4
+ $Y2=1.68
r155 1 27 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.475 $Y=1.335
+ $X2=1.475 $Y2=1.26
r156 1 39 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.475 $Y=1.335
+ $X2=1.475 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%C 3 5 6 9 13 15 19 23 25 26 29 32 33 36 37 38
+ 39 40 41 50
c105 15 0 1.58468e-19 $X=2.85 $Y=1.62
c106 3 0 8.39251e-20 $X=2.005 $Y=2.4
r107 50 51 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.31
+ $Y=0.505 $X2=5.31 $Y2=0.505
r108 47 50 237.811 $w=3.3e-07 $l=1.36e-06 $layer=POLY_cond $X=3.95 $Y=0.505
+ $X2=5.31 $Y2=0.505
r109 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=0.505 $X2=3.95 $Y2=0.505
r110 41 51 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.52 $Y=0.505
+ $X2=5.31 $Y2=0.505
r111 40 51 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.04 $Y=0.505
+ $X2=5.31 $Y2=0.505
r112 39 40 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=0.505
+ $X2=5.04 $Y2=0.505
r113 38 39 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=0.505
+ $X2=4.56 $Y2=0.505
r114 38 48 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=0.505
+ $X2=3.95 $Y2=0.505
r115 37 47 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.905 $Y=0.505
+ $X2=3.95 $Y2=0.505
r116 32 36 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.83 $Y=1.545
+ $X2=3.815 $Y2=1.62
r117 31 37 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.83 $Y=0.67
+ $X2=3.905 $Y2=0.505
r118 31 32 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.83 $Y=0.67
+ $X2=3.83 $Y2=1.545
r119 27 36 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.815 $Y=1.695
+ $X2=3.815 $Y2=1.62
r120 27 29 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=3.815 $Y=1.695
+ $X2=3.815 $Y2=2.4
r121 25 36 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.725 $Y=1.62
+ $X2=3.815 $Y2=1.62
r122 25 26 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.725 $Y=1.62
+ $X2=3.305 $Y2=1.62
r123 21 26 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.215 $Y=1.62
+ $X2=3.305 $Y2=1.62
r124 21 34 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.215 $Y=1.62
+ $X2=2.925 $Y2=1.62
r125 21 23 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=3.215 $Y=1.695
+ $X2=3.215 $Y2=2.4
r126 17 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.925 $Y=1.545
+ $X2=2.925 $Y2=1.62
r127 17 19 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.925 $Y=1.545
+ $X2=2.925 $Y2=0.74
r128 16 33 13.2179 $w=1.5e-07 $l=1.38e-07 $layer=POLY_cond $X=2.695 $Y=1.62
+ $X2=2.557 $Y2=1.62
r129 15 34 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.85 $Y=1.62
+ $X2=2.925 $Y2=1.62
r130 15 16 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.85 $Y=1.62
+ $X2=2.695 $Y2=1.62
r131 11 33 10.9219 $w=1.8e-07 $l=9.60469e-08 $layer=POLY_cond $X=2.605 $Y=1.695
+ $X2=2.557 $Y2=1.62
r132 11 13 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=2.605 $Y=1.695
+ $X2=2.605 $Y2=2.4
r133 7 33 10.9219 $w=1.5e-07 $l=1.01366e-07 $layer=POLY_cond $X=2.495 $Y=1.545
+ $X2=2.557 $Y2=1.62
r134 7 9 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.495 $Y=1.545
+ $X2=2.495 $Y2=0.74
r135 5 33 13.2179 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=2.42 $Y=1.62
+ $X2=2.557 $Y2=1.62
r136 5 6 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.42 $Y=1.62
+ $X2=2.095 $Y2=1.62
r137 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.005 $Y=1.695
+ $X2=2.095 $Y2=1.62
r138 1 3 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=2.005 $Y=1.695
+ $X2=2.005 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%A_27_368# 1 2 3 4 5 18 22 24 28 30 32 36 38
+ 42 46 48 51 53 60 61
c86 30 0 4.80254e-20 $X=4.485 $Y=2.595
c87 28 0 2.37388e-19 $X=1.175 $Y=2.815
r88 56 57 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=4.61 $Y=2.545 $X2=4.61
+ $Y2=2.595
r89 53 56 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=4.61 $Y=2.445 $X2=4.61
+ $Y2=2.545
r90 51 52 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.215 $Y=2.425
+ $X2=1.215 $Y2=2.595
r91 44 61 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=2.53 $X2=6.49
+ $Y2=2.445
r92 44 46 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.49 $Y=2.53
+ $X2=6.49 $Y2=2.815
r93 40 61 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=2.36 $X2=6.49
+ $Y2=2.445
r94 40 42 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=6.49 $Y=2.36
+ $X2=6.49 $Y2=1.985
r95 39 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=2.445
+ $X2=5.55 $Y2=2.445
r96 38 61 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.365 $Y=2.445
+ $X2=6.49 $Y2=2.445
r97 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.365 $Y=2.445
+ $X2=5.635 $Y2=2.445
r98 34 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=2.53 $X2=5.55
+ $Y2=2.445
r99 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.55 $Y=2.53
+ $X2=5.55 $Y2=2.835
r100 33 53 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.735 $Y=2.445
+ $X2=4.61 $Y2=2.445
r101 32 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=2.445
+ $X2=5.55 $Y2=2.445
r102 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.465 $Y=2.445
+ $X2=4.735 $Y2=2.445
r103 31 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=2.595
+ $X2=1.215 $Y2=2.595
r104 30 57 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.485 $Y=2.595
+ $X2=4.61 $Y2=2.595
r105 30 31 205.182 $w=1.68e-07 $l=3.145e-06 $layer=LI1_cond $X=4.485 $Y=2.595
+ $X2=1.34 $Y2=2.595
r106 26 52 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.68
+ $X2=1.215 $Y2=2.595
r107 26 28 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.215 $Y=2.68
+ $X2=1.215 $Y2=2.815
r108 25 48 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.36 $Y=2.425
+ $X2=0.235 $Y2=2.425
r109 24 51 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.09 $Y=2.425
+ $X2=1.215 $Y2=2.425
r110 24 25 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.09 $Y=2.425
+ $X2=0.36 $Y2=2.425
r111 20 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.51
+ $X2=0.235 $Y2=2.425
r112 20 22 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.235 $Y=2.51
+ $X2=0.235 $Y2=2.815
r113 16 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.34
+ $X2=0.235 $Y2=2.425
r114 16 18 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.235 $Y=2.34
+ $X2=0.235 $Y2=1.985
r115 5 46 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.315
+ $Y=1.84 $X2=6.45 $Y2=2.815
r116 5 42 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.315
+ $Y=1.84 $X2=6.45 $Y2=1.985
r117 4 60 600 $w=1.7e-07 $l=6.69104e-07 $layer=licon1_PDIFF $count=1 $X=5.415
+ $Y=1.84 $X2=5.55 $Y2=2.445
r118 4 36 600 $w=1.7e-07 $l=1.06035e-06 $layer=licon1_PDIFF $count=1 $X=5.415
+ $Y=1.84 $X2=5.55 $Y2=2.835
r119 3 56 600 $w=1.7e-07 $l=7.69545e-07 $layer=licon1_PDIFF $count=1 $X=4.515
+ $Y=1.84 $X2=4.65 $Y2=2.545
r120 2 51 600 $w=1.7e-07 $l=6.48999e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.84 $X2=1.175 $Y2=2.425
r121 2 28 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.84 $X2=1.175 $Y2=2.815
r122 1 22 600 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=2.815
r123 1 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%VPWR 1 2 9 13 15 17 22 32 33 36 39
c69 1 0 1.07767e-19 $X=0.59 $Y=1.84
r70 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r71 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r73 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r74 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33 $X2=6
+ $Y2=3.33
r75 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.48 $Y2=3.33
r76 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r77 28 29 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 25 28 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=5.52
+ $Y2=3.33
r80 25 26 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r81 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r82 23 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33 $X2=6
+ $Y2=3.33
r84 22 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r88 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r89 15 29 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 15 26 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=1.2 $Y2=3.33
r91 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6 $Y=3.245 $X2=6
+ $Y2=3.33
r92 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6 $Y=3.245 $X2=6
+ $Y2=2.8
r93 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r94 7 9 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.79
r95 2 13 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=5.865
+ $Y=1.84 $X2=6 $Y2=2.8
r96 1 9 600 $w=1.7e-07 $l=1.01526e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.725 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%A_298_368# 1 2 3 4 13 21 25
c44 23 0 1.78868e-19 $X=4.285 $Y=2.962
c45 21 0 6.80408e-20 $X=4.935 $Y=2.99
r46 25 27 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.1 $Y=2.8 $X2=5.1
+ $Y2=2.99
r47 21 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=2.99
+ $X2=5.1 $Y2=2.99
r48 21 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.935 $Y=2.99
+ $X2=4.285 $Y2=2.99
r49 18 20 61.9758 $w=2.23e-07 $l=1.21e-06 $layer=LI1_cond $X=2.91 $Y=2.962
+ $X2=4.12 $Y2=2.962
r50 15 18 61.7197 $w=2.23e-07 $l=1.205e-06 $layer=LI1_cond $X=1.705 $Y=2.962
+ $X2=2.91 $Y2=2.962
r51 13 23 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=4.173 $Y=2.962
+ $X2=4.285 $Y2=2.962
r52 13 20 2.71464 $w=2.23e-07 $l=5.3e-08 $layer=LI1_cond $X=4.173 $Y=2.962
+ $X2=4.12 $Y2=2.962
r53 4 25 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.84 $X2=5.1 $Y2=2.8
r54 3 20 600 $w=1.7e-07 $l=1.19769e-06 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.12 $Y2=2.935
r55 2 18 600 $w=1.7e-07 $l=1.19769e-06 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=1.84 $X2=2.91 $Y2=2.935
r56 1 15 600 $w=1.7e-07 $l=1.19769e-06 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.84 $X2=1.705 $Y2=2.935
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%Y 1 2 3 4 5 16 17 20 22 30 32 34 37 39 42 45
+ 46 47
c112 39 0 7.79871e-20 $X=1.71 $Y=0.925
c113 37 0 1.82358e-19 $X=5.22 $Y=1.68
c114 34 0 4.80254e-20 $X=5.135 $Y=1.765
c115 16 0 4.22428e-20 $X=1.545 $Y=1.095
r116 44 46 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=1.84
+ $X2=3.68 $Y2=1.84
r117 44 45 6.52497 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=1.84
+ $X2=3.35 $Y2=1.84
r118 39 40 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.71 $Y=0.925
+ $X2=1.71 $Y2=1.095
r119 38 47 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.515
r120 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.22 $Y=1.01
+ $X2=5.22 $Y2=1.68
r121 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.135 $Y=1.765
+ $X2=5.22 $Y2=1.68
r122 34 46 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=5.135 $Y=1.765
+ $X2=3.68 $Y2=1.765
r123 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0.925
+ $X2=2.71 $Y2=0.925
r124 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.135 $Y=0.925
+ $X2=5.22 $Y2=1.01
r125 32 33 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=5.135 $Y=0.925
+ $X2=2.875 $Y2=0.925
r126 28 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.84
+ $X2=2.71 $Y2=0.925
r127 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.71 $Y=0.84
+ $X2=2.71 $Y2=0.515
r128 26 45 48.1721 $w=2.48e-07 $l=1.045e-06 $layer=LI1_cond $X=2.305 $Y=1.875
+ $X2=3.35 $Y2=1.875
r129 23 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.925
+ $X2=1.71 $Y2=0.925
r130 22 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0.925
+ $X2=2.71 $Y2=0.925
r131 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.545 $Y=0.925
+ $X2=1.875 $Y2=0.925
r132 18 39 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.84
+ $X2=1.71 $Y2=0.925
r133 18 20 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.71 $Y=0.84
+ $X2=1.71 $Y2=0.515
r134 17 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.875 $Y=1.095
+ $X2=0.71 $Y2=1.01
r135 16 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=1.71 $Y2=1.095
r136 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=0.875 $Y2=1.095
r137 5 44 600 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.84 $X2=3.515 $Y2=1.915
r138 4 26 600 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.84 $X2=2.305 $Y2=1.915
r139 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.515
r140 2 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.71 $Y2=0.515
r141 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3_4%VGND 1 2 3 4 13 15 19 23 25 29 31 33 38 48 49
+ 55 58 61
r62 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r64 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r65 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r66 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r67 48 49 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r68 46 49 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r69 45 48 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r70 45 46 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r71 43 61 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.21
+ $Y2=0
r72 43 45 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.6
+ $Y2=0
r73 42 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r74 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r75 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r76 39 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r77 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r78 38 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.21
+ $Y2=0
r79 38 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.68
+ $Y2=0
r80 37 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r81 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r82 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r83 34 52 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r84 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r85 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r86 33 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r87 31 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r88 31 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.12
+ $Y2=0
r89 27 61 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r90 27 29 15.6137 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.505
r91 26 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.21
+ $Y2=0
r92 25 61 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.21
+ $Y2=0
r93 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.375
+ $Y2=0
r94 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r95 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.55
r96 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r97 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.675
r98 13 52 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r99 13 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.515
r100 4 29 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.14 $Y2=0.505
r101 3 23 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.21 $Y2=0.55
r102 2 19 182 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.37 $X2=1.21 $Y2=0.675
r103 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends


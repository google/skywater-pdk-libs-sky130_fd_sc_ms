* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ms__maj3_2 A B C VGND VNB VPB VPWR X
*.PININFO A:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN2 X y VGND VNB nfet_01v8_lvt m=2 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN10 y B sndNBa VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN11 sndNBa A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN20 y B sndNBc VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN21 sndNBc C VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN30 y C sndNCa VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMN31 sndNCa A VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 X y VPWR VPB pfet_01v8 m=2 w=1.12 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP10 VPWR A sndPAb VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP11 sndPAb B y VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP20 VPWR C sndPCb VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP21 sndPCb B y VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP30 VPWR A sndPAc VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP31 sndPAc C y VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ms__maj3_2

* File: sky130_fd_sc_ms__xnor3_2.pex.spice
* Created: Fri Aug 28 18:18:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_83_247# 1 2 3 4 15 19 21 24 25 26 28 29 33
+ 34 35 37 38 39 44 45 48
c131 24 0 1.07216e-19 $X=0.58 $Y=1.4
r132 48 50 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.51 $Y=2.795
+ $X2=3.51 $Y2=2.99
r133 44 45 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.35
+ $X2=3.2 $Y2=0.35
r134 38 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=3.51 $Y2=2.99
r135 38 39 128.524 $w=1.68e-07 $l=1.97e-06 $layer=LI1_cond $X=3.345 $Y=2.99
+ $X2=1.375 $Y2=2.99
r136 37 45 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=1.345 $Y=0.34
+ $X2=3.2 $Y2=0.34
r137 35 39 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.375 $Y2=2.99
r138 34 42 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.035
r139 34 35 32.3096 $w=2.78e-07 $l=7.85e-07 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.905
r140 31 33 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=1.22 $Y=1.035
+ $X2=1.22 $Y2=0.55
r141 30 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.345 $Y2=0.34
r142 30 33 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.22 $Y2=0.55
r143 28 42 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=1.235 $Y2=2.035
r144 28 29 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=0.745 $Y2=2.035
r145 27 40 1.68994 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.12
+ $X2=0.62 $Y2=1.12
r146 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.095 $Y=1.12
+ $X2=1.22 $Y2=1.035
r147 26 27 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.095 $Y=1.12
+ $X2=0.745 $Y2=1.12
r148 25 54 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.4
+ $X2=0.58 $Y2=1.565
r149 25 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.4
+ $X2=0.58 $Y2=1.235
r150 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.4 $X2=0.58 $Y2=1.4
r151 22 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.745 $Y2=2.035
r152 22 24 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.62 $Y2=1.4
r153 21 40 12.2351 $w=2.5e-07 $l=2.4e-07 $layer=LI1_cond $X=0.62 $Y=1.36
+ $X2=0.62 $Y2=1.12
r154 21 24 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=0.62 $Y=1.36 $X2=0.62
+ $Y2=1.4
r155 19 53 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.535 $Y=0.725
+ $X2=0.535 $Y2=1.235
r156 15 54 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=0.505 $Y=2.365
+ $X2=0.505 $Y2=1.565
r157 4 48 600 $w=1.7e-07 $l=1.03192e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.865 $X2=3.51 $Y2=2.795
r158 3 42 300 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.865 $X2=1.28 $Y2=2.115
r159 2 44 182 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.625 $X2=3.365 $Y2=0.36
r160 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.12
+ $Y=0.405 $X2=1.26 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A 3 7 9 12 13
c45 12 0 3.99547e-20 $X=1.12 $Y=1.54
c46 7 0 2.53685e-19 $X=1.045 $Y=0.725
c47 3 0 1.91609e-19 $X=1.045 $Y=2.365
r48 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.54
+ $X2=1.12 $Y2=1.705
r49 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.54
+ $X2=1.12 $Y2=1.375
r50 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.54 $X2=1.12 $Y2=1.54
r51 9 13 4.00154 $w=3.58e-07 $l=1.25e-07 $layer=LI1_cond $X=1.135 $Y=1.665
+ $X2=1.135 $Y2=1.54
r52 7 14 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.045 $Y=0.725
+ $X2=1.045 $Y2=1.375
r53 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.045 $Y=2.365
+ $X2=1.045 $Y2=1.705
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_397_21# 1 2 10 11 13 15 16 20 23 32 33 35
+ 37 39 42 43 44
c117 43 0 1.94615e-19 $X=3.32 $Y=1.54
c118 42 0 1.16185e-19 $X=3.32 $Y=1.54
c119 23 0 2.55111e-19 $X=3.205 $Y=2.285
c120 11 0 1.69141e-19 $X=2.195 $Y=1.49
c121 10 0 6.5827e-20 $X=2.06 $Y=1.055
r122 46 48 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.07 $Y=1.54
+ $X2=3.205 $Y2=1.54
r123 43 48 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.32 $Y=1.54
+ $X2=3.205 $Y2=1.54
r124 42 45 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=1.54
+ $X2=3.36 $Y2=1.705
r125 42 44 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=1.54
+ $X2=3.36 $Y2=1.375
r126 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.54 $X2=3.32 $Y2=1.54
r127 37 39 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=3.565 $Y=2.075
+ $X2=4.09 $Y2=2.075
r128 33 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.565 $Y=1.04
+ $X2=3.925 $Y2=1.04
r129 32 37 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.48 $Y=1.95
+ $X2=3.565 $Y2=2.075
r130 32 45 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.48 $Y=1.95
+ $X2=3.48 $Y2=1.705
r131 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.48 $Y=1.125
+ $X2=3.565 $Y2=1.04
r132 29 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.48 $Y=1.125
+ $X2=3.48 $Y2=1.375
r133 21 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.705
+ $X2=3.205 $Y2=1.54
r134 21 23 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.205 $Y=1.705
+ $X2=3.205 $Y2=2.285
r135 18 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.375
+ $X2=3.07 $Y2=1.54
r136 18 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.07 $Y=1.375
+ $X2=3.07 $Y2=0.945
r137 17 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.07 $Y=0.255
+ $X2=3.07 $Y2=0.945
r138 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.995 $Y=0.18
+ $X2=3.07 $Y2=0.255
r139 15 16 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.995 $Y=0.18
+ $X2=2.135 $Y2=0.18
r140 11 25 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.195 $Y=1.415
+ $X2=2.06 $Y2=1.415
r141 11 13 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=2.195 $Y=1.49
+ $X2=2.195 $Y2=2.185
r142 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=1.34
+ $X2=2.06 $Y2=1.415
r143 8 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.06 $Y=1.34
+ $X2=2.06 $Y2=1.055
r144 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.06 $Y=0.255
+ $X2=2.135 $Y2=0.18
r145 7 10 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.06 $Y=0.255 $X2=2.06
+ $Y2=1.055
r146 2 39 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.84 $X2=4.09 $Y2=2.115
r147 1 35 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.445 $X2=3.925 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%B 3 5 8 9 10 13 18 19 22 25 29 33 34 35 42
+ 43
c122 33 0 3.0936e-20 $X=2.625 $Y=1.655
c123 18 0 7.64129e-20 $X=2.665 $Y=2.185
c124 13 0 1.16185e-19 $X=2.57 $Y=0.945
c125 3 0 2.86506e-20 $X=1.57 $Y=0.725
r126 41 43 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.24 $Y=1.515
+ $X2=4.315 $Y2=1.515
r127 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.24
+ $Y=1.515 $X2=4.24 $Y2=1.515
r128 39 41 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.14 $Y=1.515
+ $X2=4.24 $Y2=1.515
r129 37 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.8 $Y=1.515
+ $X2=4.14 $Y2=1.515
r130 35 42 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.07 $Y=1.665
+ $X2=4.07 $Y2=1.515
r131 32 33 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.625 $Y=1.505
+ $X2=2.625 $Y2=1.655
r132 27 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.68
+ $X2=4.315 $Y2=1.515
r133 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.315 $Y=1.68
+ $X2=4.315 $Y2=2.4
r134 23 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=1.515
r135 23 25 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.14 $Y2=0.815
r136 21 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.68
+ $X2=3.8 $Y2=1.515
r137 21 22 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=3.8 $Y=1.68
+ $X2=3.8 $Y2=3.075
r138 20 34 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.755 $Y=3.15
+ $X2=2.665 $Y2=3.15
r139 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.725 $Y=3.15
+ $X2=3.8 $Y2=3.075
r140 19 20 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=3.725 $Y=3.15
+ $X2=2.755 $Y2=3.15
r141 18 33 206.016 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=2.665 $Y=2.185
+ $X2=2.665 $Y2=1.655
r142 16 34 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=3.075
+ $X2=2.665 $Y2=3.15
r143 16 18 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.665 $Y=3.075
+ $X2=2.665 $Y2=2.185
r144 13 32 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.57 $Y=0.945
+ $X2=2.57 $Y2=1.505
r145 9 34 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.575 $Y=3.15
+ $X2=2.665 $Y2=3.15
r146 9 10 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.575 $Y=3.15
+ $X2=1.675 $Y2=3.15
r147 6 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.585 $Y=3.075
+ $X2=1.675 $Y2=3.15
r148 6 8 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.585 $Y=3.075
+ $X2=1.585 $Y2=2.285
r149 5 31 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.585 $Y=1.595
+ $X2=1.585 $Y2=1.505
r150 5 8 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.585 $Y=1.595
+ $X2=1.585 $Y2=2.285
r151 3 31 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.57 $Y=0.725
+ $X2=1.57 $Y2=1.505
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_1027_48# 1 2 9 13 15 18 21 24 28 31 32
r79 33 35 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=5.21 $Y=1.64
+ $X2=5.395 $Y2=1.64
r80 28 30 3.21434 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=1.085
+ $X2=6.555 $Y2=1.17
r81 24 32 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=6.687 $Y=2.132
+ $X2=6.687 $Y2=1.95
r82 24 26 3.10849 $w=3.65e-07 $l=9.3e-08 $layer=LI1_cond $X=6.687 $Y=2.132
+ $X2=6.687 $Y2=2.225
r83 22 31 6.95506 $w=2.27e-07 $l=1.9182e-07 $layer=LI1_cond $X=6.59 $Y=1.805
+ $X2=6.532 $Y2=1.64
r84 22 32 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.59 $Y=1.805
+ $X2=6.59 $Y2=1.95
r85 21 31 6.95506 $w=2.27e-07 $l=1.65e-07 $layer=LI1_cond $X=6.532 $Y=1.475
+ $X2=6.532 $Y2=1.64
r86 21 30 12.3332 $w=2.83e-07 $l=3.05e-07 $layer=LI1_cond $X=6.532 $Y=1.475
+ $X2=6.532 $Y2=1.17
r87 18 35 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.49 $Y=1.64
+ $X2=5.395 $Y2=1.64
r88 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.64 $X2=5.49 $Y2=1.64
r89 15 31 0.0443336 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=6.39 $Y=1.64
+ $X2=6.532 $Y2=1.64
r90 15 17 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=6.39 $Y=1.64 $X2=5.49
+ $Y2=1.64
r91 11 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.805
+ $X2=5.395 $Y2=1.64
r92 11 13 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=5.395 $Y=1.805
+ $X2=5.395 $Y2=2.415
r93 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.475
+ $X2=5.21 $Y2=1.64
r94 7 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.21 $Y=1.475
+ $X2=5.21 $Y2=0.69
r95 2 26 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=6.645
+ $Y=1.84 $X2=6.785 $Y2=2.225
r96 1 28 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.41
+ $Y=0.81 $X2=6.555 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%C 1 3 4 5 6 8 12 14 17 21 24 26 27
c86 12 0 1.44369e-19 $X=6.77 $Y=1.35
c87 1 0 1.52403e-19 $X=5.71 $Y=1.085
r88 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=1.515 $X2=7.01 $Y2=1.515
r89 23 26 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=6.77 $Y=1.515
+ $X2=7.01 $Y2=1.515
r90 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.77 $Y=1.515
+ $X2=6.695 $Y2=1.515
r91 21 27 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=7.01 $Y=1.665
+ $X2=7.01 $Y2=1.515
r92 15 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.01 $Y=1.68
+ $X2=7.01 $Y2=1.515
r93 15 17 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=7.01 $Y=1.68
+ $X2=7.01 $Y2=2.16
r94 12 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.35
+ $X2=6.77 $Y2=1.515
r95 12 14 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.77 $Y=1.35 $X2=6.77
+ $Y2=1.02
r96 11 20 3.61756 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.1 $Y=1.425 $X2=6.01
+ $Y2=1.425
r97 11 24 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=6.1 $Y=1.425
+ $X2=6.695 $Y2=1.425
r98 6 20 45.2467 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.01 $Y=1.59
+ $X2=6.01 $Y2=1.425
r99 6 8 320.685 $w=1.8e-07 $l=8.25e-07 $layer=POLY_cond $X=6.01 $Y=1.59 $X2=6.01
+ $Y2=2.415
r100 4 20 82.4064 $w=1.55e-07 $l=2.65e-07 $layer=POLY_cond $X=6.01 $Y=1.16
+ $X2=6.01 $Y2=1.425
r101 4 5 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.16
+ $X2=5.785 $Y2=1.16
r102 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.71 $Y=1.085
+ $X2=5.785 $Y2=1.16
r103 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.71 $Y=1.085
+ $X2=5.71 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_1057_74# 1 2 9 11 13 14 16 18 20 23 25 26
+ 27 30 31 32 34 36 37 38 39 40 44 46 51 53
c125 51 0 1.38659e-19 $X=7.59 $Y=1.505
c126 14 0 1.44369e-19 $X=8.14 $Y=1.605
r127 56 57 4.09864 $w=2.94e-07 $l=2.5e-08 $layer=POLY_cond $X=7.69 $Y=1.505
+ $X2=7.715 $Y2=1.505
r128 52 56 16.3946 $w=2.94e-07 $l=1e-07 $layer=POLY_cond $X=7.59 $Y=1.505
+ $X2=7.69 $Y2=1.505
r129 51 54 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.582 $Y=1.505
+ $X2=7.582 $Y2=1.67
r130 51 53 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.582 $Y=1.505
+ $X2=7.582 $Y2=1.34
r131 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.59
+ $Y=1.505 $X2=7.59 $Y2=1.505
r132 46 48 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.7 $Y=2.82 $X2=5.7
+ $Y2=2.99
r133 44 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.495 $Y=1.95
+ $X2=7.495 $Y2=1.67
r134 41 53 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.495 $Y=1.18
+ $X2=7.495 $Y2=1.34
r135 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=2.035
+ $X2=7.495 $Y2=1.95
r136 39 40 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.41 $Y=2.035
+ $X2=7.21 $Y2=2.035
r137 37 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=1.095
+ $X2=7.495 $Y2=1.18
r138 37 38 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.41 $Y=1.095
+ $X2=7.06 $Y2=1.095
r139 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.125 $Y=2.12
+ $X2=7.21 $Y2=2.035
r140 35 36 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.125 $Y=2.12
+ $X2=7.125 $Y2=2.905
r141 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.975 $Y=1.01
+ $X2=7.06 $Y2=1.095
r142 33 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.975 $Y=0.83
+ $X2=6.975 $Y2=1.01
r143 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.975 $Y2=0.83
r144 31 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.89 $Y=0.745
+ $X2=6.5 $Y2=0.745
r145 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=0.66
+ $X2=6.5 $Y2=0.745
r146 29 30 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.415 $Y=0.425
+ $X2=6.415 $Y2=0.66
r147 28 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=2.99
+ $X2=5.7 $Y2=2.99
r148 27 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.04 $Y=2.99
+ $X2=7.125 $Y2=2.905
r149 27 28 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=7.04 $Y=2.99
+ $X2=5.865 $Y2=2.99
r150 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=6.415 $Y2=0.425
r151 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.33 $Y=0.34
+ $X2=5.66 $Y2=0.34
r152 21 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.66 $Y2=0.34
r153 21 23 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=5.495 $Y=0.425
+ $X2=5.495 $Y2=0.495
r154 18 59 18.4939 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.145 $Y=1.34
+ $X2=8.145 $Y2=1.505
r155 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.145 $Y=1.34
+ $X2=8.145 $Y2=0.86
r156 14 59 0.819728 $w=2.94e-07 $l=5e-09 $layer=POLY_cond $X=8.14 $Y=1.505
+ $X2=8.145 $Y2=1.505
r157 14 57 69.6769 $w=2.94e-07 $l=4.25e-07 $layer=POLY_cond $X=8.14 $Y=1.505
+ $X2=7.715 $Y2=1.505
r158 14 16 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=8.14 $Y=1.605
+ $X2=8.14 $Y2=2.4
r159 11 57 18.4939 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.715 $Y=1.34
+ $X2=7.715 $Y2=1.505
r160 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.715 $Y=1.34
+ $X2=7.715 $Y2=0.86
r161 7 56 14.2527 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.69 $Y=1.67
+ $X2=7.69 $Y2=1.505
r162 7 9 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=7.69 $Y=1.67 $X2=7.69
+ $Y2=2.4
r163 2 46 600 $w=1.7e-07 $l=9.26283e-07 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=1.995 $X2=5.7 $Y2=2.82
r164 1 23 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.495 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_27_373# 1 2 3 4 15 19 20 21 23 24 27 30 33
+ 36 40 41 44 47
c103 47 0 1.46469e-19 $X=1.68 $Y=1.295
c104 40 0 3.06279e-20 $X=1.535 $Y=1.295
c105 36 0 1.9829e-20 $X=2.275 $Y=1.11
c106 33 0 1.91609e-19 $X=0.28 $Y=2.375
c107 27 0 1.97037e-19 $X=2.44 $Y=2.01
c108 19 0 9.32687e-21 $X=1.63 $Y=1.38
r109 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.295
r110 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.295
r111 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.295
+ $X2=0.24 $Y2=1.295
r112 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.535 $Y=1.295
+ $X2=1.68 $Y2=1.295
r113 40 41 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=1.535 $Y=1.295
+ $X2=0.385 $Y2=1.295
r114 36 38 7.46783 $w=2.48e-07 $l=1.62e-07 $layer=LI1_cond $X=2.26 $Y=1.11
+ $X2=2.26 $Y2=1.272
r115 34 44 47.7784 $w=2.38e-07 $l=9.95e-07 $layer=LI1_cond $X=0.205 $Y=2.29
+ $X2=0.205 $Y2=1.295
r116 33 34 4.00454 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.375
+ $X2=0.265 $Y2=2.29
r117 30 44 11.0442 $w=2.38e-07 $l=2.3e-07 $layer=LI1_cond $X=0.205 $Y=1.065
+ $X2=0.205 $Y2=1.295
r118 25 27 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=2.44 $Y=2.565
+ $X2=2.44 $Y2=2.01
r119 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=2.65
+ $X2=2.44 $Y2=2.565
r120 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.275 $Y=2.65
+ $X2=1.715 $Y2=2.65
r121 22 48 3.05574 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=1.272
+ $X2=1.63 $Y2=1.272
r122 21 38 1.64524 $w=2.15e-07 $l=1.25e-07 $layer=LI1_cond $X=2.135 $Y=1.272
+ $X2=2.26 $Y2=1.272
r123 21 22 22.5128 $w=2.13e-07 $l=4.2e-07 $layer=LI1_cond $X=2.135 $Y=1.272
+ $X2=1.715 $Y2=1.272
r124 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.63 $Y=2.565
+ $X2=1.715 $Y2=2.65
r125 19 48 3.88258 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.63 $Y=1.38
+ $X2=1.63 $Y2=1.272
r126 19 20 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=1.63 $Y=1.38
+ $X2=1.63 $Y2=2.565
r127 13 30 6.50835 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.245 $Y=0.905
+ $X2=0.245 $Y2=1.065
r128 13 15 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=0.245 $Y=0.905
+ $X2=0.245 $Y2=0.55
r129 4 27 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.285
+ $Y=1.865 $X2=2.44 $Y2=2.01
r130 3 33 300 $w=1.7e-07 $l=5.77971e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.865 $X2=0.28 $Y2=2.375
r131 2 36 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.845 $X2=2.275 $Y2=1.11
r132 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.175
+ $Y=0.405 $X2=0.32 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%VPWR 1 2 3 4 17 21 25 27 29 33 35 43 48 54
+ 57 60 64
c84 2 0 3.71954e-20 $X=4.405 $Y=1.84
r85 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r86 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r87 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 52 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r90 52 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r91 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r92 49 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.55 $Y=3.33
+ $X2=7.465 $Y2=3.33
r93 49 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.55 $Y=3.33 $X2=7.92
+ $Y2=3.33
r94 48 63 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=8.28 $Y=3.33 $X2=8.46
+ $Y2=3.33
r95 48 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=7.92 $Y2=3.33
r96 47 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r99 44 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=4.62 $Y2=3.33
r100 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 43 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=3.33
+ $X2=7.465 $Y2=3.33
r102 43 46 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=7.38 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 39 42 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 38 41 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 38 39 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 36 54 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.785 $Y2=3.33
r109 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 35 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=3.33
+ $X2=4.62 $Y2=3.33
r111 35 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.455 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 33 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r113 33 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 29 32 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.405 $Y=1.985
+ $X2=8.405 $Y2=2.815
r115 27 63 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.46 $Y2=3.33
r116 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.405 $Y2=2.815
r117 23 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=3.245
+ $X2=7.465 $Y2=3.33
r118 23 25 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.465 $Y=3.245
+ $X2=7.465 $Y2=2.455
r119 19 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=3.245
+ $X2=4.62 $Y2=3.33
r120 19 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.62 $Y=3.245
+ $X2=4.62 $Y2=2.9
r121 15 54 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r122 15 17 29.84 $w=2.78e-07 $l=7.25e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.52
r123 4 32 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.23
+ $Y=1.84 $X2=8.365 $Y2=2.815
r124 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.23
+ $Y=1.84 $X2=8.365 $Y2=1.985
r125 3 25 300 $w=1.7e-07 $l=7.76338e-07 $layer=licon1_PDIFF $count=2 $X=7.1
+ $Y=1.84 $X2=7.465 $Y2=2.455
r126 2 21 600 $w=1.7e-07 $l=1.16254e-06 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=1.84 $X2=4.62 $Y2=2.9
r127 1 17 600 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.865 $X2=0.745 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_335_373# 1 2 3 4 15 17 18 19 20 21 25 31
+ 37 39 40 43 46
c112 43 0 1.94615e-19 $X=2.64 $Y=1.295
c113 40 0 2.00077e-19 $X=2.785 $Y=1.295
c114 17 0 5.80738e-20 $X=2.555 $Y=1.635
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r116 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.295
r117 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.295
+ $X2=2.64 $Y2=1.295
r118 39 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=5.04 $Y2=1.295
r119 39 40 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=2.785 $Y2=1.295
r120 34 37 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=5.04 $Y=2.1 $X2=5.17
+ $Y2=2.1
r121 33 43 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.655 $Y=1.55
+ $X2=2.655 $Y2=1.295
r122 28 43 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=2.655 $Y=1.285
+ $X2=2.655 $Y2=1.295
r123 27 31 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.655 $Y=1.12
+ $X2=2.8 $Y2=1.12
r124 27 28 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=1.12
+ $X2=2.655 $Y2=1.285
r125 23 25 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.995 $Y=1.135
+ $X2=5.995 $Y2=0.81
r126 22 47 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.155 $Y=1.22
+ $X2=5.04 $Y2=1.22
r127 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.83 $Y=1.22
+ $X2=5.995 $Y2=1.135
r128 21 22 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.83 $Y=1.22
+ $X2=5.155 $Y2=1.22
r129 20 34 1.2199 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=1.975
+ $X2=5.04 $Y2=2.1
r130 19 47 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=1.305
+ $X2=5.04 $Y2=1.22
r131 19 20 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.04 $Y=1.305
+ $X2=5.04 $Y2=1.975
r132 17 33 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.555 $Y=1.635
+ $X2=2.655 $Y2=1.55
r133 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.555 $Y=1.635
+ $X2=2.105 $Y2=1.635
r134 13 18 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.995 $Y=1.72
+ $X2=2.105 $Y2=1.635
r135 13 15 20.9535 $w=2.18e-07 $l=4e-07 $layer=LI1_cond $X=1.995 $Y=1.72
+ $X2=1.995 $Y2=2.12
r136 4 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.995 $X2=5.17 $Y2=2.14
r137 3 15 600 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_PDIFF $count=1 $X=1.675
+ $Y=1.865 $X2=1.97 $Y2=2.12
r138 2 25 182 $w=1.7e-07 $l=5.3479e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.37 $X2=5.995 $Y2=0.81
r139 1 31 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.625 $X2=2.8 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%A_329_81# 1 2 3 4 15 19 21 22 23 24 25 29 31
+ 36 37 41
c128 37 0 6.5827e-20 $X=2.725 $Y=0.69
c129 36 0 8.82162e-21 $X=2.555 $Y=0.69
c130 25 0 3.71954e-20 $X=6.07 $Y=2.48
c131 23 0 1.52403e-19 $X=4.67 $Y=0.965
r132 39 40 4.81237 $w=4.69e-07 $l=1.85e-07 $layer=LI1_cond $X=4.872 $Y=0.515
+ $X2=4.872 $Y2=0.7
r133 36 37 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=0.69
+ $X2=2.725 $Y2=0.69
r134 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.79 $Y=0.68
+ $X2=1.79 $Y2=0.8
r135 27 29 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.195 $Y=2.395
+ $X2=6.195 $Y2=2.14
r136 26 41 5.16603 $w=1.7e-07 $l=9.12688e-08 $layer=LI1_cond $X=4.755 $Y=2.48
+ $X2=4.67 $Y2=2.467
r137 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.07 $Y=2.48
+ $X2=6.195 $Y2=2.395
r138 25 26 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=6.07 $Y=2.48
+ $X2=4.755 $Y2=2.48
r139 24 41 1.34256 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=4.67 $Y=2.37
+ $X2=4.67 $Y2=2.467
r140 23 40 12.1197 $w=4.69e-07 $l=3.51788e-07 $layer=LI1_cond $X=4.67 $Y=0.965
+ $X2=4.872 $Y2=0.7
r141 23 24 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=4.67 $Y=0.965
+ $X2=4.67 $Y2=2.37
r142 21 41 5.16603 $w=1.7e-07 $l=9.0802e-08 $layer=LI1_cond $X=4.585 $Y=2.455
+ $X2=4.67 $Y2=2.467
r143 21 22 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.585 $Y=2.455
+ $X2=3.145 $Y2=2.455
r144 17 22 10.2712 $w=1.77e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.99 $Y=2.37
+ $X2=3.145 $Y2=2.455
r145 17 19 12.2679 $w=3.08e-07 $l=3.3e-07 $layer=LI1_cond $X=2.99 $Y=2.37
+ $X2=2.99 $Y2=2.04
r146 15 40 6.75673 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=4.585 $Y=0.7
+ $X2=4.872 $Y2=0.7
r147 15 37 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=4.585 $Y=0.7
+ $X2=2.725 $Y2=0.7
r148 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=1.79 $Y2=0.68
r149 14 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.955 $Y=0.68
+ $X2=2.555 $Y2=0.68
r150 4 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.1
+ $Y=1.995 $X2=6.235 $Y2=2.14
r151 3 19 300 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=2 $X=2.755 $Y=1.865
+ $X2=2.98 $Y2=2.04
r152 2 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.37 $X2=4.995 $Y2=0.515
r153 1 34 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.405 $X2=1.785 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%X 1 2 9 14 15 16 17 28
r34 21 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.93 $Y=1.005 $X2=7.93
+ $Y2=0.925
r35 17 30 8.39233 $w=3.28e-07 $l=1.63e-07 $layer=LI1_cond $X=7.93 $Y=1.007
+ $X2=7.93 $Y2=1.17
r36 17 21 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=7.93 $Y=1.007
+ $X2=7.93 $Y2=1.005
r37 17 28 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=7.93 $Y=0.922
+ $X2=7.93 $Y2=0.925
r38 16 17 12.8166 $w=3.28e-07 $l=3.67e-07 $layer=LI1_cond $X=7.93 $Y=0.555
+ $X2=7.93 $Y2=0.922
r39 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.01 $Y=1.84
+ $X2=8.01 $Y2=1.17
r40 14 15 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=7.922 $Y=2.005
+ $X2=7.922 $Y2=1.84
r41 7 14 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=7.922 $Y=2.012
+ $X2=7.922 $Y2=2.005
r42 7 9 26.8235 $w=3.43e-07 $l=8.03e-07 $layer=LI1_cond $X=7.922 $Y=2.012
+ $X2=7.922 $Y2=2.815
r43 2 14 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.84 $X2=7.915 $Y2=2.005
r44 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.84 $X2=7.915 $Y2=2.815
r45 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.49 $X2=7.93 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_2%VGND 1 2 3 4 15 19 21 23 25 27 29 34 42 48
+ 51 54 62
c82 54 0 1.38659e-19 $X=6.96 $Y=0
r83 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r84 55 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r85 54 59 7.08036 $w=5.6e-07 $l=3.25e-07 $layer=LI1_cond $X=7.242 $Y=0 $X2=7.242
+ $Y2=0.325
r86 54 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r87 54 55 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 52 55 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.96
+ $Y2=0
r89 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r90 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r92 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r93 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r94 43 54 7.87414 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.242
+ $Y2=0
r95 43 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.92
+ $Y2=0
r96 42 61 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=8.457
+ $Y2=0
r97 42 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=7.92
+ $Y2=0
r98 40 41 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r99 38 41 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r100 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r101 37 40 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.08
+ $Y2=0
r102 37 38 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r103 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r104 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r105 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r106 34 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r107 32 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r108 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r109 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r110 29 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r111 27 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r112 27 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r113 23 61 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.457 $Y2=0
r114 23 25 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.4 $Y2=0.635
r115 22 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r116 21 54 7.87414 $w=1.7e-07 $l=3.42e-07 $layer=LI1_cond $X=6.9 $Y=0 $X2=7.242
+ $Y2=0
r117 21 22 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.9 $Y=0 $X2=4.6
+ $Y2=0
r118 17 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r119 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.36
r120 13 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r121 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.78
r122 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.49 $X2=8.36 $Y2=0.635
r123 3 59 60.6667 $w=1.7e-07 $l=7.80705e-07 $layer=licon1_NDIFF $count=3
+ $X=6.845 $Y=0.81 $X2=7.42 $Y2=0.325
r124 2 19 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.445 $X2=4.435 $Y2=0.36
r125 1 15 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.405 $X2=0.75 $Y2=0.78
.ends


* File: sky130_fd_sc_ms__sdfxbp_1.pxi.spice
* Created: Fri Aug 28 18:14:06 2020
* 
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_31_74# N_A_31_74#_M1024_s N_A_31_74#_M1022_s
+ N_A_31_74#_M1007_g N_A_31_74#_M1032_g N_A_31_74#_c_256_n N_A_31_74#_c_257_n
+ N_A_31_74#_c_262_n N_A_31_74#_c_263_n N_A_31_74#_c_258_n N_A_31_74#_c_259_n
+ N_A_31_74#_c_265_n N_A_31_74#_c_266_n PM_SKY130_FD_SC_MS__SDFXBP_1%A_31_74#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%SCE N_SCE_c_343_n N_SCE_c_351_n N_SCE_c_352_n
+ N_SCE_M1024_g N_SCE_c_353_n N_SCE_M1022_g N_SCE_c_354_n N_SCE_c_355_n
+ N_SCE_M1018_g N_SCE_c_345_n N_SCE_M1003_g N_SCE_c_356_n SCE N_SCE_c_346_n
+ N_SCE_c_347_n N_SCE_c_348_n N_SCE_c_349_n PM_SKY130_FD_SC_MS__SDFXBP_1%SCE
x_PM_SKY130_FD_SC_MS__SDFXBP_1%D N_D_M1008_g N_D_M1028_g D N_D_c_423_n
+ N_D_c_424_n PM_SKY130_FD_SC_MS__SDFXBP_1%D
x_PM_SKY130_FD_SC_MS__SDFXBP_1%SCD N_SCD_M1027_g N_SCD_M1009_g SCD SCD
+ N_SCD_c_459_n PM_SKY130_FD_SC_MS__SDFXBP_1%SCD
x_PM_SKY130_FD_SC_MS__SDFXBP_1%CLK N_CLK_c_498_n N_CLK_M1023_g N_CLK_M1013_g CLK
+ N_CLK_c_501_n PM_SKY130_FD_SC_MS__SDFXBP_1%CLK
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_828_74# N_A_828_74#_M1015_d N_A_828_74#_M1025_d
+ N_A_828_74#_M1029_g N_A_828_74#_c_539_n N_A_828_74#_M1006_g
+ N_A_828_74#_M1010_g N_A_828_74#_M1020_g N_A_828_74#_c_561_n
+ N_A_828_74#_c_562_n N_A_828_74#_c_541_n N_A_828_74#_c_542_n
+ N_A_828_74#_c_543_n N_A_828_74#_c_544_n N_A_828_74#_c_545_n
+ N_A_828_74#_c_546_n N_A_828_74#_c_547_n N_A_828_74#_c_548_n
+ N_A_828_74#_c_614_p N_A_828_74#_c_631_p N_A_828_74#_c_549_n
+ N_A_828_74#_c_550_n N_A_828_74#_c_551_n N_A_828_74#_c_552_n
+ N_A_828_74#_c_565_n N_A_828_74#_c_566_n N_A_828_74#_c_553_n
+ N_A_828_74#_c_736_p N_A_828_74#_c_554_n N_A_828_74#_c_555_n
+ N_A_828_74#_c_556_n N_A_828_74#_c_557_n N_A_828_74#_c_558_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%A_828_74#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_612_74# N_A_612_74#_M1023_d N_A_612_74#_M1013_d
+ N_A_612_74#_M1015_g N_A_612_74#_c_738_n N_A_612_74#_c_755_n
+ N_A_612_74#_M1025_g N_A_612_74#_c_739_n N_A_612_74#_M1030_g
+ N_A_612_74#_c_741_n N_A_612_74#_M1033_g N_A_612_74#_M1000_g
+ N_A_612_74#_c_742_n N_A_612_74#_M1017_g N_A_612_74#_c_744_n
+ N_A_612_74#_c_745_n N_A_612_74#_c_746_n N_A_612_74#_c_747_n
+ N_A_612_74#_c_748_n N_A_612_74#_c_749_n N_A_612_74#_c_762_n
+ N_A_612_74#_c_750_n N_A_612_74#_c_751_n N_A_612_74#_c_765_n
+ N_A_612_74#_c_837_p N_A_612_74#_c_898_p N_A_612_74#_c_766_n
+ N_A_612_74#_c_767_n N_A_612_74#_c_768_n N_A_612_74#_c_769_n
+ N_A_612_74#_c_752_n N_A_612_74#_c_771_n N_A_612_74#_c_753_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%A_612_74#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_1243_398# N_A_1243_398#_M1011_d
+ N_A_1243_398#_M1019_d N_A_1243_398#_c_957_n N_A_1243_398#_M1031_g
+ N_A_1243_398#_M1016_g N_A_1243_398#_c_951_n N_A_1243_398#_c_952_n
+ N_A_1243_398#_c_953_n N_A_1243_398#_c_954_n N_A_1243_398#_c_955_n
+ N_A_1243_398#_c_961_n N_A_1243_398#_c_956_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%A_1243_398#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_1021_100# N_A_1021_100#_M1030_d
+ N_A_1021_100#_M1029_d N_A_1021_100#_M1019_g N_A_1021_100#_M1011_g
+ N_A_1021_100#_c_1028_n N_A_1021_100#_c_1029_n N_A_1021_100#_c_1030_n
+ N_A_1021_100#_c_1035_n N_A_1021_100#_c_1036_n N_A_1021_100#_c_1031_n
+ N_A_1021_100#_c_1032_n PM_SKY130_FD_SC_MS__SDFXBP_1%A_1021_100#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_1723_48# N_A_1723_48#_M1001_d
+ N_A_1723_48#_M1014_d N_A_1723_48#_M1021_g N_A_1723_48#_M1002_g
+ N_A_1723_48#_M1012_g N_A_1723_48#_M1005_g N_A_1723_48#_c_1115_n
+ N_A_1723_48#_M1035_g N_A_1723_48#_M1004_g N_A_1723_48#_c_1117_n
+ N_A_1723_48#_c_1118_n N_A_1723_48#_c_1119_n N_A_1723_48#_c_1129_n
+ N_A_1723_48#_c_1130_n N_A_1723_48#_c_1131_n N_A_1723_48#_c_1120_n
+ N_A_1723_48#_c_1132_n N_A_1723_48#_c_1121_n N_A_1723_48#_c_1208_p
+ N_A_1723_48#_c_1122_n N_A_1723_48#_c_1123_n N_A_1723_48#_c_1133_n
+ N_A_1723_48#_c_1134_n N_A_1723_48#_c_1124_n N_A_1723_48#_c_1125_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%A_1723_48#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_1529_74# N_A_1529_74#_M1010_d
+ N_A_1529_74#_M1000_d N_A_1529_74#_c_1251_n N_A_1529_74#_M1001_g
+ N_A_1529_74#_M1014_g N_A_1529_74#_c_1253_n N_A_1529_74#_c_1265_n
+ N_A_1529_74#_c_1266_n N_A_1529_74#_c_1267_n N_A_1529_74#_c_1268_n
+ N_A_1529_74#_c_1254_n N_A_1529_74#_c_1255_n N_A_1529_74#_c_1256_n
+ N_A_1529_74#_c_1257_n N_A_1529_74#_c_1258_n N_A_1529_74#_c_1270_n
+ N_A_1529_74#_c_1259_n N_A_1529_74#_c_1260_n N_A_1529_74#_c_1261_n
+ N_A_1529_74#_c_1262_n PM_SKY130_FD_SC_MS__SDFXBP_1%A_1529_74#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_2216_112# N_A_2216_112#_M1035_s
+ N_A_2216_112#_M1004_s N_A_2216_112#_c_1371_n N_A_2216_112#_M1034_g
+ N_A_2216_112#_c_1373_n N_A_2216_112#_M1026_g N_A_2216_112#_c_1374_n
+ N_A_2216_112#_c_1375_n N_A_2216_112#_c_1376_n N_A_2216_112#_c_1377_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%A_2216_112#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%VPWR N_VPWR_M1022_d N_VPWR_M1009_d N_VPWR_M1025_s
+ N_VPWR_M1031_d N_VPWR_M1002_d N_VPWR_M1005_s N_VPWR_M1004_d N_VPWR_c_1421_n
+ N_VPWR_c_1422_n N_VPWR_c_1423_n N_VPWR_c_1424_n N_VPWR_c_1425_n
+ N_VPWR_c_1426_n VPWR N_VPWR_c_1427_n N_VPWR_c_1428_n N_VPWR_c_1429_n
+ N_VPWR_c_1430_n N_VPWR_c_1431_n N_VPWR_c_1432_n N_VPWR_c_1433_n
+ N_VPWR_c_1420_n N_VPWR_c_1435_n N_VPWR_c_1436_n N_VPWR_c_1437_n
+ N_VPWR_c_1438_n N_VPWR_c_1439_n N_VPWR_c_1440_n N_VPWR_c_1441_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%VPWR
x_PM_SKY130_FD_SC_MS__SDFXBP_1%A_296_74# N_A_296_74#_M1008_d N_A_296_74#_M1030_s
+ N_A_296_74#_M1028_d N_A_296_74#_M1029_s N_A_296_74#_c_1574_n
+ N_A_296_74#_c_1575_n N_A_296_74#_c_1561_n N_A_296_74#_c_1562_n
+ N_A_296_74#_c_1563_n N_A_296_74#_c_1564_n N_A_296_74#_c_1569_n
+ N_A_296_74#_c_1570_n N_A_296_74#_c_1565_n N_A_296_74#_c_1566_n
+ N_A_296_74#_c_1567_n N_A_296_74#_c_1571_n N_A_296_74#_c_1625_n
+ N_A_296_74#_c_1572_n N_A_296_74#_c_1573_n N_A_296_74#_c_1679_n
+ PM_SKY130_FD_SC_MS__SDFXBP_1%A_296_74#
x_PM_SKY130_FD_SC_MS__SDFXBP_1%Q N_Q_M1012_d N_Q_M1005_d N_Q_c_1696_n
+ N_Q_c_1697_n N_Q_c_1693_n Q Q N_Q_c_1694_n Q PM_SKY130_FD_SC_MS__SDFXBP_1%Q
x_PM_SKY130_FD_SC_MS__SDFXBP_1%Q_N N_Q_N_M1026_d N_Q_N_M1034_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_MS__SDFXBP_1%Q_N
x_PM_SKY130_FD_SC_MS__SDFXBP_1%VGND N_VGND_M1024_d N_VGND_M1027_d N_VGND_M1015_s
+ N_VGND_M1016_d N_VGND_M1021_d N_VGND_M1012_s N_VGND_M1035_d N_VGND_c_1742_n
+ N_VGND_c_1743_n N_VGND_c_1744_n N_VGND_c_1745_n N_VGND_c_1746_n
+ N_VGND_c_1747_n N_VGND_c_1748_n N_VGND_c_1749_n N_VGND_c_1750_n
+ N_VGND_c_1751_n VGND N_VGND_c_1752_n N_VGND_c_1753_n N_VGND_c_1754_n
+ N_VGND_c_1755_n N_VGND_c_1756_n N_VGND_c_1757_n N_VGND_c_1758_n
+ N_VGND_c_1759_n N_VGND_c_1760_n N_VGND_c_1761_n N_VGND_c_1762_n
+ N_VGND_c_1763_n N_VGND_c_1764_n PM_SKY130_FD_SC_MS__SDFXBP_1%VGND
cc_1 VNB N_A_31_74#_M1007_g 0.0475288f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_2 VNB N_A_31_74#_c_256_n 0.017734f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.69
cc_3 VNB N_A_31_74#_c_257_n 0.0291841f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.525
cc_4 VNB N_A_31_74#_c_258_n 0.0105846f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.04
cc_5 VNB N_A_31_74#_c_259_n 0.0207058f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.565
cc_6 VNB N_SCE_c_343_n 0.0225543f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.32
cc_7 VNB N_SCE_M1024_g 0.0265269f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.525
cc_8 VNB N_SCE_c_345_n 0.0190492f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.525
cc_9 VNB N_SCE_c_346_n 0.0469821f $X=-0.19 $Y=-0.245 $X2=0.307 $Y2=1.825
cc_10 VNB N_SCE_c_347_n 0.012219f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_11 VNB N_SCE_c_348_n 0.0455055f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_12 VNB N_SCE_c_349_n 0.0162965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_M1008_g 0.0498611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_c_423_n 0.0196781f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.64
cc_15 VNB N_D_c_424_n 0.010039f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.64
cc_16 VNB N_SCD_M1027_g 0.0648667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB SCD 0.00491809f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_18 VNB N_SCD_c_459_n 0.0103114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_CLK_c_498_n 0.0219097f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.37
cc_20 VNB N_CLK_M1013_g 0.00763399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB CLK 0.00802736f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_22 VNB N_CLK_c_501_n 0.0583402f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.125
cc_23 VNB N_A_828_74#_c_539_n 0.0185816f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.125
cc_24 VNB N_A_828_74#_M1010_g 0.0216916f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_25 VNB N_A_828_74#_c_541_n 0.0094817f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.825
cc_26 VNB N_A_828_74#_c_542_n 0.0177202f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.825
cc_27 VNB N_A_828_74#_c_543_n 0.00372992f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_28 VNB N_A_828_74#_c_544_n 0.00584382f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_29 VNB N_A_828_74#_c_545_n 0.0184848f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_30 VNB N_A_828_74#_c_546_n 8.04069e-19 $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=2.04
cc_31 VNB N_A_828_74#_c_547_n 0.00304498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_828_74#_c_548_n 0.0413567f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_33 VNB N_A_828_74#_c_549_n 0.00546206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_828_74#_c_550_n 0.00244258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_828_74#_c_551_n 0.00386929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_828_74#_c_552_n 0.0249814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_828_74#_c_553_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_828_74#_c_554_n 0.00552726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_828_74#_c_555_n 0.0329659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_828_74#_c_556_n 0.00277926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_828_74#_c_557_n 0.00600252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_828_74#_c_558_n 0.00277306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_612_74#_M1015_g 0.029024f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_44 VNB N_A_612_74#_c_738_n 0.00315725f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.125
cc_45 VNB N_A_612_74#_c_739_n 0.0137968f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_46 VNB N_A_612_74#_M1030_g 0.0539353f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=2.465
cc_47 VNB N_A_612_74#_c_741_n 0.0288402f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.04
cc_48 VNB N_A_612_74#_c_742_n 0.0299913f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_49 VNB N_A_612_74#_M1017_g 0.0220815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_612_74#_c_744_n 0.00625466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_612_74#_c_745_n 9.55161e-19 $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_52 VNB N_A_612_74#_c_746_n 0.0249239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_612_74#_c_747_n 0.00836014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_612_74#_c_748_n 0.00735495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_612_74#_c_749_n 2.44598e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_612_74#_c_750_n 0.00362644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_612_74#_c_751_n 0.0311424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_612_74#_c_752_n 0.0024038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_612_74#_c_753_n 0.0109487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1243_398#_c_951_n 0.0204124f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_61 VNB N_A_1243_398#_c_952_n 0.0120695f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.525
cc_62 VNB N_A_1243_398#_c_953_n 0.0301013f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=2.465
cc_63 VNB N_A_1243_398#_c_954_n 0.0057844f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.04
cc_64 VNB N_A_1243_398#_c_955_n 0.00354476f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=2.04
cc_65 VNB N_A_1243_398#_c_956_n 0.021021f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_66 VNB N_A_1021_100#_M1011_g 0.0517822f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.64
cc_67 VNB N_A_1021_100#_c_1028_n 0.0119107f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.525
cc_68 VNB N_A_1021_100#_c_1029_n 0.0104788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1021_100#_c_1030_n 4.61231e-19 $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=2.04
cc_70 VNB N_A_1021_100#_c_1031_n 0.00360348f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.825
cc_71 VNB N_A_1021_100#_c_1032_n 0.0157658f $X=-0.19 $Y=-0.245 $X2=2.005
+ $Y2=2.04
cc_72 VNB N_A_1723_48#_M1021_g 0.024243f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_73 VNB N_A_1723_48#_M1012_g 0.02935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1723_48#_M1005_g 6.2705e-19 $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.565
cc_75 VNB N_A_1723_48#_c_1115_n 0.0643314f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=0.785
cc_76 VNB N_A_1723_48#_M1035_g 0.0241445f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_77 VNB N_A_1723_48#_c_1117_n 0.0258401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1723_48#_c_1118_n 0.00757458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1723_48#_c_1119_n 0.00412679f $X=-0.19 $Y=-0.245 $X2=2.005
+ $Y2=2.125
cc_80 VNB N_A_1723_48#_c_1120_n 0.00818639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1723_48#_c_1121_n 0.00795659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1723_48#_c_1122_n 0.0659302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1723_48#_c_1123_n 0.00861416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1723_48#_c_1124_n 0.00200882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1723_48#_c_1125_n 0.0254762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1529_74#_c_1251_n 0.0237925f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_87 VNB N_A_1529_74#_M1001_g 0.0251373f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=2.125
cc_88 VNB N_A_1529_74#_c_1253_n 0.00487183f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.525
cc_89 VNB N_A_1529_74#_c_1254_n 0.00195667f $X=-0.19 $Y=-0.245 $X2=0.307
+ $Y2=1.825
cc_90 VNB N_A_1529_74#_c_1255_n 0.00592247f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=1.825
cc_91 VNB N_A_1529_74#_c_1256_n 0.00142674f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_92 VNB N_A_1529_74#_c_1257_n 0.00337309f $X=-0.19 $Y=-0.245 $X2=2.005
+ $Y2=1.96
cc_93 VNB N_A_1529_74#_c_1258_n 0.0108965f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_94 VNB N_A_1529_74#_c_1259_n 0.0060862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1529_74#_c_1260_n 0.00558376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1529_74#_c_1261_n 0.0036429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1529_74#_c_1262_n 0.0184072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2216_112#_c_1371_n 0.0404017f $X=-0.19 $Y=-0.245 $X2=1.015
+ $Y2=1.525
cc_99 VNB N_A_2216_112#_M1034_g 0.00121087f $X=-0.19 $Y=-0.245 $X2=1.015
+ $Y2=0.58
cc_100 VNB N_A_2216_112#_c_1373_n 0.0222593f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=2.125
cc_101 VNB N_A_2216_112#_c_1374_n 0.00489156f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=0.785
cc_102 VNB N_A_2216_112#_c_1375_n 0.00116982f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=2.465
cc_103 VNB N_A_2216_112#_c_1376_n 0.00564802f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=0.565
cc_104 VNB N_A_2216_112#_c_1377_n 0.0019836f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=0.785
cc_105 VNB N_VPWR_c_1420_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_296_74#_c_1561_n 0.00692604f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.04
cc_107 VNB N_A_296_74#_c_1562_n 0.014829f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.04
cc_108 VNB N_A_296_74#_c_1563_n 0.0101071f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=0.565
cc_109 VNB N_A_296_74#_c_1564_n 0.00557634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_296_74#_c_1565_n 0.0087055f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_111 VNB N_A_296_74#_c_1566_n 0.00282848f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.69
cc_112 VNB N_A_296_74#_c_1567_n 0.0165556f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_113 VNB N_Q_c_1693_n 0.00420932f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.69
cc_114 VNB N_Q_c_1694_n 0.0108561f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.04
cc_115 VNB Q 0.00597177f $X=-0.19 $Y=-0.245 $X2=0.307 $Y2=1.825
cc_116 VNB Q_N 0.0231264f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.525
cc_117 VNB Q_N 0.0297888f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.58
cc_118 VNB Q_N 0.00654121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1742_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.565
cc_120 VNB N_VGND_c_1743_n 0.00963905f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.825
cc_121 VNB N_VGND_c_1744_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.825
cc_122 VNB N_VGND_c_1745_n 0.0129085f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.96
cc_123 VNB N_VGND_c_1746_n 0.00805174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1747_n 0.00923537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1748_n 0.0100148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1749_n 0.0134514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1750_n 0.02053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1751_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1752_n 0.0193973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1753_n 0.0455426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1754_n 0.0604741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1755_n 0.0507575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1756_n 0.0327701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1757_n 0.0190734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1758_n 0.676852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1759_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1760_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1761_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1762_n 0.00477982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1763_n 0.0125082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1764_n 0.00721303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VPB N_A_31_74#_M1032_g 0.0252813f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.64
cc_143 VPB N_A_31_74#_c_256_n 0.0224496f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.69
cc_144 VPB N_A_31_74#_c_262_n 0.0516091f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=2.465
cc_145 VPB N_A_31_74#_c_263_n 0.0184786f $X=-0.19 $Y=1.66 $X2=1.84 $Y2=2.04
cc_146 VPB N_A_31_74#_c_258_n 0.011997f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=2.04
cc_147 VPB N_A_31_74#_c_265_n 0.00569549f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_148 VPB N_A_31_74#_c_266_n 0.0334061f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_149 VPB N_SCE_c_343_n 0.0258351f $X=-0.19 $Y=1.66 $X2=0.22 $Y2=2.32
cc_150 VPB N_SCE_c_351_n 0.0111993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_SCE_c_352_n 0.0109496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_SCE_c_353_n 0.0216639f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_153 VPB N_SCE_c_354_n 0.0211699f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.64
cc_154 VPB N_SCE_c_355_n 0.0166279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_SCE_c_356_n 0.00835417f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=2.465
cc_156 VPB N_D_M1028_g 0.0442399f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.525
cc_157 VPB N_D_c_423_n 0.01299f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.64
cc_158 VPB N_D_c_424_n 0.00661974f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.64
cc_159 VPB N_SCD_M1009_g 0.0364329f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.525
cc_160 VPB SCD 0.00661602f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_161 VPB N_SCD_c_459_n 0.0283616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_CLK_M1013_g 0.027468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_828_74#_M1029_g 0.026324f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_164 VPB N_A_828_74#_M1020_g 0.0351661f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=2.465
cc_165 VPB N_A_828_74#_c_561_n 0.0181357f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=0.565
cc_166 VPB N_A_828_74#_c_562_n 0.0124151f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.565
cc_167 VPB N_A_828_74#_c_544_n 0.00143191f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_168 VPB N_A_828_74#_c_552_n 0.00590666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_828_74#_c_565_n 0.0090294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_828_74#_c_566_n 0.04579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_612_74#_c_738_n 0.00660767f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.125
cc_172 VPB N_A_612_74#_c_755_n 0.0250167f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.64
cc_173 VPB N_A_612_74#_c_739_n 0.0125862f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.785
cc_174 VPB N_A_612_74#_c_741_n 0.0201567f $X=-0.19 $Y=1.66 $X2=1.84 $Y2=2.04
cc_175 VPB N_A_612_74#_M1033_g 0.0281141f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.825
cc_176 VPB N_A_612_74#_M1000_g 0.0274469f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.69
cc_177 VPB N_A_612_74#_c_744_n 0.00171929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_612_74#_c_745_n 0.00391153f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_179 VPB N_A_612_74#_c_762_n 0.00931465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_612_74#_c_750_n 0.00136812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_612_74#_c_751_n 0.0168177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_612_74#_c_765_n 0.00525319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_612_74#_c_766_n 0.00236132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_612_74#_c_767_n 0.00707711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_612_74#_c_768_n 0.0205433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_612_74#_c_769_n 0.00444883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_612_74#_c_752_n 7.45923e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_612_74#_c_771_n 0.0159687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_612_74#_c_753_n 0.0392559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1243_398#_c_957_n 0.00626859f $X=-0.19 $Y=1.66 $X2=1.015
+ $Y2=1.525
cc_191 VPB N_A_1243_398#_M1031_g 0.0379789f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_192 VPB N_A_1243_398#_c_951_n 0.017271f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.785
cc_193 VPB N_A_1243_398#_c_955_n 0.00505656f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=2.04
cc_194 VPB N_A_1243_398#_c_961_n 0.00368866f $X=-0.19 $Y=1.66 $X2=0.275
+ $Y2=0.785
cc_195 VPB N_A_1021_100#_M1019_g 0.0305906f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_196 VPB N_A_1021_100#_c_1029_n 0.0151397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1021_100#_c_1035_n 0.00693779f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.565
cc_198 VPB N_A_1021_100#_c_1036_n 0.00863148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1021_100#_c_1031_n 0.00231038f $X=-0.19 $Y=1.66 $X2=0.17
+ $Y2=1.825
cc_200 VPB N_A_1021_100#_c_1032_n 0.0335023f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.04
cc_201 VPB N_A_1723_48#_M1002_g 0.0237989f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.64
cc_202 VPB N_A_1723_48#_M1005_g 0.030246f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=0.565
cc_203 VPB N_A_1723_48#_c_1119_n 0.00771603f $X=-0.19 $Y=1.66 $X2=2.005
+ $Y2=2.125
cc_204 VPB N_A_1723_48#_c_1129_n 0.0300599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_1723_48#_c_1130_n 0.0096416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1723_48#_c_1131_n 0.0311613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1723_48#_c_1132_n 0.00866405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1723_48#_c_1133_n 0.00999349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1723_48#_c_1134_n 0.0056542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_1723_48#_c_1125_n 0.0218285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1529_74#_M1014_g 0.0282133f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.69
cc_212 VPB N_A_1529_74#_c_1253_n 0.0135229f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.525
cc_213 VPB N_A_1529_74#_c_1265_n 0.00150872f $X=-0.19 $Y=1.66 $X2=0.365
+ $Y2=2.465
cc_214 VPB N_A_1529_74#_c_1266_n 0.00532231f $X=-0.19 $Y=1.66 $X2=1.84 $Y2=2.04
cc_215 VPB N_A_1529_74#_c_1267_n 0.0146779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1529_74#_c_1268_n 0.00242604f $X=-0.19 $Y=1.66 $X2=0.275
+ $Y2=0.785
cc_217 VPB N_A_1529_74#_c_1257_n 0.00128942f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_218 VPB N_A_1529_74#_c_1270_n 0.00321341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1529_74#_c_1261_n 0.0021202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_2216_112#_M1034_g 0.0299798f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_221 VPB N_A_2216_112#_c_1375_n 0.0183807f $X=-0.19 $Y=1.66 $X2=0.365
+ $Y2=2.465
cc_222 VPB N_VPWR_c_1421_n 0.00882483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1422_n 0.0128171f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.825
cc_224 VPB N_VPWR_c_1423_n 0.00987081f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_225 VPB N_VPWR_c_1424_n 0.00896846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1425_n 0.0185934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1426_n 0.0118539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1427_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1428_n 0.0214483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1429_n 0.0587582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1430_n 0.0592077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1431_n 0.019175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1432_n 0.0308335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1433_n 0.0189924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1420_n 0.152801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1435_n 0.0270726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1436_n 0.0167508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1437_n 0.00949386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1438_n 0.00631473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1439_n 0.0107437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1440_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1441_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_296_74#_c_1564_n 0.00374783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_296_74#_c_1569_n 0.00913235f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=0.785
cc_245 VPB N_A_296_74#_c_1570_n 8.26431e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.825
cc_246 VPB N_A_296_74#_c_1571_n 0.00881812f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.04
cc_247 VPB N_A_296_74#_c_1572_n 0.00658645f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.96
cc_248 VPB N_A_296_74#_c_1573_n 0.00471059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_Q_c_1696_n 0.00368089f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.525
cc_250 VPB N_Q_c_1697_n 0.0124404f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_251 VPB N_Q_c_1693_n 0.00291074f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.69
cc_252 VPB Q_N 0.0076353f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=0.58
cc_253 VPB Q_N 0.0503937f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=2.125
cc_254 N_A_31_74#_M1007_g N_SCE_c_343_n 0.00334293f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_255 N_A_31_74#_c_256_n N_SCE_c_343_n 0.0181178f $X=0.94 $Y=1.69 $X2=0 $Y2=0
cc_256 N_A_31_74#_c_257_n N_SCE_c_343_n 0.00903502f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_257 N_A_31_74#_c_262_n N_SCE_c_343_n 0.00996929f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A_31_74#_c_258_n N_SCE_c_343_n 0.0184949f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_259 N_A_31_74#_c_262_n N_SCE_c_351_n 0.00937675f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A_31_74#_c_262_n N_SCE_c_352_n 0.00835712f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_31_74#_M1007_g N_SCE_M1024_g 0.016521f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_262 N_A_31_74#_c_257_n N_SCE_M1024_g 0.00402581f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_263 N_A_31_74#_c_259_n N_SCE_M1024_g 0.00646213f $X=0.3 $Y=0.565 $X2=0 $Y2=0
cc_264 N_A_31_74#_c_262_n N_SCE_c_353_n 0.0110534f $X=0.365 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_31_74#_c_263_n N_SCE_c_354_n 0.0118599f $X=1.84 $Y=2.04 $X2=0 $Y2=0
cc_266 N_A_31_74#_c_258_n N_SCE_c_354_n 0.00424629f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_267 N_A_31_74#_c_262_n N_SCE_c_355_n 4.29959e-19 $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A_31_74#_c_256_n N_SCE_c_356_n 0.0283381f $X=0.94 $Y=1.69 $X2=0 $Y2=0
cc_269 N_A_31_74#_c_262_n N_SCE_c_356_n 0.00718422f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_31_74#_c_258_n N_SCE_c_356_n 0.00107844f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_271 N_A_31_74#_M1007_g N_SCE_c_346_n 0.0213603f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_272 N_A_31_74#_c_256_n N_SCE_c_346_n 0.00775549f $X=0.94 $Y=1.69 $X2=0 $Y2=0
cc_273 N_A_31_74#_c_257_n N_SCE_c_346_n 0.0109392f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_274 N_A_31_74#_c_258_n N_SCE_c_346_n 0.00778098f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_275 N_A_31_74#_c_259_n N_SCE_c_346_n 0.00484549f $X=0.3 $Y=0.565 $X2=0 $Y2=0
cc_276 N_A_31_74#_c_265_n N_SCE_c_347_n 0.00750655f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_277 N_A_31_74#_c_266_n N_SCE_c_347_n 9.67531e-19 $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_278 N_A_31_74#_c_265_n N_SCE_c_348_n 9.91346e-19 $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_279 N_A_31_74#_c_266_n N_SCE_c_348_n 0.00544003f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_280 N_A_31_74#_M1007_g N_SCE_c_349_n 0.0212279f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_281 N_A_31_74#_c_256_n N_SCE_c_349_n 0.00211101f $X=0.94 $Y=1.69 $X2=0 $Y2=0
cc_282 N_A_31_74#_c_257_n N_SCE_c_349_n 0.0256546f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_283 N_A_31_74#_c_263_n N_SCE_c_349_n 0.0110929f $X=1.84 $Y=2.04 $X2=0 $Y2=0
cc_284 N_A_31_74#_c_258_n N_SCE_c_349_n 0.0306909f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_285 N_A_31_74#_c_259_n N_SCE_c_349_n 0.00241486f $X=0.3 $Y=0.565 $X2=0 $Y2=0
cc_286 N_A_31_74#_M1007_g N_D_M1008_g 0.065468f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_287 N_A_31_74#_M1032_g N_D_M1028_g 0.0172361f $X=1.96 $Y=2.64 $X2=0 $Y2=0
cc_288 N_A_31_74#_c_256_n N_D_M1028_g 0.00305222f $X=0.94 $Y=1.69 $X2=0 $Y2=0
cc_289 N_A_31_74#_c_263_n N_D_M1028_g 0.0176642f $X=1.84 $Y=2.04 $X2=0 $Y2=0
cc_290 N_A_31_74#_c_258_n N_D_M1028_g 0.00277385f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_291 N_A_31_74#_c_265_n N_D_M1028_g 0.00116992f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_292 N_A_31_74#_c_266_n N_D_M1028_g 0.0183745f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_293 N_A_31_74#_M1007_g N_D_c_423_n 0.0214162f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_294 N_A_31_74#_c_263_n N_D_c_423_n 0.00371768f $X=1.84 $Y=2.04 $X2=0 $Y2=0
cc_295 N_A_31_74#_M1007_g N_D_c_424_n 0.00369933f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_296 N_A_31_74#_c_256_n N_D_c_424_n 0.00622556f $X=0.94 $Y=1.69 $X2=0 $Y2=0
cc_297 N_A_31_74#_c_263_n N_D_c_424_n 0.0411529f $X=1.84 $Y=2.04 $X2=0 $Y2=0
cc_298 N_A_31_74#_c_258_n N_D_c_424_n 0.0215615f $X=0.915 $Y=2.04 $X2=0 $Y2=0
cc_299 N_A_31_74#_M1032_g N_SCD_M1009_g 0.0338144f $X=1.96 $Y=2.64 $X2=0 $Y2=0
cc_300 N_A_31_74#_c_265_n N_SCD_M1009_g 2.24581e-19 $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_301 N_A_31_74#_c_266_n N_SCD_M1009_g 0.00975924f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_302 N_A_31_74#_M1032_g SCD 5.07602e-19 $X=1.96 $Y=2.64 $X2=0 $Y2=0
cc_303 N_A_31_74#_c_265_n SCD 0.0217661f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_304 N_A_31_74#_c_266_n SCD 0.00163634f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_305 N_A_31_74#_c_265_n N_SCD_c_459_n 5.05021e-19 $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_306 N_A_31_74#_c_266_n N_SCD_c_459_n 0.00883639f $X=2.005 $Y=1.96 $X2=0 $Y2=0
cc_307 N_A_31_74#_c_256_n N_VPWR_c_1421_n 9.27053e-19 $X=0.94 $Y=1.69 $X2=0
+ $Y2=0
cc_308 N_A_31_74#_c_262_n N_VPWR_c_1421_n 0.0282903f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_31_74#_c_263_n N_VPWR_c_1421_n 0.00880343f $X=1.84 $Y=2.04 $X2=0
+ $Y2=0
cc_310 N_A_31_74#_c_258_n N_VPWR_c_1421_n 0.0146916f $X=0.915 $Y=2.04 $X2=0
+ $Y2=0
cc_311 N_A_31_74#_M1032_g N_VPWR_c_1427_n 0.005209f $X=1.96 $Y=2.64 $X2=0 $Y2=0
cc_312 N_A_31_74#_M1032_g N_VPWR_c_1420_n 0.00517535f $X=1.96 $Y=2.64 $X2=0
+ $Y2=0
cc_313 N_A_31_74#_c_262_n N_VPWR_c_1420_n 0.0162216f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_31_74#_c_262_n N_VPWR_c_1435_n 0.0196804f $X=0.365 $Y=2.465 $X2=0
+ $Y2=0
cc_315 N_A_31_74#_M1032_g N_VPWR_c_1436_n 0.00128339f $X=1.96 $Y=2.64 $X2=0
+ $Y2=0
cc_316 N_A_31_74#_M1007_g N_A_296_74#_c_1574_n 6.99132e-19 $X=1.015 $Y=0.58
+ $X2=0 $Y2=0
cc_317 N_A_31_74#_M1032_g N_A_296_74#_c_1575_n 0.0105358f $X=1.96 $Y=2.64 $X2=0
+ $Y2=0
cc_318 N_A_31_74#_c_265_n N_A_296_74#_c_1575_n 0.0122883f $X=2.005 $Y=1.96 $X2=0
+ $Y2=0
cc_319 N_A_31_74#_c_266_n N_A_296_74#_c_1575_n 6.08607e-19 $X=2.005 $Y=1.96
+ $X2=0 $Y2=0
cc_320 N_A_31_74#_M1032_g N_A_296_74#_c_1573_n 0.0121629f $X=1.96 $Y=2.64 $X2=0
+ $Y2=0
cc_321 N_A_31_74#_c_263_n N_A_296_74#_c_1573_n 0.0220899f $X=1.84 $Y=2.04 $X2=0
+ $Y2=0
cc_322 N_A_31_74#_c_265_n N_A_296_74#_c_1573_n 0.00475538f $X=2.005 $Y=1.96
+ $X2=0 $Y2=0
cc_323 N_A_31_74#_c_266_n N_A_296_74#_c_1573_n 2.27493e-19 $X=2.005 $Y=1.96
+ $X2=0 $Y2=0
cc_324 N_A_31_74#_M1007_g N_VGND_c_1742_n 0.011043f $X=1.015 $Y=0.58 $X2=0 $Y2=0
cc_325 N_A_31_74#_c_259_n N_VGND_c_1742_n 0.0153602f $X=0.3 $Y=0.565 $X2=0 $Y2=0
cc_326 N_A_31_74#_c_259_n N_VGND_c_1752_n 0.0165046f $X=0.3 $Y=0.565 $X2=0 $Y2=0
cc_327 N_A_31_74#_M1007_g N_VGND_c_1753_n 0.00383152f $X=1.015 $Y=0.58 $X2=0
+ $Y2=0
cc_328 N_A_31_74#_M1007_g N_VGND_c_1758_n 0.0075725f $X=1.015 $Y=0.58 $X2=0
+ $Y2=0
cc_329 N_A_31_74#_c_259_n N_VGND_c_1758_n 0.0137323f $X=0.3 $Y=0.565 $X2=0 $Y2=0
cc_330 N_SCE_c_345_n N_D_M1008_g 0.0144151f $X=2.095 $Y=0.9 $X2=0 $Y2=0
cc_331 N_SCE_c_347_n N_D_M1008_g 0.00429476f $X=1.885 $Y=1.065 $X2=0 $Y2=0
cc_332 N_SCE_c_348_n N_D_M1008_g 0.0178081f $X=2.095 $Y=1.065 $X2=0 $Y2=0
cc_333 N_SCE_c_349_n N_D_M1008_g 0.0205821f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_334 N_SCE_c_354_n N_D_M1028_g 0.0532969f $X=1 $Y=2.17 $X2=0 $Y2=0
cc_335 N_SCE_c_349_n N_D_c_423_n 0.00458551f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_336 N_SCE_c_354_n N_D_c_424_n 4.72616e-19 $X=1 $Y=2.17 $X2=0 $Y2=0
cc_337 N_SCE_c_349_n N_D_c_424_n 0.0434752f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_338 N_SCE_c_345_n N_SCD_M1027_g 0.0474884f $X=2.095 $Y=0.9 $X2=0 $Y2=0
cc_339 N_SCE_c_347_n N_SCD_M1027_g 4.33427e-19 $X=1.885 $Y=1.065 $X2=0 $Y2=0
cc_340 N_SCE_c_353_n N_VPWR_c_1421_n 0.00351947f $X=0.59 $Y=2.245 $X2=0 $Y2=0
cc_341 N_SCE_c_354_n N_VPWR_c_1421_n 0.00323673f $X=1 $Y=2.17 $X2=0 $Y2=0
cc_342 N_SCE_c_355_n N_VPWR_c_1421_n 0.0173409f $X=1.09 $Y=2.245 $X2=0 $Y2=0
cc_343 N_SCE_c_355_n N_VPWR_c_1427_n 0.00460063f $X=1.09 $Y=2.245 $X2=0 $Y2=0
cc_344 N_SCE_c_353_n N_VPWR_c_1420_n 0.00986085f $X=0.59 $Y=2.245 $X2=0 $Y2=0
cc_345 N_SCE_c_355_n N_VPWR_c_1420_n 0.00908371f $X=1.09 $Y=2.245 $X2=0 $Y2=0
cc_346 N_SCE_c_353_n N_VPWR_c_1435_n 0.005209f $X=0.59 $Y=2.245 $X2=0 $Y2=0
cc_347 N_SCE_c_345_n N_A_296_74#_c_1574_n 0.0175259f $X=2.095 $Y=0.9 $X2=0 $Y2=0
cc_348 N_SCE_c_347_n N_A_296_74#_c_1574_n 0.0364171f $X=1.885 $Y=1.065 $X2=0
+ $Y2=0
cc_349 N_SCE_c_348_n N_A_296_74#_c_1574_n 0.00161084f $X=2.095 $Y=1.065 $X2=0
+ $Y2=0
cc_350 N_SCE_c_349_n N_A_296_74#_c_1574_n 0.00408749f $X=1.565 $Y=1.047 $X2=0
+ $Y2=0
cc_351 N_SCE_c_345_n N_A_296_74#_c_1561_n 0.00371748f $X=2.095 $Y=0.9 $X2=0
+ $Y2=0
cc_352 N_SCE_c_347_n N_A_296_74#_c_1561_n 0.0291033f $X=1.885 $Y=1.065 $X2=0
+ $Y2=0
cc_353 N_SCE_c_347_n N_A_296_74#_c_1563_n 0.00951656f $X=1.885 $Y=1.065 $X2=0
+ $Y2=0
cc_354 N_SCE_c_348_n N_A_296_74#_c_1563_n 4.32703e-19 $X=2.095 $Y=1.065 $X2=0
+ $Y2=0
cc_355 N_SCE_c_355_n N_A_296_74#_c_1573_n 0.00192554f $X=1.09 $Y=2.245 $X2=0
+ $Y2=0
cc_356 N_SCE_M1024_g N_VGND_c_1742_n 0.00513692f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_357 N_SCE_c_346_n N_VGND_c_1742_n 0.00208805f $X=0.515 $Y=1.12 $X2=0 $Y2=0
cc_358 N_SCE_c_349_n N_VGND_c_1742_n 0.0201359f $X=1.565 $Y=1.047 $X2=0 $Y2=0
cc_359 N_SCE_M1024_g N_VGND_c_1752_n 0.00434272f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_360 N_SCE_c_345_n N_VGND_c_1753_n 0.00296985f $X=2.095 $Y=0.9 $X2=0 $Y2=0
cc_361 N_SCE_M1024_g N_VGND_c_1758_n 0.00824496f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_362 N_SCE_c_345_n N_VGND_c_1758_n 0.00365767f $X=2.095 $Y=0.9 $X2=0 $Y2=0
cc_363 N_D_M1028_g N_VPWR_c_1421_n 0.00247097f $X=1.51 $Y=2.64 $X2=0 $Y2=0
cc_364 N_D_M1028_g N_VPWR_c_1427_n 0.005209f $X=1.51 $Y=2.64 $X2=0 $Y2=0
cc_365 N_D_M1028_g N_VPWR_c_1420_n 0.00983291f $X=1.51 $Y=2.64 $X2=0 $Y2=0
cc_366 N_D_M1008_g N_A_296_74#_c_1574_n 0.0094734f $X=1.405 $Y=0.58 $X2=0 $Y2=0
cc_367 N_D_M1028_g N_A_296_74#_c_1573_n 0.0137354f $X=1.51 $Y=2.64 $X2=0 $Y2=0
cc_368 N_D_M1008_g N_VGND_c_1742_n 0.00191703f $X=1.405 $Y=0.58 $X2=0 $Y2=0
cc_369 N_D_M1008_g N_VGND_c_1753_n 0.00434051f $X=1.405 $Y=0.58 $X2=0 $Y2=0
cc_370 N_D_M1008_g N_VGND_c_1758_n 0.00820179f $X=1.405 $Y=0.58 $X2=0 $Y2=0
cc_371 N_SCD_M1027_g N_CLK_c_498_n 0.0234726f $X=2.485 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_372 N_SCD_M1009_g N_CLK_M1013_g 0.0208278f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_373 N_SCD_c_459_n N_CLK_M1013_g 0.00777786f $X=2.545 $Y=1.775 $X2=0 $Y2=0
cc_374 N_SCD_M1027_g N_CLK_c_501_n 0.00333958f $X=2.485 $Y=0.58 $X2=0 $Y2=0
cc_375 N_SCD_M1027_g N_A_612_74#_c_747_n 2.01164e-19 $X=2.485 $Y=0.58 $X2=0
+ $Y2=0
cc_376 N_SCD_M1027_g N_A_612_74#_c_749_n 5.27956e-19 $X=2.485 $Y=0.58 $X2=0
+ $Y2=0
cc_377 N_SCD_M1009_g N_VPWR_c_1427_n 0.00461464f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_378 N_SCD_M1009_g N_VPWR_c_1420_n 0.00444149f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_379 N_SCD_M1009_g N_VPWR_c_1436_n 0.0152405f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_380 N_SCD_M1009_g N_A_296_74#_c_1575_n 0.0148905f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_381 SCD N_A_296_74#_c_1575_n 0.0183209f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_382 N_SCD_c_459_n N_A_296_74#_c_1575_n 4.11623e-19 $X=2.545 $Y=1.775 $X2=0
+ $Y2=0
cc_383 N_SCD_M1027_g N_A_296_74#_c_1561_n 0.00749276f $X=2.485 $Y=0.58 $X2=0
+ $Y2=0
cc_384 N_SCD_M1027_g N_A_296_74#_c_1562_n 0.0161008f $X=2.485 $Y=0.58 $X2=0
+ $Y2=0
cc_385 SCD N_A_296_74#_c_1562_n 0.0235982f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_386 N_SCD_c_459_n N_A_296_74#_c_1562_n 9.93453e-19 $X=2.545 $Y=1.775 $X2=0
+ $Y2=0
cc_387 SCD N_A_296_74#_c_1563_n 7.44219e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_388 N_SCD_M1027_g N_A_296_74#_c_1564_n 0.00391514f $X=2.485 $Y=0.58 $X2=0
+ $Y2=0
cc_389 N_SCD_M1009_g N_A_296_74#_c_1564_n 0.00528956f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_390 SCD N_A_296_74#_c_1564_n 0.0473211f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_391 N_SCD_c_459_n N_A_296_74#_c_1564_n 0.00111877f $X=2.545 $Y=1.775 $X2=0
+ $Y2=0
cc_392 N_SCD_M1009_g N_A_296_74#_c_1573_n 0.00196654f $X=2.5 $Y=2.64 $X2=0 $Y2=0
cc_393 N_SCD_M1027_g N_VGND_c_1743_n 0.00374169f $X=2.485 $Y=0.58 $X2=0 $Y2=0
cc_394 N_SCD_M1027_g N_VGND_c_1753_n 0.00461464f $X=2.485 $Y=0.58 $X2=0 $Y2=0
cc_395 N_SCD_M1027_g N_VGND_c_1758_n 0.00908754f $X=2.485 $Y=0.58 $X2=0 $Y2=0
cc_396 CLK N_A_612_74#_M1015_g 6.03388e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_397 N_CLK_c_501_n N_A_612_74#_M1015_g 0.00328824f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_398 N_CLK_c_498_n N_A_612_74#_c_747_n 0.00629682f $X=2.985 $Y=1.22 $X2=0
+ $Y2=0
cc_399 CLK N_A_612_74#_c_748_n 0.0254704f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_400 N_CLK_c_501_n N_A_612_74#_c_748_n 0.00126098f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_401 N_CLK_c_498_n N_A_612_74#_c_749_n 0.00367545f $X=2.985 $Y=1.22 $X2=0
+ $Y2=0
cc_402 CLK N_A_612_74#_c_749_n 0.0113738f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_403 N_CLK_c_501_n N_A_612_74#_c_749_n 0.00714913f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_404 CLK N_A_612_74#_c_762_n 0.00493081f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_405 N_CLK_M1013_g N_A_612_74#_c_750_n 0.00260591f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_406 CLK N_A_612_74#_c_750_n 0.0292932f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_407 N_CLK_c_501_n N_A_612_74#_c_750_n 5.13557e-19 $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_408 N_CLK_M1013_g N_A_612_74#_c_751_n 0.00604224f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_409 CLK N_A_612_74#_c_751_n 0.00137967f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_410 N_CLK_c_501_n N_A_612_74#_c_751_n 0.0125058f $X=3.21 $Y=1.385 $X2=0 $Y2=0
cc_411 N_CLK_M1013_g N_A_612_74#_c_767_n 0.00634099f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_412 CLK N_A_612_74#_c_767_n 0.0189212f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_413 N_CLK_c_501_n N_A_612_74#_c_767_n 0.00571027f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_414 N_CLK_M1013_g N_VPWR_c_1422_n 0.0097956f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_415 N_CLK_M1013_g N_VPWR_c_1428_n 0.00461464f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_416 N_CLK_M1013_g N_VPWR_c_1420_n 0.0044838f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_417 N_CLK_M1013_g N_VPWR_c_1436_n 0.0244121f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_418 N_CLK_c_498_n N_A_296_74#_c_1562_n 0.00847112f $X=2.985 $Y=1.22 $X2=0
+ $Y2=0
cc_419 CLK N_A_296_74#_c_1562_n 0.0142131f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_420 N_CLK_c_501_n N_A_296_74#_c_1562_n 0.00570301f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_421 CLK N_A_296_74#_c_1564_n 0.0152822f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_422 N_CLK_c_501_n N_A_296_74#_c_1564_n 0.0178458f $X=3.21 $Y=1.385 $X2=0
+ $Y2=0
cc_423 N_CLK_M1013_g N_A_296_74#_c_1569_n 0.0206842f $X=3.21 $Y=2.4 $X2=0 $Y2=0
cc_424 N_CLK_c_498_n N_VGND_c_1743_n 0.00336369f $X=2.985 $Y=1.22 $X2=0 $Y2=0
cc_425 N_CLK_c_498_n N_VGND_c_1744_n 0.00434272f $X=2.985 $Y=1.22 $X2=0 $Y2=0
cc_426 N_CLK_c_498_n N_VGND_c_1745_n 0.00334742f $X=2.985 $Y=1.22 $X2=0 $Y2=0
cc_427 N_CLK_c_498_n N_VGND_c_1758_n 0.00825771f $X=2.985 $Y=1.22 $X2=0 $Y2=0
cc_428 N_A_828_74#_c_541_n N_A_612_74#_M1015_g 0.0015901f $X=4.28 $Y=0.515 $X2=0
+ $Y2=0
cc_429 N_A_828_74#_c_543_n N_A_612_74#_M1015_g 0.00285142f $X=4.445 $Y=0.34
+ $X2=0 $Y2=0
cc_430 N_A_828_74#_c_541_n N_A_612_74#_c_738_n 0.00125047f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_431 N_A_828_74#_c_544_n N_A_612_74#_c_755_n 0.00156666f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_432 N_A_828_74#_c_565_n N_A_612_74#_c_755_n 7.43073e-19 $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_433 N_A_828_74#_c_566_n N_A_612_74#_c_755_n 0.00575971f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_434 N_A_828_74#_c_565_n N_A_612_74#_c_739_n 0.012686f $X=5.075 $Y=2.155 $X2=0
+ $Y2=0
cc_435 N_A_828_74#_c_566_n N_A_612_74#_c_739_n 0.0180964f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_436 N_A_828_74#_c_539_n N_A_612_74#_M1030_g 0.0134026f $X=5.71 $Y=1.03 $X2=0
+ $Y2=0
cc_437 N_A_828_74#_c_541_n N_A_612_74#_M1030_g 0.00322663f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_438 N_A_828_74#_c_542_n N_A_612_74#_M1030_g 0.00881128f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_439 N_A_828_74#_c_544_n N_A_612_74#_M1030_g 0.0301317f $X=5.155 $Y=1.82 $X2=0
+ $Y2=0
cc_440 N_A_828_74#_c_553_n N_A_612_74#_M1030_g 0.00175971f $X=5.155 $Y=0.34
+ $X2=0 $Y2=0
cc_441 N_A_828_74#_c_544_n N_A_612_74#_c_741_n 0.00848553f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_442 N_A_828_74#_c_547_n N_A_612_74#_c_741_n 2.76302e-19 $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_443 N_A_828_74#_c_548_n N_A_612_74#_c_741_n 0.0205027f $X=5.87 $Y=1.195 $X2=0
+ $Y2=0
cc_444 N_A_828_74#_c_566_n N_A_612_74#_c_741_n 0.00800603f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_445 N_A_828_74#_c_566_n N_A_612_74#_M1033_g 0.0204226f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_446 N_A_828_74#_c_562_n N_A_612_74#_M1000_g 0.0205705f $X=8.395 $Y=2.17 $X2=0
+ $Y2=0
cc_447 N_A_828_74#_c_552_n N_A_612_74#_c_742_n 0.0142778f $X=8.515 $Y=1.52 $X2=0
+ $Y2=0
cc_448 N_A_828_74#_c_554_n N_A_612_74#_c_742_n 0.00241447f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_449 N_A_828_74#_c_557_n N_A_612_74#_c_742_n 0.00614465f $X=8.05 $Y=1.43 $X2=0
+ $Y2=0
cc_450 N_A_828_74#_c_558_n N_A_612_74#_c_742_n 0.018169f $X=8.22 $Y=1.43 $X2=0
+ $Y2=0
cc_451 N_A_828_74#_M1010_g N_A_612_74#_M1017_g 0.00627384f $X=7.57 $Y=0.645
+ $X2=0 $Y2=0
cc_452 N_A_828_74#_c_549_n N_A_612_74#_M1017_g 0.00242411f $X=7.69 $Y=0.34 $X2=0
+ $Y2=0
cc_453 N_A_828_74#_c_556_n N_A_612_74#_M1017_g 0.00187705f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_454 N_A_828_74#_c_544_n N_A_612_74#_c_745_n 0.00594022f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_455 N_A_828_74#_M1010_g N_A_612_74#_c_746_n 0.00350773f $X=7.57 $Y=0.645
+ $X2=0 $Y2=0
cc_456 N_A_828_74#_c_551_n N_A_612_74#_c_746_n 0.00364871f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_457 N_A_828_74#_c_552_n N_A_612_74#_c_746_n 0.00332459f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_458 N_A_828_74#_c_555_n N_A_612_74#_c_746_n 0.0204749f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_459 N_A_828_74#_c_556_n N_A_612_74#_c_746_n 0.00225834f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_460 N_A_828_74#_c_558_n N_A_612_74#_c_746_n 0.00192158f $X=8.22 $Y=1.43 $X2=0
+ $Y2=0
cc_461 N_A_828_74#_c_541_n N_A_612_74#_c_750_n 0.0047909f $X=4.28 $Y=0.515 $X2=0
+ $Y2=0
cc_462 N_A_828_74#_c_566_n N_A_612_74#_c_768_n 0.00403509f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_463 N_A_828_74#_c_552_n N_A_612_74#_c_752_n 6.00238e-19 $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_464 N_A_828_74#_c_554_n N_A_612_74#_c_752_n 0.0203505f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_465 N_A_828_74#_c_555_n N_A_612_74#_c_752_n 2.67686e-19 $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_466 N_A_828_74#_c_557_n N_A_612_74#_c_752_n 0.00122353f $X=8.05 $Y=1.43 $X2=0
+ $Y2=0
cc_467 N_A_828_74#_c_566_n N_A_612_74#_c_771_n 0.00186306f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_468 N_A_828_74#_c_561_n N_A_612_74#_c_753_n 0.0198311f $X=8.395 $Y=2.02 $X2=0
+ $Y2=0
cc_469 N_A_828_74#_c_554_n N_A_612_74#_c_753_n 9.50416e-19 $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_470 N_A_828_74#_c_555_n N_A_612_74#_c_753_n 0.0146077f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_471 N_A_828_74#_c_557_n N_A_612_74#_c_753_n 0.00415645f $X=8.05 $Y=1.43 $X2=0
+ $Y2=0
cc_472 N_A_828_74#_c_549_n N_A_1243_398#_M1011_d 0.00181776f $X=7.69 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_473 N_A_828_74#_c_547_n N_A_1243_398#_c_952_n 0.0218583f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_474 N_A_828_74#_c_548_n N_A_1243_398#_c_952_n 0.00118201f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_475 N_A_828_74#_c_614_p N_A_1243_398#_c_952_n 0.0571895f $X=6.85 $Y=0.775
+ $X2=0 $Y2=0
cc_476 N_A_828_74#_c_549_n N_A_1243_398#_c_952_n 0.00392224f $X=7.69 $Y=0.34
+ $X2=0 $Y2=0
cc_477 N_A_828_74#_c_547_n N_A_1243_398#_c_953_n 4.15062e-19 $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_478 N_A_828_74#_c_548_n N_A_1243_398#_c_953_n 0.0210735f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_479 N_A_828_74#_c_614_p N_A_1243_398#_c_953_n 0.00391065f $X=6.85 $Y=0.775
+ $X2=0 $Y2=0
cc_480 N_A_828_74#_M1010_g N_A_1243_398#_c_954_n 0.00649287f $X=7.57 $Y=0.645
+ $X2=0 $Y2=0
cc_481 N_A_828_74#_c_549_n N_A_1243_398#_c_954_n 0.0157317f $X=7.69 $Y=0.34
+ $X2=0 $Y2=0
cc_482 N_A_828_74#_c_554_n N_A_1243_398#_c_954_n 0.0227674f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_483 N_A_828_74#_c_555_n N_A_1243_398#_c_954_n 0.00207368f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_484 N_A_828_74#_c_556_n N_A_1243_398#_c_954_n 0.00837092f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_485 N_A_828_74#_c_554_n N_A_1243_398#_c_955_n 0.00447131f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_486 N_A_828_74#_c_555_n N_A_1243_398#_c_955_n 3.97462e-19 $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_487 N_A_828_74#_c_539_n N_A_1243_398#_c_956_n 0.0135f $X=5.71 $Y=1.03 $X2=0
+ $Y2=0
cc_488 N_A_828_74#_c_545_n N_A_1243_398#_c_956_n 5.92548e-19 $X=5.75 $Y=0.34
+ $X2=0 $Y2=0
cc_489 N_A_828_74#_c_546_n N_A_1243_398#_c_956_n 0.00487885f $X=5.892 $Y=0.69
+ $X2=0 $Y2=0
cc_490 N_A_828_74#_c_547_n N_A_1243_398#_c_956_n 0.00396563f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_491 N_A_828_74#_c_614_p N_A_1243_398#_c_956_n 0.0138367f $X=6.85 $Y=0.775
+ $X2=0 $Y2=0
cc_492 N_A_828_74#_c_631_p N_A_1243_398#_c_956_n 0.00300612f $X=6.935 $Y=0.69
+ $X2=0 $Y2=0
cc_493 N_A_828_74#_c_544_n N_A_1021_100#_M1030_d 0.0042575f $X=5.155 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_494 N_A_828_74#_M1010_g N_A_1021_100#_M1011_g 0.0192422f $X=7.57 $Y=0.645
+ $X2=0 $Y2=0
cc_495 N_A_828_74#_c_549_n N_A_1021_100#_M1011_g 0.0118543f $X=7.69 $Y=0.34
+ $X2=0 $Y2=0
cc_496 N_A_828_74#_c_554_n N_A_1021_100#_M1011_g 2.8582e-19 $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_497 N_A_828_74#_c_555_n N_A_1021_100#_M1011_g 0.0171166f $X=7.615 $Y=1.255
+ $X2=0 $Y2=0
cc_498 N_A_828_74#_c_539_n N_A_1021_100#_c_1028_n 0.00496513f $X=5.71 $Y=1.03
+ $X2=0 $Y2=0
cc_499 N_A_828_74#_c_544_n N_A_1021_100#_c_1028_n 0.0694974f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_500 N_A_828_74#_c_545_n N_A_1021_100#_c_1028_n 0.012971f $X=5.75 $Y=0.34
+ $X2=0 $Y2=0
cc_501 N_A_828_74#_c_547_n N_A_1021_100#_c_1028_n 0.0347882f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_502 N_A_828_74#_c_547_n N_A_1021_100#_c_1029_n 0.0226162f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_503 N_A_828_74#_c_548_n N_A_1021_100#_c_1029_n 0.00346436f $X=5.87 $Y=1.195
+ $X2=0 $Y2=0
cc_504 N_A_828_74#_c_614_p N_A_1021_100#_c_1029_n 0.00499811f $X=6.85 $Y=0.775
+ $X2=0 $Y2=0
cc_505 N_A_828_74#_c_544_n N_A_1021_100#_c_1030_n 0.0135293f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_506 N_A_828_74#_M1029_g N_A_1021_100#_c_1035_n 0.00766532f $X=5.375 $Y=2.69
+ $X2=0 $Y2=0
cc_507 N_A_828_74#_M1029_g N_A_1021_100#_c_1036_n 0.00682306f $X=5.375 $Y=2.69
+ $X2=0 $Y2=0
cc_508 N_A_828_74#_c_544_n N_A_1021_100#_c_1036_n 0.00858845f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_509 N_A_828_74#_c_565_n N_A_1021_100#_c_1036_n 0.0369554f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_510 N_A_828_74#_c_566_n N_A_1021_100#_c_1036_n 0.00634432f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_511 N_A_828_74#_c_552_n N_A_1723_48#_c_1117_n 0.00410296f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_512 N_A_828_74#_M1020_g N_A_1723_48#_c_1130_n 6.77067e-19 $X=8.38 $Y=2.75
+ $X2=0 $Y2=0
cc_513 N_A_828_74#_M1020_g N_A_1723_48#_c_1131_n 0.0490179f $X=8.38 $Y=2.75
+ $X2=0 $Y2=0
cc_514 N_A_828_74#_c_562_n N_A_1723_48#_c_1131_n 0.00782003f $X=8.395 $Y=2.17
+ $X2=0 $Y2=0
cc_515 N_A_828_74#_c_561_n N_A_1723_48#_c_1125_n 0.0107684f $X=8.395 $Y=2.02
+ $X2=0 $Y2=0
cc_516 N_A_828_74#_c_551_n N_A_1723_48#_c_1125_n 2.93187e-19 $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_517 N_A_828_74#_c_552_n N_A_1723_48#_c_1125_n 0.0211504f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_518 N_A_828_74#_c_558_n N_A_1723_48#_c_1125_n 5.55836e-19 $X=8.22 $Y=1.43
+ $X2=0 $Y2=0
cc_519 N_A_828_74#_c_549_n N_A_1529_74#_M1010_d 6.28082e-19 $X=7.69 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_520 N_A_828_74#_c_556_n N_A_1529_74#_M1010_d 0.00812725f $X=7.695 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_521 N_A_828_74#_M1020_g N_A_1529_74#_c_1265_n 0.00674514f $X=8.38 $Y=2.75
+ $X2=0 $Y2=0
cc_522 N_A_828_74#_c_558_n N_A_1529_74#_c_1265_n 5.21567e-19 $X=8.22 $Y=1.43
+ $X2=0 $Y2=0
cc_523 N_A_828_74#_c_561_n N_A_1529_74#_c_1267_n 0.0155886f $X=8.395 $Y=2.02
+ $X2=0 $Y2=0
cc_524 N_A_828_74#_c_562_n N_A_1529_74#_c_1267_n 0.00277699f $X=8.395 $Y=2.17
+ $X2=0 $Y2=0
cc_525 N_A_828_74#_c_551_n N_A_1529_74#_c_1267_n 0.0326559f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_526 N_A_828_74#_c_552_n N_A_1529_74#_c_1267_n 0.00441003f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_527 N_A_828_74#_c_558_n N_A_1529_74#_c_1268_n 0.0144087f $X=8.22 $Y=1.43
+ $X2=0 $Y2=0
cc_528 N_A_828_74#_c_556_n N_A_1529_74#_c_1254_n 0.00498303f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_529 N_A_828_74#_c_551_n N_A_1529_74#_c_1255_n 0.0076531f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_530 N_A_828_74#_c_552_n N_A_1529_74#_c_1255_n 0.00154759f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_531 N_A_828_74#_c_551_n N_A_1529_74#_c_1256_n 0.011566f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_532 N_A_828_74#_c_552_n N_A_1529_74#_c_1256_n 0.00392698f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_533 N_A_828_74#_c_556_n N_A_1529_74#_c_1256_n 0.00577893f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_534 N_A_828_74#_c_561_n N_A_1529_74#_c_1257_n 0.00164707f $X=8.395 $Y=2.02
+ $X2=0 $Y2=0
cc_535 N_A_828_74#_c_551_n N_A_1529_74#_c_1257_n 0.0201267f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_536 N_A_828_74#_c_552_n N_A_1529_74#_c_1257_n 0.00229136f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_537 N_A_828_74#_c_561_n N_A_1529_74#_c_1270_n 0.00163108f $X=8.395 $Y=2.02
+ $X2=0 $Y2=0
cc_538 N_A_828_74#_c_562_n N_A_1529_74#_c_1270_n 0.00674514f $X=8.395 $Y=2.17
+ $X2=0 $Y2=0
cc_539 N_A_828_74#_M1010_g N_A_1529_74#_c_1259_n 9.38568e-19 $X=7.57 $Y=0.645
+ $X2=0 $Y2=0
cc_540 N_A_828_74#_c_549_n N_A_1529_74#_c_1259_n 0.00661633f $X=7.69 $Y=0.34
+ $X2=0 $Y2=0
cc_541 N_A_828_74#_c_551_n N_A_1529_74#_c_1259_n 0.00560127f $X=8.515 $Y=1.52
+ $X2=0 $Y2=0
cc_542 N_A_828_74#_c_556_n N_A_1529_74#_c_1259_n 0.0306116f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_543 N_A_828_74#_c_557_n N_A_1529_74#_c_1259_n 0.00790998f $X=8.05 $Y=1.43
+ $X2=0 $Y2=0
cc_544 N_A_828_74#_c_558_n N_A_1529_74#_c_1260_n 0.00332311f $X=8.22 $Y=1.43
+ $X2=0 $Y2=0
cc_545 N_A_828_74#_M1020_g N_VPWR_c_1424_n 0.00150721f $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_546 N_A_828_74#_M1029_g N_VPWR_c_1429_n 0.0058807f $X=5.375 $Y=2.69 $X2=0
+ $Y2=0
cc_547 N_A_828_74#_M1020_g N_VPWR_c_1430_n 0.00553757f $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_548 N_A_828_74#_M1029_g N_VPWR_c_1420_n 0.00632145f $X=5.375 $Y=2.69 $X2=0
+ $Y2=0
cc_549 N_A_828_74#_M1020_g N_VPWR_c_1420_n 0.0109043f $X=8.38 $Y=2.75 $X2=0
+ $Y2=0
cc_550 N_A_828_74#_c_565_n N_A_296_74#_c_1570_n 0.0161616f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_551 N_A_828_74#_c_566_n N_A_296_74#_c_1570_n 4.3257e-19 $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_552 N_A_828_74#_c_541_n N_A_296_74#_c_1565_n 0.00401715f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_553 N_A_828_74#_c_544_n N_A_296_74#_c_1565_n 0.0134973f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_554 N_A_828_74#_c_565_n N_A_296_74#_c_1565_n 0.0302216f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_555 N_A_828_74#_c_541_n N_A_296_74#_c_1566_n 0.00956695f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_556 N_A_828_74#_c_541_n N_A_296_74#_c_1567_n 0.0374588f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_557 N_A_828_74#_c_542_n N_A_296_74#_c_1567_n 0.0192119f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_558 N_A_828_74#_c_544_n N_A_296_74#_c_1567_n 0.0522531f $X=5.155 $Y=1.82
+ $X2=0 $Y2=0
cc_559 N_A_828_74#_M1025_d N_A_296_74#_c_1571_n 0.00298843f $X=4.485 $Y=1.84
+ $X2=0 $Y2=0
cc_560 N_A_828_74#_M1029_g N_A_296_74#_c_1571_n 7.79654e-19 $X=5.375 $Y=2.69
+ $X2=0 $Y2=0
cc_561 N_A_828_74#_c_565_n N_A_296_74#_c_1571_n 0.0406937f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_562 N_A_828_74#_c_566_n N_A_296_74#_c_1571_n 0.00774417f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_563 N_A_828_74#_M1025_d N_A_296_74#_c_1625_n 0.00538932f $X=4.485 $Y=1.84
+ $X2=0 $Y2=0
cc_564 N_A_828_74#_M1029_g N_A_296_74#_c_1625_n 0.00185506f $X=5.375 $Y=2.69
+ $X2=0 $Y2=0
cc_565 N_A_828_74#_c_565_n N_A_296_74#_c_1625_n 0.0106796f $X=5.075 $Y=2.155
+ $X2=0 $Y2=0
cc_566 N_A_828_74#_M1029_g N_A_296_74#_c_1572_n 7.62635e-19 $X=5.375 $Y=2.69
+ $X2=0 $Y2=0
cc_567 N_A_828_74#_c_614_p N_VGND_M1016_d 0.0149445f $X=6.85 $Y=0.775 $X2=0
+ $Y2=0
cc_568 N_A_828_74#_c_631_p N_VGND_M1016_d 0.00437919f $X=6.935 $Y=0.69 $X2=0
+ $Y2=0
cc_569 N_A_828_74#_c_550_n N_VGND_M1016_d 6.25492e-19 $X=7.02 $Y=0.34 $X2=0
+ $Y2=0
cc_570 N_A_828_74#_c_543_n N_VGND_c_1745_n 0.00749385f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_571 N_A_828_74#_c_545_n N_VGND_c_1746_n 0.00820472f $X=5.75 $Y=0.34 $X2=0
+ $Y2=0
cc_572 N_A_828_74#_c_546_n N_VGND_c_1746_n 0.00373972f $X=5.892 $Y=0.69 $X2=0
+ $Y2=0
cc_573 N_A_828_74#_c_614_p N_VGND_c_1746_n 0.017591f $X=6.85 $Y=0.775 $X2=0
+ $Y2=0
cc_574 N_A_828_74#_c_631_p N_VGND_c_1746_n 0.00706899f $X=6.935 $Y=0.69 $X2=0
+ $Y2=0
cc_575 N_A_828_74#_c_550_n N_VGND_c_1746_n 0.0144033f $X=7.02 $Y=0.34 $X2=0
+ $Y2=0
cc_576 N_A_828_74#_c_539_n N_VGND_c_1754_n 7.26171e-19 $X=5.71 $Y=1.03 $X2=0
+ $Y2=0
cc_577 N_A_828_74#_c_542_n N_VGND_c_1754_n 0.0402032f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_578 N_A_828_74#_c_543_n N_VGND_c_1754_n 0.0179217f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_579 N_A_828_74#_c_545_n N_VGND_c_1754_n 0.0532258f $X=5.75 $Y=0.34 $X2=0
+ $Y2=0
cc_580 N_A_828_74#_c_614_p N_VGND_c_1754_n 0.00530242f $X=6.85 $Y=0.775 $X2=0
+ $Y2=0
cc_581 N_A_828_74#_c_553_n N_VGND_c_1754_n 0.0121867f $X=5.155 $Y=0.34 $X2=0
+ $Y2=0
cc_582 N_A_828_74#_M1010_g N_VGND_c_1755_n 0.00278271f $X=7.57 $Y=0.645 $X2=0
+ $Y2=0
cc_583 N_A_828_74#_c_614_p N_VGND_c_1755_n 0.00262318f $X=6.85 $Y=0.775 $X2=0
+ $Y2=0
cc_584 N_A_828_74#_c_549_n N_VGND_c_1755_n 0.0544154f $X=7.69 $Y=0.34 $X2=0
+ $Y2=0
cc_585 N_A_828_74#_c_550_n N_VGND_c_1755_n 0.0120795f $X=7.02 $Y=0.34 $X2=0
+ $Y2=0
cc_586 N_A_828_74#_M1010_g N_VGND_c_1758_n 0.00355988f $X=7.57 $Y=0.645 $X2=0
+ $Y2=0
cc_587 N_A_828_74#_c_542_n N_VGND_c_1758_n 0.0234906f $X=5.07 $Y=0.34 $X2=0
+ $Y2=0
cc_588 N_A_828_74#_c_543_n N_VGND_c_1758_n 0.00971942f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_589 N_A_828_74#_c_545_n N_VGND_c_1758_n 0.030247f $X=5.75 $Y=0.34 $X2=0 $Y2=0
cc_590 N_A_828_74#_c_614_p N_VGND_c_1758_n 0.0163792f $X=6.85 $Y=0.775 $X2=0
+ $Y2=0
cc_591 N_A_828_74#_c_549_n N_VGND_c_1758_n 0.0304265f $X=7.69 $Y=0.34 $X2=0
+ $Y2=0
cc_592 N_A_828_74#_c_550_n N_VGND_c_1758_n 0.00658903f $X=7.02 $Y=0.34 $X2=0
+ $Y2=0
cc_593 N_A_828_74#_c_553_n N_VGND_c_1758_n 0.00660921f $X=5.155 $Y=0.34 $X2=0
+ $Y2=0
cc_594 N_A_828_74#_c_546_n A_1157_100# 0.00311414f $X=5.892 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_595 N_A_828_74#_c_547_n A_1157_100# 7.49468e-19 $X=5.87 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_596 N_A_828_74#_c_614_p A_1157_100# 0.00627545f $X=6.85 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_597 N_A_828_74#_c_736_p A_1157_100# 6.19923e-19 $X=5.892 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_598 N_A_612_74#_c_837_p N_A_1243_398#_M1019_d 0.025286f $X=7.565 $Y=2.605
+ $X2=0 $Y2=0
cc_599 N_A_612_74#_c_766_n N_A_1243_398#_M1019_d 0.0076998f $X=7.65 $Y=2.52
+ $X2=0 $Y2=0
cc_600 N_A_612_74#_c_768_n N_A_1243_398#_c_957_n 0.00621485f $X=5.84 $Y=2.035
+ $X2=0 $Y2=0
cc_601 N_A_612_74#_c_769_n N_A_1243_398#_c_957_n 0.00522333f $X=6.02 $Y=2.035
+ $X2=0 $Y2=0
cc_602 N_A_612_74#_M1033_g N_A_1243_398#_M1031_g 0.0314542f $X=5.825 $Y=2.69
+ $X2=0 $Y2=0
cc_603 N_A_612_74#_c_765_n N_A_1243_398#_M1031_g 0.00723747f $X=6.02 $Y=2.52
+ $X2=0 $Y2=0
cc_604 N_A_612_74#_c_837_p N_A_1243_398#_M1031_g 0.0190237f $X=7.565 $Y=2.605
+ $X2=0 $Y2=0
cc_605 N_A_612_74#_c_771_n N_A_1243_398#_M1031_g 0.00621485f $X=5.84 $Y=2.2
+ $X2=0 $Y2=0
cc_606 N_A_612_74#_c_741_n N_A_1243_398#_c_951_n 0.0213111f $X=5.675 $Y=1.675
+ $X2=0 $Y2=0
cc_607 N_A_612_74#_c_769_n N_A_1243_398#_c_951_n 0.00211554f $X=6.02 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_A_612_74#_c_742_n N_A_1243_398#_c_955_n 0.00445728f $X=8.065 $Y=1.63
+ $X2=0 $Y2=0
cc_609 N_A_612_74#_c_752_n N_A_1243_398#_c_955_n 0.0306852f $X=7.72 $Y=1.795
+ $X2=0 $Y2=0
cc_610 N_A_612_74#_c_753_n N_A_1243_398#_c_955_n 0.00251818f $X=7.845 $Y=1.795
+ $X2=0 $Y2=0
cc_611 N_A_612_74#_c_837_p N_A_1243_398#_c_961_n 0.0262176f $X=7.565 $Y=2.605
+ $X2=0 $Y2=0
cc_612 N_A_612_74#_c_766_n N_A_1243_398#_c_961_n 0.0194278f $X=7.65 $Y=2.52
+ $X2=0 $Y2=0
cc_613 N_A_612_74#_c_837_p N_A_1021_100#_M1019_g 0.0180279f $X=7.565 $Y=2.605
+ $X2=0 $Y2=0
cc_614 N_A_612_74#_c_766_n N_A_1021_100#_M1019_g 0.00320946f $X=7.65 $Y=2.52
+ $X2=0 $Y2=0
cc_615 N_A_612_74#_c_753_n N_A_1021_100#_M1019_g 4.29905e-19 $X=7.845 $Y=1.795
+ $X2=0 $Y2=0
cc_616 N_A_612_74#_M1030_g N_A_1021_100#_c_1028_n 0.00296701f $X=5.03 $Y=0.71
+ $X2=0 $Y2=0
cc_617 N_A_612_74#_c_741_n N_A_1021_100#_c_1029_n 0.017901f $X=5.675 $Y=1.675
+ $X2=0 $Y2=0
cc_618 N_A_612_74#_c_769_n N_A_1021_100#_c_1029_n 0.0261387f $X=6.02 $Y=2.035
+ $X2=0 $Y2=0
cc_619 N_A_612_74#_M1030_g N_A_1021_100#_c_1030_n 4.00949e-19 $X=5.03 $Y=0.71
+ $X2=0 $Y2=0
cc_620 N_A_612_74#_c_741_n N_A_1021_100#_c_1030_n 0.00714571f $X=5.675 $Y=1.675
+ $X2=0 $Y2=0
cc_621 N_A_612_74#_M1033_g N_A_1021_100#_c_1035_n 0.00921183f $X=5.825 $Y=2.69
+ $X2=0 $Y2=0
cc_622 N_A_612_74#_c_765_n N_A_1021_100#_c_1035_n 0.00299148f $X=6.02 $Y=2.52
+ $X2=0 $Y2=0
cc_623 N_A_612_74#_c_769_n N_A_1021_100#_c_1035_n 7.70348e-19 $X=6.02 $Y=2.035
+ $X2=0 $Y2=0
cc_624 N_A_612_74#_c_771_n N_A_1021_100#_c_1035_n 0.00245428f $X=5.84 $Y=2.2
+ $X2=0 $Y2=0
cc_625 N_A_612_74#_c_741_n N_A_1021_100#_c_1036_n 0.00602573f $X=5.675 $Y=1.675
+ $X2=0 $Y2=0
cc_626 N_A_612_74#_M1033_g N_A_1021_100#_c_1036_n 0.00203067f $X=5.825 $Y=2.69
+ $X2=0 $Y2=0
cc_627 N_A_612_74#_c_765_n N_A_1021_100#_c_1036_n 0.0117006f $X=6.02 $Y=2.52
+ $X2=0 $Y2=0
cc_628 N_A_612_74#_c_768_n N_A_1021_100#_c_1036_n 0.00969365f $X=5.84 $Y=2.035
+ $X2=0 $Y2=0
cc_629 N_A_612_74#_c_769_n N_A_1021_100#_c_1036_n 0.0248707f $X=6.02 $Y=2.035
+ $X2=0 $Y2=0
cc_630 N_A_612_74#_c_837_p N_A_1021_100#_c_1031_n 0.00714622f $X=7.565 $Y=2.605
+ $X2=0 $Y2=0
cc_631 N_A_612_74#_c_769_n N_A_1021_100#_c_1031_n 0.00183977f $X=6.02 $Y=2.035
+ $X2=0 $Y2=0
cc_632 N_A_612_74#_c_837_p N_A_1021_100#_c_1032_n 5.55869e-19 $X=7.565 $Y=2.605
+ $X2=0 $Y2=0
cc_633 N_A_612_74#_c_752_n N_A_1021_100#_c_1032_n 2.99208e-19 $X=7.72 $Y=1.795
+ $X2=0 $Y2=0
cc_634 N_A_612_74#_c_753_n N_A_1021_100#_c_1032_n 0.0100254f $X=7.845 $Y=1.795
+ $X2=0 $Y2=0
cc_635 N_A_612_74#_M1017_g N_A_1723_48#_M1021_g 0.0260838f $X=8.33 $Y=0.58 $X2=0
+ $Y2=0
cc_636 N_A_612_74#_c_742_n N_A_1723_48#_c_1117_n 5.66812e-19 $X=8.065 $Y=1.63
+ $X2=0 $Y2=0
cc_637 N_A_612_74#_c_746_n N_A_1723_48#_c_1117_n 0.0260838f $X=8.33 $Y=1.04
+ $X2=0 $Y2=0
cc_638 N_A_612_74#_M1000_g N_A_1529_74#_c_1265_n 0.00330427f $X=7.845 $Y=2.54
+ $X2=0 $Y2=0
cc_639 N_A_612_74#_c_753_n N_A_1529_74#_c_1265_n 0.00351335f $X=7.845 $Y=1.795
+ $X2=0 $Y2=0
cc_640 N_A_612_74#_M1000_g N_A_1529_74#_c_1266_n 0.019512f $X=7.845 $Y=2.54
+ $X2=0 $Y2=0
cc_641 N_A_612_74#_c_752_n N_A_1529_74#_c_1268_n 0.0134093f $X=7.72 $Y=1.795
+ $X2=0 $Y2=0
cc_642 N_A_612_74#_c_753_n N_A_1529_74#_c_1268_n 0.00418897f $X=7.845 $Y=1.795
+ $X2=0 $Y2=0
cc_643 N_A_612_74#_M1017_g N_A_1529_74#_c_1254_n 0.00387649f $X=8.33 $Y=0.58
+ $X2=0 $Y2=0
cc_644 N_A_612_74#_c_746_n N_A_1529_74#_c_1254_n 3.91054e-19 $X=8.33 $Y=1.04
+ $X2=0 $Y2=0
cc_645 N_A_612_74#_c_742_n N_A_1529_74#_c_1256_n 4.35709e-19 $X=8.065 $Y=1.63
+ $X2=0 $Y2=0
cc_646 N_A_612_74#_c_746_n N_A_1529_74#_c_1256_n 0.00438715f $X=8.33 $Y=1.04
+ $X2=0 $Y2=0
cc_647 N_A_612_74#_c_766_n N_A_1529_74#_c_1270_n 0.00774145f $X=7.65 $Y=2.52
+ $X2=0 $Y2=0
cc_648 N_A_612_74#_c_752_n N_A_1529_74#_c_1270_n 6.67209e-19 $X=7.72 $Y=1.795
+ $X2=0 $Y2=0
cc_649 N_A_612_74#_c_753_n N_A_1529_74#_c_1270_n 0.00159052f $X=7.845 $Y=1.795
+ $X2=0 $Y2=0
cc_650 N_A_612_74#_M1017_g N_A_1529_74#_c_1259_n 0.014391f $X=8.33 $Y=0.58 $X2=0
+ $Y2=0
cc_651 N_A_612_74#_c_746_n N_A_1529_74#_c_1259_n 0.00620238f $X=8.33 $Y=1.04
+ $X2=0 $Y2=0
cc_652 N_A_612_74#_c_762_n N_VPWR_M1025_s 0.00475059f $X=3.855 $Y=1.905 $X2=0
+ $Y2=0
cc_653 N_A_612_74#_c_837_p N_VPWR_M1031_d 0.0146731f $X=7.565 $Y=2.605 $X2=0
+ $Y2=0
cc_654 N_A_612_74#_c_755_n N_VPWR_c_1422_n 0.0211814f $X=4.395 $Y=1.75 $X2=0
+ $Y2=0
cc_655 N_A_612_74#_c_837_p N_VPWR_c_1423_n 0.0248918f $X=7.565 $Y=2.605 $X2=0
+ $Y2=0
cc_656 N_A_612_74#_c_755_n N_VPWR_c_1429_n 0.00460063f $X=4.395 $Y=1.75 $X2=0
+ $Y2=0
cc_657 N_A_612_74#_M1033_g N_VPWR_c_1429_n 0.00612719f $X=5.825 $Y=2.69 $X2=0
+ $Y2=0
cc_658 N_A_612_74#_c_837_p N_VPWR_c_1429_n 0.00488549f $X=7.565 $Y=2.605 $X2=0
+ $Y2=0
cc_659 N_A_612_74#_c_898_p N_VPWR_c_1429_n 0.00282634f $X=6.105 $Y=2.605 $X2=0
+ $Y2=0
cc_660 N_A_612_74#_M1000_g N_VPWR_c_1430_n 0.005209f $X=7.845 $Y=2.54 $X2=0
+ $Y2=0
cc_661 N_A_612_74#_c_837_p N_VPWR_c_1430_n 0.015371f $X=7.565 $Y=2.605 $X2=0
+ $Y2=0
cc_662 N_A_612_74#_c_755_n N_VPWR_c_1420_n 0.00448128f $X=4.395 $Y=1.75 $X2=0
+ $Y2=0
cc_663 N_A_612_74#_M1033_g N_VPWR_c_1420_n 0.00632145f $X=5.825 $Y=2.69 $X2=0
+ $Y2=0
cc_664 N_A_612_74#_M1000_g N_VPWR_c_1420_n 0.00989358f $X=7.845 $Y=2.54 $X2=0
+ $Y2=0
cc_665 N_A_612_74#_c_837_p N_VPWR_c_1420_n 0.0377202f $X=7.565 $Y=2.605 $X2=0
+ $Y2=0
cc_666 N_A_612_74#_c_898_p N_VPWR_c_1420_n 0.00504896f $X=6.105 $Y=2.605 $X2=0
+ $Y2=0
cc_667 N_A_612_74#_c_747_n N_A_296_74#_c_1561_n 7.94987e-19 $X=3.2 $Y=0.515
+ $X2=0 $Y2=0
cc_668 N_A_612_74#_c_749_n N_A_296_74#_c_1561_n 0.0048278f $X=3.365 $Y=0.925
+ $X2=0 $Y2=0
cc_669 N_A_612_74#_c_749_n N_A_296_74#_c_1562_n 0.00230378f $X=3.365 $Y=0.925
+ $X2=0 $Y2=0
cc_670 N_A_612_74#_c_767_n N_A_296_74#_c_1564_n 0.0135476f $X=3.435 $Y=1.905
+ $X2=0 $Y2=0
cc_671 N_A_612_74#_M1013_d N_A_296_74#_c_1569_n 0.00751229f $X=3.3 $Y=1.84 $X2=0
+ $Y2=0
cc_672 N_A_612_74#_c_762_n N_A_296_74#_c_1569_n 0.0179473f $X=3.855 $Y=1.905
+ $X2=0 $Y2=0
cc_673 N_A_612_74#_c_751_n N_A_296_74#_c_1569_n 0.00516338f $X=3.94 $Y=1.515
+ $X2=0 $Y2=0
cc_674 N_A_612_74#_c_767_n N_A_296_74#_c_1569_n 0.0210366f $X=3.435 $Y=1.905
+ $X2=0 $Y2=0
cc_675 N_A_612_74#_c_738_n N_A_296_74#_c_1570_n 0.00499927f $X=4.305 $Y=1.675
+ $X2=0 $Y2=0
cc_676 N_A_612_74#_c_755_n N_A_296_74#_c_1570_n 0.0241827f $X=4.395 $Y=1.75
+ $X2=0 $Y2=0
cc_677 N_A_612_74#_c_744_n N_A_296_74#_c_1570_n 0.00492873f $X=4.395 $Y=1.675
+ $X2=0 $Y2=0
cc_678 N_A_612_74#_c_762_n N_A_296_74#_c_1570_n 0.013382f $X=3.855 $Y=1.905
+ $X2=0 $Y2=0
cc_679 N_A_612_74#_c_750_n N_A_296_74#_c_1570_n 0.0119771f $X=3.94 $Y=1.515
+ $X2=0 $Y2=0
cc_680 N_A_612_74#_c_767_n N_A_296_74#_c_1570_n 0.00732007f $X=3.435 $Y=1.905
+ $X2=0 $Y2=0
cc_681 N_A_612_74#_c_739_n N_A_296_74#_c_1565_n 0.0157813f $X=4.955 $Y=1.675
+ $X2=0 $Y2=0
cc_682 N_A_612_74#_M1030_g N_A_296_74#_c_1565_n 0.00274293f $X=5.03 $Y=0.71
+ $X2=0 $Y2=0
cc_683 N_A_612_74#_c_744_n N_A_296_74#_c_1565_n 0.00779732f $X=4.395 $Y=1.675
+ $X2=0 $Y2=0
cc_684 N_A_612_74#_c_738_n N_A_296_74#_c_1566_n 0.00247513f $X=4.305 $Y=1.675
+ $X2=0 $Y2=0
cc_685 N_A_612_74#_c_744_n N_A_296_74#_c_1566_n 0.00128466f $X=4.395 $Y=1.675
+ $X2=0 $Y2=0
cc_686 N_A_612_74#_c_750_n N_A_296_74#_c_1566_n 0.0135314f $X=3.94 $Y=1.515
+ $X2=0 $Y2=0
cc_687 N_A_612_74#_c_751_n N_A_296_74#_c_1566_n 0.00327963f $X=3.94 $Y=1.515
+ $X2=0 $Y2=0
cc_688 N_A_612_74#_M1015_g N_A_296_74#_c_1567_n 0.00672586f $X=4.065 $Y=0.74
+ $X2=0 $Y2=0
cc_689 N_A_612_74#_M1030_g N_A_296_74#_c_1567_n 0.0124213f $X=5.03 $Y=0.71 $X2=0
+ $Y2=0
cc_690 N_A_612_74#_c_750_n N_A_296_74#_c_1567_n 0.00962885f $X=3.94 $Y=1.515
+ $X2=0 $Y2=0
cc_691 N_A_612_74#_c_755_n N_A_296_74#_c_1625_n 0.0197538f $X=4.395 $Y=1.75
+ $X2=0 $Y2=0
cc_692 N_A_612_74#_c_755_n N_A_296_74#_c_1572_n 0.0057602f $X=4.395 $Y=1.75
+ $X2=0 $Y2=0
cc_693 N_A_612_74#_c_765_n A_1183_496# 5.73081e-19 $X=6.02 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_694 N_A_612_74#_c_837_p A_1183_496# 0.00289478f $X=7.565 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_695 N_A_612_74#_c_898_p A_1183_496# 0.00298884f $X=6.105 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_696 N_A_612_74#_c_748_n N_VGND_M1015_s 0.0104039f $X=3.855 $Y=0.925 $X2=0
+ $Y2=0
cc_697 N_A_612_74#_c_750_n N_VGND_M1015_s 0.0037774f $X=3.94 $Y=1.515 $X2=0
+ $Y2=0
cc_698 N_A_612_74#_c_747_n N_VGND_c_1743_n 0.0180182f $X=3.2 $Y=0.515 $X2=0
+ $Y2=0
cc_699 N_A_612_74#_c_747_n N_VGND_c_1744_n 0.0145323f $X=3.2 $Y=0.515 $X2=0
+ $Y2=0
cc_700 N_A_612_74#_M1015_g N_VGND_c_1745_n 0.00908753f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_701 N_A_612_74#_c_747_n N_VGND_c_1745_n 0.0216229f $X=3.2 $Y=0.515 $X2=0
+ $Y2=0
cc_702 N_A_612_74#_c_748_n N_VGND_c_1745_n 0.0274963f $X=3.855 $Y=0.925 $X2=0
+ $Y2=0
cc_703 N_A_612_74#_c_751_n N_VGND_c_1745_n 3.3849e-19 $X=3.94 $Y=1.515 $X2=0
+ $Y2=0
cc_704 N_A_612_74#_M1017_g N_VGND_c_1747_n 9.27404e-19 $X=8.33 $Y=0.58 $X2=0
+ $Y2=0
cc_705 N_A_612_74#_M1015_g N_VGND_c_1754_n 0.00461464f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_706 N_A_612_74#_M1030_g N_VGND_c_1754_n 7.26171e-19 $X=5.03 $Y=0.71 $X2=0
+ $Y2=0
cc_707 N_A_612_74#_M1017_g N_VGND_c_1755_n 0.00291649f $X=8.33 $Y=0.58 $X2=0
+ $Y2=0
cc_708 N_A_612_74#_M1015_g N_VGND_c_1758_n 0.00814502f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_709 N_A_612_74#_M1017_g N_VGND_c_1758_n 0.00360937f $X=8.33 $Y=0.58 $X2=0
+ $Y2=0
cc_710 N_A_612_74#_c_747_n N_VGND_c_1758_n 0.0119861f $X=3.2 $Y=0.515 $X2=0
+ $Y2=0
cc_711 N_A_612_74#_c_748_n N_VGND_c_1758_n 0.0124019f $X=3.855 $Y=0.925 $X2=0
+ $Y2=0
cc_712 N_A_1243_398#_c_951_n N_A_1021_100#_M1019_g 0.032189f $X=6.305 $Y=1.99
+ $X2=0 $Y2=0
cc_713 N_A_1243_398#_c_955_n N_A_1021_100#_M1019_g 0.00555975f $X=7.275 $Y=2.1
+ $X2=0 $Y2=0
cc_714 N_A_1243_398#_c_961_n N_A_1021_100#_M1019_g 0.00671668f $X=7.275 $Y=2.225
+ $X2=0 $Y2=0
cc_715 N_A_1243_398#_c_951_n N_A_1021_100#_M1011_g 0.00455773f $X=6.305 $Y=1.99
+ $X2=0 $Y2=0
cc_716 N_A_1243_398#_c_952_n N_A_1021_100#_M1011_g 0.0191626f $X=7.19 $Y=1.195
+ $X2=0 $Y2=0
cc_717 N_A_1243_398#_c_953_n N_A_1021_100#_M1011_g 0.00674159f $X=6.41 $Y=1.195
+ $X2=0 $Y2=0
cc_718 N_A_1243_398#_c_954_n N_A_1021_100#_M1011_g 0.0137575f $X=7.275 $Y=1.36
+ $X2=0 $Y2=0
cc_719 N_A_1243_398#_c_955_n N_A_1021_100#_M1011_g 0.0109379f $X=7.275 $Y=2.1
+ $X2=0 $Y2=0
cc_720 N_A_1243_398#_c_956_n N_A_1021_100#_M1011_g 0.00866418f $X=6.41 $Y=1.03
+ $X2=0 $Y2=0
cc_721 N_A_1243_398#_c_953_n N_A_1021_100#_c_1028_n 0.00347455f $X=6.41 $Y=1.195
+ $X2=0 $Y2=0
cc_722 N_A_1243_398#_c_957_n N_A_1021_100#_c_1029_n 0.00109522f $X=6.305 $Y=2.08
+ $X2=0 $Y2=0
cc_723 N_A_1243_398#_c_951_n N_A_1021_100#_c_1029_n 0.0160739f $X=6.305 $Y=1.99
+ $X2=0 $Y2=0
cc_724 N_A_1243_398#_c_952_n N_A_1021_100#_c_1029_n 0.0333579f $X=7.19 $Y=1.195
+ $X2=0 $Y2=0
cc_725 N_A_1243_398#_c_953_n N_A_1021_100#_c_1029_n 0.0040357f $X=6.41 $Y=1.195
+ $X2=0 $Y2=0
cc_726 N_A_1243_398#_M1031_g N_A_1021_100#_c_1035_n 0.0012163f $X=6.305 $Y=2.69
+ $X2=0 $Y2=0
cc_727 N_A_1243_398#_c_951_n N_A_1021_100#_c_1031_n 0.00145248f $X=6.305 $Y=1.99
+ $X2=0 $Y2=0
cc_728 N_A_1243_398#_c_952_n N_A_1021_100#_c_1031_n 0.0278385f $X=7.19 $Y=1.195
+ $X2=0 $Y2=0
cc_729 N_A_1243_398#_c_955_n N_A_1021_100#_c_1031_n 0.0288169f $X=7.275 $Y=2.1
+ $X2=0 $Y2=0
cc_730 N_A_1243_398#_c_961_n N_A_1021_100#_c_1031_n 0.00256538f $X=7.275
+ $Y=2.225 $X2=0 $Y2=0
cc_731 N_A_1243_398#_c_951_n N_A_1021_100#_c_1032_n 0.0147992f $X=6.305 $Y=1.99
+ $X2=0 $Y2=0
cc_732 N_A_1243_398#_c_952_n N_A_1021_100#_c_1032_n 0.00354312f $X=7.19 $Y=1.195
+ $X2=0 $Y2=0
cc_733 N_A_1243_398#_c_955_n N_A_1021_100#_c_1032_n 0.00861106f $X=7.275 $Y=2.1
+ $X2=0 $Y2=0
cc_734 N_A_1243_398#_c_961_n N_A_1021_100#_c_1032_n 0.0073456f $X=7.275 $Y=2.225
+ $X2=0 $Y2=0
cc_735 N_A_1243_398#_M1031_g N_VPWR_c_1423_n 0.00404978f $X=6.305 $Y=2.69 $X2=0
+ $Y2=0
cc_736 N_A_1243_398#_M1031_g N_VPWR_c_1429_n 0.00492183f $X=6.305 $Y=2.69 $X2=0
+ $Y2=0
cc_737 N_A_1243_398#_M1031_g N_VPWR_c_1420_n 0.00632145f $X=6.305 $Y=2.69 $X2=0
+ $Y2=0
cc_738 N_A_1243_398#_c_956_n N_VGND_c_1746_n 0.0021844f $X=6.41 $Y=1.03 $X2=0
+ $Y2=0
cc_739 N_A_1243_398#_c_956_n N_VGND_c_1754_n 0.00378853f $X=6.41 $Y=1.03 $X2=0
+ $Y2=0
cc_740 N_A_1243_398#_c_956_n N_VGND_c_1758_n 0.00505379f $X=6.41 $Y=1.03 $X2=0
+ $Y2=0
cc_741 N_A_1021_100#_M1019_g N_VPWR_c_1423_n 0.00520853f $X=6.925 $Y=2.54 $X2=0
+ $Y2=0
cc_742 N_A_1021_100#_c_1035_n N_VPWR_c_1429_n 0.0122756f $X=5.6 $Y=2.69 $X2=0
+ $Y2=0
cc_743 N_A_1021_100#_M1019_g N_VPWR_c_1430_n 0.00392086f $X=6.925 $Y=2.54 $X2=0
+ $Y2=0
cc_744 N_A_1021_100#_M1019_g N_VPWR_c_1420_n 0.00505743f $X=6.925 $Y=2.54 $X2=0
+ $Y2=0
cc_745 N_A_1021_100#_c_1035_n N_VPWR_c_1420_n 0.0123853f $X=5.6 $Y=2.69 $X2=0
+ $Y2=0
cc_746 N_A_1021_100#_c_1035_n N_A_296_74#_c_1571_n 0.00719893f $X=5.6 $Y=2.69
+ $X2=0 $Y2=0
cc_747 N_A_1021_100#_c_1035_n N_A_296_74#_c_1572_n 0.0114934f $X=5.6 $Y=2.69
+ $X2=0 $Y2=0
cc_748 N_A_1021_100#_M1011_g N_VGND_c_1746_n 0.00121343f $X=7.135 $Y=0.645 $X2=0
+ $Y2=0
cc_749 N_A_1021_100#_M1011_g N_VGND_c_1755_n 0.00278271f $X=7.135 $Y=0.645 $X2=0
+ $Y2=0
cc_750 N_A_1021_100#_M1011_g N_VGND_c_1758_n 0.00358571f $X=7.135 $Y=0.645 $X2=0
+ $Y2=0
cc_751 N_A_1723_48#_c_1122_n N_A_1529_74#_c_1251_n 0.0145987f $X=10.41 $Y=1.485
+ $X2=0 $Y2=0
cc_752 N_A_1723_48#_c_1124_n N_A_1529_74#_c_1251_n 0.00241371f $X=9.865 $Y=1.485
+ $X2=0 $Y2=0
cc_753 N_A_1723_48#_c_1125_n N_A_1529_74#_c_1251_n 0.0169561f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_754 N_A_1723_48#_M1021_g N_A_1529_74#_M1001_g 0.00661561f $X=8.69 $Y=0.58
+ $X2=0 $Y2=0
cc_755 N_A_1723_48#_c_1117_n N_A_1529_74#_M1001_g 0.004134f $X=8.965 $Y=1.07
+ $X2=0 $Y2=0
cc_756 N_A_1723_48#_c_1120_n N_A_1529_74#_M1001_g 0.00391579f $X=9.77 $Y=0.75
+ $X2=0 $Y2=0
cc_757 N_A_1723_48#_c_1121_n N_A_1529_74#_M1001_g 0.00533837f $X=9.865 $Y=1.32
+ $X2=0 $Y2=0
cc_758 N_A_1723_48#_M1002_g N_A_1529_74#_M1014_g 0.0135875f $X=8.8 $Y=2.75 $X2=0
+ $Y2=0
cc_759 N_A_1723_48#_c_1130_n N_A_1529_74#_M1014_g 0.0174492f $X=9.6 $Y=2.235
+ $X2=0 $Y2=0
cc_760 N_A_1723_48#_c_1132_n N_A_1529_74#_M1014_g 0.0171617f $X=9.765 $Y=2.815
+ $X2=0 $Y2=0
cc_761 N_A_1723_48#_c_1133_n N_A_1529_74#_M1014_g 0.00674839f $X=9.765 $Y=2.105
+ $X2=0 $Y2=0
cc_762 N_A_1723_48#_c_1125_n N_A_1529_74#_M1014_g 0.0180446f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_763 N_A_1723_48#_c_1130_n N_A_1529_74#_c_1253_n 8.63567e-19 $X=9.6 $Y=2.235
+ $X2=0 $Y2=0
cc_764 N_A_1723_48#_c_1134_n N_A_1529_74#_c_1253_n 0.00882211f $X=9.775 $Y=1.94
+ $X2=0 $Y2=0
cc_765 N_A_1723_48#_c_1117_n N_A_1529_74#_c_1267_n 8.34571e-19 $X=8.965 $Y=1.07
+ $X2=0 $Y2=0
cc_766 N_A_1723_48#_c_1130_n N_A_1529_74#_c_1267_n 0.0235169f $X=9.6 $Y=2.235
+ $X2=0 $Y2=0
cc_767 N_A_1723_48#_c_1131_n N_A_1529_74#_c_1267_n 0.00518345f $X=8.875 $Y=2.215
+ $X2=0 $Y2=0
cc_768 N_A_1723_48#_c_1133_n N_A_1529_74#_c_1267_n 2.90376e-19 $X=9.765 $Y=2.105
+ $X2=0 $Y2=0
cc_769 N_A_1723_48#_c_1125_n N_A_1529_74#_c_1267_n 0.00941005f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_770 N_A_1723_48#_M1021_g N_A_1529_74#_c_1254_n 0.00387486f $X=8.69 $Y=0.58
+ $X2=0 $Y2=0
cc_771 N_A_1723_48#_M1021_g N_A_1529_74#_c_1255_n 0.00634929f $X=8.69 $Y=0.58
+ $X2=0 $Y2=0
cc_772 N_A_1723_48#_c_1117_n N_A_1529_74#_c_1255_n 0.00917885f $X=8.965 $Y=1.07
+ $X2=0 $Y2=0
cc_773 N_A_1723_48#_c_1125_n N_A_1529_74#_c_1257_n 0.0124128f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_774 N_A_1723_48#_c_1117_n N_A_1529_74#_c_1258_n 8.97248e-19 $X=8.965 $Y=1.07
+ $X2=0 $Y2=0
cc_775 N_A_1723_48#_c_1125_n N_A_1529_74#_c_1258_n 0.00274661f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_776 N_A_1723_48#_c_1130_n N_A_1529_74#_c_1270_n 0.00872496f $X=9.6 $Y=2.235
+ $X2=0 $Y2=0
cc_777 N_A_1723_48#_M1021_g N_A_1529_74#_c_1259_n 0.00162923f $X=8.69 $Y=0.58
+ $X2=0 $Y2=0
cc_778 N_A_1723_48#_c_1117_n N_A_1529_74#_c_1260_n 0.00772788f $X=8.965 $Y=1.07
+ $X2=0 $Y2=0
cc_779 N_A_1723_48#_c_1125_n N_A_1529_74#_c_1260_n 0.00369631f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_780 N_A_1723_48#_c_1130_n N_A_1529_74#_c_1261_n 0.0129935f $X=9.6 $Y=2.235
+ $X2=0 $Y2=0
cc_781 N_A_1723_48#_c_1121_n N_A_1529_74#_c_1261_n 0.0170792f $X=9.865 $Y=1.32
+ $X2=0 $Y2=0
cc_782 N_A_1723_48#_c_1122_n N_A_1529_74#_c_1261_n 3.22361e-19 $X=10.41 $Y=1.485
+ $X2=0 $Y2=0
cc_783 N_A_1723_48#_c_1123_n N_A_1529_74#_c_1261_n 0.00167119f $X=9.77 $Y=0.93
+ $X2=0 $Y2=0
cc_784 N_A_1723_48#_c_1133_n N_A_1529_74#_c_1261_n 6.76444e-19 $X=9.765 $Y=2.105
+ $X2=0 $Y2=0
cc_785 N_A_1723_48#_c_1134_n N_A_1529_74#_c_1261_n 0.00898092f $X=9.775 $Y=1.94
+ $X2=0 $Y2=0
cc_786 N_A_1723_48#_c_1124_n N_A_1529_74#_c_1261_n 0.0277915f $X=9.865 $Y=1.485
+ $X2=0 $Y2=0
cc_787 N_A_1723_48#_c_1125_n N_A_1529_74#_c_1261_n 0.00161269f $X=8.875 $Y=2.05
+ $X2=0 $Y2=0
cc_788 N_A_1723_48#_c_1117_n N_A_1529_74#_c_1262_n 0.0169561f $X=8.965 $Y=1.07
+ $X2=0 $Y2=0
cc_789 N_A_1723_48#_c_1121_n N_A_1529_74#_c_1262_n 0.00508573f $X=9.865 $Y=1.32
+ $X2=0 $Y2=0
cc_790 N_A_1723_48#_c_1123_n N_A_1529_74#_c_1262_n 0.00109024f $X=9.77 $Y=0.93
+ $X2=0 $Y2=0
cc_791 N_A_1723_48#_M1035_g N_A_2216_112#_c_1371_n 0.0214307f $X=11.44 $Y=0.835
+ $X2=0 $Y2=0
cc_792 N_A_1723_48#_c_1118_n N_A_2216_112#_c_1371_n 0.00369421f $X=11.44
+ $Y=1.455 $X2=0 $Y2=0
cc_793 N_A_1723_48#_c_1119_n N_A_2216_112#_M1034_g 0.00369421f $X=11.467 $Y=1.79
+ $X2=0 $Y2=0
cc_794 N_A_1723_48#_c_1129_n N_A_2216_112#_M1034_g 0.0162374f $X=11.467 $Y=1.94
+ $X2=0 $Y2=0
cc_795 N_A_1723_48#_M1035_g N_A_2216_112#_c_1373_n 0.0116936f $X=11.44 $Y=0.835
+ $X2=0 $Y2=0
cc_796 N_A_1723_48#_M1012_g N_A_2216_112#_c_1374_n 8.54002e-19 $X=10.45 $Y=0.74
+ $X2=0 $Y2=0
cc_797 N_A_1723_48#_M1035_g N_A_2216_112#_c_1374_n 0.00786691f $X=11.44 $Y=0.835
+ $X2=0 $Y2=0
cc_798 N_A_1723_48#_c_1115_n N_A_2216_112#_c_1375_n 0.00666886f $X=11.365
+ $Y=1.455 $X2=0 $Y2=0
cc_799 N_A_1723_48#_c_1119_n N_A_2216_112#_c_1375_n 0.0148816f $X=11.467 $Y=1.79
+ $X2=0 $Y2=0
cc_800 N_A_1723_48#_c_1129_n N_A_2216_112#_c_1375_n 0.00642329f $X=11.467
+ $Y=1.94 $X2=0 $Y2=0
cc_801 N_A_1723_48#_c_1115_n N_A_2216_112#_c_1376_n 0.00159431f $X=11.365
+ $Y=1.455 $X2=0 $Y2=0
cc_802 N_A_1723_48#_M1035_g N_A_2216_112#_c_1376_n 0.0105795f $X=11.44 $Y=0.835
+ $X2=0 $Y2=0
cc_803 N_A_1723_48#_c_1118_n N_A_2216_112#_c_1376_n 0.0124075f $X=11.44 $Y=1.455
+ $X2=0 $Y2=0
cc_804 N_A_1723_48#_c_1129_n N_A_2216_112#_c_1376_n 0.00187208f $X=11.467
+ $Y=1.94 $X2=0 $Y2=0
cc_805 N_A_1723_48#_c_1115_n N_A_2216_112#_c_1377_n 0.0133125f $X=11.365
+ $Y=1.455 $X2=0 $Y2=0
cc_806 N_A_1723_48#_c_1130_n N_VPWR_M1002_d 0.00790346f $X=9.6 $Y=2.235 $X2=0
+ $Y2=0
cc_807 N_A_1723_48#_M1002_g N_VPWR_c_1424_n 0.0178964f $X=8.8 $Y=2.75 $X2=0
+ $Y2=0
cc_808 N_A_1723_48#_c_1130_n N_VPWR_c_1424_n 0.0270838f $X=9.6 $Y=2.235 $X2=0
+ $Y2=0
cc_809 N_A_1723_48#_c_1131_n N_VPWR_c_1424_n 0.00365262f $X=8.875 $Y=2.215 $X2=0
+ $Y2=0
cc_810 N_A_1723_48#_c_1132_n N_VPWR_c_1424_n 0.0133529f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_811 N_A_1723_48#_M1005_g N_VPWR_c_1425_n 0.0242874f $X=10.51 $Y=2.4 $X2=0
+ $Y2=0
cc_812 N_A_1723_48#_c_1208_p N_VPWR_c_1425_n 0.0274929f $X=10.41 $Y=1.485 $X2=0
+ $Y2=0
cc_813 N_A_1723_48#_c_1122_n N_VPWR_c_1425_n 0.00712264f $X=10.41 $Y=1.485 $X2=0
+ $Y2=0
cc_814 N_A_1723_48#_c_1134_n N_VPWR_c_1425_n 0.0964204f $X=9.775 $Y=1.94 $X2=0
+ $Y2=0
cc_815 N_A_1723_48#_c_1129_n N_VPWR_c_1426_n 0.0182757f $X=11.467 $Y=1.94 $X2=0
+ $Y2=0
cc_816 N_A_1723_48#_M1002_g N_VPWR_c_1430_n 0.00460063f $X=8.8 $Y=2.75 $X2=0
+ $Y2=0
cc_817 N_A_1723_48#_c_1132_n N_VPWR_c_1431_n 0.0154414f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_818 N_A_1723_48#_M1005_g N_VPWR_c_1432_n 0.00460063f $X=10.51 $Y=2.4 $X2=0
+ $Y2=0
cc_819 N_A_1723_48#_c_1129_n N_VPWR_c_1432_n 0.00502645f $X=11.467 $Y=1.94 $X2=0
+ $Y2=0
cc_820 N_A_1723_48#_M1002_g N_VPWR_c_1420_n 0.00908371f $X=8.8 $Y=2.75 $X2=0
+ $Y2=0
cc_821 N_A_1723_48#_M1005_g N_VPWR_c_1420_n 0.00913687f $X=10.51 $Y=2.4 $X2=0
+ $Y2=0
cc_822 N_A_1723_48#_c_1129_n N_VPWR_c_1420_n 0.00516335f $X=11.467 $Y=1.94 $X2=0
+ $Y2=0
cc_823 N_A_1723_48#_c_1132_n N_VPWR_c_1420_n 0.0127129f $X=9.765 $Y=2.815 $X2=0
+ $Y2=0
cc_824 N_A_1723_48#_M1005_g N_Q_c_1696_n 0.00194411f $X=10.51 $Y=2.4 $X2=0 $Y2=0
cc_825 N_A_1723_48#_c_1115_n N_Q_c_1696_n 0.00224485f $X=11.365 $Y=1.455 $X2=0
+ $Y2=0
cc_826 N_A_1723_48#_c_1129_n N_Q_c_1696_n 0.00312869f $X=11.467 $Y=1.94 $X2=0
+ $Y2=0
cc_827 N_A_1723_48#_M1012_g N_Q_c_1693_n 0.00613182f $X=10.45 $Y=0.74 $X2=0
+ $Y2=0
cc_828 N_A_1723_48#_c_1115_n N_Q_c_1693_n 0.0198946f $X=11.365 $Y=1.455 $X2=0
+ $Y2=0
cc_829 N_A_1723_48#_M1035_g N_Q_c_1693_n 3.80806e-19 $X=11.44 $Y=0.835 $X2=0
+ $Y2=0
cc_830 N_A_1723_48#_c_1208_p N_Q_c_1693_n 0.025206f $X=10.41 $Y=1.485 $X2=0
+ $Y2=0
cc_831 N_A_1723_48#_c_1122_n N_Q_c_1693_n 0.00770035f $X=10.41 $Y=1.485 $X2=0
+ $Y2=0
cc_832 N_A_1723_48#_M1012_g N_Q_c_1694_n 0.00817254f $X=10.45 $Y=0.74 $X2=0
+ $Y2=0
cc_833 N_A_1723_48#_M1035_g N_Q_c_1694_n 0.00300585f $X=11.44 $Y=0.835 $X2=0
+ $Y2=0
cc_834 N_A_1723_48#_M1012_g Q 0.00303502f $X=10.45 $Y=0.74 $X2=0 $Y2=0
cc_835 N_A_1723_48#_c_1115_n Q 0.00589477f $X=11.365 $Y=1.455 $X2=0 $Y2=0
cc_836 N_A_1723_48#_c_1208_p Q 0.0056311f $X=10.41 $Y=1.485 $X2=0 $Y2=0
cc_837 N_A_1723_48#_M1035_g Q_N 2.58792e-19 $X=11.44 $Y=0.835 $X2=0 $Y2=0
cc_838 N_A_1723_48#_c_1129_n Q_N 0.00119087f $X=11.467 $Y=1.94 $X2=0 $Y2=0
cc_839 N_A_1723_48#_M1021_g N_VGND_c_1747_n 0.0111294f $X=8.69 $Y=0.58 $X2=0
+ $Y2=0
cc_840 N_A_1723_48#_c_1117_n N_VGND_c_1747_n 0.00254075f $X=8.965 $Y=1.07 $X2=0
+ $Y2=0
cc_841 N_A_1723_48#_c_1120_n N_VGND_c_1747_n 0.019141f $X=9.77 $Y=0.75 $X2=0
+ $Y2=0
cc_842 N_A_1723_48#_M1012_g N_VGND_c_1748_n 0.00626792f $X=10.45 $Y=0.74 $X2=0
+ $Y2=0
cc_843 N_A_1723_48#_c_1120_n N_VGND_c_1748_n 0.0536441f $X=9.77 $Y=0.75 $X2=0
+ $Y2=0
cc_844 N_A_1723_48#_c_1208_p N_VGND_c_1748_n 0.0130317f $X=10.41 $Y=1.485 $X2=0
+ $Y2=0
cc_845 N_A_1723_48#_c_1122_n N_VGND_c_1748_n 0.00387455f $X=10.41 $Y=1.485 $X2=0
+ $Y2=0
cc_846 N_A_1723_48#_M1035_g N_VGND_c_1749_n 0.0123472f $X=11.44 $Y=0.835 $X2=0
+ $Y2=0
cc_847 N_A_1723_48#_c_1120_n N_VGND_c_1750_n 0.0158774f $X=9.77 $Y=0.75 $X2=0
+ $Y2=0
cc_848 N_A_1723_48#_M1021_g N_VGND_c_1755_n 0.00383152f $X=8.69 $Y=0.58 $X2=0
+ $Y2=0
cc_849 N_A_1723_48#_M1012_g N_VGND_c_1756_n 0.00434272f $X=10.45 $Y=0.74 $X2=0
+ $Y2=0
cc_850 N_A_1723_48#_M1035_g N_VGND_c_1756_n 0.00375057f $X=11.44 $Y=0.835 $X2=0
+ $Y2=0
cc_851 N_A_1723_48#_M1021_g N_VGND_c_1758_n 0.0075694f $X=8.69 $Y=0.58 $X2=0
+ $Y2=0
cc_852 N_A_1723_48#_M1012_g N_VGND_c_1758_n 0.00830282f $X=10.45 $Y=0.74 $X2=0
+ $Y2=0
cc_853 N_A_1723_48#_M1035_g N_VGND_c_1758_n 0.00409726f $X=11.44 $Y=0.835 $X2=0
+ $Y2=0
cc_854 N_A_1723_48#_c_1120_n N_VGND_c_1758_n 0.0131847f $X=9.77 $Y=0.75 $X2=0
+ $Y2=0
cc_855 N_A_1529_74#_M1014_g N_VPWR_c_1424_n 0.00668659f $X=9.54 $Y=2.46 $X2=0
+ $Y2=0
cc_856 N_A_1529_74#_c_1266_n N_VPWR_c_1424_n 0.00487611f $X=8.07 $Y=2.815 $X2=0
+ $Y2=0
cc_857 N_A_1529_74#_M1014_g N_VPWR_c_1425_n 0.00448333f $X=9.54 $Y=2.46 $X2=0
+ $Y2=0
cc_858 N_A_1529_74#_c_1266_n N_VPWR_c_1430_n 0.014549f $X=8.07 $Y=2.815 $X2=0
+ $Y2=0
cc_859 N_A_1529_74#_M1014_g N_VPWR_c_1431_n 0.005209f $X=9.54 $Y=2.46 $X2=0
+ $Y2=0
cc_860 N_A_1529_74#_M1014_g N_VPWR_c_1420_n 0.00988987f $X=9.54 $Y=2.46 $X2=0
+ $Y2=0
cc_861 N_A_1529_74#_c_1266_n N_VPWR_c_1420_n 0.0119743f $X=8.07 $Y=2.815 $X2=0
+ $Y2=0
cc_862 N_A_1529_74#_M1001_g N_VGND_c_1747_n 0.0145549f $X=9.46 $Y=0.645 $X2=0
+ $Y2=0
cc_863 N_A_1529_74#_c_1255_n N_VGND_c_1747_n 0.0090058f $X=8.85 $Y=1.065 $X2=0
+ $Y2=0
cc_864 N_A_1529_74#_c_1258_n N_VGND_c_1747_n 0.0146855f $X=9.28 $Y=1.185 $X2=0
+ $Y2=0
cc_865 N_A_1529_74#_c_1259_n N_VGND_c_1747_n 0.0199258f $X=8.475 $Y=0.58 $X2=0
+ $Y2=0
cc_866 N_A_1529_74#_c_1260_n N_VGND_c_1747_n 0.0157382f $X=8.935 $Y=1.065 $X2=0
+ $Y2=0
cc_867 N_A_1529_74#_c_1261_n N_VGND_c_1747_n 0.00565625f $X=9.445 $Y=1.265 $X2=0
+ $Y2=0
cc_868 N_A_1529_74#_c_1262_n N_VGND_c_1747_n 5.47931e-19 $X=9.445 $Y=1.265 $X2=0
+ $Y2=0
cc_869 N_A_1529_74#_M1001_g N_VGND_c_1748_n 0.00318791f $X=9.46 $Y=0.645 $X2=0
+ $Y2=0
cc_870 N_A_1529_74#_M1001_g N_VGND_c_1750_n 0.00383152f $X=9.46 $Y=0.645 $X2=0
+ $Y2=0
cc_871 N_A_1529_74#_c_1259_n N_VGND_c_1755_n 0.0224701f $X=8.475 $Y=0.58 $X2=0
+ $Y2=0
cc_872 N_A_1529_74#_M1001_g N_VGND_c_1758_n 0.00762539f $X=9.46 $Y=0.645 $X2=0
+ $Y2=0
cc_873 N_A_1529_74#_c_1259_n N_VGND_c_1758_n 0.0185858f $X=8.475 $Y=0.58 $X2=0
+ $Y2=0
cc_874 N_A_2216_112#_c_1371_n N_VPWR_c_1426_n 0.00267634f $X=11.985 $Y=1.64
+ $X2=0 $Y2=0
cc_875 N_A_2216_112#_M1034_g N_VPWR_c_1426_n 0.00607682f $X=11.985 $Y=2.4 $X2=0
+ $Y2=0
cc_876 N_A_2216_112#_c_1375_n N_VPWR_c_1426_n 0.030344f $X=11.255 $Y=2.16 $X2=0
+ $Y2=0
cc_877 N_A_2216_112#_c_1376_n N_VPWR_c_1426_n 0.0130288f $X=11.89 $Y=1.385 $X2=0
+ $Y2=0
cc_878 N_A_2216_112#_c_1375_n N_VPWR_c_1432_n 0.00775887f $X=11.255 $Y=2.16
+ $X2=0 $Y2=0
cc_879 N_A_2216_112#_M1034_g N_VPWR_c_1433_n 0.005209f $X=11.985 $Y=2.4 $X2=0
+ $Y2=0
cc_880 N_A_2216_112#_M1034_g N_VPWR_c_1420_n 0.00990545f $X=11.985 $Y=2.4 $X2=0
+ $Y2=0
cc_881 N_A_2216_112#_c_1375_n N_VPWR_c_1420_n 0.00855956f $X=11.255 $Y=2.16
+ $X2=0 $Y2=0
cc_882 N_A_2216_112#_c_1375_n N_Q_c_1693_n 0.10299f $X=11.255 $Y=2.16 $X2=0
+ $Y2=0
cc_883 N_A_2216_112#_c_1377_n N_Q_c_1693_n 0.0253889f $X=11.215 $Y=1.385 $X2=0
+ $Y2=0
cc_884 N_A_2216_112#_c_1374_n N_Q_c_1694_n 0.0534224f $X=11.225 $Y=0.835 $X2=0
+ $Y2=0
cc_885 N_A_2216_112#_c_1373_n Q_N 0.00609353f $X=11.985 $Y=1.22 $X2=0 $Y2=0
cc_886 N_A_2216_112#_c_1371_n Q_N 0.00871962f $X=11.985 $Y=1.64 $X2=0 $Y2=0
cc_887 N_A_2216_112#_c_1373_n Q_N 0.0127686f $X=11.985 $Y=1.22 $X2=0 $Y2=0
cc_888 N_A_2216_112#_c_1376_n Q_N 0.0267051f $X=11.89 $Y=1.385 $X2=0 $Y2=0
cc_889 N_A_2216_112#_M1034_g Q_N 0.0181768f $X=11.985 $Y=2.4 $X2=0 $Y2=0
cc_890 N_A_2216_112#_c_1373_n Q_N 0.00323868f $X=11.985 $Y=1.22 $X2=0 $Y2=0
cc_891 N_A_2216_112#_c_1371_n N_VGND_c_1749_n 0.0031522f $X=11.985 $Y=1.64 $X2=0
+ $Y2=0
cc_892 N_A_2216_112#_c_1373_n N_VGND_c_1749_n 0.00695589f $X=11.985 $Y=1.22
+ $X2=0 $Y2=0
cc_893 N_A_2216_112#_c_1374_n N_VGND_c_1749_n 0.0182577f $X=11.225 $Y=0.835
+ $X2=0 $Y2=0
cc_894 N_A_2216_112#_c_1376_n N_VGND_c_1749_n 0.0252425f $X=11.89 $Y=1.385 $X2=0
+ $Y2=0
cc_895 N_A_2216_112#_c_1374_n N_VGND_c_1756_n 0.0054549f $X=11.225 $Y=0.835
+ $X2=0 $Y2=0
cc_896 N_A_2216_112#_c_1373_n N_VGND_c_1757_n 0.00434272f $X=11.985 $Y=1.22
+ $X2=0 $Y2=0
cc_897 N_A_2216_112#_c_1373_n N_VGND_c_1758_n 0.00828717f $X=11.985 $Y=1.22
+ $X2=0 $Y2=0
cc_898 N_A_2216_112#_c_1374_n N_VGND_c_1758_n 0.00708918f $X=11.225 $Y=0.835
+ $X2=0 $Y2=0
cc_899 N_VPWR_M1009_d N_A_296_74#_c_1575_n 0.0110613f $X=2.59 $Y=2.32 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1420_n N_A_296_74#_c_1575_n 0.0232759f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1436_n N_A_296_74#_c_1575_n 0.0217273f $X=2.855 $Y=2.815 $X2=0
+ $Y2=0
cc_902 N_VPWR_M1009_d N_A_296_74#_c_1564_n 0.00964217f $X=2.59 $Y=2.32 $X2=0
+ $Y2=0
cc_903 N_VPWR_M1025_s N_A_296_74#_c_1569_n 0.0115547f $X=3.85 $Y=1.84 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1422_n N_A_296_74#_c_1569_n 0.0288112f $X=4.08 $Y=2.815 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1420_n N_A_296_74#_c_1569_n 0.0255591f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1436_n N_A_296_74#_c_1569_n 0.00214766f $X=2.855 $Y=2.815 $X2=0
+ $Y2=0
cc_907 N_VPWR_M1025_s N_A_296_74#_c_1570_n 0.0125907f $X=3.85 $Y=1.84 $X2=0
+ $Y2=0
cc_908 N_VPWR_c_1429_n N_A_296_74#_c_1571_n 0.00487697f $X=6.45 $Y=3.33 $X2=0
+ $Y2=0
cc_909 N_VPWR_c_1420_n N_A_296_74#_c_1571_n 0.00841085f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_910 N_VPWR_M1025_s N_A_296_74#_c_1625_n 5.64071e-19 $X=3.85 $Y=1.84 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1422_n N_A_296_74#_c_1625_n 0.00696805f $X=4.08 $Y=2.815 $X2=0
+ $Y2=0
cc_912 N_VPWR_c_1429_n N_A_296_74#_c_1625_n 0.00238305f $X=6.45 $Y=3.33 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1420_n N_A_296_74#_c_1625_n 0.0105802f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1422_n N_A_296_74#_c_1572_n 0.00545691f $X=4.08 $Y=2.815 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1429_n N_A_296_74#_c_1572_n 0.0086639f $X=6.45 $Y=3.33 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1420_n N_A_296_74#_c_1572_n 0.00869469f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1421_n N_A_296_74#_c_1573_n 0.0200631f $X=0.865 $Y=2.465 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1427_n N_A_296_74#_c_1573_n 0.0144623f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1420_n N_A_296_74#_c_1573_n 0.0118344f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1436_n N_A_296_74#_c_1573_n 0.00632485f $X=2.855 $Y=2.815 $X2=0
+ $Y2=0
cc_921 N_VPWR_M1009_d N_A_296_74#_c_1679_n 0.00223497f $X=2.59 $Y=2.32 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1420_n N_A_296_74#_c_1679_n 6.82232e-19 $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1436_n N_A_296_74#_c_1679_n 0.0146376f $X=2.855 $Y=2.815 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1425_n N_Q_c_1696_n 0.0395806f $X=10.285 $Y=1.985 $X2=0 $Y2=0
cc_925 N_VPWR_c_1426_n N_Q_c_1697_n 0.00304034f $X=11.705 $Y=2.16 $X2=0 $Y2=0
cc_926 N_VPWR_c_1432_n N_Q_c_1697_n 0.0117353f $X=11.54 $Y=3.33 $X2=0 $Y2=0
cc_927 N_VPWR_c_1420_n N_Q_c_1697_n 0.00971347f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_928 N_VPWR_c_1426_n Q_N 0.0368843f $X=11.705 $Y=2.16 $X2=0 $Y2=0
cc_929 N_VPWR_c_1433_n Q_N 0.014549f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_930 N_VPWR_c_1420_n Q_N 0.0119743f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_931 N_A_296_74#_c_1575_n A_410_464# 0.0123094f $X=2.895 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_932 N_A_296_74#_c_1574_n N_VGND_c_1742_n 0.00833256f $X=2.22 $Y=0.515 $X2=0
+ $Y2=0
cc_933 N_A_296_74#_c_1561_n N_VGND_c_1743_n 0.00120995f $X=2.305 $Y=1.18 $X2=0
+ $Y2=0
cc_934 N_A_296_74#_c_1562_n N_VGND_c_1743_n 0.0115398f $X=2.895 $Y=1.265 $X2=0
+ $Y2=0
cc_935 N_A_296_74#_c_1574_n N_VGND_c_1753_n 0.0294503f $X=2.22 $Y=0.515 $X2=0
+ $Y2=0
cc_936 N_A_296_74#_c_1574_n N_VGND_c_1758_n 0.0318847f $X=2.22 $Y=0.515 $X2=0
+ $Y2=0
cc_937 N_A_296_74#_c_1574_n A_434_74# 0.00164902f $X=2.22 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_938 N_Q_c_1694_n N_VGND_c_1748_n 0.0302899f $X=10.665 $Y=0.515 $X2=0 $Y2=0
cc_939 N_Q_c_1694_n N_VGND_c_1749_n 0.00650919f $X=10.665 $Y=0.515 $X2=0 $Y2=0
cc_940 N_Q_c_1694_n N_VGND_c_1756_n 0.0183567f $X=10.665 $Y=0.515 $X2=0 $Y2=0
cc_941 N_Q_c_1694_n N_VGND_c_1758_n 0.0151377f $X=10.665 $Y=0.515 $X2=0 $Y2=0
cc_942 Q_N N_VGND_c_1749_n 0.0260234f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_943 Q_N N_VGND_c_1757_n 0.0150211f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_944 Q_N N_VGND_c_1758_n 0.0123721f $X=12.155 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__or4b_2.pxi.spice
* Created: Wed Sep  2 12:29:17 2020
* 
x_PM_SKY130_FD_SC_MS__OR4B_2%D_N N_D_N_c_84_n N_D_N_M1003_g N_D_N_M1010_g D_N
+ N_D_N_c_86_n PM_SKY130_FD_SC_MS__OR4B_2%D_N
x_PM_SKY130_FD_SC_MS__OR4B_2%A_190_48# N_A_190_48#_M1004_d N_A_190_48#_M1002_d
+ N_A_190_48#_M1006_d N_A_190_48#_M1005_g N_A_190_48#_M1009_g
+ N_A_190_48#_c_113_n N_A_190_48#_M1013_g N_A_190_48#_M1012_g
+ N_A_190_48#_c_116_n N_A_190_48#_c_117_n N_A_190_48#_c_118_n
+ N_A_190_48#_c_200_p N_A_190_48#_c_119_n N_A_190_48#_c_120_n
+ N_A_190_48#_c_121_n N_A_190_48#_c_130_n N_A_190_48#_c_122_n
+ N_A_190_48#_c_123_n N_A_190_48#_c_124_n N_A_190_48#_c_125_n
+ N_A_190_48#_c_131_n N_A_190_48#_c_126_n N_A_190_48#_c_127_n
+ PM_SKY130_FD_SC_MS__OR4B_2%A_190_48#
x_PM_SKY130_FD_SC_MS__OR4B_2%A N_A_M1004_g N_A_M1000_g A A N_A_c_239_n
+ N_A_c_240_n PM_SKY130_FD_SC_MS__OR4B_2%A
x_PM_SKY130_FD_SC_MS__OR4B_2%B N_B_M1007_g N_B_M1008_g B B N_B_c_287_n
+ PM_SKY130_FD_SC_MS__OR4B_2%B
x_PM_SKY130_FD_SC_MS__OR4B_2%C N_C_M1001_g N_C_M1002_g C C C N_C_c_326_n
+ PM_SKY130_FD_SC_MS__OR4B_2%C
x_PM_SKY130_FD_SC_MS__OR4B_2%A_27_368# N_A_27_368#_M1010_s N_A_27_368#_M1003_s
+ N_A_27_368#_M1006_g N_A_27_368#_M1011_g N_A_27_368#_c_361_n
+ N_A_27_368#_c_362_n N_A_27_368#_c_363_n N_A_27_368#_c_364_n
+ N_A_27_368#_c_394_n N_A_27_368#_c_369_n N_A_27_368#_c_398_n
+ N_A_27_368#_c_432_p N_A_27_368#_c_370_n N_A_27_368#_c_365_n
+ N_A_27_368#_c_366_n PM_SKY130_FD_SC_MS__OR4B_2%A_27_368#
x_PM_SKY130_FD_SC_MS__OR4B_2%VPWR N_VPWR_M1003_d N_VPWR_M1012_s N_VPWR_c_459_n
+ VPWR N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_458_n N_VPWR_c_463_n
+ N_VPWR_c_464_n PM_SKY130_FD_SC_MS__OR4B_2%VPWR
x_PM_SKY130_FD_SC_MS__OR4B_2%X N_X_M1005_d N_X_M1009_d N_X_c_502_n N_X_c_503_n X
+ N_X_c_504_n PM_SKY130_FD_SC_MS__OR4B_2%X
x_PM_SKY130_FD_SC_MS__OR4B_2%VGND N_VGND_M1010_d N_VGND_M1013_s N_VGND_M1008_d
+ N_VGND_M1011_d N_VGND_c_547_n N_VGND_c_548_n N_VGND_c_549_n N_VGND_c_550_n
+ N_VGND_c_551_n VGND N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n
+ N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n
+ PM_SKY130_FD_SC_MS__OR4B_2%VGND
cc_1 VNB N_D_N_c_84_n 0.0339332f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.77
cc_2 VNB N_D_N_M1010_g 0.0335586f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.835
cc_3 VNB N_D_N_c_86_n 0.0147527f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_190_48#_M1005_g 0.0217322f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_5 VNB N_A_190_48#_M1009_g 0.0110629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_190_48#_c_113_n 0.0134199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_190_48#_M1013_g 0.0229022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_190_48#_M1012_g 0.00168498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_190_48#_c_116_n 0.00626877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_190_48#_c_117_n 0.00305584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_190_48#_c_118_n 0.00740858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_190_48#_c_119_n 0.00379109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_190_48#_c_120_n 0.00326291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_190_48#_c_121_n 0.0126446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_190_48#_c_122_n 0.00293951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_190_48#_c_123_n 0.00951601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_190_48#_c_124_n 0.0103969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_190_48#_c_125_n 0.00809499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_190_48#_c_126_n 0.0186681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_190_48#_c_127_n 0.031148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_M1004_g 0.0266404f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_22 VNB N_A_c_239_n 0.0268394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_240_n 0.00183238f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_24 VNB N_B_M1008_g 0.0350429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB B 0.00220385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_287_n 0.0180468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_M1002_g 0.0343028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB C 0.00367115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C_c_326_n 0.0168455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_368#_M1011_g 0.0311486f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_31 VNB N_A_27_368#_c_361_n 0.0214174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_368#_c_362_n 0.00510302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_368#_c_363_n 0.00942464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_368#_c_364_n 0.0086419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_368#_c_365_n 0.00386761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_368#_c_366_n 0.0207748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_458_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_502_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_503_n 0.00434772f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_40 VNB N_X_c_504_n 0.00226257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_547_n 0.0157056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_548_n 0.0117064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_549_n 0.0147881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_550_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_551_n 0.0366542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_552_n 0.0190549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_553_n 0.0197882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_554_n 0.0191517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_555_n 0.0255552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_556_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_557_n 0.0100021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_558_n 0.265964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_D_N_c_84_n 0.0366557f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.77
cc_54 VPB N_D_N_c_86_n 0.00730023f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_55 VPB N_A_190_48#_M1009_g 0.0238834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_190_48#_M1012_g 0.0243326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_190_48#_c_130_n 0.0377236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_190_48#_c_131_n 0.010431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_190_48#_c_126_n 0.013323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_M1000_g 0.0290868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_c_239_n 0.00574133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_c_240_n 0.0031429f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_63 VPB N_B_M1007_g 0.0208594f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_64 VPB B 0.00207778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B_c_287_n 0.0137801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_C_M1001_g 0.0221952f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_67 VPB C 0.0029589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_C_c_326_n 0.0128841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_368#_M1006_g 0.0282981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_368#_c_364_n 0.00320434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_368#_c_369_n 0.0349325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_368#_c_370_n 0.0013256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_368#_c_365_n 0.00178662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_27_368#_c_366_n 0.0153136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_459_n 0.0162527f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_76 VPB N_VPWR_c_460_n 0.0177898f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_77 VPB N_VPWR_c_461_n 0.0603644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_458_n 0.070198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_463_n 0.0274712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_464_n 0.0156038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB X 0.00206185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_X_c_504_n 0.00105576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 N_D_N_M1010_g N_A_190_48#_M1005_g 0.0140885f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_84 N_D_N_c_84_n N_A_190_48#_M1009_g 0.0302802f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_85 N_D_N_c_84_n N_A_190_48#_c_116_n 0.0140885f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_86 N_D_N_M1010_g N_A_27_368#_c_361_n 0.00872945f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_87 N_D_N_c_84_n N_A_27_368#_c_362_n 2.93656e-19 $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_88 N_D_N_M1010_g N_A_27_368#_c_362_n 0.0120739f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_89 N_D_N_c_86_n N_A_27_368#_c_362_n 0.00649299f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_90 N_D_N_c_84_n N_A_27_368#_c_363_n 0.00168251f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_91 N_D_N_M1010_g N_A_27_368#_c_363_n 0.00377477f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_92 N_D_N_c_86_n N_A_27_368#_c_363_n 0.0286137f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_93 N_D_N_c_84_n N_A_27_368#_c_364_n 0.00457725f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_94 N_D_N_M1010_g N_A_27_368#_c_364_n 0.00640717f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_95 N_D_N_c_86_n N_A_27_368#_c_364_n 0.0329135f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_96 N_D_N_c_84_n N_A_27_368#_c_369_n 0.030358f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_97 N_D_N_c_86_n N_A_27_368#_c_369_n 0.0338794f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_98 N_D_N_c_84_n N_VPWR_c_459_n 0.00339971f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_99 N_D_N_c_84_n N_VPWR_c_458_n 0.00555093f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_100 N_D_N_c_84_n N_VPWR_c_463_n 0.0046462f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_101 N_D_N_M1010_g N_X_c_502_n 6.35749e-19 $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_102 N_D_N_M1010_g N_VGND_c_547_n 0.00459404f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_103 N_D_N_M1010_g N_VGND_c_555_n 0.0043356f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_104 N_D_N_M1010_g N_VGND_c_558_n 0.00487769f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_105 N_A_190_48#_M1013_g N_A_M1004_g 0.0160656f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_190_48#_c_117_n N_A_M1004_g 0.00351998f $X=1.66 $Y=1.3 $X2=0 $Y2=0
cc_107 N_A_190_48#_c_118_n N_A_M1004_g 0.0156668f $X=2.175 $Y=1.045 $X2=0 $Y2=0
cc_108 N_A_190_48#_c_119_n N_A_M1004_g 0.00321875f $X=2.34 $Y=0.615 $X2=0 $Y2=0
cc_109 N_A_190_48#_c_122_n N_A_M1004_g 0.00107033f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_110 N_A_190_48#_c_127_n N_A_M1004_g 0.00252021f $X=1.555 $Y=1.375 $X2=0 $Y2=0
cc_111 N_A_190_48#_M1012_g N_A_M1000_g 0.0302142f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_190_48#_M1012_g N_A_c_239_n 0.00181814f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_190_48#_c_118_n N_A_c_239_n 5.20343e-19 $X=2.175 $Y=1.045 $X2=0 $Y2=0
cc_114 N_A_190_48#_c_122_n N_A_c_239_n 0.00161664f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A_190_48#_c_123_n N_A_c_239_n 7.46556e-19 $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_116 N_A_190_48#_c_127_n N_A_c_239_n 0.0171073f $X=1.555 $Y=1.375 $X2=0 $Y2=0
cc_117 N_A_190_48#_M1012_g N_A_c_240_n 0.00610477f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_190_48#_c_118_n N_A_c_240_n 0.0144509f $X=2.175 $Y=1.045 $X2=0 $Y2=0
cc_119 N_A_190_48#_c_122_n N_A_c_240_n 0.0197025f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_120 N_A_190_48#_c_123_n N_A_c_240_n 0.00726462f $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_121 N_A_190_48#_c_127_n N_A_c_240_n 3.4058e-19 $X=1.555 $Y=1.375 $X2=0 $Y2=0
cc_122 N_A_190_48#_c_119_n N_B_M1008_g 0.00321875f $X=2.34 $Y=0.615 $X2=0 $Y2=0
cc_123 N_A_190_48#_c_124_n N_B_M1008_g 0.016738f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_124 N_A_190_48#_c_123_n B 0.00100747f $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_125 N_A_190_48#_c_124_n B 0.0140616f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_126 N_A_190_48#_c_124_n N_B_c_287_n 9.60242e-19 $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_127 N_A_190_48#_c_124_n N_C_M1002_g 0.0148482f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_128 N_A_190_48#_c_125_n N_C_M1002_g 0.00468012f $X=3.705 $Y=1.115 $X2=0 $Y2=0
cc_129 N_A_190_48#_c_124_n C 0.0160291f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_130 N_A_190_48#_c_124_n N_C_c_326_n 0.00108269f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_131 N_A_190_48#_c_131_n N_A_27_368#_M1006_g 0.024632f $X=4.03 $Y=2.105 $X2=0
+ $Y2=0
cc_132 N_A_190_48#_c_126_n N_A_27_368#_M1006_g 0.00309918f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_133 N_A_190_48#_c_120_n N_A_27_368#_M1011_g 0.00700031f $X=3.54 $Y=0.615
+ $X2=0 $Y2=0
cc_134 N_A_190_48#_c_121_n N_A_27_368#_M1011_g 0.0127639f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_135 N_A_190_48#_c_125_n N_A_27_368#_M1011_g 0.0092772f $X=3.705 $Y=1.115
+ $X2=0 $Y2=0
cc_136 N_A_190_48#_c_126_n N_A_27_368#_M1011_g 0.00539566f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_137 N_A_190_48#_M1005_g N_A_27_368#_c_361_n 5.93853e-19 $X=1.025 $Y=0.74
+ $X2=0 $Y2=0
cc_138 N_A_190_48#_M1005_g N_A_27_368#_c_362_n 0.0015418f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_190_48#_M1005_g N_A_27_368#_c_364_n 0.00655019f $X=1.025 $Y=0.74
+ $X2=0 $Y2=0
cc_140 N_A_190_48#_M1009_g N_A_27_368#_c_394_n 0.016896f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_141 N_A_190_48#_M1012_g N_A_27_368#_c_394_n 0.0188375f $X=1.49 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_190_48#_c_127_n N_A_27_368#_c_394_n 0.0027222f $X=1.555 $Y=1.375
+ $X2=0 $Y2=0
cc_143 N_A_190_48#_M1009_g N_A_27_368#_c_369_n 0.00798707f $X=1.04 $Y=2.4 $X2=0
+ $Y2=0
cc_144 N_A_190_48#_c_130_n N_A_27_368#_c_398_n 0.0141265f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_145 N_A_190_48#_c_131_n N_A_27_368#_c_370_n 0.0559687f $X=4.03 $Y=2.105 $X2=0
+ $Y2=0
cc_146 N_A_190_48#_c_126_n N_A_27_368#_c_370_n 0.00677874f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_147 N_A_190_48#_c_125_n N_A_27_368#_c_365_n 0.0280161f $X=3.705 $Y=1.115
+ $X2=0 $Y2=0
cc_148 N_A_190_48#_c_131_n N_A_27_368#_c_365_n 0.00244567f $X=4.03 $Y=2.105
+ $X2=0 $Y2=0
cc_149 N_A_190_48#_c_126_n N_A_27_368#_c_365_n 0.0249903f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_150 N_A_190_48#_c_121_n N_A_27_368#_c_366_n 0.00145734f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_151 N_A_190_48#_c_125_n N_A_27_368#_c_366_n 0.00306887f $X=3.705 $Y=1.115
+ $X2=0 $Y2=0
cc_152 N_A_190_48#_c_131_n N_A_27_368#_c_366_n 6.75574e-19 $X=4.03 $Y=2.105
+ $X2=0 $Y2=0
cc_153 N_A_190_48#_c_126_n N_A_27_368#_c_366_n 0.00231223f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_154 N_A_190_48#_M1009_g N_VPWR_c_459_n 0.0118162f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_190_48#_M1012_g N_VPWR_c_459_n 0.00138681f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_190_48#_M1009_g N_VPWR_c_460_n 0.00460063f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_190_48#_M1012_g N_VPWR_c_460_n 0.00461464f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_190_48#_c_130_n N_VPWR_c_461_n 0.0164205f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_159 N_A_190_48#_M1009_g N_VPWR_c_458_n 0.0046086f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_190_48#_M1012_g N_VPWR_c_458_n 0.0046086f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_190_48#_c_130_n N_VPWR_c_458_n 0.0135915f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_162 N_A_190_48#_M1009_g N_VPWR_c_464_n 0.00105016f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_190_48#_M1012_g N_VPWR_c_464_n 0.0144568f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_190_48#_M1005_g N_X_c_502_n 0.00922867f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_190_48#_M1013_g N_X_c_502_n 0.00930665f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_190_48#_M1005_g N_X_c_503_n 0.0026107f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_190_48#_c_113_n N_X_c_503_n 0.00246648f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_168 N_A_190_48#_M1013_g N_X_c_503_n 0.00294637f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_190_48#_c_200_p N_X_c_503_n 0.00733863f $X=1.745 $Y=1.045 $X2=0 $Y2=0
cc_170 N_A_190_48#_M1009_g X 0.00584623f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_190_48#_c_113_n X 0.00501807f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_172 N_A_190_48#_M1012_g X 0.00739803f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A_190_48#_c_122_n X 0.00200011f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_174 N_A_190_48#_c_127_n X 8.69852e-19 $X=1.555 $Y=1.375 $X2=0 $Y2=0
cc_175 N_A_190_48#_M1005_g N_X_c_504_n 0.00330399f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_190_48#_M1009_g N_X_c_504_n 0.00755278f $X=1.04 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_190_48#_c_113_n N_X_c_504_n 0.00668903f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_178 N_A_190_48#_M1013_g N_X_c_504_n 9.29964e-19 $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_190_48#_M1012_g N_X_c_504_n 0.00289597f $X=1.49 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_190_48#_c_116_n N_X_c_504_n 0.00212694f $X=1.04 $Y=1.375 $X2=0 $Y2=0
cc_181 N_A_190_48#_c_117_n N_X_c_504_n 0.00551929f $X=1.66 $Y=1.3 $X2=0 $Y2=0
cc_182 N_A_190_48#_c_122_n N_X_c_504_n 0.0242992f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_183 N_A_190_48#_c_127_n N_X_c_504_n 0.00110944f $X=1.555 $Y=1.375 $X2=0 $Y2=0
cc_184 N_A_190_48#_c_118_n N_VGND_M1013_s 0.00218122f $X=2.175 $Y=1.045 $X2=0
+ $Y2=0
cc_185 N_A_190_48#_c_200_p N_VGND_M1013_s 0.00305443f $X=1.745 $Y=1.045 $X2=0
+ $Y2=0
cc_186 N_A_190_48#_c_124_n N_VGND_M1008_d 0.00526182f $X=3.375 $Y=1.115 $X2=0
+ $Y2=0
cc_187 N_A_190_48#_c_121_n N_VGND_M1011_d 0.00330281f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_188 N_A_190_48#_M1005_g N_VGND_c_547_n 0.00709895f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_190_48#_M1013_g N_VGND_c_548_n 0.00743057f $X=1.455 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_190_48#_c_118_n N_VGND_c_548_n 0.0147668f $X=2.175 $Y=1.045 $X2=0
+ $Y2=0
cc_191 N_A_190_48#_c_200_p N_VGND_c_548_n 0.0129834f $X=1.745 $Y=1.045 $X2=0
+ $Y2=0
cc_192 N_A_190_48#_c_119_n N_VGND_c_548_n 0.0130314f $X=2.34 $Y=0.615 $X2=0
+ $Y2=0
cc_193 N_A_190_48#_c_127_n N_VGND_c_548_n 5.79689e-19 $X=1.555 $Y=1.375 $X2=0
+ $Y2=0
cc_194 N_A_190_48#_c_119_n N_VGND_c_549_n 0.0134386f $X=2.34 $Y=0.615 $X2=0
+ $Y2=0
cc_195 N_A_190_48#_c_120_n N_VGND_c_549_n 0.00163718f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_196 N_A_190_48#_c_124_n N_VGND_c_549_n 0.0314461f $X=3.375 $Y=1.115 $X2=0
+ $Y2=0
cc_197 N_A_190_48#_c_120_n N_VGND_c_551_n 0.0188012f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_198 N_A_190_48#_c_121_n N_VGND_c_551_n 0.027045f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_199 N_A_190_48#_M1005_g N_VGND_c_552_n 0.00417277f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_200 N_A_190_48#_M1013_g N_VGND_c_552_n 0.00434272f $X=1.455 $Y=0.74 $X2=0
+ $Y2=0
cc_201 N_A_190_48#_c_119_n N_VGND_c_553_n 0.010412f $X=2.34 $Y=0.615 $X2=0 $Y2=0
cc_202 N_A_190_48#_c_120_n N_VGND_c_554_n 0.010139f $X=3.54 $Y=0.615 $X2=0 $Y2=0
cc_203 N_A_190_48#_M1005_g N_VGND_c_558_n 0.00770365f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_204 N_A_190_48#_M1013_g N_VGND_c_558_n 0.00825059f $X=1.455 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_190_48#_c_119_n N_VGND_c_558_n 0.0113592f $X=2.34 $Y=0.615 $X2=0
+ $Y2=0
cc_206 N_A_190_48#_c_120_n N_VGND_c_558_n 0.0112086f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_207 N_A_M1000_g N_B_M1007_g 0.0664f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_208 N_A_c_240_n N_B_M1007_g 4.25461e-19 $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_209 N_A_M1004_g N_B_M1008_g 0.0230804f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_210 N_A_c_239_n N_B_M1008_g 0.00559311f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_211 N_A_c_240_n N_B_M1008_g 7.46398e-19 $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_212 N_A_M1000_g B 0.00143696f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_213 N_A_c_239_n B 0.00110276f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_214 N_A_c_240_n B 0.0376777f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A_c_239_n N_B_c_287_n 0.0197624f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A_c_240_n N_B_c_287_n 0.00114872f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_M1000_g N_A_27_368#_c_394_n 0.0134763f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_218 N_A_c_239_n N_A_27_368#_c_394_n 3.5167e-19 $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A_c_240_n N_A_27_368#_c_394_n 0.0211204f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_220 N_A_c_240_n N_VPWR_M1012_s 0.00384934f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_221 N_A_M1000_g N_VPWR_c_461_n 0.00461464f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_222 N_A_M1000_g N_VPWR_c_458_n 0.00460677f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_223 N_A_M1000_g N_VPWR_c_464_n 0.0135675f $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_224 N_A_M1004_g N_X_c_502_n 8.75421e-19 $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_225 N_A_M1000_g X 2.76706e-19 $X=2.185 $Y=2.46 $X2=0 $Y2=0
cc_226 N_A_c_240_n X 0.0111395f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A_M1004_g N_VGND_c_548_n 0.00862467f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_228 N_A_M1004_g N_VGND_c_549_n 5.59444e-19 $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_229 N_A_M1004_g N_VGND_c_553_n 0.00421418f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_230 N_A_M1004_g N_VGND_c_558_n 0.00432128f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_231 N_B_M1007_g N_C_M1001_g 0.0487255f $X=2.605 $Y=2.46 $X2=0 $Y2=0
cc_232 B N_C_M1001_g 0.00125169f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B_M1008_g N_C_M1002_g 0.0250853f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_234 N_B_M1007_g C 5.8851e-19 $X=2.605 $Y=2.46 $X2=0 $Y2=0
cc_235 B C 0.0434887f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B_c_287_n C 0.00188716f $X=2.65 $Y=1.635 $X2=0 $Y2=0
cc_237 B N_C_c_326_n 3.99347e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B_c_287_n N_C_c_326_n 0.0206935f $X=2.65 $Y=1.635 $X2=0 $Y2=0
cc_239 N_B_M1007_g N_A_27_368#_c_398_n 0.0138361f $X=2.605 $Y=2.46 $X2=0 $Y2=0
cc_240 B N_A_27_368#_c_398_n 0.00742996f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B_M1007_g N_VPWR_c_461_n 0.00368591f $X=2.605 $Y=2.46 $X2=0 $Y2=0
cc_242 N_B_M1007_g N_VPWR_c_458_n 0.00451809f $X=2.605 $Y=2.46 $X2=0 $Y2=0
cc_243 N_B_M1007_g N_VPWR_c_464_n 0.00120517f $X=2.605 $Y=2.46 $X2=0 $Y2=0
cc_244 B A_539_392# 0.00294111f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_245 N_B_M1008_g N_VGND_c_548_n 5.60991e-19 $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_246 N_B_M1008_g N_VGND_c_549_n 0.0142125f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_247 N_B_M1008_g N_VGND_c_553_n 0.00421418f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_248 N_B_M1008_g N_VGND_c_558_n 0.00432128f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_249 N_C_M1001_g N_A_27_368#_M1006_g 0.0429408f $X=3.115 $Y=2.46 $X2=0 $Y2=0
cc_250 C N_A_27_368#_M1006_g 0.00250531f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_251 N_C_c_326_n N_A_27_368#_M1006_g 0.0111791f $X=3.19 $Y=1.635 $X2=0 $Y2=0
cc_252 N_C_M1002_g N_A_27_368#_M1011_g 0.0173114f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_253 N_C_M1001_g N_A_27_368#_c_398_n 0.0127032f $X=3.115 $Y=2.46 $X2=0 $Y2=0
cc_254 C N_A_27_368#_c_398_n 0.0205527f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_255 N_C_M1001_g N_A_27_368#_c_370_n 7.79231e-19 $X=3.115 $Y=2.46 $X2=0 $Y2=0
cc_256 C N_A_27_368#_c_370_n 0.0376258f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_257 N_C_M1002_g N_A_27_368#_c_365_n 0.00238017f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_258 C N_A_27_368#_c_365_n 0.0240984f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_259 N_C_M1002_g N_A_27_368#_c_366_n 0.0111791f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_260 C N_A_27_368#_c_366_n 3.43837e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_261 N_C_M1001_g N_VPWR_c_461_n 0.00368591f $X=3.115 $Y=2.46 $X2=0 $Y2=0
cc_262 N_C_M1001_g N_VPWR_c_458_n 0.00452895f $X=3.115 $Y=2.46 $X2=0 $Y2=0
cc_263 C A_641_392# 0.0058651f $X=3.035 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_264 N_C_M1002_g N_VGND_c_549_n 0.00481242f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_265 N_C_M1002_g N_VGND_c_554_n 0.00505936f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_266 N_C_M1002_g N_VGND_c_558_n 0.00514438f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_267 N_A_27_368#_c_364_n N_VPWR_M1003_d 0.00275776f $X=0.805 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_27_368#_c_369_n N_VPWR_M1003_d 0.0105812f $X=0.89 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_27_368#_c_394_n N_VPWR_M1012_s 0.0171418f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_270 N_A_27_368#_c_394_n N_VPWR_c_459_n 0.00225335f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_271 N_A_27_368#_c_369_n N_VPWR_c_459_n 0.0227941f $X=0.89 $Y=2.405 $X2=0
+ $Y2=0
cc_272 N_A_27_368#_M1006_g N_VPWR_c_461_n 0.00419919f $X=3.655 $Y=2.46 $X2=0
+ $Y2=0
cc_273 N_A_27_368#_c_398_n N_VPWR_c_461_n 0.0290273f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_274 N_A_27_368#_c_432_p N_VPWR_c_461_n 0.00426915f $X=2.465 $Y=2.775 $X2=0
+ $Y2=0
cc_275 N_A_27_368#_M1006_g N_VPWR_c_458_n 0.00633599f $X=3.655 $Y=2.46 $X2=0
+ $Y2=0
cc_276 N_A_27_368#_c_394_n N_VPWR_c_458_n 0.0247941f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_277 N_A_27_368#_c_369_n N_VPWR_c_458_n 0.0182424f $X=0.89 $Y=2.405 $X2=0
+ $Y2=0
cc_278 N_A_27_368#_c_398_n N_VPWR_c_458_n 0.0377243f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_279 N_A_27_368#_c_432_p N_VPWR_c_458_n 0.00575379f $X=2.465 $Y=2.775 $X2=0
+ $Y2=0
cc_280 N_A_27_368#_c_369_n N_VPWR_c_463_n 0.006683f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_281 N_A_27_368#_c_394_n N_VPWR_c_464_n 0.0271244f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_282 N_A_27_368#_c_394_n N_X_M1009_d 0.00479467f $X=2.295 $Y=2.405 $X2=0 $Y2=0
cc_283 N_A_27_368#_c_361_n N_X_c_502_n 0.00448258f $X=0.295 $Y=0.835 $X2=0 $Y2=0
cc_284 N_A_27_368#_c_362_n N_X_c_503_n 0.0143703f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_285 N_A_27_368#_c_394_n X 0.0194343f $X=2.295 $Y=2.405 $X2=0 $Y2=0
cc_286 N_A_27_368#_c_369_n X 0.016649f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_287 N_A_27_368#_c_364_n N_X_c_504_n 0.0556985f $X=0.805 $Y=1.95 $X2=0 $Y2=0
cc_288 N_A_27_368#_c_394_n A_455_392# 0.00555572f $X=2.295 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_27_368#_c_432_p A_455_392# 0.00185043f $X=2.465 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_290 N_A_27_368#_c_398_n A_539_392# 0.0100529f $X=3.525 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_27_368#_c_398_n A_641_392# 0.0102834f $X=3.525 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_27_368#_c_362_n N_VGND_M1010_d 0.0041785f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A_27_368#_c_361_n N_VGND_c_547_n 0.0114804f $X=0.295 $Y=0.835 $X2=0
+ $Y2=0
cc_294 N_A_27_368#_c_362_n N_VGND_c_547_n 0.0215468f $X=0.72 $Y=1.095 $X2=0
+ $Y2=0
cc_295 N_A_27_368#_M1011_g N_VGND_c_551_n 0.0126413f $X=3.755 $Y=0.79 $X2=0
+ $Y2=0
cc_296 N_A_27_368#_M1011_g N_VGND_c_554_n 0.00485498f $X=3.755 $Y=0.79 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_361_n N_VGND_c_555_n 0.00811255f $X=0.295 $Y=0.835 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_M1011_g N_VGND_c_558_n 0.00514438f $X=3.755 $Y=0.79 $X2=0
+ $Y2=0
cc_299 N_A_27_368#_c_361_n N_VGND_c_558_n 0.0106114f $X=0.295 $Y=0.835 $X2=0
+ $Y2=0
cc_300 N_X_c_502_n N_VGND_c_547_n 0.0373918f $X=1.24 $Y=0.515 $X2=0 $Y2=0
cc_301 N_X_c_502_n N_VGND_c_548_n 0.0170646f $X=1.24 $Y=0.515 $X2=0 $Y2=0
cc_302 N_X_c_502_n N_VGND_c_552_n 0.0151167f $X=1.24 $Y=0.515 $X2=0 $Y2=0
cc_303 N_X_c_502_n N_VGND_c_558_n 0.0123643f $X=1.24 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dlymetal6s6s_1.pex.spice
* Created: Wed Sep  2 12:07:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%A 3 7 9 12 13
c32 3 0 5.46905e-20 $X=0.49 $Y=2.05
r33 12 15 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.44
+ $X2=0.402 $Y2=1.605
r34 12 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.44
+ $X2=0.402 $Y2=1.275
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.39
+ $Y=1.44 $X2=0.39 $Y2=1.44
r36 9 13 5.98039 $w=4.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.33 $Y=1.665
+ $X2=0.33 $Y2=1.44
r37 7 14 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.48 $Y=0.9 $X2=0.48
+ $Y2=1.275
r38 3 15 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=0.49 $Y=2.05
+ $X2=0.49 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%A_28_138# 1 2 9 13 15 17 19 20 22 29
+ 33
c66 19 0 1.94125e-19 $X=0.81 $Y=1.605
r67 33 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.44
+ $X2=0.955 $Y2=1.605
r68 33 35 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.955 $Y=1.44
+ $X2=0.955 $Y2=1.26
r69 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.955
+ $Y=1.44 $X2=0.955 $Y2=1.44
r70 30 32 18.9224 $w=2.45e-07 $l=3.8e-07 $layer=LI1_cond $X=0.882 $Y=1.06
+ $X2=0.882 $Y2=1.44
r71 27 29 7.56208 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.08
+ $X2=0.43 $Y2=2.08
r72 22 24 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=0.247 $Y=0.865
+ $X2=0.247 $Y2=1.06
r73 19 32 9.37148 $w=2.45e-07 $l=1.9775e-07 $layer=LI1_cond $X=0.81 $Y=1.605
+ $X2=0.882 $Y2=1.44
r74 19 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.81 $Y=1.605
+ $X2=0.81 $Y2=1.935
r75 17 20 6.89401 $w=2.05e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.725 $Y=2.037
+ $X2=0.81 $Y2=1.935
r76 17 29 15.9601 $w=2.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.725 $Y=2.037
+ $X2=0.43 $Y2=2.037
r77 16 24 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.395 $Y=1.06
+ $X2=0.247 $Y2=1.06
r78 15 30 2.87745 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.725 $Y=1.06
+ $X2=0.882 $Y2=1.06
r79 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.725 $Y=1.06
+ $X2=0.395 $Y2=1.06
r80 13 36 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=1.005 $Y=2.4
+ $X2=1.005 $Y2=1.605
r81 9 35 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.97 $Y=0.74 $X2=0.97
+ $Y2=1.26
r82 2 27 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.265 $Y2=2.06
r83 1 22 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.69 $X2=0.265 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%A_209_74# 1 2 9 13 17 20 25 26 28 29
+ 30 31 41
c69 41 0 5.46905e-20 $X=1.23 $Y=2
c70 26 0 1.94125e-19 $X=1.83 $Y=1.44
c71 13 0 5.55505e-20 $X=1.975 $Y=2.05
r72 41 43 29.8172 $w=3.13e-07 $l=8.15e-07 $layer=LI1_cond $X=1.222 $Y=2
+ $X2=1.222 $Y2=2.815
r73 28 41 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=1.222 $Y=1.992
+ $X2=1.222 $Y2=2
r74 28 29 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=1.222 $Y=1.992
+ $X2=1.222 $Y2=1.835
r75 26 39 39.9775 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.44
+ $X2=1.865 $Y2=1.605
r76 26 38 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.44
+ $X2=1.865 $Y2=1.275
r77 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.44 $X2=1.83 $Y2=1.44
r78 23 31 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=1.46
+ $X2=1.295 $Y2=1.46
r79 23 25 17.8827 $w=2.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.38 $Y=1.46
+ $X2=1.83 $Y2=1.46
r80 21 31 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.295 $Y=1.605
+ $X2=1.295 $Y2=1.46
r81 21 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.295 $Y=1.605
+ $X2=1.295 $Y2=1.835
r82 20 31 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.295 $Y=1.315
+ $X2=1.295 $Y2=1.46
r83 20 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.295 $Y=1.315
+ $X2=1.295 $Y2=1.075
r84 15 30 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.235 $Y=0.93
+ $X2=1.235 $Y2=1.075
r85 15 17 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.235 $Y=0.93
+ $X2=1.235 $Y2=0.57
r86 13 39 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=1.975 $Y=2.05
+ $X2=1.975 $Y2=1.605
r87 9 38 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.92 $Y=0.9 $X2=1.92
+ $Y2=1.275
r88 2 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.815
r89 2 41 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2
r90 1 17 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%A_316_138# 1 2 9 13 15 17 19 20 22 29
+ 33
c69 33 0 3.02239e-19 $X=2.44 $Y=1.44
r70 33 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.44 $Y=1.44
+ $X2=2.44 $Y2=1.605
r71 33 35 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.44 $Y=1.44
+ $X2=2.44 $Y2=1.26
r72 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.44 $X2=2.44 $Y2=1.44
r73 27 29 4.97949 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.75 $Y=2.06
+ $X2=1.87 $Y2=2.06
r74 22 24 7.88514 $w=2.83e-07 $l=1.95e-07 $layer=LI1_cond $X=1.692 $Y=0.865
+ $X2=1.692 $Y2=1.06
r75 19 32 9.12826 $w=2.69e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.25 $Y=1.605
+ $X2=2.345 $Y2=1.44
r76 19 20 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.25 $Y=1.605
+ $X2=2.25 $Y2=1.895
r77 17 20 7.11011 $w=2.45e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.165 $Y=2.017
+ $X2=2.25 $Y2=1.895
r78 17 29 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=2.165 $Y=2.017
+ $X2=1.87 $Y2=2.017
r79 16 24 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.835 $Y=1.06
+ $X2=1.692 $Y2=1.06
r80 15 32 17.2342 $w=2.69e-07 $l=4.61302e-07 $layer=LI1_cond $X=2.165 $Y=1.06
+ $X2=2.345 $Y2=1.44
r81 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.165 $Y=1.06
+ $X2=1.835 $Y2=1.06
r82 13 36 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=2.49 $Y=2.4
+ $X2=2.49 $Y2=1.605
r83 9 35 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.41 $Y=0.74 $X2=2.41
+ $Y2=1.26
r84 2 27 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.84 $X2=1.75 $Y2=2.06
r85 1 22 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.69 $X2=1.705 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%A_497_74# 1 2 9 13 17 21 24 29 32 33
+ 42 45 46
c70 45 0 5.55505e-20 $X=2.715 $Y=2
c71 9 0 1.48579e-19 $X=3.36 $Y=0.9
r72 45 47 5.47606 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=2.685 $Y=2 $X2=2.685
+ $Y2=2.16
r73 45 46 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2
+ $X2=2.685 $Y2=1.835
r74 41 42 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.36 $Y=1.44 $X2=3.46
+ $Y2=1.44
r75 30 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.27 $Y=1.44 $X2=3.36
+ $Y2=1.44
r76 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.44 $X2=3.27 $Y2=1.44
r77 27 33 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.46
+ $X2=2.78 $Y2=1.46
r78 27 29 16.0945 $w=2.88e-07 $l=4.05e-07 $layer=LI1_cond $X=2.865 $Y=1.46
+ $X2=3.27 $Y2=1.46
r79 25 33 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.78 $Y=1.605
+ $X2=2.78 $Y2=1.46
r80 25 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.78 $Y=1.605
+ $X2=2.78 $Y2=1.835
r81 24 33 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.78 $Y=1.315
+ $X2=2.78 $Y2=1.46
r82 24 32 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.78 $Y=1.315
+ $X2=2.78 $Y2=1.075
r83 21 47 25.1617 $w=2.98e-07 $l=6.55e-07 $layer=LI1_cond $X=2.715 $Y=2.815
+ $X2=2.715 $Y2=2.16
r84 15 32 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=2.697 $Y=0.908
+ $X2=2.697 $Y2=1.075
r85 15 17 11.6276 $w=3.33e-07 $l=3.38e-07 $layer=LI1_cond $X=2.697 $Y=0.908
+ $X2=2.697 $Y2=0.57
r86 11 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.46 $Y=1.605
+ $X2=3.46 $Y2=1.44
r87 11 13 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=3.46 $Y=1.605
+ $X2=3.46 $Y2=2.05
r88 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=1.275
+ $X2=3.36 $Y2=1.44
r89 7 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.36 $Y=1.275
+ $X2=3.36 $Y2=0.9
r90 2 45 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.84 $X2=2.715 $Y2=2
r91 2 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.84 $X2=2.715 $Y2=2.815
r92 1 17 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.37 $X2=2.625 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%A_604_138# 1 2 9 13 17 19 20 21 22 24
+ 29
r66 29 32 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=1.44
+ $X2=3.925 $Y2=1.605
r67 29 31 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.925 $Y=1.44
+ $X2=3.925 $Y2=1.26
r68 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.44 $X2=3.925 $Y2=1.44
r69 24 25 20.2615 $w=2.83e-07 $l=4.7e-07 $layer=LI1_cond $X=3.235 $Y=2.06
+ $X2=3.705 $Y2=2.06
r70 22 25 2.77065 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=1.895
+ $X2=3.705 $Y2=2.06
r71 21 28 8.10771 $w=2.93e-07 $l=2.09893e-07 $layer=LI1_cond $X=3.705 $Y=1.605
+ $X2=3.807 $Y2=1.44
r72 21 22 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.705 $Y=1.605
+ $X2=3.705 $Y2=1.895
r73 19 28 15.8225 $w=2.93e-07 $l=4.70277e-07 $layer=LI1_cond $X=3.605 $Y=1.06
+ $X2=3.807 $Y2=1.44
r74 19 20 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.605 $Y=1.06
+ $X2=3.275 $Y2=1.06
r75 15 20 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=3.167 $Y=0.975
+ $X2=3.275 $Y2=1.06
r76 15 17 5.89622 $w=2.13e-07 $l=1.1e-07 $layer=LI1_cond $X=3.167 $Y=0.975
+ $X2=3.167 $Y2=0.865
r77 13 32 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=3.98 $Y=2.4
+ $X2=3.98 $Y2=1.605
r78 9 31 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.85 $Y=0.74 $X2=3.85
+ $Y2=1.26
r79 2 24 600 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=1.84 $X2=3.235 $Y2=2.06
r80 1 17 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.69 $X2=3.145 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%VPWR 1 2 3 12 16 20 22 24 29 34 41 42
+ 45 48 51 58
r49 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 49 58 0.0655027 $w=4.9e-07 $l=2.35e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.925 $Y2=3.33
r51 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r55 39 51 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=3.732 $Y2=3.33
r56 39 41 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 38 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 35 48 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.247 $Y2=3.33
r60 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 34 51 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=3.732 $Y2=3.33
r62 34 37 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.585 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 33 58 0.202083 $w=4.9e-07 $l=7.25e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.925 $Y2=3.33
r64 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 30 45 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.737 $Y2=3.33
r67 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 29 48 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.1 $Y=3.33
+ $X2=2.247 $Y2=3.33
r69 29 32 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 24 45 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.737 $Y2=3.33
r73 24 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 22 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 22 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 18 51 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.732 $Y=3.245
+ $X2=3.732 $Y2=3.33
r77 18 20 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=3.732 $Y=3.245
+ $X2=3.732 $Y2=2.475
r78 14 48 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.247 $Y=3.245
+ $X2=2.247 $Y2=3.33
r79 14 16 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=2.247 $Y=3.245
+ $X2=2.247 $Y2=2.475
r80 10 45 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=3.245
+ $X2=0.737 $Y2=3.33
r81 10 12 30.0807 $w=2.93e-07 $l=7.7e-07 $layer=LI1_cond $X=0.737 $Y=3.245
+ $X2=0.737 $Y2=2.475
r82 3 20 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=3.55
+ $Y=1.84 $X2=3.75 $Y2=2.475
r83 2 16 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=2.065
+ $Y=1.84 $X2=2.265 $Y2=2.475
r84 1 12 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%X 1 2 9 13 17 18 23 24 26 28 32
r52 28 32 1.20842 $w=1.7e-07 $l=1.255e-06 $layer=MET1_cond $X=3.845 $Y=2.405
+ $X2=2.59 $Y2=2.405
r53 23 27 5.41124 $w=3.73e-07 $l=1.6e-07 $layer=LI1_cond $X=4.162 $Y=2 $X2=4.162
+ $Y2=2.16
r54 23 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r55 23 24 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.162 $Y=2
+ $X2=4.162 $Y2=1.835
r56 18 28 0.0580243 $w=1.7e-07 $l=1.9e-07 $layer=MET1_cond $X=4.035 $Y=2.405
+ $X2=3.845 $Y2=2.405
r57 18 26 0.081654 $w=7.45e-07 $l=2.85e-07 $layer=MET1_cond $X=4.035 $Y=2.32
+ $X2=4.035 $Y2=2.035
r58 18 32 0.178133 $w=1.7e-07 $l=1.85e-07 $layer=MET1_cond $X=2.405 $Y=2.405
+ $X2=2.59 $Y2=2.405
r59 17 24 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.265 $Y=1.075
+ $X2=4.265 $Y2=1.835
r60 13 27 25.1617 $w=2.98e-07 $l=6.55e-07 $layer=LI1_cond $X=4.2 $Y=2.815
+ $X2=4.2 $Y2=2.16
r61 7 17 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=4.16 $Y=0.885
+ $X2=4.16 $Y2=1.075
r62 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.16 $Y=0.885
+ $X2=4.16 $Y2=0.57
r63 2 23 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=4.07
+ $Y=1.84 $X2=4.205 $Y2=2
r64 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.07
+ $Y=1.84 $X2=4.205 $Y2=2.815
r65 1 9 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=3.925
+ $Y=0.37 $X2=4.065 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__DLYMETAL6S6S_1%VGND 1 2 3 12 16 20 22 24 29 34 41 42
+ 45 48 51 58
c59 16 0 1.5366e-19 $X=2.195 $Y=0.72
r60 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 49 58 0.0655027 $w=4.9e-07 $l=2.35e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.925 $Y2=0
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 42 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r65 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.635
+ $Y2=0
r67 39 41 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=4.56
+ $Y2=0
r68 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.195
+ $Y2=0
r71 35 37 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=3.12
+ $Y2=0
r72 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.635
+ $Y2=0
r73 34 37 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.12
+ $Y2=0
r74 33 58 0.06829 $w=4.9e-07 $l=2.45e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.925
+ $Y2=0
r75 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r76 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r77 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=0.755
+ $Y2=0
r78 30 32 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=0.92 $Y=0 $X2=1.68
+ $Y2=0
r79 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.195
+ $Y2=0
r80 29 32 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.68
+ $Y2=0
r81 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r82 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.755
+ $Y2=0
r84 24 26 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.24
+ $Y2=0
r85 22 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r86 22 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r87 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0.085
+ $X2=3.635 $Y2=0
r88 18 20 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.635 $Y=0.085
+ $X2=3.635 $Y2=0.72
r89 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r90 14 16 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.72
r91 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r92 10 12 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.72
r93 3 20 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=3.435
+ $Y=0.69 $X2=3.635 $Y2=0.72
r94 2 16 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.69 $X2=2.195 $Y2=0.72
r95 1 12 182 $w=1.7e-07 $l=2.14476e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.69 $X2=0.755 $Y2=0.72
.ends


* NGSPICE file created from sky130_fd_sc_ms__mux2i_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
M1000 Y A1 a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=1.0767e+12p pd=1.031e+07u as=8.917e+11p ps=8.33e+06u
M1001 a_481_368# A0 Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.3104e+12p pd=1.13e+07u as=1.6576e+12p ps=1.416e+07u
M1002 VPWR a_1030_268# a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.387e+12p pd=1.732e+07u as=1.2992e+12p ps=1.128e+07u
M1003 a_481_368# S VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR S a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_114_85# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR S a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_475_85# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=8.806e+11p pd=8.3e+06u as=0p ps=0u
M1008 a_119_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_114_85# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.795e+12p ps=1.331e+07u
M1011 a_119_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_119_368# a_1030_268# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_475_85# a_1030_268# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_1030_268# a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A0 a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_114_85# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A0 a_481_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_481_368# A0 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1030_268# a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_119_368# a_1030_268# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_114_85# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A1 a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1030_268# S VGND VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1025 VGND S a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_1030_268# a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1030_268# S VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1028 VGND S a_114_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_475_85# a_1030_268# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y A0 a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A0 a_475_85# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_481_368# S VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR S a_1030_268# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_475_85# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


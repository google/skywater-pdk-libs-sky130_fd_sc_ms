* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_1333_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_861_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 Y A3 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_1333_368# A2 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_861_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 VPWR A1 a_1333_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 a_861_368# A2 a_1333_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X27 a_1333_368# A2 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 a_861_368# A2 a_1333_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 VPWR A1 a_1333_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X33 Y A3 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X34 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 a_1333_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X38 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__einvn_1.pxi.spice
* Created: Wed Sep  2 12:08:12 2020
* 
x_PM_SKY130_FD_SC_MS__EINVN_1%TE_B N_TE_B_M1004_g N_TE_B_c_44_n N_TE_B_M1005_g
+ N_TE_B_c_45_n N_TE_B_c_51_n N_TE_B_M1000_g TE_B N_TE_B_c_47_n N_TE_B_c_48_n
+ PM_SKY130_FD_SC_MS__EINVN_1%TE_B
x_PM_SKY130_FD_SC_MS__EINVN_1%A_22_46# N_A_22_46#_M1005_s N_A_22_46#_M1004_s
+ N_A_22_46#_c_91_n N_A_22_46#_c_92_n N_A_22_46#_M1002_g N_A_22_46#_c_93_n
+ N_A_22_46#_c_94_n N_A_22_46#_c_126_p N_A_22_46#_c_95_n N_A_22_46#_c_96_n
+ N_A_22_46#_c_99_n N_A_22_46#_c_97_n PM_SKY130_FD_SC_MS__EINVN_1%A_22_46#
x_PM_SKY130_FD_SC_MS__EINVN_1%A N_A_M1003_g N_A_M1001_g A N_A_c_136_n
+ N_A_c_137_n N_A_c_138_n PM_SKY130_FD_SC_MS__EINVN_1%A
x_PM_SKY130_FD_SC_MS__EINVN_1%VPWR N_VPWR_M1004_d N_VPWR_c_170_n VPWR
+ N_VPWR_c_171_n N_VPWR_c_172_n N_VPWR_c_169_n N_VPWR_c_174_n
+ PM_SKY130_FD_SC_MS__EINVN_1%VPWR
x_PM_SKY130_FD_SC_MS__EINVN_1%Z N_Z_M1003_d N_Z_M1001_d N_Z_c_195_n N_Z_c_193_n
+ N_Z_c_194_n Z Z PM_SKY130_FD_SC_MS__EINVN_1%Z
x_PM_SKY130_FD_SC_MS__EINVN_1%VGND N_VGND_M1005_d N_VGND_c_217_n VGND
+ N_VGND_c_218_n N_VGND_c_219_n N_VGND_c_220_n N_VGND_c_221_n
+ PM_SKY130_FD_SC_MS__EINVN_1%VGND
cc_1 VNB N_TE_B_c_44_n 0.019244f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.43
cc_2 VNB N_TE_B_c_45_n 0.0161612f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.685
cc_3 VNB TE_B 0.00343606f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_TE_B_c_47_n 0.0295513f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.595
cc_5 VNB N_TE_B_c_48_n 0.00549215f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.605
cc_6 VNB N_A_22_46#_c_91_n 0.0464381f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.685
cc_7 VNB N_A_22_46#_c_92_n 0.0137421f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.4
cc_8 VNB N_A_22_46#_c_93_n 0.0189997f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.595
cc_9 VNB N_A_22_46#_c_94_n 0.0201391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_22_46#_c_95_n 0.066973f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.595
cc_11 VNB N_A_22_46#_c_96_n 0.0247124f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.605
cc_12 VNB N_A_22_46#_c_97_n 0.0199392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_c_136_n 0.0311378f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.4
cc_14 VNB N_A_c_137_n 0.00786651f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.4
cc_15 VNB N_A_c_138_n 0.0207146f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.595
cc_16 VNB N_VPWR_c_169_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.595
cc_17 VNB N_Z_c_193_n 0.0228045f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.4
cc_18 VNB N_Z_c_194_n 0.0420195f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.595
cc_19 VNB N_VGND_c_217_n 0.0100327f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.11
cc_20 VNB N_VGND_c_218_n 0.0257484f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.4
cc_21 VNB N_VGND_c_219_n 0.0344986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_220_n 0.169809f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.595
cc_23 VNB N_VGND_c_221_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.595
cc_24 VPB N_TE_B_M1004_g 0.0276251f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=2.24
cc_25 VPB N_TE_B_c_45_n 0.0114606f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.685
cc_26 VPB N_TE_B_c_51_n 0.0188129f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.76
cc_27 VPB TE_B 0.00149535f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_28 VPB N_TE_B_c_47_n 0.0131742f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.595
cc_29 VPB N_TE_B_c_48_n 9.38834e-19 $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.605
cc_30 VPB N_A_22_46#_c_94_n 0.0140006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_A_22_46#_c_99_n 0.0460708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A_M1001_g 0.0261966f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.11
cc_33 VPB N_A_c_136_n 0.00567549f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=2.4
cc_34 VPB N_A_c_137_n 0.00617913f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=2.4
cc_35 VPB N_VPWR_c_170_n 0.0214828f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.11
cc_36 VPB N_VPWR_c_171_n 0.0304179f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=2.4
cc_37 VPB N_VPWR_c_172_n 0.0341405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_169_n 0.0784328f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.595
cc_39 VPB N_VPWR_c_174_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.595
cc_40 VPB N_Z_c_195_n 0.0146645f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=2.4
cc_41 VPB N_Z_c_193_n 0.0140507f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=2.4
cc_42 VPB Z 0.0400096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 N_TE_B_c_44_n N_A_22_46#_c_91_n 0.00493939f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_44 N_TE_B_c_44_n N_A_22_46#_c_92_n 0.0115742f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_45 N_TE_B_c_45_n N_A_22_46#_c_92_n 0.00997937f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_46 TE_B N_A_22_46#_c_92_n 0.00122005f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_47 N_TE_B_c_44_n N_A_22_46#_c_93_n 0.00482005f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_48 N_TE_B_M1004_g N_A_22_46#_c_94_n 0.00445973f $X=0.78 $Y=2.24 $X2=0 $Y2=0
cc_49 N_TE_B_c_44_n N_A_22_46#_c_94_n 0.00404556f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_50 N_TE_B_c_47_n N_A_22_46#_c_94_n 0.00227767f $X=0.895 $Y=1.595 $X2=0 $Y2=0
cc_51 N_TE_B_c_48_n N_A_22_46#_c_94_n 0.0256401f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_52 N_TE_B_c_44_n N_A_22_46#_c_96_n 0.00379808f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_53 N_TE_B_c_47_n N_A_22_46#_c_96_n 0.00675751f $X=0.895 $Y=1.595 $X2=0 $Y2=0
cc_54 N_TE_B_c_48_n N_A_22_46#_c_96_n 0.022249f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_55 N_TE_B_M1004_g N_A_22_46#_c_99_n 0.00972944f $X=0.78 $Y=2.24 $X2=0 $Y2=0
cc_56 N_TE_B_c_47_n N_A_22_46#_c_99_n 0.00514378f $X=0.895 $Y=1.595 $X2=0 $Y2=0
cc_57 N_TE_B_c_48_n N_A_22_46#_c_99_n 0.0173903f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_58 N_TE_B_c_44_n N_A_22_46#_c_97_n 0.0023126f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_59 N_TE_B_c_51_n N_A_M1001_g 0.0385618f $X=1.315 $Y=1.76 $X2=0 $Y2=0
cc_60 N_TE_B_c_45_n N_A_c_136_n 0.0385618f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_61 TE_B N_A_c_136_n 0.00130594f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_62 N_TE_B_c_44_n N_A_c_137_n 0.001417f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_63 N_TE_B_c_45_n N_A_c_137_n 0.00137165f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_64 TE_B N_A_c_137_n 0.0229496f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_65 N_TE_B_c_47_n N_A_c_137_n 5.88986e-19 $X=0.895 $Y=1.595 $X2=0 $Y2=0
cc_66 N_TE_B_M1004_g N_VPWR_c_170_n 0.00657963f $X=0.78 $Y=2.24 $X2=0 $Y2=0
cc_67 N_TE_B_c_45_n N_VPWR_c_170_n 0.00285467f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_68 N_TE_B_c_51_n N_VPWR_c_170_n 0.024249f $X=1.315 $Y=1.76 $X2=0 $Y2=0
cc_69 TE_B N_VPWR_c_170_n 0.0119134f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_70 N_TE_B_c_48_n N_VPWR_c_170_n 0.0119721f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_71 N_TE_B_M1004_g N_VPWR_c_171_n 0.00402065f $X=0.78 $Y=2.24 $X2=0 $Y2=0
cc_72 N_TE_B_c_51_n N_VPWR_c_172_n 0.00460063f $X=1.315 $Y=1.76 $X2=0 $Y2=0
cc_73 N_TE_B_M1004_g N_VPWR_c_169_n 0.00517376f $X=0.78 $Y=2.24 $X2=0 $Y2=0
cc_74 N_TE_B_c_51_n N_VPWR_c_169_n 0.00908371f $X=1.315 $Y=1.76 $X2=0 $Y2=0
cc_75 N_TE_B_c_51_n N_Z_c_195_n 0.00305188f $X=1.315 $Y=1.76 $X2=0 $Y2=0
cc_76 N_TE_B_c_44_n N_VGND_c_217_n 0.00300331f $X=0.82 $Y=1.43 $X2=0 $Y2=0
cc_77 N_TE_B_c_45_n N_VGND_c_217_n 0.00160902f $X=1.225 $Y=1.685 $X2=0 $Y2=0
cc_78 N_TE_B_c_48_n N_VGND_c_217_n 0.0285478f $X=1.085 $Y=1.605 $X2=0 $Y2=0
cc_79 N_A_22_46#_c_92_n N_A_c_136_n 0.0253488f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_80 N_A_22_46#_c_92_n N_A_c_137_n 4.88499e-19 $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_81 N_A_22_46#_c_91_n N_A_c_138_n 0.0253488f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_82 N_A_22_46#_c_99_n N_VPWR_c_170_n 0.0161981f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_83 N_A_22_46#_c_99_n N_VPWR_c_171_n 0.00510886f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_84 N_A_22_46#_c_99_n N_VPWR_c_169_n 0.00894968f $X=0.555 $Y=2.075 $X2=0 $Y2=0
cc_85 N_A_22_46#_c_92_n N_Z_c_194_n 0.0019742f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_86 N_A_22_46#_c_91_n N_VGND_c_217_n 0.0256607f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_87 N_A_22_46#_c_92_n N_VGND_c_217_n 0.016172f $X=1.33 $Y=0.425 $X2=0 $Y2=0
cc_88 N_A_22_46#_c_93_n N_VGND_c_217_n 0.0419197f $X=0.44 $Y=0.92 $X2=0 $Y2=0
cc_89 N_A_22_46#_c_126_p N_VGND_c_217_n 0.0248316f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_90 N_A_22_46#_c_97_n N_VGND_c_217_n 0.00277657f $X=0.78 $Y=0.395 $X2=0 $Y2=0
cc_91 N_A_22_46#_c_91_n N_VGND_c_218_n 0.00502076f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_92 N_A_22_46#_c_126_p N_VGND_c_218_n 0.0454726f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_93 N_A_22_46#_c_95_n N_VGND_c_218_n 0.0116198f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_94 N_A_22_46#_c_91_n N_VGND_c_219_n 0.0045897f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_95 N_A_22_46#_c_91_n N_VGND_c_220_n 0.0093352f $X=1.255 $Y=0.35 $X2=0 $Y2=0
cc_96 N_A_22_46#_c_126_p N_VGND_c_220_n 0.0228727f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_97 N_A_22_46#_c_95_n N_VGND_c_220_n 0.0114391f $X=0.615 $Y=0.395 $X2=0 $Y2=0
cc_98 N_A_22_46#_c_97_n N_VGND_c_220_n 0.00394079f $X=0.78 $Y=0.395 $X2=0 $Y2=0
cc_99 N_A_M1001_g N_VPWR_c_170_n 0.00342385f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_M1001_g N_VPWR_c_172_n 0.0048691f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_M1001_g N_VPWR_c_169_n 0.00877303f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_M1001_g N_Z_c_195_n 0.00635975f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_c_136_n N_Z_c_195_n 7.74224e-19 $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A_c_137_n N_Z_c_195_n 0.0154469f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A_M1001_g N_Z_c_193_n 0.00316404f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_c_136_n N_Z_c_193_n 0.00739878f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A_c_137_n N_Z_c_193_n 0.0332868f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_c_138_n N_Z_c_193_n 0.00337861f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_c_136_n N_Z_c_194_n 0.0012388f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A_c_137_n N_Z_c_194_n 0.0145144f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A_c_138_n N_Z_c_194_n 0.0126824f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_112 N_A_M1001_g Z 0.0161483f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_c_138_n N_VGND_c_217_n 0.00292024f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_114 N_A_c_138_n N_VGND_c_219_n 0.00467453f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_115 N_A_c_138_n N_VGND_c_220_n 0.00505379f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_116 N_VPWR_c_170_n N_Z_c_195_n 0.0327712f $X=1.09 $Y=2.115 $X2=0 $Y2=0
cc_117 N_VPWR_c_172_n Z 0.0242759f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_118 N_VPWR_c_169_n Z 0.0199549f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_119 N_Z_c_194_n N_VGND_c_217_n 0.0230605f $X=1.935 $Y=0.645 $X2=0 $Y2=0
cc_120 N_Z_c_194_n N_VGND_c_219_n 0.0157999f $X=1.935 $Y=0.645 $X2=0 $Y2=0
cc_121 N_Z_c_194_n N_VGND_c_220_n 0.0184123f $X=1.935 $Y=0.645 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__inv_16.pex.spice
* Created: Wed Sep  2 12:10:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__INV_16%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 129 133 135 137 140
+ 148 155 161 167 174 181 219 227
c337 91 0 1.79483e-19 $X=5.575 $Y=0.74
c338 75 0 1.75317e-19 $X=4.645 $Y=0.74
r339 214 219 0.638396 $w=2.3e-07 $l=9.95e-07 $layer=MET1_cond $X=5.93 $Y=1.665
+ $X2=6.925 $Y2=1.665
r340 209 214 0.638396 $w=2.3e-07 $l=9.95e-07 $layer=MET1_cond $X=4.935 $Y=1.665
+ $X2=5.93 $Y2=1.665
r341 209 227 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=4.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r342 194 199 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=2.17 $Y=1.665
+ $X2=3.11 $Y2=1.665
r343 189 194 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=1.23 $Y=1.665
+ $X2=2.17 $Y2=1.665
r344 184 185 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.575 $Y=1.515
+ $X2=6.655 $Y2=1.515
r345 183 184 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=6.205 $Y=1.515
+ $X2=6.575 $Y2=1.515
r346 182 183 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.145 $Y=1.515
+ $X2=6.205 $Y2=1.515
r347 181 214 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.93 $Y=1.665
+ $X2=5.93 $Y2=1.665
r348 180 182 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.93 $Y=1.515
+ $X2=6.145 $Y2=1.515
r349 180 181 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.93
+ $Y=1.515 $X2=5.93 $Y2=1.515
r350 178 180 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=5.655 $Y=1.515
+ $X2=5.93 $Y2=1.515
r351 177 178 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.575 $Y=1.515
+ $X2=5.655 $Y2=1.515
r352 176 177 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=5.175 $Y=1.515
+ $X2=5.575 $Y2=1.515
r353 175 176 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.145 $Y=1.515
+ $X2=5.175 $Y2=1.515
r354 174 209 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.935 $Y=1.665
+ $X2=4.935 $Y2=1.665
r355 173 175 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.935 $Y=1.515
+ $X2=5.145 $Y2=1.515
r356 173 174 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.515 $X2=4.935 $Y2=1.515
r357 171 173 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=4.705 $Y=1.515
+ $X2=4.935 $Y2=1.515
r358 170 171 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.645 $Y=1.515
+ $X2=4.705 $Y2=1.515
r359 169 170 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.255 $Y=1.515
+ $X2=4.645 $Y2=1.515
r360 168 169 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.215 $Y=1.515
+ $X2=4.255 $Y2=1.515
r361 166 168 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.025 $Y=1.515
+ $X2=4.215 $Y2=1.515
r362 166 167 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.515 $X2=4.025 $Y2=1.515
r363 164 166 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.805 $Y=1.515
+ $X2=4.025 $Y2=1.515
r364 163 164 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.785 $Y=1.515
+ $X2=3.805 $Y2=1.515
r365 162 163 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.355 $Y=1.515
+ $X2=3.785 $Y2=1.515
r366 161 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.11 $Y=1.665
+ $X2=3.11 $Y2=1.665
r367 160 162 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=3.11 $Y=1.515
+ $X2=3.355 $Y2=1.515
r368 160 161 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.515 $X2=3.11 $Y2=1.515
r369 158 160 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=2.855 $Y=1.515
+ $X2=3.11 $Y2=1.515
r370 157 158 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.425 $Y=1.515
+ $X2=2.855 $Y2=1.515
r371 156 157 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.405 $Y=1.515
+ $X2=2.425 $Y2=1.515
r372 155 194 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=1.665
r373 154 156 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.17 $Y=1.515
+ $X2=2.405 $Y2=1.515
r374 154 155 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.515 $X2=2.17 $Y2=1.515
r375 152 154 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.925 $Y=1.515
+ $X2=2.17 $Y2=1.515
r376 151 152 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.905 $Y=1.515
+ $X2=1.925 $Y2=1.515
r377 150 151 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.495 $Y=1.515
+ $X2=1.905 $Y2=1.515
r378 149 150 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.455 $Y=1.515
+ $X2=1.495 $Y2=1.515
r379 148 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=1.665
r380 147 149 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.23 $Y=1.515
+ $X2=1.455 $Y2=1.515
r381 147 148 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.515 $X2=1.23 $Y2=1.515
r382 145 147 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.995 $Y=1.515
+ $X2=1.23 $Y2=1.515
r383 144 145 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.515
+ $X2=0.995 $Y2=1.515
r384 143 144 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=0.565 $Y=1.515
+ $X2=0.955 $Y2=1.515
r385 141 143 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.565 $Y2=1.515
r386 140 219 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.925 $Y=1.665
+ $X2=6.925 $Y2=1.665
r387 139 140 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.925
+ $Y=1.515 $X2=6.925 $Y2=1.515
r388 137 185 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.745 $Y=1.515
+ $X2=6.655 $Y2=1.515
r389 137 139 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.745 $Y=1.515
+ $X2=6.925 $Y2=1.515
r390 135 227 0.0352882 $w=2.3e-07 $l=5.5e-08 $layer=MET1_cond $X=4.025 $Y=1.665
+ $X2=4.08 $Y2=1.665
r391 135 199 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=4.025 $Y=1.665
+ $X2=3.11 $Y2=1.665
r392 135 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.025 $Y=1.665
+ $X2=4.025 $Y2=1.665
r393 132 133 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=7.595 $Y=1.515
+ $X2=7.655 $Y2=1.515
r394 131 132 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=7.205 $Y=1.515
+ $X2=7.595 $Y2=1.515
r395 130 131 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=7.165 $Y=1.515
+ $X2=7.205 $Y2=1.515
r396 129 139 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.515
+ $X2=6.925 $Y2=1.515
r397 129 130 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.09 $Y=1.515
+ $X2=7.165 $Y2=1.515
r398 125 133 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.68
+ $X2=7.655 $Y2=1.515
r399 125 127 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.655 $Y=1.68
+ $X2=7.655 $Y2=2.4
r400 121 132 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.595 $Y=1.35
+ $X2=7.595 $Y2=1.515
r401 121 123 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.595 $Y=1.35
+ $X2=7.595 $Y2=0.74
r402 117 131 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=1.68
+ $X2=7.205 $Y2=1.515
r403 117 119 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.205 $Y=1.68
+ $X2=7.205 $Y2=2.4
r404 113 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.35
+ $X2=7.165 $Y2=1.515
r405 113 115 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.165 $Y=1.35
+ $X2=7.165 $Y2=0.74
r406 109 185 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.655 $Y=1.68
+ $X2=6.655 $Y2=1.515
r407 109 111 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.655 $Y=1.68
+ $X2=6.655 $Y2=2.4
r408 105 184 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.575 $Y=1.35
+ $X2=6.575 $Y2=1.515
r409 105 107 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.575 $Y=1.35
+ $X2=6.575 $Y2=0.74
r410 101 183 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.68
+ $X2=6.205 $Y2=1.515
r411 101 103 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.205 $Y=1.68
+ $X2=6.205 $Y2=2.4
r412 97 182 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.145 $Y=1.35
+ $X2=6.145 $Y2=1.515
r413 97 99 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.145 $Y=1.35
+ $X2=6.145 $Y2=0.74
r414 93 178 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.68
+ $X2=5.655 $Y2=1.515
r415 93 95 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.655 $Y=1.68
+ $X2=5.655 $Y2=2.4
r416 89 177 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.35
+ $X2=5.575 $Y2=1.515
r417 89 91 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.575 $Y=1.35
+ $X2=5.575 $Y2=0.74
r418 85 176 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.68
+ $X2=5.175 $Y2=1.515
r419 85 87 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.175 $Y=1.68
+ $X2=5.175 $Y2=2.4
r420 81 175 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.35
+ $X2=5.145 $Y2=1.515
r421 81 83 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.145 $Y=1.35
+ $X2=5.145 $Y2=0.74
r422 77 171 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.68
+ $X2=4.705 $Y2=1.515
r423 77 79 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.705 $Y=1.68
+ $X2=4.705 $Y2=2.4
r424 73 170 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.645 $Y=1.35
+ $X2=4.645 $Y2=1.515
r425 73 75 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.645 $Y=1.35
+ $X2=4.645 $Y2=0.74
r426 69 169 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=1.68
+ $X2=4.255 $Y2=1.515
r427 69 71 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.255 $Y=1.68
+ $X2=4.255 $Y2=2.4
r428 65 168 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.215 $Y=1.35
+ $X2=4.215 $Y2=1.515
r429 65 67 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.215 $Y=1.35
+ $X2=4.215 $Y2=0.74
r430 61 164 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.68
+ $X2=3.805 $Y2=1.515
r431 61 63 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.805 $Y=1.68
+ $X2=3.805 $Y2=2.4
r432 57 163 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.35
+ $X2=3.785 $Y2=1.515
r433 57 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.785 $Y=1.35
+ $X2=3.785 $Y2=0.74
r434 53 162 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=1.515
r435 53 55 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=0.74
r436 49 162 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.68
+ $X2=3.355 $Y2=1.515
r437 49 51 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.355 $Y=1.68
+ $X2=3.355 $Y2=2.4
r438 45 158 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=1.515
r439 45 47 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=0.74
r440 41 158 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.855 $Y2=1.515
r441 41 43 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.855 $Y2=2.4
r442 37 157 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=1.515
r443 37 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=0.74
r444 33 156 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=1.515
r445 33 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=2.4
r446 29 152 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.515
r447 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.74
r448 25 151 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=1.515
r449 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=2.4
r450 21 150 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.515
r451 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r452 17 149 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.515
r453 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r454 13 145 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r455 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r456 9 144 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.515
r457 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r458 5 143 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=1.515
r459 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.565 $Y=1.35
+ $X2=0.565 $Y2=0.74
r460 1 141 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.515
r461 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__INV_16%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 42 48 54 60
+ 66 72 76 78 83 84 86 87 88 90 95 100 112 116 121 130 133 136 139 142 146
r147 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r150 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r151 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r154 125 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r155 125 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r156 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 122 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=6.93 $Y2=3.33
r158 122 124 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=7.44 $Y2=3.33
r159 121 145 4.55093 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.947 $Y2=3.33
r160 121 124 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.44 $Y2=3.33
r161 120 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r162 120 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r163 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r164 117 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=5.93 $Y2=3.33
r165 117 119 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.48 $Y2=3.33
r166 116 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.93 $Y2=3.33
r167 116 119 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 115 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r169 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r170 112 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.93 $Y2=3.33
r171 112 114 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.52 $Y2=3.33
r172 111 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r173 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r174 108 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r175 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r176 105 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.12 $Y2=3.33
r177 105 107 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.6 $Y2=3.33
r178 104 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r179 104 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r181 101 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.17 $Y2=3.33
r182 101 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r183 100 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.12 $Y2=3.33
r184 100 103 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r185 99 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r186 99 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r187 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r188 96 130 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.2 $Y2=3.33
r189 96 98 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 95 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.17 $Y2=3.33
r191 95 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r192 94 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 94 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r194 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 91 127 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r196 91 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r197 90 130 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 90 93 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r199 88 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r200 88 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r201 86 110 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.81 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 86 87 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.81 $Y=3.33
+ $X2=4.952 $Y2=3.33
r203 85 114 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=5.52 $Y2=3.33
r204 85 87 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=4.952 $Y2=3.33
r205 83 107 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 83 84 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=4.032 $Y2=3.33
r207 82 110 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.56 $Y2=3.33
r208 82 84 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.032 $Y2=3.33
r209 78 81 30.8557 $w=3.08e-07 $l=8.3e-07 $layer=LI1_cond $X=7.89 $Y=1.985
+ $X2=7.89 $Y2=2.815
r210 76 145 3.04826 $w=3.1e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.947 $Y2=3.33
r211 76 81 15.9855 $w=3.08e-07 $l=4.3e-07 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.89 $Y2=2.815
r212 72 75 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.93 $Y=2.105
+ $X2=6.93 $Y2=2.815
r213 70 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=3.33
r214 70 75 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.93 $Y=3.245
+ $X2=6.93 $Y2=2.815
r215 66 69 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.93 $Y=2.105
+ $X2=5.93 $Y2=2.815
r216 64 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=3.245
+ $X2=5.93 $Y2=3.33
r217 64 69 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.93 $Y=3.245
+ $X2=5.93 $Y2=2.815
r218 60 63 28.71 $w=2.83e-07 $l=7.1e-07 $layer=LI1_cond $X=4.952 $Y=2.105
+ $X2=4.952 $Y2=2.815
r219 58 87 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.952 $Y=3.245
+ $X2=4.952 $Y2=3.33
r220 58 63 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=4.952 $Y=3.245
+ $X2=4.952 $Y2=2.815
r221 54 57 34.8185 $w=2.33e-07 $l=7.1e-07 $layer=LI1_cond $X=4.032 $Y=2.105
+ $X2=4.032 $Y2=2.815
r222 52 84 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.032 $Y=3.245
+ $X2=4.032 $Y2=3.33
r223 52 57 21.0873 $w=2.33e-07 $l=4.3e-07 $layer=LI1_cond $X=4.032 $Y=3.245
+ $X2=4.032 $Y2=2.815
r224 48 51 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=3.12 $Y=2.105
+ $X2=3.12 $Y2=2.815
r225 46 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=3.33
r226 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.12 $Y2=2.815
r227 42 45 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.17 $Y=2.105
+ $X2=2.17 $Y2=2.815
r228 40 133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r229 40 45 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.815
r230 36 39 28.215 $w=2.88e-07 $l=7.1e-07 $layer=LI1_cond $X=1.2 $Y=2.105 $X2=1.2
+ $Y2=2.815
r231 34 130 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245
+ $X2=1.2 $Y2=3.33
r232 34 39 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=3.245
+ $X2=1.2 $Y2=2.815
r233 30 33 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r234 28 127 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r235 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r236 9 81 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=2.815
r237 9 78 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=1.985
r238 8 75 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.93 $Y2=2.815
r239 8 72 400 $w=1.7e-07 $l=3.45326e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.93 $Y2=2.105
r240 7 69 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.84 $X2=5.93 $Y2=2.815
r241 7 66 400 $w=1.7e-07 $l=3.45326e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.84 $X2=5.93 $Y2=2.105
r242 6 63 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.84 $X2=4.93 $Y2=2.815
r243 6 60 400 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.84 $X2=4.93 $Y2=2.105
r244 5 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.84 $X2=4.03 $Y2=2.815
r245 5 54 400 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.84 $X2=4.03 $Y2=2.105
r246 4 51 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.815
r247 4 48 400 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.105
r248 3 45 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.84 $X2=2.13 $Y2=2.815
r249 3 42 400 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.84 $X2=2.13 $Y2=2.105
r250 2 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r251 2 36 400 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.105
r252 1 33 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r253 1 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__INV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 51
+ 57 61 65 69 73 77 79 81 83 85 89 91 92 93 97 98 101 108 118 125 132 134 139
+ 144 149
c248 91 0 1.71499e-19 $X=0.725 $Y=1.49
c249 83 0 1.79483e-19 $X=6.36 $Y=1.015
c250 79 0 1.75317e-19 $X=5.37 $Y=1.025
r251 149 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.48 $Y=2.035
+ $X2=4.48 $Y2=2.035
r252 149 150 1.98543 $w=2.88e-07 $l=4.5e-08 $layer=LI1_cond $X=4.485 $Y=1.985
+ $X2=4.485 $Y2=1.94
r253 144 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.63 $Y=2.035
+ $X2=2.63 $Y2=2.035
r254 144 145 1.62839 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.63 $Y=1.985
+ $X2=2.63 $Y2=1.94
r255 142 147 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=1.68 $Y=2.035
+ $X2=2.63 $Y2=2.035
r256 139 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.035
r257 139 140 3.16711 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.025
+ $X2=1.68 $Y2=1.94
r258 132 136 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=7.405 $Y=1.985
+ $X2=7.405 $Y2=2.815
r259 132 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.43 $Y=2.035
+ $X2=7.43 $Y2=2.035
r260 127 134 0.641604 $w=2.3e-07 $l=1e-06 $layer=MET1_cond $X=6.43 $Y=2.035
+ $X2=7.43 $Y2=2.035
r261 125 129 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.43 $Y=1.985
+ $X2=6.43 $Y2=2.815
r262 125 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.43 $Y=2.035
+ $X2=6.43 $Y2=2.035
r263 120 127 0.641604 $w=2.3e-07 $l=1e-06 $layer=MET1_cond $X=5.43 $Y=2.035
+ $X2=6.43 $Y2=2.035
r264 120 152 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=5.43 $Y=2.035
+ $X2=4.48 $Y2=2.035
r265 118 122 30.366 $w=3.13e-07 $l=8.3e-07 $layer=LI1_cond $X=5.422 $Y=1.985
+ $X2=5.422 $Y2=2.815
r266 118 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.43 $Y=2.035
+ $X2=5.43 $Y2=2.035
r267 113 147 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=3.58 $Y=2.035
+ $X2=2.63 $Y2=2.035
r268 111 115 32.4247 $w=2.93e-07 $l=8.3e-07 $layer=LI1_cond $X=3.562 $Y=1.985
+ $X2=3.562 $Y2=2.815
r269 111 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.58 $Y=2.035
+ $X2=3.58 $Y2=2.035
r270 108 111 57.4268 $w=2.93e-07 $l=1.47e-06 $layer=LI1_cond $X=3.562 $Y=0.515
+ $X2=3.562 $Y2=1.985
r271 103 142 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=0.73 $Y=2.035
+ $X2=1.68 $Y2=2.035
r272 101 105 29.8915 $w=3.18e-07 $l=8.3e-07 $layer=LI1_cond $X=0.725 $Y=1.985
+ $X2=0.725 $Y2=2.815
r273 101 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=2.035
+ $X2=0.73 $Y2=2.035
r274 98 152 0.256642 $w=2.3e-07 $l=4e-07 $layer=MET1_cond $X=4.08 $Y=2.035
+ $X2=4.48 $Y2=2.035
r275 98 113 0.320802 $w=2.3e-07 $l=5e-07 $layer=MET1_cond $X=4.08 $Y=2.035
+ $X2=3.58 $Y2=2.035
r276 97 132 35.1907 $w=2.78e-07 $l=8.55e-07 $layer=LI1_cond $X=7.405 $Y=1.13
+ $X2=7.405 $Y2=1.985
r277 95 125 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=6.43 $Y=1.45
+ $X2=6.43 $Y2=1.985
r278 94 118 19.8659 $w=3.13e-07 $l=5.43e-07 $layer=LI1_cond $X=5.422 $Y=1.442
+ $X2=5.422 $Y2=1.985
r279 92 93 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=0.75 $Y=1.33 $X2=0.75
+ $Y2=1.13
r280 91 101 17.8269 $w=3.18e-07 $l=4.95e-07 $layer=LI1_cond $X=0.725 $Y=1.49
+ $X2=0.725 $Y2=1.985
r281 91 92 6.07707 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.725 $Y=1.49
+ $X2=0.725 $Y2=1.33
r282 87 97 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=0.965
+ $X2=7.38 $Y2=1.13
r283 87 89 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.38 $Y=0.965
+ $X2=7.38 $Y2=0.515
r284 83 95 16.9553 $w=3.13e-07 $l=4.68695e-07 $layer=LI1_cond $X=6.36 $Y=1.015
+ $X2=6.43 $Y2=1.45
r285 83 85 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.36 $Y=1.015
+ $X2=6.36 $Y2=0.515
r286 79 94 17.0147 $w=2.99e-07 $l=4.42236e-07 $layer=LI1_cond $X=5.37 $Y=1.025
+ $X2=5.422 $Y2=1.442
r287 79 81 18.9595 $w=3.08e-07 $l=5.1e-07 $layer=LI1_cond $X=5.37 $Y=1.025
+ $X2=5.37 $Y2=0.515
r288 75 149 3.97394 $w=2.88e-07 $l=1e-07 $layer=LI1_cond $X=4.485 $Y=2.085
+ $X2=4.485 $Y2=1.985
r289 75 77 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=4.485 $Y=2.085
+ $X2=4.485 $Y2=2.4
r290 73 150 64.4012 $w=2.53e-07 $l=1.425e-06 $layer=LI1_cond $X=4.467 $Y=0.515
+ $X2=4.467 $Y2=1.94
r291 69 145 52.9752 $w=3.08e-07 $l=1.425e-06 $layer=LI1_cond $X=2.64 $Y=0.515
+ $X2=2.64 $Y2=1.94
r292 63 144 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.63 $Y=2.105
+ $X2=2.63 $Y2=1.985
r293 63 65 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.63 $Y=2.105
+ $X2=2.63 $Y2=2.815
r294 61 140 56.6287 $w=2.88e-07 $l=1.425e-06 $layer=LI1_cond $X=1.7 $Y=0.515
+ $X2=1.7 $Y2=1.94
r295 55 139 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=2.105
+ $X2=1.68 $Y2=2.025
r296 55 57 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.68 $Y=2.105
+ $X2=1.68 $Y2=2.815
r297 49 93 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=1.13
r298 49 51 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=0.515
r299 16 136 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.43 $Y2=2.815
r300 16 132 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.84 $X2=7.43 $Y2=1.985
r301 15 129 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.815
r302 15 125 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=1.985
r303 14 122 400 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.84 $X2=5.43 $Y2=2.815
r304 14 118 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.84 $X2=5.43 $Y2=1.985
r305 13 149 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.84 $X2=4.48 $Y2=1.985
r306 13 77 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.84 $X2=4.48 $Y2=2.4
r307 12 115 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.58 $Y2=2.815
r308 12 111 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.58 $Y2=1.985
r309 11 144 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=1.985
r310 11 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.815
r311 10 139 400 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.025
r312 10 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.815
r313 9 105 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r314 9 101 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r315 8 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.37 $X2=7.38 $Y2=0.515
r316 7 85 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.22
+ $Y=0.37 $X2=6.36 $Y2=0.515
r317 6 81 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.37 $X2=5.36 $Y2=0.515
r318 5 73 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.29
+ $Y=0.37 $X2=4.43 $Y2=0.515
r319 4 108 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.37 $X2=3.57 $Y2=0.515
r320 3 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.5
+ $Y=0.37 $X2=2.64 $Y2=0.515
r321 2 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.71 $Y2=0.515
r322 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__INV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 58 60 62 65 66 68 69 71 72 73 75 80 85 100 104 113 116 119 122 126
r136 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r137 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r138 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r139 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r140 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r141 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r142 108 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r143 108 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r144 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r145 105 122 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=6.875 $Y2=0
r146 105 107 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=7.44 $Y2=0
r147 104 125 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.937 $Y2=0
r148 104 107 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.44 $Y2=0
r149 103 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r150 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r151 100 122 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.875 $Y2=0
r152 100 102 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.48 $Y2=0
r153 99 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r154 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r155 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r156 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r157 93 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r158 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r159 90 119 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.245 $Y=0
+ $X2=3.11 $Y2=0
r160 90 92 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.6
+ $Y2=0
r161 89 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r162 89 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r163 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r164 86 116 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.165
+ $Y2=0
r165 86 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.64 $Y2=0
r166 85 119 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=3.11 $Y2=0
r167 85 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0
+ $X2=2.64 $Y2=0
r168 84 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r169 84 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r170 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r171 81 113 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.245 $Y2=0
r172 81 83 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r173 80 116 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.165
+ $Y2=0
r174 80 83 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.68
+ $Y2=0
r175 79 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r176 79 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r177 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r178 76 110 4.01078 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r179 76 78 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r180 75 113 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=1.245 $Y2=0
r181 75 78 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r182 73 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r183 73 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r184 71 98 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.705 $Y=0
+ $X2=5.52 $Y2=0
r185 71 72 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=5.865
+ $Y2=0
r186 70 102 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.025 $Y=0
+ $X2=6.48 $Y2=0
r187 70 72 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.025 $Y=0 $X2=5.865
+ $Y2=0
r188 68 95 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r189 68 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.895
+ $Y2=0
r190 67 98 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=5.52 $Y2=0
r191 67 69 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.025 $Y=0 $X2=4.895
+ $Y2=0
r192 65 92 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.6
+ $Y2=0
r193 65 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.02
+ $Y2=0
r194 64 95 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.15 $Y=0 $X2=4.56
+ $Y2=0
r195 64 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.15 $Y=0 $X2=4.02
+ $Y2=0
r196 60 125 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.937 $Y2=0
r197 60 62 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.515
r198 56 122 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=0.085
+ $X2=6.875 $Y2=0
r199 56 58 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=6.875 $Y=0.085
+ $X2=6.875 $Y2=0.53
r200 52 72 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.865 $Y=0.085
+ $X2=5.865 $Y2=0
r201 52 54 16.0262 $w=3.18e-07 $l=4.45e-07 $layer=LI1_cond $X=5.865 $Y=0.085
+ $X2=5.865 $Y2=0.53
r202 48 69 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0.085
+ $X2=4.895 $Y2=0
r203 48 50 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=4.895 $Y=0.085
+ $X2=4.895 $Y2=0.53
r204 44 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r205 44 46 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.515
r206 40 119 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0
r207 40 42 18.3537 $w=2.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0.515
r208 36 116 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r209 36 38 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.515
r210 32 113 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r211 32 34 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.515
r212 28 110 3.20143 $w=2.6e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.222 $Y2=0
r213 28 30 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.315 $Y2=0.515
r214 9 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.67
+ $Y=0.37 $X2=7.81 $Y2=0.515
r215 8 58 91 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=2 $X=6.65
+ $Y=0.37 $X2=6.87 $Y2=0.53
r216 7 54 91 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=2 $X=5.65
+ $Y=0.37 $X2=5.86 $Y2=0.53
r217 6 50 91 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_NDIFF $count=2 $X=4.72
+ $Y=0.37 $X2=4.895 $Y2=0.53
r218 5 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.37 $X2=4 $Y2=0.515
r219 4 42 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.93
+ $Y=0.37 $X2=3.12 $Y2=0.515
r220 3 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r221 2 34 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r222 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends


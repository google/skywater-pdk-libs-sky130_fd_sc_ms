* File: sky130_fd_sc_ms__or3b_2.pex.spice
* Created: Fri Aug 28 18:08:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR3B_2%C_N 1 3 6 8 12
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r26 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r27 4 11 39.4323 $w=3.92e-07 $l=2.62857e-07 $layer=POLY_cond $X=0.565 $Y=1.3
+ $X2=0.372 $Y2=1.465
r28 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.565 $Y=1.3
+ $X2=0.565 $Y2=0.835
r29 1 11 52.9661 $w=3.92e-07 $l=3.75659e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.372 $Y2=1.465
r30 1 3 128.533 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%A_190_260# 1 2 3 12 16 18 22 26 28 29 30 33
+ 35 39 47 49 50 52
r114 49 50 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.375
+ $X2=3.495 $Y2=2.29
r115 46 56 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.567 $Y=1.465
+ $X2=1.567 $Y2=1.63
r116 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.465 $X2=1.57 $Y2=1.465
r117 41 52 3.27229 $w=2.87e-07 $l=1.54771e-07 $layer=LI1_cond $X=3.67 $Y=1.18
+ $X2=3.552 $Y2=1.095
r118 41 50 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.67 $Y=1.18
+ $X2=3.67 $Y2=2.29
r119 37 52 3.27229 $w=2.87e-07 $l=8.5e-08 $layer=LI1_cond $X=3.552 $Y=1.01
+ $X2=3.552 $Y2=1.095
r120 37 39 11.2399 $w=4.03e-07 $l=3.95e-07 $layer=LI1_cond $X=3.552 $Y=1.01
+ $X2=3.552 $Y2=0.615
r121 36 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=1.095
+ $X2=2.515 $Y2=1.095
r122 35 52 3.2872 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=3.35 $Y=1.095
+ $X2=3.552 $Y2=1.095
r123 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.35 $Y=1.095
+ $X2=2.68 $Y2=1.095
r124 31 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.515 $Y2=1.095
r125 31 33 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.515 $Y2=0.615
r126 30 45 15.7282 $w=2.87e-07 $l=4.5722e-07 $layer=LI1_cond $X=1.795 $Y=1.095
+ $X2=1.6 $Y2=1.465
r127 29 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=2.515 $Y2=1.095
r128 29 30 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.35 $Y=1.095
+ $X2=1.795 $Y2=1.095
r129 26 54 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.505 $Y=0.74
+ $X2=1.505 $Y2=1.3
r130 22 56 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.49 $Y=2.4
+ $X2=1.49 $Y2=1.63
r131 19 28 6.66866 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.15 $Y=1.375
+ $X2=1.05 $Y2=1.375
r132 18 46 15.5026 $w=3.35e-07 $l=9e-08 $layer=POLY_cond $X=1.567 $Y=1.375
+ $X2=1.567 $Y2=1.465
r133 18 54 30.7523 $w=3.35e-07 $l=7.5e-08 $layer=POLY_cond $X=1.567 $Y=1.375
+ $X2=1.567 $Y2=1.3
r134 18 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.4 $Y=1.375
+ $X2=1.15 $Y2=1.375
r135 14 28 18.8402 $w=1.65e-07 $l=8.66025e-08 $layer=POLY_cond $X=1.075 $Y=1.3
+ $X2=1.05 $Y2=1.375
r136 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.075 $Y=1.3
+ $X2=1.075 $Y2=0.74
r137 10 28 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=1.04 $Y=1.45
+ $X2=1.05 $Y2=1.375
r138 10 12 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=1.04 $Y=1.45
+ $X2=1.04 $Y2=2.4
r139 3 49 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=1.84 $X2=3.4 $Y2=2.375
r140 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.375
+ $Y=0.47 $X2=3.515 $Y2=0.615
r141 1 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.47 $X2=2.515 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%A 3 7 9 10 14 15
r44 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.515
+ $X2=2.14 $Y2=1.68
r45 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.515
+ $X2=2.14 $Y2=1.35
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.515 $X2=2.14 $Y2=1.515
r47 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=2.035
r48 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.515
r49 7 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.23 $Y=0.79 $X2=2.23
+ $Y2=1.35
r50 3 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.215 $Y=2.34
+ $X2=2.215 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%B 3 7 9 12 13
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.515
+ $X2=2.68 $Y2=1.68
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.515
+ $X2=2.68 $Y2=1.35
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.515 $X2=2.68 $Y2=1.515
r45 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.68 $Y=1.665
+ $X2=2.68 $Y2=1.515
r46 7 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.73 $Y=0.79 $X2=2.73
+ $Y2=1.35
r47 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.635 $Y=2.34
+ $X2=2.635 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%A_27_368# 1 2 9 12 15 16 19 20 21 24 25 28 31
+ 35
r95 28 29 6.23986 $w=5.67e-07 $l=2.9e-07 $layer=LI1_cond $X=0.445 $Y=2.115
+ $X2=0.445 $Y2=2.405
r96 25 35 48.5591 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.25 $Y=1.515
+ $X2=3.25 $Y2=1.725
r97 25 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.515
+ $X2=3.25 $Y2=1.35
r98 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.515 $X2=3.25 $Y2=1.515
r99 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.25 $Y=1.95
+ $X2=3.25 $Y2=1.515
r100 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=3.25 $Y2=1.95
r101 20 21 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=2.645 $Y2=2.035
r102 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=2.12
+ $X2=2.645 $Y2=2.035
r103 18 19 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.56 $Y=2.12 $X2=2.56
+ $Y2=2.32
r104 17 29 7.95352 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=0.775 $Y=2.405
+ $X2=0.445 $Y2=2.405
r105 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=2.405
+ $X2=2.56 $Y2=2.32
r106 16 17 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.475 $Y=2.405
+ $X2=0.775 $Y2=2.405
r107 15 28 10.1404 $w=5.67e-07 $l=3.16938e-07 $layer=LI1_cond $X=0.69 $Y=1.95
+ $X2=0.445 $Y2=2.115
r108 14 31 8.86325 $w=4.68e-07 $l=4.6465e-07 $layer=LI1_cond $X=0.69 $Y=1.13
+ $X2=0.35 $Y2=0.835
r109 14 15 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.69 $Y=1.13
+ $X2=0.69 $Y2=1.95
r110 12 34 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.3 $Y=0.79 $X2=3.3
+ $Y2=1.35
r111 9 35 164.683 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=3.175 $Y=2.34
+ $X2=3.175 $Y2=1.725
r112 2 28 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r113 1 31 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.56 $X2=0.35 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%VPWR 1 2 11 13 17 19 26 27 30 33
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 24 27 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 23 26 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 21 33 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.852 $Y2=3.33
r47 21 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=3.33 $X2=2.16
+ $Y2=3.33
r48 19 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 19 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 15 33 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.852 $Y=3.245
+ $X2=1.852 $Y2=3.33
r51 15 17 11.127 $w=4.33e-07 $l=4.2e-07 $layer=LI1_cond $X=1.852 $Y=3.245
+ $X2=1.852 $Y2=2.825
r52 14 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r53 13 33 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=1.852 $Y2=3.33
r54 13 14 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=0.98 $Y2=3.33
r55 9 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r56 9 11 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.78
r57 2 17 600 $w=1.7e-07 $l=1.11183e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.85 $Y2=2.825
r58 1 11 600 $w=1.7e-07 $l=1.04422e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%X 1 2 8 11 14 15 16
r37 15 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=1.985
+ $X2=1.235 $Y2=1.985
r38 15 16 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=1.985
+ $X2=1.68 $Y2=1.985
r39 15 20 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.26 $Y=1.985
+ $X2=1.235 $Y2=1.985
r40 13 14 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.26 $Y=0.96
+ $X2=1.26 $Y2=1.13
r41 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.29 $Y=0.515
+ $X2=1.29 $Y2=0.96
r42 8 15 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=1.82 $X2=1.15
+ $Y2=1.985
r43 8 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.15 $Y=1.82 $X2=1.15
+ $Y2=1.13
r44 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.265 $Y2=1.985
r45 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.37 $X2=1.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_2%VGND 1 2 3 12 14 18 22 24 25 27 28 29 40 41
+ 44
r51 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r54 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r55 35 44 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.135 $Y=0 $X2=1.88
+ $Y2=0
r56 35 37 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.64
+ $Y2=0
r57 33 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r58 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r59 29 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 29 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r61 27 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.64
+ $Y2=0
r62 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.015
+ $Y2=0
r63 26 40 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.6
+ $Y2=0
r64 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.015
+ $Y2=0
r65 24 32 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.72
+ $Y2=0
r66 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.86
+ $Y2=0
r67 20 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0
r68 20 22 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.645
r69 16 44 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=0.085
+ $X2=1.88 $Y2=0
r70 16 18 13.2507 $w=5.08e-07 $l=5.65e-07 $layer=LI1_cond $X=1.88 $Y=0.085
+ $X2=1.88 $Y2=0.65
r71 15 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.86
+ $Y2=0
r72 14 44 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.88
+ $Y2=0
r73 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=0.945
+ $Y2=0
r74 10 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0
r75 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0.57
r76 3 22 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.47 $X2=3.015 $Y2=0.645
r77 2 18 182 $w=1.7e-07 $l=4.38178e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.37 $X2=1.9 $Y2=0.65
r78 1 12 182 $w=1.7e-07 $l=2.24944e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.56 $X2=0.86 $Y2=0.57
.ends


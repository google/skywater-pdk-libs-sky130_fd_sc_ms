* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_27_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_1235_74# A3 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_325_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_325_74# A2 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_852_74# A2 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_325_74# A2 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1235_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 Y A1 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_852_74# A3 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 Y A1 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_1235_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND A4 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR A4 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 a_325_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X27 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 a_852_74# A3 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 a_852_74# A2 a_325_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND A4 a_1235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 a_27_368# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 a_1235_74# A3 a_852_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

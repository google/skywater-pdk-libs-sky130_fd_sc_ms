* File: sky130_fd_sc_ms__sedfxbp_2.spice
* Created: Wed Sep  2 12:32:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sedfxbp_2.pex.spice"
.subckt sky130_fd_sc_ms__sedfxbp_2  VNB VPB D DE SCD SCE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1001 A_141_74# N_D_M1001_g N_A_32_74#_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1659 PD=0.66 PS=1.63 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1042 N_VGND_M1042_d N_DE_M1042_g A_141_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_DE_M1020_g N_A_183_290#_M1020_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1021 A_527_113# N_A_183_290#_M1021_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_A_32_74#_M1005_d N_A_575_87#_M1005_g A_527_113# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_691_113#_M1009_d N_A_661_87#_M1009_g N_A_32_74#_M1005_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_SCE_M1037_g N_A_661_87#_M1037_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1017 A_1091_125# N_SCD_M1017_g N_VGND_M1037_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_691_113#_M1033_d N_SCE_M1033_g A_1091_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_1377_368#_M1029_d N_CLK_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_1586_74#_M1004_d N_A_1377_368#_M1004_g N_VGND_M1004_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_1784_97#_M1035_d N_A_1377_368#_M1035_g N_A_691_113#_M1035_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1038 A_1920_97# N_A_1586_74#_M1038_g N_A_1784_97#_M1035_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.09765 AS=0.1113 PD=0.885 PS=0.95 NRD=50.712 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_2013_71#_M1025_g A_1920_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.136292 AS=0.09765 PD=0.990566 PS=0.885 NRD=24.276 NRS=50.712 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1018 N_A_2013_71#_M1018_d N_A_1784_97#_M1018_g N_VGND_M1025_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.207683 PD=1.85 PS=1.50943 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 A_2417_74# N_A_2013_71#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1010 N_A_2489_74#_M1010_d N_A_1586_74#_M1010_g A_2417_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1011 A_2591_74# N_A_1377_368#_M1011_g N_A_2489_74#_M1010_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_575_87#_M1022_g A_2591_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.199681 AS=0.0504 PD=1.28534 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_A_575_87#_M1012_d N_A_2489_74#_M1012_g N_VGND_M1022_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.351819 PD=2.05 PS=2.26466 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_Q_M1026_d N_A_2489_74#_M1026_g N_VGND_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1047 N_Q_M1026_d N_A_2489_74#_M1047_g N_VGND_M1047_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1023 N_Q_N_M1023_d N_A_575_87#_M1023_g N_VGND_M1047_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1041 N_Q_N_M1023_d N_A_575_87#_M1041_g N_VGND_M1041_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 A_135_464# N_D_M1027_g N_A_32_74#_M1027_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1792 PD=0.88 PS=1.84 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1003 N_VPWR_M1003_d N_A_183_290#_M1003_g A_135_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.0768 PD=1.84 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90000.6
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1013 N_VPWR_M1013_d N_DE_M1013_g N_A_183_290#_M1013_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.14 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1045 A_581_462# N_DE_M1045_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=0.64 AD=0.0672
+ AS=0.16 PD=0.85 PS=1.14 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.9 SB=90001
+ A=0.1152 P=1.64 MULT=1
MM1024 N_A_32_74#_M1024_d N_A_575_87#_M1024_g A_581_462# VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.3 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1028 N_A_691_113#_M1028_d N_SCE_M1028_g N_A_32_74#_M1024_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.0864 PD=1.84 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90001.7 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1014 N_VPWR_M1014_d N_SCE_M1014_g N_A_661_87#_M1014_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1632 AS=0.1856 PD=1.15 PS=1.86 NRD=69.2455 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1031 A_1091_453# N_SCD_M1031_g N_VPWR_M1014_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1632 PD=0.88 PS=1.15 NRD=19.9955 NRS=1.5366 M=1 R=3.55556
+ SA=90000.9 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1040 N_A_691_113#_M1040_d N_A_661_87#_M1040_g A_1091_453# VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.0768 PD=1.84 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556
+ SA=90001.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1000 N_A_1377_368#_M1000_d N_CLK_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1008 N_A_1586_74#_M1008_d N_A_1377_368#_M1008_g N_VPWR_M1008_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1015 N_A_1784_97#_M1015_d N_A_1586_74#_M1015_g N_A_691_113#_M1015_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1019 A_1947_508# N_A_1377_368#_M1019_g N_A_1784_97#_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0693 AS=0.0567 PD=0.75 PS=0.69 NRD=51.5943 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1016 N_VPWR_M1016_d N_A_2013_71#_M1016_g A_1947_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0936833 AS=0.0693 PD=0.89 PS=0.75 NRD=2.3443 NRS=51.5943 M=1 R=2.33333
+ SA=90001.1 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1032 N_A_2013_71#_M1032_d N_A_1784_97#_M1032_g N_VPWR_M1016_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.187367 PD=2.24 PS=1.78 NRD=0 NRS=19.9167 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1043 A_2377_392# N_A_2013_71#_M1043_g N_VPWR_M1043_s VPB PSHORT L=0.18 W=1
+ AD=0.3875 AS=0.3882 PD=1.775 PS=2.89 NRD=65.4828 NRS=16.7253 M=1 R=5.55556
+ SA=90000.3 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1034 N_A_2489_74#_M1034_d N_A_1377_368#_M1034_g A_2377_392# VPB PSHORT L=0.18
+ W=1 AD=0.219366 AS=0.3875 PD=1.90845 PS=1.775 NRD=0 NRS=65.4828 M=1 R=5.55556
+ SA=90001.2 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1030 A_2675_508# N_A_1586_74#_M1030_g N_A_2489_74#_M1034_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0921338 PD=0.66 PS=0.801549 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90001.8 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_575_87#_M1006_g A_2675_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.108436 AS=0.0504 PD=0.9 PS=0.66 NRD=46.886 NRS=30.4759 M=1 R=2.33333
+ SA=90002.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1044 N_A_575_87#_M1044_d N_A_2489_74#_M1044_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.289164 PD=2.8 PS=2.4 NRD=0 NRS=26.3783 M=1 R=6.22222
+ SA=90001.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1036 N_Q_M1036_d N_A_2489_74#_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1039 N_Q_M1036_d N_A_2489_74#_M1039_g N_VPWR_M1039_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1039_s N_A_575_87#_M1002_g N_Q_N_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1046 N_VPWR_M1046_d N_A_575_87#_M1046_g N_Q_N_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX48_noxref VNB VPB NWDIODE A=32.8476 P=39.04
c_188 VNB 0 1.45871e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sedfxbp_2.pxi.spice"
*
.ends
*
*

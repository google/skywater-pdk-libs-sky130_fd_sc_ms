* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2b_4 A B_N VGND VNB VPB VPWR X
M1000 a_81_296# A VGND VNB nlowvt w=640000u l=150000u
+  ad=4.672e+11p pd=4.02e+06u as=1.1509e+12p ps=1.032e+07u
M1001 a_81_296# a_676_48# a_492_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=8.2e+11p ps=7.64e+06u
M1002 a_492_392# a_676_48# a_81_296# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_492_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.5272e+12p ps=1.358e+07u
M1004 VPWR A a_492_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_81_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1006 a_81_296# a_676_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_81_296# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_81_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1009 VPWR a_81_296# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_81_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_81_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_81_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_81_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_676_48# B_N VGND VNB nlowvt w=640000u l=150000u
+  ad=6.272e+11p pd=3.24e+06u as=0p ps=0u
M1015 a_676_48# B_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1016 VPWR a_81_296# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_676_48# a_81_296# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

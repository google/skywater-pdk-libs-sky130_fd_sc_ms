* File: sky130_fd_sc_ms__and4bb_2.pex.spice
* Created: Wed Sep  2 11:59:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4BB_2%A_N 3 5 7 8 12
c31 12 0 1.82461e-19 $X=0.385 $Y=1.615
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r33 8 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r34 5 11 45.7042 $w=3.84e-07 $l=3.19374e-07 $layer=POLY_cond $X=0.6 $Y=1.87
+ $X2=0.455 $Y2=1.615
r35 5 7 136.567 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=0.6 $Y=1.87 $X2=0.6
+ $Y2=2.38
r36 1 11 39.2873 $w=3.84e-07 $l=1.83916e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.455 $Y2=1.615
r37 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%A_27_74# 1 2 9 13 17 21 22 23 25 26 28 34
c66 34 0 1.82461e-19 $X=1.17 $Y=1.505
c67 13 0 1.77462e-19 $X=1.485 $Y=0.78
r68 32 34 14.8156 $w=2.44e-07 $l=7.5e-08 $layer=POLY_cond $X=1.095 $Y=1.505
+ $X2=1.17 $Y2=1.505
r69 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.505 $X2=1.095 $Y2=1.505
r70 25 31 9.01265 $w=3.61e-07 $l=2.32282e-07 $layer=LI1_cond $X=0.85 $Y=1.67
+ $X2=1.012 $Y2=1.505
r71 25 26 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.85 $Y=1.67
+ $X2=0.85 $Y2=1.95
r72 24 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=2.035
+ $X2=0.375 $Y2=2.035
r73 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.85 $Y2=1.95
r74 23 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.54 $Y2=2.035
r75 21 31 10.4765 $w=3.61e-07 $l=4.15536e-07 $layer=LI1_cond $X=0.765 $Y=1.195
+ $X2=1.012 $Y2=1.505
r76 21 22 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.765 $Y=1.195
+ $X2=0.365 $Y2=1.195
r77 15 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.365 $Y2=1.195
r78 15 17 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.24 $Y2=0.645
r79 11 34 62.2254 $w=2.44e-07 $l=3.88844e-07 $layer=POLY_cond $X=1.485 $Y=1.34
+ $X2=1.17 $Y2=1.505
r80 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.485 $Y=1.34
+ $X2=1.485 $Y2=0.78
r81 7 34 9.95785 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.67
+ $X2=1.17 $Y2=1.505
r82 7 9 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.17 $Y=1.67 $X2=1.17
+ $Y2=2.46
r83 2 28 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.23
+ $Y=1.96 $X2=0.375 $Y2=2.115
r84 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%A_354_252# 1 2 9 12 16 17 19 20 22 23 24 26
+ 27 29 30 33 35 36 42
c114 36 0 1.65552e-19 $X=5 $Y=0.665
c115 20 0 2.96366e-19 $X=2.1 $Y=1.085
r116 36 39 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=5 $Y=0.665 $X2=5
+ $Y2=0.795
r117 31 33 1.83723 $w=3.43e-07 $l=5.5e-08 $layer=LI1_cond $X=4.992 $Y=1.93
+ $X2=4.992 $Y2=1.985
r118 29 31 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=4.82 $Y=1.845
+ $X2=4.992 $Y2=1.93
r119 29 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.82 $Y=1.845
+ $X2=4.535 $Y2=1.845
r120 28 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=0.665
+ $X2=4.45 $Y2=0.665
r121 27 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.665
+ $X2=5 $Y2=0.665
r122 27 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.835 $Y=0.665
+ $X2=4.535 $Y2=0.665
r123 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=1.76
+ $X2=4.535 $Y2=1.845
r124 25 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.665
r125 25 26 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=1.76
r126 23 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0.665
+ $X2=4.45 $Y2=0.665
r127 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.365 $Y=0.665
+ $X2=3.645 $Y2=0.665
r128 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=0.75
+ $X2=3.645 $Y2=0.665
r129 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.56 $Y=0.75
+ $X2=3.56 $Y2=1
r130 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.475 $Y=1.085
+ $X2=3.56 $Y2=1
r131 19 20 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=3.475 $Y=1.085
+ $X2=2.1 $Y2=1.085
r132 17 43 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.425
+ $X2=1.935 $Y2=1.59
r133 17 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.425
+ $X2=1.935 $Y2=1.26
r134 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.425 $X2=1.935 $Y2=1.425
r135 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.935 $Y=1.17
+ $X2=2.1 $Y2=1.085
r136 14 16 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=1.17
+ $X2=1.935 $Y2=1.425
r137 12 43 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=1.89 $Y=2.46
+ $X2=1.89 $Y2=1.59
r138 9 42 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.875 $Y=0.78
+ $X2=1.875 $Y2=1.26
r139 2 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.85
+ $Y=1.84 $X2=4.99 $Y2=1.985
r140 1 39 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.6 $X2=5 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%C 3 7 9 12
c37 9 0 1.78968e-19 $X=2.64 $Y=1.665
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.475 $Y=1.585
+ $X2=2.475 $Y2=1.75
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.475 $Y=1.585
+ $X2=2.475 $Y2=1.42
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.475
+ $Y=1.585 $X2=2.475 $Y2=1.585
r41 9 13 5.28203 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.6
+ $X2=2.475 $Y2=1.6
r42 7 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=2.55 $Y=2.46 $X2=2.55
+ $Y2=1.75
r43 3 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.415 $Y=0.78
+ $X2=2.415 $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%D 3 7 9 12
c41 7 0 1.78968e-19 $X=3 $Y=2.46
r42 12 15 40.0728 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.052 $Y=1.585
+ $X2=3.052 $Y2=1.75
r43 12 14 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.052 $Y=1.585
+ $X2=3.052 $Y2=1.42
r44 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.585 $X2=3.09 $Y2=1.585
r45 7 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=3 $Y=2.46 $X2=3
+ $Y2=1.75
r46 3 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.925 $Y=0.78
+ $X2=2.925 $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%A_225_82# 1 2 3 12 16 20 24 28 31 34 36 40
+ 42 45 46 48 50 54 62
c129 54 0 1.46091e-19 $X=3.69 $Y=1.505
c130 20 0 1.65552e-19 $X=4.195 $Y=0.78
r131 61 62 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.195 $Y=1.505
+ $X2=4.225 $Y2=1.505
r132 60 61 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.775 $Y=1.505
+ $X2=4.195 $Y2=1.505
r133 59 60 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.765 $Y=1.505
+ $X2=3.775 $Y2=1.505
r134 55 59 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=1.505
+ $X2=3.765 $Y2=1.505
r135 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.69
+ $Y=1.505 $X2=3.69 $Y2=1.505
r136 51 54 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.58 $Y=1.505
+ $X2=3.69 $Y2=1.505
r137 44 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=1.67
+ $X2=3.58 $Y2=1.505
r138 44 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.58 $Y=1.67
+ $X2=3.58 $Y2=1.95
r139 43 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.94 $Y=2.035
+ $X2=2.775 $Y2=2.035
r140 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.495 $Y=2.035
+ $X2=3.58 $Y2=1.95
r141 42 43 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.495 $Y=2.035
+ $X2=2.94 $Y2=2.035
r142 38 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=2.12
+ $X2=2.775 $Y2=2.035
r143 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.775 $Y=2.12
+ $X2=2.775 $Y2=2.815
r144 37 48 2.76166 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.76 $Y=2.035
+ $X2=1.595 $Y2=2.03
r145 36 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=2.035
+ $X2=2.775 $Y2=2.035
r146 36 37 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.61 $Y=2.035
+ $X2=1.76 $Y2=2.035
r147 32 48 3.70735 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.595 $Y=2.12
+ $X2=1.595 $Y2=2.03
r148 32 34 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.595 $Y=2.12
+ $X2=1.595 $Y2=2.815
r149 31 48 3.70735 $w=2.5e-07 $l=1.23693e-07 $layer=LI1_cond $X=1.515 $Y=1.94
+ $X2=1.595 $Y2=2.03
r150 31 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.515 $Y=1.94
+ $X2=1.515 $Y2=1.17
r151 26 46 11.4679 $w=4.93e-07 $l=2.47e-07 $layer=LI1_cond $X=1.352 $Y=0.923
+ $X2=1.352 $Y2=1.17
r152 26 28 8.89206 $w=4.93e-07 $l=3.68e-07 $layer=LI1_cond $X=1.352 $Y=0.923
+ $X2=1.352 $Y2=0.555
r153 22 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.225 $Y=1.67
+ $X2=4.225 $Y2=1.505
r154 22 24 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=4.225 $Y=1.67
+ $X2=4.225 $Y2=2.4
r155 18 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=1.34
+ $X2=4.195 $Y2=1.505
r156 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.195 $Y=1.34
+ $X2=4.195 $Y2=0.78
r157 14 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.34
+ $X2=3.765 $Y2=1.505
r158 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.765 $Y=1.34
+ $X2=3.765 $Y2=0.78
r159 10 60 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=1.67
+ $X2=3.775 $Y2=1.505
r160 10 12 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=3.775 $Y=1.67
+ $X2=3.775 $Y2=2.4
r161 3 50 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.96 $X2=2.775 $Y2=2.115
r162 3 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.96 $X2=2.775 $Y2=2.815
r163 2 48 400 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.96 $X2=1.595 $Y2=2.105
r164 2 34 400 $w=1.7e-07 $l=1.00869e-06 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.96 $X2=1.595 $Y2=2.815
r165 1 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.41 $X2=1.27 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%B_N 3 5 7 8 14
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.425 $X2=4.99 $Y2=1.425
r29 12 14 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.785 $Y=1.425
+ $X2=4.99 $Y2=1.425
r30 10 12 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=4.76 $Y=1.425
+ $X2=4.785 $Y2=1.425
r31 8 15 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.99 $Y=1.295
+ $X2=4.99 $Y2=1.425
r32 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.26
+ $X2=4.785 $Y2=1.425
r33 5 7 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.785 $Y=1.26
+ $X2=4.785 $Y2=0.875
r34 1 10 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.76 $Y=1.59
+ $X2=4.76 $Y2=1.425
r35 1 3 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=4.76 $Y=1.59 $X2=4.76
+ $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%VPWR 1 2 3 4 15 21 25 29 34 35 37 38 40 41
+ 42 48 60 61 64
r71 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r73 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r74 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r75 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r77 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r78 52 54 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r82 48 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 46 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r86 42 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r87 40 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.49 $Y2=3.33
r89 39 60 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.615 $Y=3.33
+ $X2=5.04 $Y2=3.33
r90 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.615 $Y=3.33
+ $X2=4.49 $Y2=3.33
r91 37 54 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.2 $Y=3.33 $X2=3.12
+ $Y2=3.33
r92 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=3.33
+ $X2=3.365 $Y2=3.33
r93 36 57 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.53 $Y=3.33
+ $X2=4.08 $Y2=3.33
r94 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=3.33
+ $X2=3.365 $Y2=3.33
r95 34 45 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.78 $Y=3.33 $X2=0.72
+ $Y2=3.33
r96 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=0.945 $Y2=3.33
r97 33 50 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.11 $Y=3.33
+ $X2=1.68 $Y2=3.33
r98 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=3.33
+ $X2=0.945 $Y2=3.33
r99 29 32 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=4.49 $Y=2.265
+ $X2=4.49 $Y2=2.815
r100 27 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=3.245
+ $X2=4.49 $Y2=3.33
r101 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.49 $Y=3.245
+ $X2=4.49 $Y2=2.815
r102 23 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=3.245
+ $X2=3.365 $Y2=3.33
r103 23 25 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.365 $Y=3.245
+ $X2=3.365 $Y2=2.405
r104 19 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r105 19 21 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.41
r106 15 18 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.815
r107 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=3.245
+ $X2=0.945 $Y2=3.33
r108 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.945 $Y=3.245
+ $X2=0.945 $Y2=2.815
r109 4 32 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.84 $X2=4.45 $Y2=2.815
r110 4 29 600 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.84 $X2=4.45 $Y2=2.265
r111 3 25 300 $w=1.7e-07 $l=5.66039e-07 $layer=licon1_PDIFF $count=2 $X=3.09
+ $Y=1.96 $X2=3.365 $Y2=2.405
r112 2 21 300 $w=1.7e-07 $l=5.61249e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.96 $X2=2.23 $Y2=2.41
r113 1 18 600 $w=1.7e-07 $l=9.74192e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.96 $X2=0.945 $Y2=2.815
r114 1 15 600 $w=1.7e-07 $l=5.27304e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.96 $X2=0.945 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%X 1 2 12 14 15 16 23 32
r35 21 23 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=4.015 $Y=2.02
+ $X2=4.015 $Y2=2.035
r36 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=4.015 $Y=2.405
+ $X2=4.015 $Y2=2.775
r37 14 21 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.015 $Y=1.985
+ $X2=4.015 $Y2=2.02
r38 14 32 7.87078 $w=3.58e-07 $l=1.45e-07 $layer=LI1_cond $X=4.015 $Y=1.985
+ $X2=4.015 $Y2=1.84
r39 14 15 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=4.015 $Y=2.07
+ $X2=4.015 $Y2=2.405
r40 14 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.015 $Y=2.07
+ $X2=4.015 $Y2=2.035
r41 10 12 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=3.98 $Y=1.045
+ $X2=4.11 $Y2=1.045
r42 7 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.11 $Y=1.17 $X2=4.11
+ $Y2=1.045
r43 7 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.11 $Y=1.17 $X2=4.11
+ $Y2=1.84
r44 2 14 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.84 $X2=4 $Y2=2.005
r45 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.84 $X2=4 $Y2=2.815
r46 1 10 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.84
+ $Y=0.41 $X2=3.98 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_2%VGND 1 2 3 12 16 18 20 25 33 40 41 44 47 51
r62 51 54 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=4.49
+ $Y2=0.325
r63 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r64 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r65 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r67 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r68 38 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.49
+ $Y2=0
r69 38 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=5.04
+ $Y2=0
r70 37 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r71 37 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r72 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r73 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r74 34 36 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=4.08
+ $Y2=0
r75 33 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.49
+ $Y2=0
r76 33 36 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.08
+ $Y2=0
r77 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r78 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r79 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r80 26 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r81 26 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r82 25 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r83 25 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.64
+ $Y2=0
r84 23 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r85 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r86 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r87 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r88 18 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r89 18 29 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r90 18 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r91 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r92 14 16 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.665
r93 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r94 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.645
r95 3 54 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.41 $X2=4.49 $Y2=0.325
r96 2 16 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3 $Y=0.41
+ $X2=3.14 $Y2=0.665
r97 1 12 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.645
.ends


* File: sky130_fd_sc_ms__clkinv_2.spice
* Created: Wed Sep  2 12:01:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkinv_2.pex.spice"
.subckt sky130_fd_sc_ms__clkinv_2  VNB VPB A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.1638 PD=1.41 PS=1.2 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.1638 PD=1.41 PS=1.2 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90001.1
+ A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1000_d N_A_M1001_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX5_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ms__clkinv_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfstp_2.spice
* Created: Fri Aug 28 17:24:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfstp_2.pex.spice"
.subckt sky130_fd_sc_ms__dfstp_2  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_D_M1031_g N_A_27_74#_M1031_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_225_74#_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_A_398_74#_M1015_d N_A_225_74#_M1015_g N_VGND_M1033_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_612_74#_M1018_d N_A_225_74#_M1018_g N_A_27_74#_M1018_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.14595 AS=0.18665 PD=1.115 PS=1.8 NRD=71.424 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 A_781_74# N_A_398_74#_M1012_g N_A_612_74#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.14595 PD=0.66 PS=1.115 NRD=18.564 NRS=47.136 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_767_384#_M1024_g A_781_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1057_118# N_A_612_74#_M1002_g N_A_767_384#_M1002_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_1057_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.120611 AS=0.0504 PD=0.954906 PS=0.66 NRD=38.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1000 A_1278_74# N_A_612_74#_M1000_g N_VGND_M1022_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.183789 PD=0.88 PS=1.45509 NRD=12.18 NRS=28.584 M=1 R=4.26667
+ SA=75000.9 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_1356_74#_M1001_d N_A_398_74#_M1001_g A_1278_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.163804 AS=0.0768 PD=1.39472 PS=0.88 NRD=21.552 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1008 A_1489_118# N_A_225_74#_M1008_g N_A_1356_74#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08085 AS=0.107496 PD=0.805 PS=0.915283 NRD=39.276 NRS=34.284 M=1
+ R=2.8 SA=75002.4 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1030 A_1596_118# N_A_1566_92#_M1030_g A_1489_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.08085 PD=0.84 PS=0.805 NRD=44.28 NRS=39.276 M=1 R=2.8
+ SA=75002.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SET_B_M1004_g A_1596_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.17955 AS=0.0882 PD=1.275 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75003.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1027 N_A_1566_92#_M1027_d N_A_1356_74#_M1027_g N_VGND_M1004_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.17955 PD=1.41 PS=1.275 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75004.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1356_74#_M1013_g N_A_2022_94#_M1013_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.144093 AS=0.1824 PD=1.08522 PS=1.85 NRD=15.468 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1013_d N_A_2022_94#_M1005_g N_Q_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.1036 PD=1.25478 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_A_2022_94#_M1025_g N_Q_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2294 AS=0.1036 PD=2.1 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_D_M1020_g N_A_27_74#_M1020_s VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1014 N_VPWR_M1014_d N_CLK_M1014_g N_A_225_74#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1017 N_A_398_74#_M1017_d N_A_225_74#_M1017_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1023 N_A_612_74#_M1023_d N_A_398_74#_M1023_g N_A_27_74#_M1023_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90004.6 A=0.0756 P=1.2 MULT=1
MM1021 A_719_456# N_A_225_74#_M1021_g N_A_612_74#_M1023_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0672 PD=0.66 PS=0.74 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90004.1 A=0.0756 P=1.2 MULT=1
MM1032 N_VPWR_M1032_d N_A_767_384#_M1032_g A_719_456# VPB PSHORT L=0.18 W=0.42
+ AD=0.240525 AS=0.0504 PD=1.545 PS=0.66 NRD=79.7259 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1009 N_A_767_384#_M1009_d N_A_612_74#_M1009_g N_VPWR_M1032_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.240525 PD=0.69 PS=1.545 NRD=0 NRS=242.802 M=1 R=2.33333
+ SA=90002.2 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1016 N_VPWR_M1016_d N_SET_B_M1016_g N_A_767_384#_M1009_d VPB PSHORT L=0.18
+ W=0.42 AD=0.13846 AS=0.0567 PD=1.09437 PS=0.69 NRD=128.818 NRS=0 M=1 R=2.33333
+ SA=90002.7 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1011 A_1269_341# N_A_612_74#_M1011_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=1
+ AD=0.184812 AS=0.329665 PD=1.58 PS=2.60563 NRD=25.5706 NRS=54.0962 M=1
+ R=5.55556 SA=90001.5 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1003 N_A_1356_74#_M1003_d N_A_225_74#_M1003_g A_1269_341# VPB PSHORT L=0.18
+ W=1 AD=0.288873 AS=0.184812 PD=2.23944 PS=1.58 NRD=20.0152 NRS=25.5706 M=1
+ R=5.55556 SA=90001.9 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1010 A_1524_508# N_A_398_74#_M1010_g N_A_1356_74#_M1003_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.121327 PD=0.66 PS=0.940563 NRD=30.4759 NRS=73.875 M=1
+ R=2.33333 SA=90002.4 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1028 N_VPWR_M1028_d N_A_1566_92#_M1028_g A_1524_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=39.8531 NRS=30.4759 M=1 R=2.33333
+ SA=90002.8 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1007 N_A_1356_74#_M1007_d N_SET_B_M1007_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0756 PD=1.4 PS=0.78 NRD=0 NRS=0 M=1 R=2.33333 SA=90003.3
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1019 N_A_1566_92#_M1019_d N_A_1356_74#_M1019_g N_VPWR_M1019_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_1356_74#_M1006_g N_A_2022_94#_M1006_s VPB PSHORT
+ L=0.18 W=1 AD=0.183302 AS=0.28 PD=1.39151 PS=2.56 NRD=16.2525 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1026 N_Q_M1026_d N_A_2022_94#_M1026_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.205298 PD=1.39 PS=1.55849 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1029 N_Q_M1026_d N_A_2022_94#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.4057 P=28.75
c_1623 A_719_456# 0 2.15866e-20 $X=3.595 $Y=2.28
*
.include "sky130_fd_sc_ms__dfstp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlxbn_1.spice
* Created: Fri Aug 28 17:28:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlxbn_1.pex.spice"
.subckt sky130_fd_sc_ms__dlxbn_1  VNB VPB D GATE_N VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_D_M1020_g N_A_27_120#_M1020_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.161184 AS=0.15675 PD=1.20233 PS=1.67 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_A_232_82#_M1003_d N_GATE_N_M1003_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_232_82#_M1008_g N_A_343_80#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.193727 AS=0.3182 PD=1.49072 PS=2.34 NRD=33.528 NRS=1.62 M=1
+ R=4.93333 SA=75000.4 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1013 A_575_79# N_A_27_120#_M1013_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.167548 PD=0.88 PS=1.28928 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75000.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1012 N_A_653_79#_M1012_d N_A_232_82#_M1012_g A_575_79# VNB NLOWVT L=0.15
+ W=0.64 AD=0.247487 AS=0.0768 PD=1.79321 PS=0.88 NRD=18.744 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1010 A_852_123# N_A_343_80#_M1010_g N_A_653_79#_M1012_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.162413 PD=0.66 PS=1.17679 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_863_294#_M1004_g A_852_123# VNB NLOWVT L=0.15 W=0.42
+ AD=0.101262 AS=0.0504 PD=0.84 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_863_294#_M1005_d N_A_653_79#_M1005_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2183 AS=0.178413 PD=2.07 PS=1.48 NRD=1.62 NRS=9.72 M=1 R=4.93333
+ SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_863_294#_M1009_g N_Q_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.140829 AS=0.2109 PD=1.26202 PS=2.05 NRD=7.296 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_1350_424#_M1017_d N_A_863_294#_M1017_g N_VGND_M1009_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.104671 PD=1.67 PS=0.937984 NRD=0 NRS=7.632 M=1
+ R=3.66667 SA=75000.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1007 N_Q_N_M1007_d N_A_1350_424#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_120#_M1000_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2814 PD=1.16 PS=2.35 NRD=0 NRS=15.2281 M=1 R=4.66667 SA=90000.2
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1001 N_A_232_82#_M1001_d N_GATE_N_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1344 PD=2.24 PS=1.16 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1021 N_VPWR_M1021_d N_A_232_82#_M1021_g N_A_343_80#_M1021_s VPB PSHORT L=0.18
+ W=0.84 AD=0.161152 AS=0.2352 PD=1.2463 PS=2.24 NRD=19.9167 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1002 A_574_392# N_A_27_120#_M1002_g N_VPWR_M1021_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.191848 PD=1.24 PS=1.4837 NRD=12.7853 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1014 N_A_653_79#_M1014_d N_A_343_80#_M1014_g A_574_392# VPB PSHORT L=0.18 W=1
+ AD=0.270704 AS=0.12 PD=2.21127 PS=1.24 NRD=19.7 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90001 A=0.18 P=2.36 MULT=1
MM1006 A_808_392# N_A_232_82#_M1006_g N_A_653_79#_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.06405 AS=0.113696 PD=0.725 PS=0.928732 NRD=45.7237 NRS=89.1031 M=1
+ R=2.33333 SA=90001.9 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_863_294#_M1011_g A_808_392# VPB PSHORT L=0.18 W=0.42
+ AD=0.115064 AS=0.06405 PD=0.908182 PS=0.725 NRD=39.8531 NRS=45.7237 M=1
+ R=2.33333 SA=90002.4 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1015 N_A_863_294#_M1015_d N_A_653_79#_M1015_g N_VPWR_M1011_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.306836 PD=2.77 PS=2.42182 NRD=0 NRS=15.3857 M=1
+ R=6.22222 SA=90001.3 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1019_d N_A_863_294#_M1019_g N_Q_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.196 AS=0.2968 PD=1.65143 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1016 N_A_1350_424#_M1016_d N_A_863_294#_M1016_g N_VPWR_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.147 PD=2.24 PS=1.23857 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1018 N_Q_N_M1018_d N_A_1350_424#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.2968 PD=2.8 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.97 P=20.96
*
.include "sky130_fd_sc_ms__dlxbn_1.pxi.spice"
*
.ends
*
*

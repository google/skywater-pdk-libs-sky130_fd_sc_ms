* File: sky130_fd_sc_ms__nand2b_2.pex.spice
* Created: Fri Aug 28 17:42:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND2B_2%A_N 1 3 6 8 12
c28 12 0 1.50161e-19 $X=0.405 $Y=1.515
c29 1 0 1.52201e-19 $X=0.505 $Y=1.8
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.515 $X2=0.405 $Y2=1.515
r31 8 12 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.405 $Y2=1.565
r32 4 11 38.6342 $w=2.88e-07 $l=2.00237e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.417 $Y2=1.515
r33 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.69
r34 1 11 54.4391 $w=2.88e-07 $l=3.26044e-07 $layer=POLY_cond $X=0.505 $Y=1.8
+ $X2=0.417 $Y2=1.515
r35 1 3 144.6 $w=1.8e-07 $l=5.4e-07 $layer=POLY_cond $X=0.505 $Y=1.8 $X2=0.505
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_2%A_27_74# 1 2 7 11 15 17 21 25 27 28 31 35
+ 36 37 39 40 42 46
c93 46 0 1.50161e-19 $X=0.97 $Y=1.305
c94 39 0 3.18194e-19 $X=0.89 $Y=1.47
c95 28 0 2.31616e-19 $X=1.97 $Y=1.395
c96 11 0 1.49852e-19 $X=1.505 $Y=2.4
r97 46 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.97 $Y=1.305 $X2=0.97
+ $Y2=1.395
r98 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.305 $X2=0.97 $Y2=1.305
r99 43 45 9.02113 $w=2.84e-07 $l=2.1e-07 $layer=LI1_cond $X=0.97 $Y=1.095
+ $X2=0.97 $Y2=1.305
r100 39 45 9.03839 $w=2.84e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.89 $Y=1.47
+ $X2=0.97 $Y2=1.305
r101 39 40 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.89 $Y=1.47
+ $X2=0.89 $Y2=1.95
r102 38 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r103 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.89 $Y2=1.95
r104 37 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.445 $Y2=2.035
r105 35 43 3.73949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.095
+ $X2=0.97 $Y2=1.095
r106 35 36 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.805 $Y=1.095
+ $X2=0.445 $Y2=1.095
r107 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r108 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r109 23 28 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=2 $Y=1.32
+ $X2=1.97 $Y2=1.395
r110 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2 $Y=1.32 $X2=2
+ $Y2=0.74
r111 19 28 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.955 $Y=1.47
+ $X2=1.97 $Y2=1.395
r112 19 21 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=1.955 $Y=1.47
+ $X2=1.955 $Y2=2.4
r113 18 27 13.2179 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.645 $Y=1.395
+ $X2=1.53 $Y2=1.395
r114 17 28 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=1.865 $Y=1.395
+ $X2=1.97 $Y2=1.395
r115 17 18 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.865 $Y=1.395
+ $X2=1.645 $Y2=1.395
r116 13 27 10.9219 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=1.57 $Y=1.32
+ $X2=1.53 $Y2=1.395
r117 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.57 $Y=1.32
+ $X2=1.57 $Y2=0.74
r118 9 27 10.9219 $w=1.8e-07 $l=8.66025e-08 $layer=POLY_cond $X=1.505 $Y=1.47
+ $X2=1.53 $Y2=1.395
r119 9 11 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=1.505 $Y=1.47
+ $X2=1.505 $Y2=2.4
r120 8 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.395
+ $X2=0.97 $Y2=1.395
r121 7 27 13.2179 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.415 $Y=1.395
+ $X2=1.53 $Y2=1.395
r122 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.415 $Y=1.395
+ $X2=1.135 $Y2=1.395
r123 2 42 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r124 1 31 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_2%B 3 7 11 15 17 24 26
c47 24 0 8.98252e-20 $X=2.61 $Y=1.515
r48 25 26 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.855 $Y=1.515
+ $X2=2.865 $Y2=1.515
r49 23 25 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.61 $Y=1.515
+ $X2=2.855 $Y2=1.515
r50 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r51 21 23 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.43 $Y=1.515
+ $X2=2.61 $Y2=1.515
r52 19 21 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.405 $Y=1.515
+ $X2=2.43 $Y2=1.515
r53 17 24 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.515
r54 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=2.865 $Y2=1.515
r55 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=2.865 $Y2=0.74
r56 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.855 $Y2=1.515
r57 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.855 $Y2=2.4
r58 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.35
+ $X2=2.43 $Y2=1.515
r59 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.43 $Y=1.35 $X2=2.43
+ $Y2=0.74
r60 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=1.515
r61 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_2%VPWR 1 2 3 12 16 18 20 23 24 25 31 35 41 45
r47 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 39 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r53 36 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 35 44 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r55 35 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 31 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r57 31 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 25 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 25 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 23 28 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 23 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.91 $Y2=3.33
r64 22 33 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 22 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.91 $Y2=3.33
r66 18 44 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r67 18 20 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.805
r68 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r69 14 16 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.805
r70 10 24 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=3.245
+ $X2=0.91 $Y2=3.33
r71 10 12 26.1636 $w=3.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.91 $Y=3.245
+ $X2=0.91 $Y2=2.405
r72 3 20 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.805
r73 2 16 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.84 $X2=2.18 $Y2=2.805
r74 1 12 300 $w=1.7e-07 $l=7.07124e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.915 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_2%Y 1 2 3 10 16 18 19 22 25 26
c41 26 0 1.91337e-19 $X=2.16 $Y=2.035
c42 19 0 1.41791e-19 $X=1.87 $Y=1.305
c43 10 0 1.49852e-19 $X=2.045 $Y=2.01
r44 26 29 2.49594 $w=2.3e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=2.01 $X2=2.16
+ $Y2=1.82
r45 25 29 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.82
r46 24 25 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=1.39
+ $X2=2.16 $Y2=1.665
r47 20 26 3.9473 $w=3.15e-07 $l=1.43875e-07 $layer=LI1_cond $X=2.275 $Y=2.075
+ $X2=2.16 $Y2=2.01
r48 20 22 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=2.275 $Y=2.075
+ $X2=2.63 $Y2=2.075
r49 18 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=1.305
+ $X2=2.16 $Y2=1.39
r50 18 19 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.045 $Y=1.305
+ $X2=1.87 $Y2=1.305
r51 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.785 $Y=1.22
+ $X2=1.87 $Y2=1.305
r52 14 16 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.785 $Y=1.22
+ $X2=1.785 $Y2=0.825
r53 10 26 3.9473 $w=3.15e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=2.01
+ $X2=2.16 $Y2=2.01
r54 10 12 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.045 $Y=2.01
+ $X2=1.73 $Y2=2.01
r55 3 22 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.115
r56 2 12 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.73 $Y2=2.01
r57 1 16 182 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.37 $X2=1.785 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_2%VGND 1 2 9 13 15 17 22 29 30 33 36
c40 1 0 1.65994e-19 $X=0.57 $Y=0.37
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r44 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.645
+ $Y2=0
r46 27 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=3.12
+ $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.745
+ $Y2=0
r50 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.645
+ $Y2=0
r52 22 25 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=0 $X2=1.2
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.745
+ $Y2=0
r56 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r58 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0
r60 11 13 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0.515
r61 7 33 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r62 7 9 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.675
r63 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.505
+ $Y=0.37 $X2=2.645 $Y2=0.515
r64 1 9 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2B_2%A_242_74# 1 2 3 13 15 16 17 18 19 22 26 29
+ 30 31
r77 29 31 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.16 $Y=2.37
+ $X2=3.16 $Y2=1.13
r78 24 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0.965
+ $X2=3.08 $Y2=1.13
r79 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.08 $Y=0.965
+ $X2=3.08 $Y2=0.515
r80 20 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.215 $Y=0.425
+ $X2=2.215 $Y2=0.515
r81 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.05 $Y=0.34
+ $X2=2.215 $Y2=0.425
r82 18 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.05 $Y=0.34
+ $X2=1.52 $Y2=0.34
r83 16 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.455
+ $X2=3.16 $Y2=2.37
r84 16 17 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=3.075 $Y=2.455
+ $X2=1.475 $Y2=2.455
r85 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.39 $Y=2.37
+ $X2=1.475 $Y2=2.455
r86 15 30 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.39 $Y=2.37
+ $X2=1.39 $Y2=0.97
r87 11 30 7.49019 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.805
+ $X2=1.355 $Y2=0.97
r88 11 13 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.355 $Y=0.805
+ $X2=1.355 $Y2=0.515
r89 10 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=0.425
+ $X2=1.52 $Y2=0.34
r90 10 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.355 $Y=0.425
+ $X2=1.355 $Y2=0.515
r91 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
r92 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.075
+ $Y=0.37 $X2=2.215 $Y2=0.515
r93 1 13 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.21
+ $Y=0.37 $X2=1.355 $Y2=0.515
.ends


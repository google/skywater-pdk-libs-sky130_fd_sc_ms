* File: sky130_fd_sc_ms__o31ai_1.pex.spice
* Created: Wed Sep  2 12:25:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O31AI_1%A1 1 3 6 8 13
c23 8 0 1.68631e-19 $X=0.24 $Y=1.295
r24 13 14 3.8254 $w=3.15e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.52 $Y2=1.385
r25 11 13 34.4286 $w=3.15e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.385
+ $X2=0.495 $Y2=1.385
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r27 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r28 4 14 15.85 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.55 $X2=0.52
+ $Y2=1.385
r29 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.52 $Y=1.55 $X2=0.52
+ $Y2=2.4
r30 1 13 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r31 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%A2 3 7 9 10 11 12 18 19
c40 18 0 1.68631e-19 $X=1.015 $Y=1.465
r41 18 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.465
+ $X2=1.015 $Y2=1.63
r42 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.465
+ $X2=1.015 $Y2=1.3
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.465 $X2=1.015 $Y2=1.465
r44 11 12 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.892 $Y=2.405
+ $X2=0.892 $Y2=2.775
r45 10 11 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.892 $Y=2.035
+ $X2=0.892 $Y2=2.405
r46 9 10 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.892 $Y=1.665
+ $X2=0.892 $Y2=2.035
r47 9 19 4.16027 $w=5.73e-07 $l=2e-07 $layer=LI1_cond $X=0.892 $Y=1.665
+ $X2=0.892 $Y2=1.465
r48 7 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.94 $Y=2.4 $X2=0.94
+ $Y2=1.63
r49 3 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=0.74
+ $X2=0.925 $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%A3 3 7 9 13
c34 13 0 1.76087e-19 $X=1.855 $Y=1.515
r35 13 15 5.80723 $w=2.49e-07 $l=3e-08 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.885 $Y2=1.515
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.515 $X2=1.855 $Y2=1.515
r37 9 14 8.1743 $w=4.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.855 $Y2=1.565
r38 5 15 14.627 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.35
+ $X2=1.885 $Y2=1.515
r39 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.885 $Y=1.35
+ $X2=1.885 $Y2=0.74
r40 1 13 66.7831 $w=2.49e-07 $l=4.19464e-07 $layer=POLY_cond $X=1.51 $Y=1.68
+ $X2=1.855 $Y2=1.515
r41 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.51 $Y=1.68 $X2=1.51
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%B1 3 7 9 15 16
c26 16 0 1.76087e-19 $X=2.61 $Y=1.465
c27 3 0 1.49438e-20 $X=2.335 $Y=0.74
r28 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.465 $X2=2.61 $Y2=1.465
r29 13 15 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=2.35 $Y=1.465
+ $X2=2.61 $Y2=1.465
r30 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.335 $Y=1.465
+ $X2=2.35 $Y2=1.465
r31 9 16 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.61 $Y=1.665 $X2=2.61
+ $Y2=1.465
r32 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.63
+ $X2=2.35 $Y2=1.465
r33 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.35 $Y=1.63 $X2=2.35
+ $Y2=2.4
r34 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.3
+ $X2=2.335 $Y2=1.465
r35 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.335 $Y=1.3 $X2=2.335
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%VPWR 1 2 7 9 13 15 19 21 34
r27 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 22 30 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33 $X2=0.19
+ $Y2=3.33
r35 22 24 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 21 33 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.645 $Y2=3.33
r37 21 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 19 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 19 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.575 $Y=2.115
+ $X2=2.575 $Y2=2.815
r41 13 33 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.645 $Y2=3.33
r42 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=2.815
r43 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.255 $Y=1.985
+ $X2=0.255 $Y2=2.815
r44 7 30 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.19 $Y2=3.33
r45 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r46 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.84 $X2=2.575 $Y2=2.815
r47 2 15 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.84 $X2=2.575 $Y2=2.115
r48 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.815
r49 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%Y 1 2 9 10 13 15 16 20 21
r42 20 21 12.1537 $w=8.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=2.115
+ $X2=1.79 $Y2=1.95
r43 15 16 5.12955 $w=8.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=1.79 $Y2=2.775
r44 15 20 4.02045 $w=8.78e-07 $l=2.9e-07 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=1.79 $Y2=2.115
r45 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.6 $Y=0.96 $X2=2.6
+ $Y2=0.515
r46 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.435 $Y=1.045
+ $X2=2.6 $Y2=0.96
r47 9 10 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.435 $Y=1.045
+ $X2=1.52 $Y2=1.045
r48 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.435 $Y=1.13
+ $X2=1.52 $Y2=1.045
r49 7 21 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.435 $Y=1.13
+ $X2=1.435 $Y2=1.95
r50 2 16 200 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=3 $X=1.6
+ $Y=1.84 $X2=1.735 $Y2=2.815
r51 2 20 200 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=3 $X=1.6
+ $Y=1.84 $X2=1.735 $Y2=2.115
r52 1 13 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.41
+ $Y=0.37 $X2=2.6 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%VGND 1 2 7 9 11 20 21 29 35
r36 33 35 7.72401 $w=5.33e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=0.182
+ $X2=1.755 $Y2=0.182
r37 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r38 31 33 2.01209 $w=5.33e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=0.182 $X2=1.68
+ $Y2=0.182
r39 27 31 8.71908 $w=5.33e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=0.182
+ $X2=1.59 $Y2=0.182
r40 27 29 9.28897 $w=5.33e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=0.182
+ $X2=1.055 $Y2=0.182
r41 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 21 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r44 20 35 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=1.755
+ $Y2=0
r45 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r47 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r48 16 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.055
+ $Y2=0
r49 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 14 24 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r51 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r52 11 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r53 11 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r54 7 24 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r55 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r56 2 31 91 $w=1.7e-07 $l=5.92495e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.59 $Y2=0.365
r57 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31AI_1%A_114_74# 1 2 9 12 14 16
c31 9 0 1.49438e-20 $X=1.935 $Y=0.705
r32 16 18 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.1 $Y=0.57 $X2=2.1
+ $Y2=0.705
r33 12 14 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.75 $Y=0.515
+ $X2=0.75 $Y2=0.705
r34 10 14 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0.705
+ $X2=0.75 $Y2=0.705
r35 9 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0.705
+ $X2=2.1 $Y2=0.705
r36 9 10 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.935 $Y=0.705
+ $X2=0.875 $Y2=0.705
r37 2 16 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.37 $X2=2.1 $Y2=0.57
r38 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends


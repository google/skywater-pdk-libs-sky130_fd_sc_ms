* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
M1000 Y a_231_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.2544e+12p pd=1.12e+07u as=2.8737e+12p ps=1.85e+07u
M1001 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_373_74# a_231_74# a_678_74# VNB nlowvt w=740000u l=150000u
+  ad=8.504e+11p pd=6.86e+06u as=4.662e+11p ps=4.22e+06u
M1003 Y a_27_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_231_74# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_231_74# B_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=5.278e+11p ps=4.3e+06u
M1006 a_886_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=0p ps=0u
M1007 VPWR a_27_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y D VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_886_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A_N a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_373_74# a_27_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.257e+11p ps=2.09e+06u
M1013 a_886_74# C a_678_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR D Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_678_74# a_231_74# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_27_368# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_231_74# B_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.8e+11p pd=2.76e+06u as=0p ps=0u
M1018 VGND A_N a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1019 a_678_74# C a_886_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

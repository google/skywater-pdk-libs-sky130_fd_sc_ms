* File: sky130_fd_sc_ms__o211ai_2.pxi.spice
* Created: Fri Aug 28 17:53:22 2020
* 
x_PM_SKY130_FD_SC_MS__O211AI_2%C1 N_C1_M1001_g N_C1_M1008_g N_C1_M1002_g
+ N_C1_M1009_g C1 N_C1_c_90_n N_C1_c_91_n PM_SKY130_FD_SC_MS__O211AI_2%C1
x_PM_SKY130_FD_SC_MS__O211AI_2%B1 N_B1_M1011_g N_B1_M1000_g N_B1_M1014_g
+ N_B1_M1015_g B1 B1 N_B1_c_135_n N_B1_c_136_n PM_SKY130_FD_SC_MS__O211AI_2%B1
x_PM_SKY130_FD_SC_MS__O211AI_2%A2 N_A2_M1007_g N_A2_M1003_g N_A2_M1010_g
+ N_A2_M1005_g A2 A2 N_A2_c_190_n N_A2_c_191_n N_A2_c_192_n
+ PM_SKY130_FD_SC_MS__O211AI_2%A2
x_PM_SKY130_FD_SC_MS__O211AI_2%A1 N_A1_M1012_g N_A1_M1004_g N_A1_M1006_g
+ N_A1_M1013_g A1 N_A1_c_248_n N_A1_c_249_n PM_SKY130_FD_SC_MS__O211AI_2%A1
x_PM_SKY130_FD_SC_MS__O211AI_2%VPWR N_VPWR_M1008_s N_VPWR_M1009_s N_VPWR_M1014_s
+ N_VPWR_M1012_s N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n
+ N_VPWR_c_296_n N_VPWR_c_297_n VPWR N_VPWR_c_298_n N_VPWR_c_299_n
+ N_VPWR_c_300_n N_VPWR_c_291_n N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n
+ PM_SKY130_FD_SC_MS__O211AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O211AI_2%Y N_Y_M1001_s N_Y_M1008_d N_Y_M1011_d N_Y_M1007_d
+ N_Y_c_360_n N_Y_c_354_n N_Y_c_367_n N_Y_c_357_n N_Y_c_358_n N_Y_c_355_n
+ N_Y_c_372_n N_Y_c_384_n N_Y_c_392_n Y Y PM_SKY130_FD_SC_MS__O211AI_2%Y
x_PM_SKY130_FD_SC_MS__O211AI_2%A_505_368# N_A_505_368#_M1007_s
+ N_A_505_368#_M1010_s N_A_505_368#_M1013_d N_A_505_368#_c_417_n
+ N_A_505_368#_c_418_n N_A_505_368#_c_419_n N_A_505_368#_c_420_n
+ N_A_505_368#_c_421_n N_A_505_368#_c_422_n N_A_505_368#_c_423_n
+ PM_SKY130_FD_SC_MS__O211AI_2%A_505_368#
x_PM_SKY130_FD_SC_MS__O211AI_2%A_30_84# N_A_30_84#_M1001_d N_A_30_84#_M1002_d
+ N_A_30_84#_M1015_s N_A_30_84#_c_455_n N_A_30_84#_c_456_n N_A_30_84#_c_457_n
+ N_A_30_84#_c_458_n N_A_30_84#_c_459_n PM_SKY130_FD_SC_MS__O211AI_2%A_30_84#
x_PM_SKY130_FD_SC_MS__O211AI_2%A_303_84# N_A_303_84#_M1000_d N_A_303_84#_M1003_s
+ N_A_303_84#_M1004_d N_A_303_84#_c_493_n N_A_303_84#_c_494_n
+ N_A_303_84#_c_495_n N_A_303_84#_c_496_n N_A_303_84#_c_497_n
+ N_A_303_84#_c_498_n PM_SKY130_FD_SC_MS__O211AI_2%A_303_84#
x_PM_SKY130_FD_SC_MS__O211AI_2%VGND N_VGND_M1003_d N_VGND_M1005_d N_VGND_M1006_s
+ N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n VGND
+ N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n
+ N_VGND_c_549_n PM_SKY130_FD_SC_MS__O211AI_2%VGND
cc_1 VNB N_C1_M1001_g 0.0263047f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.79
cc_2 VNB N_C1_M1002_g 0.0196764f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_3 VNB N_C1_M1009_g 0.00157753f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_4 VNB N_C1_c_90_n 0.0165723f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_5 VNB N_C1_c_91_n 0.0557289f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.515
cc_6 VNB N_B1_M1000_g 0.0212084f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_7 VNB N_B1_M1015_g 0.0270227f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_8 VNB N_B1_c_135_n 0.00829772f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_9 VNB N_B1_c_136_n 0.0365174f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_10 VNB N_A2_M1007_g 5.45338e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.79
cc_11 VNB N_A2_M1003_g 0.0288139f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_12 VNB N_A2_M1010_g 4.92613e-19 $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_13 VNB N_A2_M1005_g 0.0215493f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_14 VNB A2 0.00374074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_190_n 0.0383468f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_16 VNB N_A2_c_191_n 0.0334943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_192_n 0.00344733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1012_g 5.13153e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.79
cc_19 VNB N_A1_M1004_g 0.0211184f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_20 VNB N_A1_M1006_g 0.0256402f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_21 VNB N_A1_M1013_g 7.75396e-19 $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_22 VNB A1 0.0263416f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_23 VNB N_A1_c_248_n 0.0780743f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_24 VNB N_A1_c_249_n 0.00232983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_291_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_354_n 0.00148201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_355_n 0.00410134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_30_84#_c_455_n 0.0296889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_30_84#_c_456_n 0.00482743f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_30 VNB N_A_30_84#_c_457_n 0.00951014f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_31 VNB N_A_30_84#_c_458_n 0.0119635f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_32 VNB N_A_30_84#_c_459_n 0.00572319f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.515
cc_33 VNB N_A_303_84#_c_493_n 0.0174175f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.79
cc_34 VNB N_A_303_84#_c_494_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.4
cc_35 VNB N_A_303_84#_c_495_n 0.00814736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_303_84#_c_496_n 0.00229554f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_37 VNB N_A_303_84#_c_497_n 0.00243322f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.515
cc_38 VNB N_A_303_84#_c_498_n 0.00126893f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_39 VNB N_VGND_c_540_n 0.0103499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_541_n 0.00257504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_542_n 0.0125081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_543_n 0.0342758f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_43 VNB N_VGND_c_544_n 0.0629405f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.515
cc_44 VNB N_VGND_c_545_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_546_n 0.016335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_547_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_548_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_549_n 0.289293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_C1_M1008_g 0.0249926f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_50 VPB N_C1_M1009_g 0.0228982f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_51 VPB N_C1_c_90_n 0.00965371f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_52 VPB N_C1_c_91_n 0.00819868f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.515
cc_53 VPB N_B1_M1011_g 0.0208406f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.79
cc_54 VPB N_B1_M1014_g 0.0246451f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.79
cc_55 VPB N_B1_c_135_n 0.00800118f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.515
cc_56 VPB N_B1_c_136_n 0.00596533f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_57 VPB N_A2_M1007_g 0.0263624f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.79
cc_58 VPB N_A2_M1010_g 0.0218935f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=0.79
cc_59 VPB A2 0.00342514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A2_c_192_n 0.00482195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A1_M1012_g 0.0227456f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.79
cc_62 VPB N_A1_M1013_g 0.0317389f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_63 VPB N_VPWR_c_292_n 0.0116091f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.63
cc_64 VPB N_VPWR_c_293_n 0.0495763f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_65 VPB N_VPWR_c_294_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_66 VPB N_VPWR_c_295_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.515
cc_67 VPB N_VPWR_c_296_n 0.0149195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_297_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_298_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_299_n 0.0389588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_300_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_291_n 0.0792231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_302_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_303_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_304_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_Y_c_354_n 0.00250791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_Y_c_357_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.515
cc_78 VPB N_Y_c_358_n 0.0167585f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.515
cc_79 VPB Y 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_505_368#_c_417_n 0.0055433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_505_368#_c_418_n 0.00473643f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_82 VPB N_A_505_368#_c_419_n 0.00376758f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=2.4
cc_83 VPB N_A_505_368#_c_420_n 0.00316801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_505_368#_c_421_n 0.00310192f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_85 VPB N_A_505_368#_c_422_n 0.00898246f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.515
cc_86 VPB N_A_505_368#_c_423_n 0.0401925f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.515
cc_87 N_C1_M1009_g N_B1_M1011_g 0.0235602f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_88 N_C1_M1002_g N_B1_M1000_g 0.0214079f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_89 N_C1_c_91_n N_B1_c_135_n 0.0045463f $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_90 N_C1_c_91_n N_B1_c_136_n 0.0235602f $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_91 N_C1_M1008_g N_VPWR_c_293_n 0.00501904f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_92 N_C1_c_90_n N_VPWR_c_293_n 0.0217879f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_93 N_C1_c_91_n N_VPWR_c_293_n 0.0010552f $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_94 N_C1_M1008_g N_VPWR_c_294_n 0.005209f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_95 N_C1_M1009_g N_VPWR_c_294_n 0.005209f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_96 N_C1_M1009_g N_VPWR_c_295_n 0.0027763f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_97 N_C1_M1008_g N_VPWR_c_291_n 0.00986107f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_98 N_C1_M1009_g N_VPWR_c_291_n 0.00982376f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_99 N_C1_M1001_g N_Y_c_360_n 0.00489796f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_100 N_C1_M1002_g N_Y_c_360_n 0.00460661f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_101 N_C1_M1001_g N_Y_c_354_n 0.002587f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_102 N_C1_M1002_g N_Y_c_354_n 0.00463156f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_103 N_C1_M1009_g N_Y_c_354_n 0.00313006f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_104 N_C1_c_90_n N_Y_c_354_n 0.0318657f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_105 N_C1_c_91_n N_Y_c_354_n 0.0181656f $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_106 N_C1_M1009_g N_Y_c_367_n 0.017337f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_107 N_C1_M1009_g N_Y_c_357_n 6.50516e-19 $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_108 N_C1_M1001_g N_Y_c_355_n 0.00325382f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_109 N_C1_M1002_g N_Y_c_355_n 0.00190678f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_110 N_C1_c_91_n N_Y_c_355_n 0.00210354f $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_111 N_C1_M1008_g N_Y_c_372_n 0.00364186f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_112 N_C1_M1009_g N_Y_c_372_n 0.00196977f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_113 N_C1_M1008_g Y 0.0112644f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_114 N_C1_M1009_g Y 0.0119382f $X=0.985 $Y=2.4 $X2=0 $Y2=0
cc_115 N_C1_M1001_g N_A_30_84#_c_455_n 0.00159319f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_116 N_C1_c_90_n N_A_30_84#_c_455_n 0.0217837f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_117 N_C1_c_91_n N_A_30_84#_c_455_n 0.00125844f $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_118 N_C1_M1001_g N_A_30_84#_c_456_n 0.0141481f $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_119 N_C1_M1002_g N_A_30_84#_c_456_n 0.0134522f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_120 N_C1_M1002_g N_A_30_84#_c_459_n 0.00240868f $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_121 N_C1_c_91_n N_A_30_84#_c_459_n 6.77396e-19 $X=0.94 $Y=1.515 $X2=0 $Y2=0
cc_122 N_C1_M1001_g N_VGND_c_544_n 8.76084e-19 $X=0.51 $Y=0.79 $X2=0 $Y2=0
cc_123 N_C1_M1002_g N_VGND_c_544_n 8.76084e-19 $X=0.94 $Y=0.79 $X2=0 $Y2=0
cc_124 N_B1_M1015_g N_A2_c_190_n 0.00856729f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_125 N_B1_c_135_n N_A2_c_190_n 3.61578e-19 $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_126 N_B1_M1014_g N_A2_c_192_n 6.44754e-19 $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B1_c_135_n N_A2_c_192_n 0.0184224f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_128 N_B1_c_136_n N_A2_c_192_n 5.69806e-19 $X=1.94 $Y=1.515 $X2=0 $Y2=0
cc_129 N_B1_M1011_g N_VPWR_c_295_n 0.0027763f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_130 N_B1_M1014_g N_VPWR_c_296_n 0.00501904f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_131 N_B1_M1011_g N_VPWR_c_298_n 0.005209f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_132 N_B1_M1014_g N_VPWR_c_298_n 0.005209f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_133 N_B1_M1011_g N_VPWR_c_291_n 0.00982376f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_134 N_B1_M1014_g N_VPWR_c_291_n 0.00987399f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_135 N_B1_M1000_g N_Y_c_354_n 7.9877e-19 $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_136 N_B1_c_135_n N_Y_c_354_n 0.0317179f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_137 N_B1_M1011_g N_Y_c_367_n 0.0128923f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_138 N_B1_c_135_n N_Y_c_367_n 0.027843f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_139 N_B1_M1011_g N_Y_c_357_n 0.0119382f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B1_M1014_g N_Y_c_357_n 0.0166062f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_141 N_B1_M1014_g N_Y_c_358_n 0.0150541f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_142 N_B1_c_135_n N_Y_c_358_n 0.012644f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B1_M1011_g N_Y_c_384_n 8.84614e-19 $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_144 N_B1_M1014_g N_Y_c_384_n 8.84614e-19 $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_145 N_B1_c_135_n N_Y_c_384_n 0.0235495f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_146 N_B1_c_136_n N_Y_c_384_n 5.54777e-19 $X=1.94 $Y=1.515 $X2=0 $Y2=0
cc_147 N_B1_M1011_g Y 6.50516e-19 $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_148 N_B1_M1000_g N_A_30_84#_c_458_n 0.0168204f $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_149 N_B1_M1015_g N_A_30_84#_c_458_n 0.0198009f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_150 N_B1_c_135_n N_A_30_84#_c_458_n 0.00395247f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_151 N_B1_M1000_g N_A_30_84#_c_459_n 0.0105901f $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_152 N_B1_M1015_g N_A_30_84#_c_459_n 6.5477e-19 $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_153 N_B1_c_135_n N_A_30_84#_c_459_n 0.0271148f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_154 N_B1_c_136_n N_A_30_84#_c_459_n 5.44797e-19 $X=1.94 $Y=1.515 $X2=0 $Y2=0
cc_155 N_B1_M1015_g N_A_303_84#_c_493_n 0.00994167f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_156 N_B1_c_135_n N_A_303_84#_c_493_n 0.00797813f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_157 N_B1_M1000_g N_A_303_84#_c_497_n 0.0015116f $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_158 N_B1_M1015_g N_A_303_84#_c_497_n 0.00598046f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_159 N_B1_c_135_n N_A_303_84#_c_497_n 0.0261926f $X=1.85 $Y=1.515 $X2=0 $Y2=0
cc_160 N_B1_c_136_n N_A_303_84#_c_497_n 0.0041721f $X=1.94 $Y=1.515 $X2=0 $Y2=0
cc_161 N_B1_M1015_g N_VGND_c_540_n 0.0023272f $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_162 N_B1_M1000_g N_VGND_c_544_n 8.94875e-19 $X=1.44 $Y=0.79 $X2=0 $Y2=0
cc_163 N_B1_M1015_g N_VGND_c_544_n 8.76084e-19 $X=1.94 $Y=0.79 $X2=0 $Y2=0
cc_164 N_A2_M1010_g N_A1_M1012_g 0.0169146f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A2_M1005_g N_A1_M1004_g 0.0299183f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A2_M1005_g N_A1_c_248_n 0.0196111f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_167 A2 N_A1_c_248_n 4.12017e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_168 A2 N_A1_c_249_n 0.0210188f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A2_c_191_n N_A1_c_249_n 4.12009e-19 $X=3.37 $Y=1.485 $X2=0 $Y2=0
cc_170 N_A2_M1007_g N_VPWR_c_296_n 8.64401e-19 $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A2_M1007_g N_VPWR_c_299_n 0.00333926f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A2_M1010_g N_VPWR_c_299_n 0.00333926f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A2_M1007_g N_VPWR_c_291_n 0.0042782f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A2_M1010_g N_VPWR_c_291_n 0.00422798f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A2_M1007_g N_Y_c_358_n 0.0150541f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A2_c_190_n N_Y_c_358_n 0.00178623f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_177 N_A2_c_192_n N_Y_c_358_n 0.0386558f $X=3.005 $Y=1.55 $X2=0 $Y2=0
cc_178 N_A2_M1007_g N_Y_c_392_n 0.0150733f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A2_M1010_g N_Y_c_392_n 0.0110375f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_180 A2 N_Y_c_392_n 0.0191677f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A2_c_191_n N_Y_c_392_n 5.16252e-19 $X=3.37 $Y=1.485 $X2=0 $Y2=0
cc_182 N_A2_c_192_n N_Y_c_392_n 0.00324682f $X=3.005 $Y=1.55 $X2=0 $Y2=0
cc_183 N_A2_M1007_g N_A_505_368#_c_418_n 0.01495f $X=2.895 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A2_M1010_g N_A_505_368#_c_418_n 0.0137017f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A2_M1010_g N_A_505_368#_c_420_n 6.10014e-19 $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A2_M1003_g N_A_30_84#_c_458_n 0.00137242f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A2_M1003_g N_A_303_84#_c_493_n 0.0147855f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_188 A2 N_A_303_84#_c_493_n 0.00496209f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_c_190_n N_A_303_84#_c_493_n 0.009857f $X=2.805 $Y=1.485 $X2=0 $Y2=0
cc_190 N_A2_c_192_n N_A_303_84#_c_493_n 0.0433508f $X=3.005 $Y=1.55 $X2=0 $Y2=0
cc_191 N_A2_M1003_g N_A_303_84#_c_494_n 3.92313e-19 $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A2_M1005_g N_A_303_84#_c_494_n 3.92313e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A2_M1005_g N_A_303_84#_c_495_n 0.0127221f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_194 A2 N_A_303_84#_c_495_n 0.0148851f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_195 A2 N_A_303_84#_c_498_n 0.0147323f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A2_c_191_n N_A_303_84#_c_498_n 7.87695e-19 $X=3.37 $Y=1.485 $X2=0 $Y2=0
cc_197 N_A2_M1003_g N_VGND_c_540_n 0.0112914f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_M1005_g N_VGND_c_540_n 4.58208e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A2_M1003_g N_VGND_c_541_n 4.58208e-19 $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_M1005_g N_VGND_c_541_n 0.0096639f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_M1003_g N_VGND_c_545_n 0.00383152f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A2_M1005_g N_VGND_c_545_n 0.00383152f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_M1003_g N_VGND_c_549_n 0.0075754f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A2_M1005_g N_VGND_c_549_n 0.0075754f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_M1012_g N_VPWR_c_297_n 0.0147538f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A1_M1013_g N_VPWR_c_297_n 0.00387724f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A1_M1012_g N_VPWR_c_299_n 0.00460063f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A1_M1013_g N_VPWR_c_300_n 0.005209f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_M1012_g N_VPWR_c_291_n 0.00908665f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A1_M1013_g N_VPWR_c_291_n 0.00985824f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A1_M1012_g N_A_505_368#_c_418_n 0.00101073f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_M1012_g N_A_505_368#_c_421_n 0.0147251f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A1_M1013_g N_A_505_368#_c_421_n 0.0132272f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A1_c_248_n N_A_505_368#_c_421_n 0.00363102f $X=4.295 $Y=1.475 $X2=0
+ $Y2=0
cc_215 N_A1_c_249_n N_A_505_368#_c_421_n 0.0490884f $X=4.365 $Y=1.415 $X2=0
+ $Y2=0
cc_216 N_A1_M1013_g N_A_505_368#_c_422_n 0.0012834f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A1_c_248_n N_A_505_368#_c_422_n 0.00225013f $X=4.295 $Y=1.475 $X2=0
+ $Y2=0
cc_218 N_A1_c_249_n N_A_505_368#_c_422_n 0.0296207f $X=4.365 $Y=1.415 $X2=0
+ $Y2=0
cc_219 N_A1_M1012_g N_A_505_368#_c_423_n 9.71985e-19 $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A1_M1013_g N_A_505_368#_c_423_n 0.0142717f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A1_M1004_g N_A_303_84#_c_495_n 0.0128457f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1006_g N_A_303_84#_c_495_n 0.00127757f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_c_248_n N_A_303_84#_c_495_n 0.00465862f $X=4.295 $Y=1.475 $X2=0
+ $Y2=0
cc_224 N_A1_c_249_n N_A_303_84#_c_495_n 0.0371669f $X=4.365 $Y=1.415 $X2=0 $Y2=0
cc_225 N_A1_M1004_g N_A_303_84#_c_496_n 4.44262e-19 $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1006_g N_A_303_84#_c_496_n 4.4892e-19 $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1004_g N_VGND_c_541_n 0.00949565f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1006_g N_VGND_c_541_n 4.51649e-19 $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1004_g N_VGND_c_543_n 4.93565e-19 $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1006_g N_VGND_c_543_n 0.0124427f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_231 A1 N_VGND_c_543_n 0.0263105f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_232 N_A1_c_248_n N_VGND_c_543_n 0.00176634f $X=4.295 $Y=1.475 $X2=0 $Y2=0
cc_233 N_A1_c_249_n N_VGND_c_543_n 0.00136555f $X=4.365 $Y=1.415 $X2=0 $Y2=0
cc_234 N_A1_M1004_g N_VGND_c_546_n 0.00398535f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1006_g N_VGND_c_546_n 0.00383152f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1004_g N_VGND_c_549_n 0.00787968f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1006_g N_VGND_c_549_n 0.00757973f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_238 N_VPWR_M1009_s N_Y_c_367_n 0.00332066f $X=1.075 $Y=1.84 $X2=0 $Y2=0
cc_239 N_VPWR_c_295_n N_Y_c_367_n 0.0126919f $X=1.21 $Y=2.455 $X2=0 $Y2=0
cc_240 N_VPWR_c_295_n N_Y_c_357_n 0.0233699f $X=1.21 $Y=2.455 $X2=0 $Y2=0
cc_241 N_VPWR_c_296_n N_Y_c_357_n 0.0234083f $X=2.11 $Y=2.455 $X2=0 $Y2=0
cc_242 N_VPWR_c_298_n N_Y_c_357_n 0.0144623f $X=2.025 $Y=3.33 $X2=0 $Y2=0
cc_243 N_VPWR_c_291_n N_Y_c_357_n 0.0118344f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_M1014_s N_Y_c_358_n 0.0118091f $X=1.975 $Y=1.84 $X2=0 $Y2=0
cc_245 N_VPWR_c_296_n N_Y_c_358_n 0.0197477f $X=2.11 $Y=2.455 $X2=0 $Y2=0
cc_246 N_VPWR_c_293_n Y 0.0289761f $X=0.31 $Y=2.115 $X2=0 $Y2=0
cc_247 N_VPWR_c_294_n Y 0.0144623f $X=1.125 $Y=3.33 $X2=0 $Y2=0
cc_248 N_VPWR_c_295_n Y 0.0233699f $X=1.21 $Y=2.455 $X2=0 $Y2=0
cc_249 N_VPWR_c_291_n Y 0.0118344f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_250 N_VPWR_c_296_n N_A_505_368#_c_417_n 0.0397231f $X=2.11 $Y=2.455 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_297_n N_A_505_368#_c_418_n 0.0103602f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_299_n N_A_505_368#_c_418_n 0.0581059f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_291_n N_A_505_368#_c_418_n 0.0324093f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_296_n N_A_505_368#_c_419_n 0.011925f $X=2.11 $Y=2.455 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_299_n N_A_505_368#_c_419_n 0.0179217f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_291_n N_A_505_368#_c_419_n 0.00971942f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_M1012_s N_A_505_368#_c_421_n 0.00218982f $X=3.885 $Y=1.84 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_297_n N_A_505_368#_c_421_n 0.0189268f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_297_n N_A_505_368#_c_423_n 0.0315588f $X=4.02 $Y=2.325 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_300_n N_A_505_368#_c_423_n 0.014549f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_291_n N_A_505_368#_c_423_n 0.0119743f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_Y_c_358_n N_A_505_368#_M1007_s 0.00526196f $X=2.955 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_263 N_Y_c_358_n N_A_505_368#_c_417_n 0.0197477f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_264 N_Y_M1007_d N_A_505_368#_c_418_n 0.00165831f $X=2.985 $Y=1.84 $X2=0 $Y2=0
cc_265 N_Y_c_392_n N_A_505_368#_c_418_n 0.0159318f $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_266 N_Y_c_360_n N_A_30_84#_c_455_n 0.0216593f $X=0.725 $Y=0.68 $X2=0 $Y2=0
cc_267 N_Y_M1001_s N_A_30_84#_c_456_n 0.00176461f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_268 N_Y_c_360_n N_A_30_84#_c_456_n 0.0158928f $X=0.725 $Y=0.68 $X2=0 $Y2=0
cc_269 N_Y_c_360_n N_A_30_84#_c_459_n 0.017638f $X=0.725 $Y=0.68 $X2=0 $Y2=0
cc_270 N_A_505_368#_c_420_n N_A_303_84#_c_495_n 0.00549175f $X=3.57 $Y=1.99
+ $X2=0 $Y2=0
cc_271 N_A_505_368#_c_421_n N_A_303_84#_c_495_n 8.52231e-19 $X=4.355 $Y=1.905
+ $X2=0 $Y2=0
cc_272 N_A_30_84#_c_458_n N_A_303_84#_M1000_d 0.00244396f $X=2.16 $Y=0.565
+ $X2=-0.19 $Y2=-0.245
cc_273 N_A_30_84#_M1015_s N_A_303_84#_c_493_n 0.0131383f $X=2.015 $Y=0.42 $X2=0
+ $Y2=0
cc_274 N_A_30_84#_c_458_n N_A_303_84#_c_493_n 0.0220402f $X=2.16 $Y=0.565 $X2=0
+ $Y2=0
cc_275 N_A_30_84#_c_458_n N_A_303_84#_c_497_n 0.0210984f $X=2.16 $Y=0.565 $X2=0
+ $Y2=0
cc_276 N_A_30_84#_c_459_n N_A_303_84#_c_497_n 0.0112335f $X=1.225 $Y=0.565 $X2=0
+ $Y2=0
cc_277 N_A_30_84#_c_458_n N_VGND_c_540_n 0.0338381f $X=2.16 $Y=0.565 $X2=0 $Y2=0
cc_278 N_A_30_84#_c_456_n N_VGND_c_544_n 0.0437462f $X=1.06 $Y=0.34 $X2=0 $Y2=0
cc_279 N_A_30_84#_c_457_n N_VGND_c_544_n 0.0179217f $X=0.38 $Y=0.34 $X2=0 $Y2=0
cc_280 N_A_30_84#_c_458_n N_VGND_c_544_n 0.065133f $X=2.16 $Y=0.565 $X2=0 $Y2=0
cc_281 N_A_30_84#_c_459_n N_VGND_c_544_n 0.0236566f $X=1.225 $Y=0.565 $X2=0
+ $Y2=0
cc_282 N_A_30_84#_c_456_n N_VGND_c_549_n 0.0255585f $X=1.06 $Y=0.34 $X2=0 $Y2=0
cc_283 N_A_30_84#_c_457_n N_VGND_c_549_n 0.00971942f $X=0.38 $Y=0.34 $X2=0 $Y2=0
cc_284 N_A_30_84#_c_458_n N_VGND_c_549_n 0.0361835f $X=2.16 $Y=0.565 $X2=0 $Y2=0
cc_285 N_A_30_84#_c_459_n N_VGND_c_549_n 0.0128296f $X=1.225 $Y=0.565 $X2=0
+ $Y2=0
cc_286 N_A_303_84#_c_493_n N_VGND_M1003_d 0.00326148f $X=3.07 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_303_84#_c_495_n N_VGND_M1005_d 0.00188382f $X=3.935 $Y=1.065 $X2=0
+ $Y2=0
cc_288 N_A_303_84#_c_493_n N_VGND_c_540_n 0.0205937f $X=3.07 $Y=1.065 $X2=0
+ $Y2=0
cc_289 N_A_303_84#_c_494_n N_VGND_c_540_n 0.016636f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_290 N_A_303_84#_c_494_n N_VGND_c_541_n 0.016636f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_291 N_A_303_84#_c_495_n N_VGND_c_541_n 0.0160414f $X=3.935 $Y=1.065 $X2=0
+ $Y2=0
cc_292 N_A_303_84#_c_496_n N_VGND_c_541_n 0.0163061f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
cc_293 N_A_303_84#_c_496_n N_VGND_c_543_n 0.0246508f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
cc_294 N_A_303_84#_c_494_n N_VGND_c_545_n 0.00749631f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_295 N_A_303_84#_c_496_n N_VGND_c_546_n 0.00995046f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0
cc_296 N_A_303_84#_c_494_n N_VGND_c_549_n 0.0062048f $X=3.155 $Y=0.515 $X2=0
+ $Y2=0
cc_297 N_A_303_84#_c_496_n N_VGND_c_549_n 0.00823613f $X=4.02 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__nand4b_2.spice
* Created: Wed Sep  2 12:14:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4b_2.pex.spice"
.subckt sky130_fd_sc_ms__nand4b_2  VNB VPB A_N B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_N_M1010_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1726 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_225_74#_M1002_d N_A_27_74#_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1962 AS=0.1147 PD=2.05 PS=1.05 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1015 N_A_225_74#_M1015_d N_A_27_74#_M1015_g N_Y_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1147 PD=1.02 PS=1.05 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_225_74#_M1015_d N_B_M1001_g N_A_490_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1773 PD=1.02 PS=1.28 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_A_225_74#_M1007_d N_B_M1007_g N_A_490_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.197775 AS=0.1773 PD=2.05 PS=1.28 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_719_123#_M1000_d N_C_M1000_g N_A_490_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.204075 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1006 N_A_719_123#_M1006_d N_C_M1006_g N_A_490_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 N_A_719_123#_M1006_d N_D_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1005 N_A_719_123#_M1005_d N_D_M1005_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.111 PD=2.05 PS=1.04 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A_N_M1008_g N_A_27_74#_M1008_s VPB PSHORT L=0.18 W=1
+ AD=0.185943 AS=0.28 PD=1.39623 PS=2.56 NRD=16.0752 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1011 N_Y_M1011_d N_A_27_74#_M1011_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.208257 PD=1.39 PS=1.56377 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90004 A=0.2016 P=2.6 MULT=1
MM1016 N_Y_M1011_d N_A_27_74#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3556 PD=1.39 PS=1.755 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90003.6 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1012_d N_B_M1012_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3556 PD=1.39 PS=1.755 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.9 SB=90002.7
+ A=0.2016 P=2.6 MULT=1
MM1017 N_Y_M1012_d N_B_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.4 SB=90002.3
+ A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_C_M1009_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.9 SB=90001.7
+ A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1009_d N_C_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2632 PD=1.39 PS=1.59 NRD=0 NRS=18.4589 M=1 R=6.22222 SA=90003.4
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2632 PD=1.39 PS=1.59 NRD=0 NRS=14.9326 M=1 R=6.22222 SA=90004 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1013 N_Y_M1004_d N_D_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3192 PD=1.39 PS=2.81 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.5 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__nand4b_2.pxi.spice"
*
.ends
*
*

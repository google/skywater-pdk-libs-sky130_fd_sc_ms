* File: sky130_fd_sc_ms__xnor2_1.pxi.spice
* Created: Wed Sep  2 12:33:17 2020
* 
x_PM_SKY130_FD_SC_MS__XNOR2_1%B N_B_c_63_n N_B_M1002_g N_B_c_64_n N_B_M1001_g
+ N_B_M1005_g N_B_M1008_g N_B_c_72_n N_B_c_87_p N_B_c_129_p N_B_c_73_n
+ N_B_c_66_n N_B_c_67_n B N_B_c_68_n PM_SKY130_FD_SC_MS__XNOR2_1%B
x_PM_SKY130_FD_SC_MS__XNOR2_1%A N_A_M1006_g N_A_c_163_n N_A_M1007_g N_A_c_157_n
+ N_A_c_158_n N_A_M1003_g N_A_M1000_g A N_A_c_160_n N_A_c_161_n
+ PM_SKY130_FD_SC_MS__XNOR2_1%A
x_PM_SKY130_FD_SC_MS__XNOR2_1%A_141_385# N_A_141_385#_M1002_d
+ N_A_141_385#_M1007_d N_A_141_385#_M1009_g N_A_141_385#_M1004_g
+ N_A_141_385#_c_223_n N_A_141_385#_c_224_n N_A_141_385#_c_225_n
+ N_A_141_385#_c_230_n N_A_141_385#_c_226_n N_A_141_385#_c_227_n
+ N_A_141_385#_c_228_n PM_SKY130_FD_SC_MS__XNOR2_1%A_141_385#
x_PM_SKY130_FD_SC_MS__XNOR2_1%VPWR N_VPWR_M1007_s N_VPWR_M1001_d N_VPWR_M1009_d
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_315_n VPWR N_VPWR_c_316_n N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_308_n PM_SKY130_FD_SC_MS__XNOR2_1%VPWR
x_PM_SKY130_FD_SC_MS__XNOR2_1%Y N_Y_M1004_d N_Y_M1005_d N_Y_c_364_n N_Y_c_361_n
+ N_Y_c_358_n N_Y_c_359_n N_Y_c_360_n Y N_Y_c_363_n
+ PM_SKY130_FD_SC_MS__XNOR2_1%Y
x_PM_SKY130_FD_SC_MS__XNOR2_1%VGND N_VGND_M1006_s N_VGND_M1000_d N_VGND_c_395_n
+ N_VGND_c_396_n N_VGND_c_397_n VGND N_VGND_c_398_n N_VGND_c_399_n
+ N_VGND_c_400_n N_VGND_c_401_n PM_SKY130_FD_SC_MS__XNOR2_1%VGND
x_PM_SKY130_FD_SC_MS__XNOR2_1%A_293_74# N_A_293_74#_M1000_s N_A_293_74#_M1008_d
+ N_A_293_74#_c_434_n N_A_293_74#_c_433_n N_A_293_74#_c_437_n
+ PM_SKY130_FD_SC_MS__XNOR2_1%A_293_74#
cc_1 VNB N_B_c_63_n 0.0162445f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.31
cc_2 VNB N_B_c_64_n 0.0403713f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.765
cc_3 VNB N_B_M1008_g 0.0257826f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.74
cc_4 VNB N_B_c_66_n 0.0050024f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_5 VNB N_B_c_67_n 0.0223387f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_6 VNB N_B_c_68_n 0.00348558f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.607
cc_7 VNB N_A_M1006_g 0.0615073f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.765
cc_8 VNB N_A_c_157_n 0.10165f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.68
cc_9 VNB N_A_c_158_n 0.011606f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_10 VNB N_A_M1000_g 0.0193389f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.95
cc_11 VNB N_A_c_160_n 0.0301021f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_12 VNB N_A_c_161_n 0.00208705f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_13 VNB N_A_141_385#_M1009_g 0.00174221f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_14 VNB N_A_141_385#_M1004_g 0.0249763f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.74
cc_15 VNB N_A_141_385#_c_223_n 0.00745634f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.95
cc_16 VNB N_A_141_385#_c_224_n 0.0267453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_141_385#_c_225_n 0.00354512f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_18 VNB N_A_141_385#_c_226_n 0.00494238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_141_385#_c_227_n 0.00608349f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.6
cc_20 VNB N_A_141_385#_c_228_n 0.0325947f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.35
cc_21 VNB N_VPWR_c_308_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_358_n 0.027697f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.74
cc_23 VNB N_Y_c_359_n 0.0247615f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.78
cc_24 VNB N_Y_c_360_n 0.0105427f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.035
cc_25 VNB N_VGND_c_395_n 0.0106846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_396_n 0.0498887f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_27 VNB N_VGND_c_397_n 0.00813052f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.74
cc_28 VNB N_VGND_c_398_n 0.0423941f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.95
cc_29 VNB N_VGND_c_399_n 0.0320561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_400_n 0.196578f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_31 VNB N_VGND_c_401_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.35
cc_32 VNB N_A_293_74#_c_433_n 0.00381723f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_33 VPB N_B_c_64_n 0.0112213f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.765
cc_34 VPB N_B_M1001_g 0.0238141f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.345
cc_35 VPB N_B_M1005_g 0.0221369f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=2.4
cc_36 VPB N_B_c_72_n 0.0029942f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.95
cc_37 VPB N_B_c_73_n 0.00144869f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.95
cc_38 VPB N_B_c_66_n 6.49643e-19 $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_39 VPB N_B_c_67_n 0.00544473f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_40 VPB N_B_c_68_n 0.00310203f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.607
cc_41 VPB N_A_M1006_g 0.00332562f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.765
cc_42 VPB N_A_c_163_n 0.0418111f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.345
cc_43 VPB N_A_M1003_g 0.0237232f $X=-0.19 $Y=1.66 $X2=2.39 $Y2=1.35
cc_44 VPB N_A_c_160_n 0.00719193f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_45 VPB N_A_c_161_n 0.00248204f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_46 VPB N_A_141_385#_M1009_g 0.0267699f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=2.4
cc_47 VPB N_A_141_385#_c_230_n 0.00316304f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_48 VPB N_A_141_385#_c_226_n 0.00206422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_309_n 0.0185196f $X=-0.19 $Y=1.66 $X2=2.39 $Y2=1.35
cc_50 VPB N_VPWR_c_310_n 0.00626527f $X=-0.19 $Y=1.66 $X2=2.39 $Y2=0.74
cc_51 VPB N_VPWR_c_311_n 0.0141048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_312_n 0.0417722f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.95
cc_53 VPB N_VPWR_c_313_n 0.0138995f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.68
cc_54 VPB N_VPWR_c_314_n 0.0139106f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_55 VPB N_VPWR_c_315_n 0.0393536f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_56 VPB N_VPWR_c_316_n 0.0271489f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.6
cc_57 VPB N_VPWR_c_317_n 0.0299529f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.607
cc_58 VPB N_VPWR_c_318_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_308_n 0.0804683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_Y_c_361_n 0.0114589f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=2.4
cc_61 VPB N_Y_c_359_n 0.00939072f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.78
cc_62 VPB N_Y_c_363_n 0.00432573f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_63 N_B_c_63_n N_A_M1006_g 0.0574491f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_64 N_B_c_64_n N_A_M1006_g 0.00613719f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_65 N_B_c_64_n N_A_c_163_n 0.00357319f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_66 N_B_M1001_g N_A_c_163_n 0.018872f $X=1.065 $Y=2.345 $X2=0 $Y2=0
cc_67 N_B_c_63_n N_A_c_157_n 0.0103003f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_68 N_B_M1008_g N_A_c_157_n 0.0302512f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_69 N_B_c_64_n N_A_M1003_g 0.00202528f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_70 N_B_M1001_g N_A_M1003_g 0.0128184f $X=1.065 $Y=2.345 $X2=0 $Y2=0
cc_71 N_B_M1005_g N_A_M1003_g 0.0451984f $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_72 N_B_c_72_n N_A_M1003_g 0.00159306f $X=1.26 $Y=1.95 $X2=0 $Y2=0
cc_73 N_B_c_87_p N_A_M1003_g 0.0186908f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_74 N_B_c_73_n N_A_M1003_g 0.00246204f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_75 N_B_c_68_n N_A_M1003_g 2.55756e-19 $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_76 N_B_c_64_n N_A_c_160_n 0.0182538f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B_c_87_p N_A_c_160_n 9.80789e-19 $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_78 N_B_c_66_n N_A_c_160_n 0.0022979f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B_c_67_n N_A_c_160_n 0.0451984f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_80 N_B_c_68_n N_A_c_160_n 0.00152861f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_81 N_B_c_64_n N_A_c_161_n 0.00117724f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_82 N_B_c_87_p N_A_c_161_n 0.0233058f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_83 N_B_c_73_n N_A_c_161_n 0.00747764f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_84 N_B_c_66_n N_A_c_161_n 0.0267388f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B_c_67_n N_A_c_161_n 3.06344e-19 $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B_c_68_n N_A_c_161_n 0.028107f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_87 N_B_M1005_g N_A_141_385#_M1009_g 0.0244077f $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_88 N_B_c_73_n N_A_141_385#_M1009_g 7.77809e-19 $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_89 N_B_c_67_n N_A_141_385#_M1009_g 0.00254364f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B_M1008_g N_A_141_385#_M1004_g 0.0296051f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B_c_63_n N_A_141_385#_c_223_n 0.00760958f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_92 N_B_c_64_n N_A_141_385#_c_224_n 0.00130476f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B_M1008_g N_A_141_385#_c_224_n 0.0111001f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B_c_66_n N_A_141_385#_c_224_n 0.0337543f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_95 N_B_c_67_n N_A_141_385#_c_224_n 0.00474488f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B_c_68_n N_A_141_385#_c_224_n 0.00695518f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_97 N_B_c_63_n N_A_141_385#_c_225_n 0.0161471f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_98 N_B_c_64_n N_A_141_385#_c_225_n 0.00968723f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B_c_68_n N_A_141_385#_c_225_n 0.0226832f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_100 N_B_c_64_n N_A_141_385#_c_230_n 0.00528172f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B_M1001_g N_A_141_385#_c_230_n 0.0206323f $X=1.065 $Y=2.345 $X2=0 $Y2=0
cc_102 N_B_c_68_n N_A_141_385#_c_230_n 0.00354299f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_103 N_B_c_63_n N_A_141_385#_c_226_n 3.17485e-19 $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_104 N_B_c_64_n N_A_141_385#_c_226_n 0.00757095f $X=1.065 $Y=1.765 $X2=0 $Y2=0
cc_105 N_B_M1001_g N_A_141_385#_c_226_n 9.73898e-19 $X=1.065 $Y=2.345 $X2=0
+ $Y2=0
cc_106 N_B_c_72_n N_A_141_385#_c_226_n 0.00497962f $X=1.26 $Y=1.95 $X2=0 $Y2=0
cc_107 N_B_c_68_n N_A_141_385#_c_226_n 0.0262595f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_108 N_B_M1008_g N_A_141_385#_c_227_n 0.00363004f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B_c_66_n N_A_141_385#_c_227_n 0.0226425f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_110 N_B_c_67_n N_A_141_385#_c_227_n 9.00083e-19 $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B_M1008_g N_A_141_385#_c_228_n 0.0210954f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B_c_66_n N_A_141_385#_c_228_n 3.20341e-19 $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_113 N_B_c_72_n N_VPWR_M1001_d 3.71142e-19 $X=1.26 $Y=1.95 $X2=0 $Y2=0
cc_114 N_B_c_87_p N_VPWR_M1001_d 0.0147186f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_115 N_B_c_129_p N_VPWR_M1001_d 0.00667044f $X=1.345 $Y=2.035 $X2=0 $Y2=0
cc_116 N_B_M1001_g N_VPWR_c_313_n 0.00757726f $X=1.065 $Y=2.345 $X2=0 $Y2=0
cc_117 N_B_M1005_g N_VPWR_c_313_n 0.00116997f $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_118 N_B_c_87_p N_VPWR_c_313_n 0.0218557f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_119 N_B_M1005_g N_VPWR_c_315_n 9.75459e-19 $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_120 N_B_M1001_g N_VPWR_c_316_n 0.00516889f $X=1.065 $Y=2.345 $X2=0 $Y2=0
cc_121 N_B_M1005_g N_VPWR_c_317_n 0.00349978f $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B_M1001_g N_VPWR_c_308_n 0.00583598f $X=1.065 $Y=2.345 $X2=0 $Y2=0
cc_123 N_B_M1005_g N_VPWR_c_308_n 0.00430474f $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B_c_87_p A_379_368# 0.00633429f $X=2.015 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_125 N_B_c_73_n A_379_368# 0.00150072f $X=2.1 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_126 N_B_c_66_n N_Y_c_364_n 0.00805994f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_127 N_B_c_67_n N_Y_c_364_n 0.00291447f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_128 N_B_c_66_n N_Y_c_359_n 0.00136308f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_129 N_B_M1005_g N_Y_c_363_n 0.0307534f $X=2.225 $Y=2.4 $X2=0 $Y2=0
cc_130 N_B_c_87_p N_Y_c_363_n 0.00691392f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_131 N_B_c_66_n N_Y_c_363_n 0.00412171f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_132 N_B_c_67_n N_Y_c_363_n 6.13299e-19 $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_133 N_B_c_63_n N_VGND_c_396_n 0.00207013f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_134 N_B_M1008_g N_VGND_c_397_n 0.00452091f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B_M1008_g N_VGND_c_399_n 0.00327917f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_136 N_B_c_63_n N_VGND_c_400_n 9.39239e-19 $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_137 N_B_M1008_g N_VGND_c_400_n 0.00415199f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B_M1008_g N_A_293_74#_c_434_n 0.00969414f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_139 N_B_c_63_n N_A_293_74#_c_433_n 0.00216277f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_140 N_B_M1008_g N_A_293_74#_c_433_n 5.82005e-19 $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_141 N_B_M1008_g N_A_293_74#_c_437_n 0.00488999f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_M1006_g N_A_141_385#_c_223_n 0.00118315f $X=0.485 $Y=0.915 $X2=0
+ $Y2=0
cc_143 N_A_c_157_n N_A_141_385#_c_223_n 0.00622038f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_A_141_385#_c_223_n 0.0040271f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_A_141_385#_c_224_n 0.0145878f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_c_160_n N_A_141_385#_c_224_n 0.00178426f $X=1.68 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A_c_161_n N_A_141_385#_c_224_n 0.0248926f $X=1.68 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_M1006_g N_A_141_385#_c_225_n 8.41489e-19 $X=0.485 $Y=0.915 $X2=0
+ $Y2=0
cc_149 N_A_M1000_g N_A_141_385#_c_225_n 0.00210586f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_c_163_n N_A_141_385#_c_230_n 0.0165343f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_A_141_385#_c_226_n 0.0112389f $X=0.485 $Y=0.915 $X2=0 $Y2=0
cc_152 N_A_c_163_n N_A_141_385#_c_226_n 0.0140571f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_153 N_A_c_163_n N_VPWR_c_309_n 0.00269596f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_154 N_A_c_163_n N_VPWR_c_310_n 0.00221999f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_155 N_A_c_163_n N_VPWR_c_312_n 0.00714651f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_156 N_A_M1003_g N_VPWR_c_313_n 0.015493f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_c_163_n N_VPWR_c_316_n 0.00516889f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_VPWR_c_317_n 0.00460063f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_c_163_n N_VPWR_c_308_n 0.00583598f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_160 N_A_M1003_g N_VPWR_c_308_n 0.00908371f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_M1003_g N_Y_c_363_n 0.00572801f $X=1.805 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_M1006_g N_VGND_c_396_n 0.0288731f $X=0.485 $Y=0.915 $X2=0 $Y2=0
cc_163 N_A_c_158_n N_VGND_c_396_n 0.00763335f $X=0.56 $Y=0.18 $X2=0 $Y2=0
cc_164 N_A_c_157_n N_VGND_c_397_n 0.0100525f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_165 N_A_c_158_n N_VGND_c_398_n 0.0440575f $X=0.56 $Y=0.18 $X2=0 $Y2=0
cc_166 N_A_c_157_n N_VGND_c_400_n 0.0504593f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_167 N_A_c_158_n N_VGND_c_400_n 0.00749832f $X=0.56 $Y=0.18 $X2=0 $Y2=0
cc_168 N_A_M1000_g N_A_293_74#_c_434_n 0.00987582f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_c_157_n N_A_293_74#_c_433_n 0.00435764f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_170 N_A_M1000_g N_A_293_74#_c_433_n 0.00493339f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_M1000_g N_A_293_74#_c_437_n 5.82005e-19 $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_141_385#_c_230_n N_VPWR_c_309_n 0.00955198f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_173 N_A_141_385#_c_226_n N_VPWR_c_309_n 0.0159936f $X=0.805 $Y=1.95 $X2=0
+ $Y2=0
cc_174 N_A_141_385#_c_230_n N_VPWR_c_312_n 0.0193641f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_175 N_A_141_385#_c_230_n N_VPWR_c_313_n 0.019537f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_176 N_A_141_385#_M1009_g N_VPWR_c_315_n 0.0174069f $X=2.795 $Y=2.4 $X2=0
+ $Y2=0
cc_177 N_A_141_385#_c_230_n N_VPWR_c_316_n 0.00796853f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_178 N_A_141_385#_M1009_g N_VPWR_c_317_n 0.00460063f $X=2.795 $Y=2.4 $X2=0
+ $Y2=0
cc_179 N_A_141_385#_M1009_g N_VPWR_c_308_n 0.00909693f $X=2.795 $Y=2.4 $X2=0
+ $Y2=0
cc_180 N_A_141_385#_c_230_n N_VPWR_c_308_n 0.0105631f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_181 N_A_141_385#_c_224_n N_Y_c_364_n 0.00498172f $X=2.635 $Y=1.095 $X2=0
+ $Y2=0
cc_182 N_A_141_385#_c_227_n N_Y_c_364_n 0.00233195f $X=2.785 $Y=1.095 $X2=0
+ $Y2=0
cc_183 N_A_141_385#_M1009_g N_Y_c_361_n 0.0162523f $X=2.795 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_141_385#_c_227_n N_Y_c_361_n 0.0129931f $X=2.785 $Y=1.095 $X2=0 $Y2=0
cc_185 N_A_141_385#_c_228_n N_Y_c_361_n 0.00237689f $X=2.84 $Y=1.465 $X2=0 $Y2=0
cc_186 N_A_141_385#_M1004_g N_Y_c_358_n 0.0105687f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_141_385#_M1009_g N_Y_c_359_n 0.00675616f $X=2.795 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_141_385#_M1004_g N_Y_c_359_n 0.00330707f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_141_385#_c_227_n N_Y_c_359_n 0.0329445f $X=2.785 $Y=1.095 $X2=0 $Y2=0
cc_190 N_A_141_385#_c_228_n N_Y_c_359_n 0.00803238f $X=2.84 $Y=1.465 $X2=0 $Y2=0
cc_191 N_A_141_385#_c_227_n N_Y_c_360_n 0.00984957f $X=2.785 $Y=1.095 $X2=0
+ $Y2=0
cc_192 N_A_141_385#_c_228_n N_Y_c_360_n 0.0012888f $X=2.84 $Y=1.465 $X2=0 $Y2=0
cc_193 N_A_141_385#_M1009_g N_Y_c_363_n 2.54997e-19 $X=2.795 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_141_385#_c_224_n N_VGND_M1000_d 0.00367023f $X=2.635 $Y=1.095 $X2=0
+ $Y2=0
cc_195 N_A_141_385#_c_223_n N_VGND_c_396_n 0.0145372f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_141_385#_c_225_n N_VGND_c_396_n 0.00994413f $X=1.225 $Y=1.095 $X2=0
+ $Y2=0
cc_197 N_A_141_385#_c_223_n N_VGND_c_398_n 0.00749462f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_198 N_A_141_385#_M1004_g N_VGND_c_399_n 0.00437532f $X=2.82 $Y=0.74 $X2=0
+ $Y2=0
cc_199 N_A_141_385#_M1004_g N_VGND_c_400_n 0.00829339f $X=2.82 $Y=0.74 $X2=0
+ $Y2=0
cc_200 N_A_141_385#_c_223_n N_VGND_c_400_n 0.00907254f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_201 N_A_141_385#_c_225_n A_112_119# 0.00433061f $X=1.225 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_141_385#_c_224_n N_A_293_74#_M1000_s 0.00283795f $X=2.635 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_203 N_A_141_385#_c_224_n N_A_293_74#_M1008_d 0.00119058f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_204 N_A_141_385#_c_227_n N_A_293_74#_M1008_d 5.84861e-19 $X=2.785 $Y=1.095
+ $X2=0 $Y2=0
cc_205 N_A_141_385#_c_224_n N_A_293_74#_c_434_n 0.039534f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_206 N_A_141_385#_c_223_n N_A_293_74#_c_433_n 0.0190291f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_141_385#_c_224_n N_A_293_74#_c_433_n 0.0207364f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_208 N_A_141_385#_M1004_g N_A_293_74#_c_437_n 0.00452712f $X=2.82 $Y=0.74
+ $X2=0 $Y2=0
cc_209 N_A_141_385#_c_224_n N_A_293_74#_c_437_n 0.0103265f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_210 N_A_141_385#_c_227_n N_A_293_74#_c_437_n 0.00637681f $X=2.785 $Y=1.095
+ $X2=0 $Y2=0
cc_211 N_VPWR_M1009_d N_Y_c_361_n 0.00783725f $X=2.885 $Y=1.84 $X2=0 $Y2=0
cc_212 N_VPWR_c_315_n N_Y_c_361_n 0.0225368f $X=3.02 $Y=2.3 $X2=0 $Y2=0
cc_213 N_VPWR_c_313_n N_Y_c_363_n 0.036577f $X=1.58 $Y=2.415 $X2=0 $Y2=0
cc_214 N_VPWR_c_315_n N_Y_c_363_n 0.0267695f $X=3.02 $Y=2.3 $X2=0 $Y2=0
cc_215 N_VPWR_c_317_n N_Y_c_363_n 0.0279296f $X=2.855 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_308_n N_Y_c_363_n 0.022764f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_c_309_n N_VGND_c_396_n 0.00899431f $X=0.34 $Y=2.07 $X2=0 $Y2=0
cc_218 A_379_368# N_Y_c_363_n 0.0076621f $X=1.895 $Y=1.84 $X2=2.3 $Y2=1.515
cc_219 N_Y_c_358_n N_VGND_c_399_n 0.013297f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_220 N_Y_c_358_n N_VGND_c_400_n 0.0110061f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_221 N_Y_c_358_n N_A_293_74#_c_437_n 0.0220168f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_222 N_VGND_M1000_d N_A_293_74#_c_434_n 0.00697375f $X=1.89 $Y=0.37 $X2=0
+ $Y2=0
cc_223 N_VGND_c_397_n N_A_293_74#_c_434_n 0.0239631f $X=2.1 $Y=0.37 $X2=0 $Y2=0
cc_224 N_VGND_c_398_n N_A_293_74#_c_434_n 0.00227739f $X=1.935 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_399_n N_A_293_74#_c_434_n 0.00232204f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_400_n N_A_293_74#_c_434_n 0.00980247f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_398_n N_A_293_74#_c_433_n 0.00745853f $X=1.935 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_400_n N_A_293_74#_c_433_n 0.00921561f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_399_n N_A_293_74#_c_437_n 0.00677194f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_400_n N_A_293_74#_c_437_n 0.0103183f $X=3.12 $Y=0 $X2=0 $Y2=0

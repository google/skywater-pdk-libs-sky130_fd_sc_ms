* File: sky130_fd_sc_ms__sdlclkp_4.pxi.spice
* Created: Wed Sep  2 12:32:16 2020
* 
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%SCE N_SCE_M1025_g N_SCE_M1023_g SCE
+ N_SCE_c_181_n N_SCE_c_182_n PM_SKY130_FD_SC_MS__SDLCLKP_4%SCE
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%GATE N_GATE_M1001_g N_GATE_M1026_g GATE
+ N_GATE_c_208_n PM_SKY130_FD_SC_MS__SDLCLKP_4%GATE
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%A_354_105# N_A_354_105#_M1021_d
+ N_A_354_105#_M1004_d N_A_354_105#_M1005_g N_A_354_105#_c_241_n
+ N_A_354_105#_M1017_g N_A_354_105#_c_243_n N_A_354_105#_c_244_n
+ N_A_354_105#_c_245_n N_A_354_105#_c_253_n N_A_354_105#_c_246_n
+ N_A_354_105#_c_247_n N_A_354_105#_c_248_n N_A_354_105#_c_249_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%A_354_105#
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%A_324_79# N_A_324_79#_M1013_s
+ N_A_324_79#_M1002_s N_A_324_79#_c_319_n N_A_324_79#_M1021_g
+ N_A_324_79#_c_320_n N_A_324_79#_c_321_n N_A_324_79#_M1004_g
+ N_A_324_79#_c_339_n N_A_324_79#_c_340_n N_A_324_79#_c_323_n
+ N_A_324_79#_c_324_n N_A_324_79#_M1024_g N_A_324_79#_M1008_g
+ N_A_324_79#_c_325_n N_A_324_79#_c_326_n N_A_324_79#_c_327_n
+ N_A_324_79#_c_328_n N_A_324_79#_c_329_n N_A_324_79#_c_330_n
+ N_A_324_79#_c_331_n N_A_324_79#_c_379_p N_A_324_79#_c_332_n
+ N_A_324_79#_c_333_n N_A_324_79#_c_334_n N_A_324_79#_c_367_n
+ N_A_324_79#_c_342_n N_A_324_79#_c_335_n N_A_324_79#_c_336_n
+ N_A_324_79#_c_337_n PM_SKY130_FD_SC_MS__SDLCLKP_4%A_324_79#
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%A_792_48# N_A_792_48#_M1006_d
+ N_A_792_48#_M1022_d N_A_792_48#_M1007_g N_A_792_48#_M1014_g
+ N_A_792_48#_M1012_g N_A_792_48#_M1019_g N_A_792_48#_c_484_n
+ N_A_792_48#_c_485_n N_A_792_48#_c_486_n N_A_792_48#_c_476_n
+ N_A_792_48#_c_488_n N_A_792_48#_c_507_n N_A_792_48#_c_509_n
+ N_A_792_48#_c_477_n N_A_792_48#_c_478_n N_A_792_48#_c_490_n
+ N_A_792_48#_c_491_n N_A_792_48#_c_479_n N_A_792_48#_c_480_n
+ N_A_792_48#_c_481_n PM_SKY130_FD_SC_MS__SDLCLKP_4%A_792_48#
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%A_634_74# N_A_634_74#_M1024_d
+ N_A_634_74#_M1005_d N_A_634_74#_M1022_g N_A_634_74#_M1006_g
+ N_A_634_74#_c_603_n N_A_634_74#_c_604_n N_A_634_74#_c_605_n
+ N_A_634_74#_c_606_n N_A_634_74#_c_607_n N_A_634_74#_c_608_n
+ N_A_634_74#_c_609_n N_A_634_74#_c_610_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%A_634_74#
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%CLK N_CLK_M1002_g N_CLK_c_681_n N_CLK_M1013_g
+ N_CLK_M1020_g N_CLK_c_683_n N_CLK_M1011_g CLK N_CLK_c_685_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%CLK
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%A_1292_368# N_A_1292_368#_M1012_d
+ N_A_1292_368#_M1020_d N_A_1292_368#_M1009_g N_A_1292_368#_M1000_g
+ N_A_1292_368#_M1010_g N_A_1292_368#_M1003_g N_A_1292_368#_M1016_g
+ N_A_1292_368#_M1015_g N_A_1292_368#_M1018_g N_A_1292_368#_M1027_g
+ N_A_1292_368#_c_754_n N_A_1292_368#_c_743_n N_A_1292_368#_c_755_n
+ N_A_1292_368#_c_756_n N_A_1292_368#_c_744_n N_A_1292_368#_c_745_n
+ N_A_1292_368#_c_746_n N_A_1292_368#_c_747_n N_A_1292_368#_c_809_p
+ N_A_1292_368#_c_748_n N_A_1292_368#_c_749_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%A_1292_368#
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%VPWR N_VPWR_M1025_s N_VPWR_M1004_s
+ N_VPWR_M1014_d N_VPWR_M1002_d N_VPWR_M1019_d N_VPWR_M1010_s N_VPWR_M1018_s
+ N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n N_VPWR_c_866_n N_VPWR_c_867_n
+ N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_871_n N_VPWR_c_872_n
+ VPWR N_VPWR_c_873_n N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n
+ N_VPWR_c_877_n N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n
+ N_VPWR_c_862_n PM_SKY130_FD_SC_MS__SDLCLKP_4%VPWR
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%A_119_143# N_A_119_143#_M1023_d
+ N_A_119_143#_M1024_s N_A_119_143#_M1001_d N_A_119_143#_M1005_s
+ N_A_119_143#_c_967_n N_A_119_143#_c_968_n N_A_119_143#_c_969_n
+ N_A_119_143#_c_970_n N_A_119_143#_c_974_n N_A_119_143#_c_975_n
+ N_A_119_143#_c_976_n N_A_119_143#_c_977_n N_A_119_143#_c_1021_n
+ N_A_119_143#_c_971_n N_A_119_143#_c_972_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%A_119_143#
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%GCLK N_GCLK_M1000_s N_GCLK_M1015_s
+ N_GCLK_M1009_d N_GCLK_M1016_d N_GCLK_c_1067_n N_GCLK_c_1062_n N_GCLK_c_1068_n
+ N_GCLK_c_1069_n N_GCLK_c_1063_n N_GCLK_c_1064_n N_GCLK_c_1070_n
+ N_GCLK_c_1065_n N_GCLK_c_1066_n N_GCLK_c_1072_n GCLK N_GCLK_c_1106_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%GCLK
x_PM_SKY130_FD_SC_MS__SDLCLKP_4%VGND N_VGND_M1023_s N_VGND_M1026_d
+ N_VGND_M1007_d N_VGND_M1013_d N_VGND_M1000_d N_VGND_M1003_d N_VGND_M1027_d
+ N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n
+ N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n
+ N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n N_VGND_c_1143_n
+ N_VGND_c_1144_n VGND N_VGND_c_1145_n N_VGND_c_1146_n N_VGND_c_1147_n
+ N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_4%VGND
cc_1 VNB N_SCE_M1023_g 0.0277275f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.99
cc_2 VNB N_SCE_c_181_n 0.0231115f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_3 VNB N_SCE_c_182_n 0.00872743f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_4 VNB N_GATE_M1026_g 0.0240981f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.99
cc_5 VNB GATE 0.0059014f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_GATE_c_208_n 0.0205209f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_7 VNB N_A_354_105#_c_241_n 0.0221071f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.62
cc_8 VNB N_A_354_105#_M1017_g 0.0437828f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.785
cc_9 VNB N_A_354_105#_c_243_n 0.00699887f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_10 VNB N_A_354_105#_c_244_n 8.06639e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_354_105#_c_245_n 6.67232e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_354_105#_c_246_n 0.00206511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_354_105#_c_247_n 0.00282247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_354_105#_c_248_n 0.00353693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_354_105#_c_249_n 0.0329462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_324_79#_c_319_n 0.0191913f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.99
cc_17 VNB N_A_324_79#_c_320_n 0.0223453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_324_79#_c_321_n 0.0128593f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.62
cc_19 VNB N_A_324_79#_M1004_g 0.00886371f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.785
cc_20 VNB N_A_324_79#_c_323_n 0.0422786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_324_79#_c_324_n 0.0210931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_324_79#_c_325_n 0.00491788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_324_79#_c_326_n 0.00525298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_324_79#_c_327_n 0.00566241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_324_79#_c_328_n 0.00487706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_324_79#_c_329_n 0.00149564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_324_79#_c_330_n 0.0141001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_324_79#_c_331_n 0.00262393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_324_79#_c_332_n 0.0149264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_324_79#_c_333_n 0.00222644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_324_79#_c_334_n 0.00452749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_324_79#_c_335_n 0.012119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_324_79#_c_336_n 0.0019697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_324_79#_c_337_n 0.0569887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_792_48#_M1007_g 0.0571831f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_A_792_48#_M1012_g 0.0248678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_792_48#_M1019_g 0.00188561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_792_48#_c_476_n 0.00941361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_792_48#_c_477_n 0.0157893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_792_48#_c_478_n 0.00166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_792_48#_c_479_n 0.00395206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_792_48#_c_480_n 0.0115363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_792_48#_c_481_n 0.0371752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_634_74#_M1022_g 6.47399e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_45 VNB N_A_634_74#_c_603_n 0.00321093f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.785
cc_46 VNB N_A_634_74#_c_604_n 0.00131206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_634_74#_c_605_n 0.0213092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_634_74#_c_606_n 0.0035258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_634_74#_c_607_n 0.00692367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_634_74#_c_608_n 0.00462435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_634_74#_c_609_n 0.0399923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_634_74#_c_610_n 0.0228989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_CLK_M1002_g 0.00671413f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.395
cc_54 VNB N_CLK_c_681_n 0.0200962f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.455
cc_55 VNB N_CLK_M1020_g 0.00597977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_CLK_c_683_n 0.0171643f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_57 VNB CLK 0.0075037f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.785
cc_58 VNB N_CLK_c_685_n 0.0496165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1292_368#_M1009_g 0.00162616f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_60 VNB N_A_1292_368#_M1000_g 0.0233521f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.62
cc_61 VNB N_A_1292_368#_M1010_g 0.00174205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1292_368#_M1003_g 0.0209649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1292_368#_M1016_g 0.00164311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1292_368#_M1015_g 0.0202297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1292_368#_M1018_g 0.00248079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1292_368#_M1027_g 0.0260342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1292_368#_c_743_n 0.00912363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1292_368#_c_744_n 0.0130086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1292_368#_c_745_n 0.00269775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1292_368#_c_746_n 0.00378119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1292_368#_c_747_n 2.98518e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1292_368#_c_748_n 0.00266677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1292_368#_c_749_n 0.11703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VPWR_c_862_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_119_143#_c_967_n 0.00958489f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.785
cc_76 VNB N_A_119_143#_c_968_n 8.44192e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_119_143#_c_969_n 0.00496514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_119_143#_c_970_n 0.00458561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_119_143#_c_971_n 0.0096811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_119_143#_c_972_n 0.00838916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_GCLK_c_1062_n 0.00254365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_GCLK_c_1063_n 0.00351355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_GCLK_c_1064_n 0.00205014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_GCLK_c_1065_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_GCLK_c_1066_n 5.71281e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1132_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1133_n 0.067074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1134_n 0.0192463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1135_n 0.00644324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1136_n 0.00600048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1137_n 0.0126279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1138_n 0.00503707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1139_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1140_n 0.0505914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1141_n 0.0643337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1142_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1143_n 0.0380624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1144_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1145_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1146_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1147_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1148_n 0.028177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1149_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1150_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1151_n 0.535277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VPB N_SCE_M1025_g 0.0291858f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.395
cc_107 VPB N_SCE_c_181_n 0.0154497f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.62
cc_108 VPB N_SCE_c_182_n 0.00565041f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.62
cc_109 VPB N_GATE_M1001_g 0.0259131f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.395
cc_110 VPB GATE 0.00348266f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_111 VPB N_GATE_c_208_n 0.0130964f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.62
cc_112 VPB N_A_354_105#_M1005_g 0.0261831f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_113 VPB N_A_354_105#_c_244_n 0.00167859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_354_105#_c_245_n 0.00497365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_354_105#_c_253_n 0.00934855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_354_105#_c_246_n 0.00371457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_354_105#_c_247_n 6.44492e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_354_105#_c_248_n 0.00276779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_354_105#_c_249_n 0.0171087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_324_79#_M1004_g 0.0390951f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.785
cc_121 VPB N_A_324_79#_c_339_n 0.11926f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.62
cc_122 VPB N_A_324_79#_c_340_n 0.0130767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_324_79#_M1008_g 0.0479025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_324_79#_c_342_n 0.00695691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_324_79#_c_335_n 0.00294593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_792_48#_M1014_g 0.0375464f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.62
cc_127 VPB N_A_792_48#_M1019_g 0.0255355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_792_48#_c_484_n 0.00622092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_792_48#_c_485_n 0.00449717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_792_48#_c_486_n 0.0138111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_792_48#_c_476_n 0.00315538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_792_48#_c_488_n 0.0136815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_792_48#_c_478_n 0.00816786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_792_48#_c_490_n 0.00430204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_792_48#_c_491_n 5.03018e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_792_48#_c_480_n 0.0338369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_634_74#_M1022_g 0.0279138f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_138 VPB N_A_634_74#_c_604_n 0.0134653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_CLK_M1002_g 0.0259205f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.395
cc_140 VPB N_CLK_M1020_g 0.0270494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1292_368#_M1009_g 0.0231906f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_142 VPB N_A_1292_368#_M1010_g 0.0241486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1292_368#_M1016_g 0.0231739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_1292_368#_M1018_g 0.0295324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1292_368#_c_754_n 0.00280241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_1292_368#_c_755_n 0.00393707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1292_368#_c_756_n 0.00245802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1292_368#_c_747_n 0.00143083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_863_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_864_n 0.0571167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_865_n 0.0185736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_866_n 0.0169956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_867_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_868_n 0.0081889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_869_n 0.0120013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_870_n 0.0651854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_871_n 0.023151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_872_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_873_n 0.0330329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_874_n 0.0681025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_875_n 0.0387399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_876_n 0.0220372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_877_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_878_n 0.0264107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_879_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_880_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_881_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_862_n 0.138477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_119_143#_c_970_n 0.00859518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_119_143#_c_974_n 0.0141086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_119_143#_c_975_n 0.00497553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_119_143#_c_976_n 0.0118392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_119_143#_c_977_n 0.022588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_GCLK_c_1067_n 0.002787f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.785
cc_175 VPB N_GCLK_c_1068_n 0.00291589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_GCLK_c_1069_n 0.00249343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_GCLK_c_1070_n 0.00275653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_GCLK_c_1066_n 0.00264693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_GCLK_c_1072_n 0.00105536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 N_SCE_M1025_g N_GATE_M1001_g 0.0391586f $X=0.505 $Y=2.395 $X2=0 $Y2=0
cc_181 N_SCE_M1023_g N_GATE_M1026_g 0.0177982f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_182 N_SCE_c_181_n GATE 0.00127121f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_183 N_SCE_c_182_n GATE 0.0171967f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_184 N_SCE_c_181_n N_GATE_c_208_n 0.0391586f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_185 N_SCE_c_182_n N_GATE_c_208_n 3.90315e-19 $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_186 N_SCE_M1025_g N_VPWR_c_864_n 0.0255967f $X=0.505 $Y=2.395 $X2=0 $Y2=0
cc_187 N_SCE_c_181_n N_VPWR_c_864_n 0.00454265f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_188 N_SCE_c_182_n N_VPWR_c_864_n 0.0271638f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_189 N_SCE_M1025_g N_VPWR_c_873_n 0.00477175f $X=0.505 $Y=2.395 $X2=0 $Y2=0
cc_190 N_SCE_M1025_g N_VPWR_c_862_n 0.00504253f $X=0.505 $Y=2.395 $X2=0 $Y2=0
cc_191 N_SCE_M1023_g N_A_119_143#_c_967_n 6.33101e-19 $X=0.52 $Y=0.99 $X2=0
+ $Y2=0
cc_192 N_SCE_M1023_g N_A_119_143#_c_969_n 0.00128972f $X=0.52 $Y=0.99 $X2=0
+ $Y2=0
cc_193 N_SCE_M1025_g N_A_119_143#_c_976_n 0.00100651f $X=0.505 $Y=2.395 $X2=0
+ $Y2=0
cc_194 N_SCE_M1025_g N_A_119_143#_c_977_n 0.00147726f $X=0.505 $Y=2.395 $X2=0
+ $Y2=0
cc_195 N_SCE_M1023_g N_VGND_c_1133_n 0.00746819f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_196 N_SCE_c_181_n N_VGND_c_1133_n 0.00533261f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_197 N_SCE_c_182_n N_VGND_c_1133_n 0.0272945f $X=0.385 $Y=1.62 $X2=0 $Y2=0
cc_198 N_SCE_M1023_g N_VGND_c_1134_n 0.00370133f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_199 N_SCE_M1023_g N_VGND_c_1151_n 0.00445256f $X=0.52 $Y=0.99 $X2=0 $Y2=0
cc_200 N_GATE_M1026_g N_A_324_79#_c_319_n 0.0141001f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_201 N_GATE_c_208_n N_A_324_79#_c_321_n 8.07007e-19 $X=1 $Y=1.62 $X2=0 $Y2=0
cc_202 N_GATE_M1001_g N_VPWR_c_864_n 0.0030268f $X=0.925 $Y=2.395 $X2=0 $Y2=0
cc_203 N_GATE_M1001_g N_VPWR_c_873_n 0.0055029f $X=0.925 $Y=2.395 $X2=0 $Y2=0
cc_204 N_GATE_M1001_g N_VPWR_c_878_n 0.00350614f $X=0.925 $Y=2.395 $X2=0 $Y2=0
cc_205 N_GATE_M1001_g N_VPWR_c_862_n 0.00601096f $X=0.925 $Y=2.395 $X2=0 $Y2=0
cc_206 N_GATE_M1026_g N_A_119_143#_c_967_n 0.0109495f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_207 GATE N_A_119_143#_c_967_n 0.00907303f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_208 N_GATE_c_208_n N_A_119_143#_c_967_n 0.00231117f $X=1 $Y=1.62 $X2=0 $Y2=0
cc_209 N_GATE_M1026_g N_A_119_143#_c_968_n 0.0103937f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_210 GATE N_A_119_143#_c_968_n 0.00878437f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_211 N_GATE_c_208_n N_A_119_143#_c_968_n 0.00126549f $X=1 $Y=1.62 $X2=0 $Y2=0
cc_212 N_GATE_M1026_g N_A_119_143#_c_969_n 0.00269077f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_213 N_GATE_M1001_g N_A_119_143#_c_970_n 0.00432161f $X=0.925 $Y=2.395 $X2=0
+ $Y2=0
cc_214 N_GATE_M1026_g N_A_119_143#_c_970_n 0.00678895f $X=0.995 $Y=0.99 $X2=0
+ $Y2=0
cc_215 GATE N_A_119_143#_c_970_n 0.0269205f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_216 N_GATE_c_208_n N_A_119_143#_c_970_n 0.00151897f $X=1 $Y=1.62 $X2=0 $Y2=0
cc_217 N_GATE_M1001_g N_A_119_143#_c_976_n 0.00743333f $X=0.925 $Y=2.395 $X2=0
+ $Y2=0
cc_218 N_GATE_M1001_g N_A_119_143#_c_977_n 0.0146287f $X=0.925 $Y=2.395 $X2=0
+ $Y2=0
cc_219 GATE N_A_119_143#_c_977_n 0.0276031f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_220 N_GATE_c_208_n N_A_119_143#_c_977_n 0.00367709f $X=1 $Y=1.62 $X2=0 $Y2=0
cc_221 N_GATE_M1026_g N_VGND_c_1134_n 0.00287494f $X=0.995 $Y=0.99 $X2=0 $Y2=0
cc_222 N_GATE_M1026_g N_VGND_c_1151_n 0.00445256f $X=0.995 $Y=0.99 $X2=0 $Y2=0
cc_223 N_A_354_105#_c_243_n N_A_324_79#_c_319_n 6.11846e-19 $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_224 N_A_354_105#_c_243_n N_A_324_79#_c_320_n 0.0190885f $X=1.91 $Y=1.12 $X2=0
+ $Y2=0
cc_225 N_A_354_105#_c_244_n N_A_324_79#_c_320_n 0.00248561f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_226 N_A_354_105#_c_243_n N_A_324_79#_M1004_g 0.00361705f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_227 N_A_354_105#_c_244_n N_A_324_79#_M1004_g 0.0198003f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_228 N_A_354_105#_c_253_n N_A_324_79#_M1004_g 0.0168571f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_229 N_A_354_105#_c_249_n N_A_324_79#_M1004_g 0.00202336f $X=3.405 $Y=1.57
+ $X2=0 $Y2=0
cc_230 N_A_354_105#_M1005_g N_A_324_79#_c_339_n 0.0123546f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_231 N_A_354_105#_c_246_n N_A_324_79#_c_323_n 0.00132308f $X=2.925 $Y=1.65
+ $X2=0 $Y2=0
cc_232 N_A_354_105#_c_247_n N_A_324_79#_c_323_n 7.91151e-19 $X=2.53 $Y=1.65
+ $X2=0 $Y2=0
cc_233 N_A_354_105#_c_248_n N_A_324_79#_c_323_n 0.00143623f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_234 N_A_354_105#_c_249_n N_A_324_79#_c_323_n 0.015893f $X=3.405 $Y=1.57 $X2=0
+ $Y2=0
cc_235 N_A_354_105#_M1017_g N_A_324_79#_c_324_n 0.0217463f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_236 N_A_354_105#_M1005_g N_A_324_79#_M1008_g 0.0142498f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_237 N_A_354_105#_M1017_g N_A_324_79#_c_325_n 3.16786e-19 $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_238 N_A_354_105#_c_246_n N_A_324_79#_c_325_n 0.0115741f $X=2.925 $Y=1.65
+ $X2=0 $Y2=0
cc_239 N_A_354_105#_c_247_n N_A_324_79#_c_325_n 0.0063017f $X=2.53 $Y=1.65 $X2=0
+ $Y2=0
cc_240 N_A_354_105#_c_248_n N_A_324_79#_c_325_n 0.00415249f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_241 N_A_354_105#_M1017_g N_A_324_79#_c_327_n 0.0129965f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_242 N_A_354_105#_M1017_g N_A_324_79#_c_329_n 0.00199569f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_243 N_A_354_105#_M1017_g N_A_324_79#_c_331_n 0.00133148f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_244 N_A_354_105#_c_243_n N_A_324_79#_c_367_n 0.0253307f $X=1.91 $Y=1.12 $X2=0
+ $Y2=0
cc_245 N_A_354_105#_c_244_n N_A_324_79#_c_367_n 0.00871007f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_246 N_A_354_105#_c_247_n N_A_324_79#_c_367_n 0.0174669f $X=2.53 $Y=1.65 $X2=0
+ $Y2=0
cc_247 N_A_354_105#_c_243_n N_A_324_79#_c_337_n 0.00335921f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_248 N_A_354_105#_c_244_n N_A_324_79#_c_337_n 0.00146387f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_249 N_A_354_105#_c_247_n N_A_324_79#_c_337_n 0.00579073f $X=2.53 $Y=1.65
+ $X2=0 $Y2=0
cc_250 N_A_354_105#_c_248_n N_A_324_79#_c_337_n 6.1217e-19 $X=3.09 $Y=1.57 $X2=0
+ $Y2=0
cc_251 N_A_354_105#_c_249_n N_A_324_79#_c_337_n 0.00379557f $X=3.405 $Y=1.57
+ $X2=0 $Y2=0
cc_252 N_A_354_105#_M1017_g N_A_792_48#_M1007_g 0.0653275f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_253 N_A_354_105#_c_249_n N_A_792_48#_M1007_g 0.00247769f $X=3.405 $Y=1.57
+ $X2=0 $Y2=0
cc_254 N_A_354_105#_M1005_g N_A_792_48#_c_480_n 0.00247769f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_255 N_A_354_105#_M1017_g N_A_634_74#_c_603_n 0.00730232f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_256 N_A_354_105#_c_241_n N_A_634_74#_c_604_n 0.0147699f $X=3.57 $Y=1.48 $X2=0
+ $Y2=0
cc_257 N_A_354_105#_c_248_n N_A_634_74#_c_604_n 0.0251391f $X=3.09 $Y=1.57 $X2=0
+ $Y2=0
cc_258 N_A_354_105#_c_249_n N_A_634_74#_c_604_n 0.00837301f $X=3.405 $Y=1.57
+ $X2=0 $Y2=0
cc_259 N_A_354_105#_M1017_g N_A_634_74#_c_605_n 0.00308854f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_260 N_A_354_105#_c_241_n N_A_634_74#_c_606_n 3.55064e-19 $X=3.57 $Y=1.48
+ $X2=0 $Y2=0
cc_261 N_A_354_105#_M1017_g N_A_634_74#_c_606_n 0.00876954f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_262 N_A_354_105#_c_248_n N_A_634_74#_c_606_n 0.00397264f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_263 N_A_354_105#_c_249_n N_A_634_74#_c_606_n 0.00597586f $X=3.405 $Y=1.57
+ $X2=0 $Y2=0
cc_264 N_A_354_105#_c_241_n N_A_634_74#_c_607_n 0.00317399f $X=3.57 $Y=1.48
+ $X2=0 $Y2=0
cc_265 N_A_354_105#_M1017_g N_A_634_74#_c_607_n 0.0107752f $X=3.645 $Y=0.58
+ $X2=0 $Y2=0
cc_266 N_A_354_105#_M1005_g N_VPWR_c_862_n 0.00112709f $X=3.315 $Y=2.315 $X2=0
+ $Y2=0
cc_267 N_A_354_105#_c_243_n N_A_119_143#_c_970_n 0.0322212f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_268 N_A_354_105#_c_245_n N_A_119_143#_c_970_n 0.0143581f $X=2.075 $Y=1.65
+ $X2=0 $Y2=0
cc_269 N_A_354_105#_M1004_d N_A_119_143#_c_974_n 0.00810352f $X=2.31 $Y=2.12
+ $X2=0 $Y2=0
cc_270 N_A_354_105#_M1005_g N_A_119_143#_c_974_n 0.00789033f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_271 N_A_354_105#_c_244_n N_A_119_143#_c_974_n 0.00621497f $X=2.365 $Y=1.65
+ $X2=0 $Y2=0
cc_272 N_A_354_105#_c_245_n N_A_119_143#_c_974_n 0.00862623f $X=2.075 $Y=1.65
+ $X2=0 $Y2=0
cc_273 N_A_354_105#_c_253_n N_A_119_143#_c_974_n 0.0263015f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_274 N_A_354_105#_c_246_n N_A_119_143#_c_974_n 0.00740026f $X=2.925 $Y=1.65
+ $X2=0 $Y2=0
cc_275 N_A_354_105#_M1005_g N_A_119_143#_c_975_n 0.00596902f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_276 N_A_354_105#_c_253_n N_A_119_143#_c_975_n 0.0158435f $X=2.53 $Y=1.975
+ $X2=0 $Y2=0
cc_277 N_A_354_105#_c_248_n N_A_119_143#_c_975_n 0.0245639f $X=3.09 $Y=1.57
+ $X2=0 $Y2=0
cc_278 N_A_354_105#_c_249_n N_A_119_143#_c_975_n 0.00219377f $X=3.405 $Y=1.57
+ $X2=0 $Y2=0
cc_279 N_A_354_105#_M1021_d N_A_119_143#_c_972_n 0.00709289f $X=1.77 $Y=0.525
+ $X2=0 $Y2=0
cc_280 N_A_354_105#_c_243_n N_A_119_143#_c_972_n 0.0201545f $X=1.91 $Y=1.12
+ $X2=0 $Y2=0
cc_281 N_A_354_105#_M1017_g N_VGND_c_1135_n 3.67768e-19 $X=3.645 $Y=0.58 $X2=0
+ $Y2=0
cc_282 N_A_354_105#_M1017_g N_VGND_c_1141_n 0.00280452f $X=3.645 $Y=0.58 $X2=0
+ $Y2=0
cc_283 N_A_354_105#_M1017_g N_VGND_c_1151_n 0.00354535f $X=3.645 $Y=0.58 $X2=0
+ $Y2=0
cc_284 N_A_324_79#_c_332_n N_A_792_48#_M1006_d 0.00273752f $X=5.445 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_285 N_A_324_79#_c_327_n N_A_792_48#_M1007_g 0.00107336f $X=3.765 $Y=0.355
+ $X2=0 $Y2=0
cc_286 N_A_324_79#_c_329_n N_A_792_48#_M1007_g 0.00274065f $X=3.85 $Y=0.895
+ $X2=0 $Y2=0
cc_287 N_A_324_79#_c_330_n N_A_792_48#_M1007_g 0.0153072f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_288 N_A_324_79#_c_379_p N_A_792_48#_M1007_g 0.00137341f $X=4.69 $Y=0.895
+ $X2=0 $Y2=0
cc_289 N_A_324_79#_c_333_n N_A_792_48#_M1007_g 3.77334e-19 $X=4.775 $Y=0.34
+ $X2=0 $Y2=0
cc_290 N_A_324_79#_M1008_g N_A_792_48#_M1014_g 0.035737f $X=3.85 $Y=2.485 $X2=0
+ $Y2=0
cc_291 N_A_324_79#_c_342_n N_A_792_48#_c_485_n 0.013888f $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_292 N_A_324_79#_c_335_n N_A_792_48#_c_476_n 0.0502011f $X=5.607 $Y=1.82 $X2=0
+ $Y2=0
cc_293 N_A_324_79#_M1002_s N_A_792_48#_c_488_n 0.0120995f $X=5.46 $Y=1.84 $X2=0
+ $Y2=0
cc_294 N_A_324_79#_c_342_n N_A_792_48#_c_488_n 0.021703f $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A_324_79#_c_342_n N_A_792_48#_c_507_n 0.00728723f $X=5.605 $Y=1.985
+ $X2=0 $Y2=0
cc_296 N_A_324_79#_c_335_n N_A_792_48#_c_507_n 0.00347829f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_297 N_A_324_79#_c_335_n N_A_792_48#_c_509_n 0.00218713f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_298 N_A_324_79#_c_342_n N_A_792_48#_c_490_n 0.0075272f $X=5.605 $Y=1.985
+ $X2=0 $Y2=0
cc_299 N_A_324_79#_c_335_n N_A_792_48#_c_490_n 0.00742029f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_300 N_A_324_79#_c_332_n N_A_792_48#_c_479_n 0.0203619f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_301 N_A_324_79#_c_334_n N_A_792_48#_c_479_n 0.0397103f $X=5.67 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_324_79#_c_327_n N_A_634_74#_M1024_d 0.00320041f $X=3.765 $Y=0.355
+ $X2=-0.19 $Y2=-0.245
cc_303 N_A_324_79#_c_335_n N_A_634_74#_M1022_g 9.59979e-19 $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_304 N_A_324_79#_c_324_n N_A_634_74#_c_603_n 0.00236682f $X=3.095 $Y=1.045
+ $X2=0 $Y2=0
cc_305 N_A_324_79#_c_325_n N_A_634_74#_c_603_n 0.00641233f $X=2.805 $Y=1.15
+ $X2=0 $Y2=0
cc_306 N_A_324_79#_c_326_n N_A_634_74#_c_603_n 0.00468717f $X=2.89 $Y=1.065
+ $X2=0 $Y2=0
cc_307 N_A_324_79#_c_331_n N_A_634_74#_c_603_n 0.0100839f $X=3.935 $Y=0.98 $X2=0
+ $Y2=0
cc_308 N_A_324_79#_c_339_n N_A_634_74#_c_604_n 0.00495646f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_309 N_A_324_79#_M1008_g N_A_634_74#_c_604_n 0.00743278f $X=3.85 $Y=2.485
+ $X2=0 $Y2=0
cc_310 N_A_324_79#_c_330_n N_A_634_74#_c_605_n 0.0488693f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_311 N_A_324_79#_c_331_n N_A_634_74#_c_605_n 0.0143583f $X=3.935 $Y=0.98 $X2=0
+ $Y2=0
cc_312 N_A_324_79#_c_324_n N_A_634_74#_c_606_n 0.00454113f $X=3.095 $Y=1.045
+ $X2=0 $Y2=0
cc_313 N_A_324_79#_c_326_n N_A_634_74#_c_606_n 0.0136555f $X=2.89 $Y=1.065 $X2=0
+ $Y2=0
cc_314 N_A_324_79#_c_327_n N_A_634_74#_c_606_n 0.0238927f $X=3.765 $Y=0.355
+ $X2=0 $Y2=0
cc_315 N_A_324_79#_c_329_n N_A_634_74#_c_606_n 0.0151262f $X=3.85 $Y=0.895 $X2=0
+ $Y2=0
cc_316 N_A_324_79#_c_331_n N_A_634_74#_c_606_n 0.00380883f $X=3.935 $Y=0.98
+ $X2=0 $Y2=0
cc_317 N_A_324_79#_c_330_n N_A_634_74#_c_608_n 0.0135682f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_318 N_A_324_79#_c_330_n N_A_634_74#_c_609_n 0.00130489f $X=4.605 $Y=0.98
+ $X2=0 $Y2=0
cc_319 N_A_324_79#_c_332_n N_A_634_74#_c_610_n 0.0156771f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_320 N_A_324_79#_c_334_n N_A_634_74#_c_610_n 0.00385526f $X=5.67 $Y=0.515
+ $X2=0 $Y2=0
cc_321 N_A_324_79#_c_335_n N_A_634_74#_c_610_n 0.00125296f $X=5.607 $Y=1.82
+ $X2=0 $Y2=0
cc_322 N_A_324_79#_c_342_n N_CLK_M1002_g 0.00670381f $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_324_79#_c_332_n N_CLK_c_681_n 0.00462516f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_324 N_A_324_79#_c_334_n N_CLK_c_681_n 0.0043874f $X=5.67 $Y=0.515 $X2=0 $Y2=0
cc_325 N_A_324_79#_c_335_n N_CLK_c_681_n 0.00343873f $X=5.607 $Y=1.82 $X2=0
+ $Y2=0
cc_326 N_A_324_79#_c_336_n N_CLK_c_681_n 0.00232496f $X=5.64 $Y=1.01 $X2=0 $Y2=0
cc_327 N_A_324_79#_c_342_n N_CLK_M1020_g 7.35762e-19 $X=5.605 $Y=1.985 $X2=0
+ $Y2=0
cc_328 N_A_324_79#_c_335_n CLK 0.0279712f $X=5.607 $Y=1.82 $X2=0 $Y2=0
cc_329 N_A_324_79#_c_336_n CLK 0.0029255f $X=5.64 $Y=1.01 $X2=0 $Y2=0
cc_330 N_A_324_79#_c_335_n N_CLK_c_685_n 0.0148131f $X=5.607 $Y=1.82 $X2=0 $Y2=0
cc_331 N_A_324_79#_c_336_n N_CLK_c_685_n 0.00113546f $X=5.64 $Y=1.01 $X2=0 $Y2=0
cc_332 N_A_324_79#_M1008_g N_VPWR_c_865_n 0.0104158f $X=3.85 $Y=2.485 $X2=0
+ $Y2=0
cc_333 N_A_324_79#_c_340_n N_VPWR_c_874_n 0.0578172f $X=2.31 $Y=3.15 $X2=0 $Y2=0
cc_334 N_A_324_79#_M1004_g N_VPWR_c_878_n 0.0236672f $X=2.22 $Y=2.54 $X2=0 $Y2=0
cc_335 N_A_324_79#_c_340_n N_VPWR_c_878_n 0.00826345f $X=2.31 $Y=3.15 $X2=0
+ $Y2=0
cc_336 N_A_324_79#_c_339_n N_VPWR_c_862_n 0.0571785f $X=3.76 $Y=3.15 $X2=0 $Y2=0
cc_337 N_A_324_79#_c_340_n N_VPWR_c_862_n 0.00459104f $X=2.31 $Y=3.15 $X2=0
+ $Y2=0
cc_338 N_A_324_79#_c_326_n N_A_119_143#_M1024_s 0.00828024f $X=2.89 $Y=1.065
+ $X2=0 $Y2=0
cc_339 N_A_324_79#_c_328_n N_A_119_143#_M1024_s 9.10245e-19 $X=2.975 $Y=0.355
+ $X2=0 $Y2=0
cc_340 N_A_324_79#_c_319_n N_A_119_143#_c_967_n 4.34451e-19 $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_341 N_A_324_79#_c_319_n N_A_119_143#_c_970_n 0.0157986f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_342 N_A_324_79#_c_321_n N_A_119_143#_c_970_n 0.005009f $X=1.77 $Y=1.415 $X2=0
+ $Y2=0
cc_343 N_A_324_79#_M1004_g N_A_119_143#_c_970_n 0.00632018f $X=2.22 $Y=2.54
+ $X2=0 $Y2=0
cc_344 N_A_324_79#_M1004_g N_A_119_143#_c_974_n 0.0264121f $X=2.22 $Y=2.54 $X2=0
+ $Y2=0
cc_345 N_A_324_79#_c_339_n N_A_119_143#_c_974_n 0.0177273f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_346 N_A_324_79#_M1004_g N_A_119_143#_c_975_n 0.0043978f $X=2.22 $Y=2.54 $X2=0
+ $Y2=0
cc_347 N_A_324_79#_M1004_g N_A_119_143#_c_977_n 0.0106436f $X=2.22 $Y=2.54 $X2=0
+ $Y2=0
cc_348 N_A_324_79#_c_319_n N_A_119_143#_c_1021_n 0.00435069f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_349 N_A_324_79#_c_319_n N_A_119_143#_c_971_n 0.00731619f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_350 N_A_324_79#_c_324_n N_A_119_143#_c_971_n 0.00124433f $X=3.095 $Y=1.045
+ $X2=0 $Y2=0
cc_351 N_A_324_79#_c_325_n N_A_119_143#_c_971_n 0.00459251f $X=2.805 $Y=1.15
+ $X2=0 $Y2=0
cc_352 N_A_324_79#_c_326_n N_A_119_143#_c_971_n 0.0356041f $X=2.89 $Y=1.065
+ $X2=0 $Y2=0
cc_353 N_A_324_79#_c_328_n N_A_119_143#_c_971_n 0.00767896f $X=2.975 $Y=0.355
+ $X2=0 $Y2=0
cc_354 N_A_324_79#_c_367_n N_A_119_143#_c_971_n 0.0218607f $X=2.41 $Y=1.15 $X2=0
+ $Y2=0
cc_355 N_A_324_79#_c_337_n N_A_119_143#_c_971_n 0.00799329f $X=2.352 $Y=1.12
+ $X2=0 $Y2=0
cc_356 N_A_324_79#_c_319_n N_A_119_143#_c_972_n 0.0129997f $X=1.695 $Y=1.34
+ $X2=0 $Y2=0
cc_357 N_A_324_79#_c_320_n N_A_119_143#_c_972_n 5.7542e-19 $X=2.13 $Y=1.415
+ $X2=0 $Y2=0
cc_358 N_A_324_79#_c_367_n N_A_119_143#_c_972_n 0.00303811f $X=2.41 $Y=1.15
+ $X2=0 $Y2=0
cc_359 N_A_324_79#_c_337_n N_A_119_143#_c_972_n 0.00583436f $X=2.352 $Y=1.12
+ $X2=0 $Y2=0
cc_360 N_A_324_79#_c_330_n N_VGND_M1007_d 0.00468885f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_361 N_A_324_79#_c_379_p N_VGND_M1007_d 0.00845472f $X=4.69 $Y=0.895 $X2=0
+ $Y2=0
cc_362 N_A_324_79#_c_333_n N_VGND_M1007_d 6.47853e-19 $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_363 N_A_324_79#_c_327_n N_VGND_c_1135_n 0.0110244f $X=3.765 $Y=0.355 $X2=0
+ $Y2=0
cc_364 N_A_324_79#_c_330_n N_VGND_c_1135_n 0.0244958f $X=4.605 $Y=0.98 $X2=0
+ $Y2=0
cc_365 N_A_324_79#_c_379_p N_VGND_c_1135_n 0.0228902f $X=4.69 $Y=0.895 $X2=0
+ $Y2=0
cc_366 N_A_324_79#_c_333_n N_VGND_c_1135_n 0.0148567f $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_367 N_A_324_79#_c_332_n N_VGND_c_1136_n 0.011924f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_368 N_A_324_79#_c_319_n N_VGND_c_1141_n 0.00361406f $X=1.695 $Y=1.34 $X2=0
+ $Y2=0
cc_369 N_A_324_79#_c_324_n N_VGND_c_1141_n 0.00280452f $X=3.095 $Y=1.045 $X2=0
+ $Y2=0
cc_370 N_A_324_79#_c_327_n N_VGND_c_1141_n 0.056759f $X=3.765 $Y=0.355 $X2=0
+ $Y2=0
cc_371 N_A_324_79#_c_328_n N_VGND_c_1141_n 0.0111306f $X=2.975 $Y=0.355 $X2=0
+ $Y2=0
cc_372 N_A_324_79#_c_332_n N_VGND_c_1143_n 0.0705353f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_373 N_A_324_79#_c_333_n N_VGND_c_1143_n 0.0121867f $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_374 N_A_324_79#_c_319_n N_VGND_c_1148_n 0.00218072f $X=1.695 $Y=1.34 $X2=0
+ $Y2=0
cc_375 N_A_324_79#_c_319_n N_VGND_c_1151_n 0.0049796f $X=1.695 $Y=1.34 $X2=0
+ $Y2=0
cc_376 N_A_324_79#_c_324_n N_VGND_c_1151_n 0.00359824f $X=3.095 $Y=1.045 $X2=0
+ $Y2=0
cc_377 N_A_324_79#_c_327_n N_VGND_c_1151_n 0.0346109f $X=3.765 $Y=0.355 $X2=0
+ $Y2=0
cc_378 N_A_324_79#_c_328_n N_VGND_c_1151_n 0.00656177f $X=2.975 $Y=0.355 $X2=0
+ $Y2=0
cc_379 N_A_324_79#_c_332_n N_VGND_c_1151_n 0.0395478f $X=5.445 $Y=0.34 $X2=0
+ $Y2=0
cc_380 N_A_324_79#_c_333_n N_VGND_c_1151_n 0.00660921f $X=4.775 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_324_79#_c_329_n A_744_74# 7.18336e-19 $X=3.85 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_792_48#_M1007_g N_A_634_74#_M1022_g 2.22928e-19 $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_383 N_A_792_48#_c_484_n N_A_634_74#_M1022_g 0.0134232f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_384 N_A_792_48#_c_485_n N_A_634_74#_M1022_g 0.00604334f $X=5.075 $Y=2.24
+ $X2=0 $Y2=0
cc_385 N_A_792_48#_c_486_n N_A_634_74#_M1022_g 0.00714115f $X=5.045 $Y=2.73
+ $X2=0 $Y2=0
cc_386 N_A_792_48#_c_476_n N_A_634_74#_M1022_g 0.00408775f $X=5.185 $Y=1.735
+ $X2=0 $Y2=0
cc_387 N_A_792_48#_c_478_n N_A_634_74#_M1022_g 9.37036e-19 $X=4.125 $Y=1.74
+ $X2=0 $Y2=0
cc_388 N_A_792_48#_c_490_n N_A_634_74#_M1022_g 0.00129846f $X=5.045 $Y=1.9 $X2=0
+ $Y2=0
cc_389 N_A_792_48#_c_491_n N_A_634_74#_M1022_g 0.00205775f $X=5.075 $Y=2.325
+ $X2=0 $Y2=0
cc_390 N_A_792_48#_c_480_n N_A_634_74#_M1022_g 0.0268379f $X=4.27 $Y=1.74 $X2=0
+ $Y2=0
cc_391 N_A_792_48#_M1007_g N_A_634_74#_c_603_n 9.44671e-19 $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_392 N_A_792_48#_M1007_g N_A_634_74#_c_604_n 0.00449852f $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_393 N_A_792_48#_M1014_g N_A_634_74#_c_604_n 0.00749833f $X=4.27 $Y=2.485
+ $X2=0 $Y2=0
cc_394 N_A_792_48#_c_478_n N_A_634_74#_c_604_n 0.0190551f $X=4.125 $Y=1.74 $X2=0
+ $Y2=0
cc_395 N_A_792_48#_M1007_g N_A_634_74#_c_605_n 0.0109782f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_396 N_A_792_48#_c_484_n N_A_634_74#_c_605_n 0.0144756f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_397 N_A_792_48#_c_478_n N_A_634_74#_c_605_n 0.0242156f $X=4.125 $Y=1.74 $X2=0
+ $Y2=0
cc_398 N_A_792_48#_c_480_n N_A_634_74#_c_605_n 0.00326369f $X=4.27 $Y=1.74 $X2=0
+ $Y2=0
cc_399 N_A_792_48#_M1007_g N_A_634_74#_c_608_n 9.69453e-19 $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_400 N_A_792_48#_c_484_n N_A_634_74#_c_608_n 0.0204769f $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_401 N_A_792_48#_c_476_n N_A_634_74#_c_608_n 0.0248004f $X=5.185 $Y=1.735
+ $X2=0 $Y2=0
cc_402 N_A_792_48#_c_490_n N_A_634_74#_c_608_n 0.00401739f $X=5.045 $Y=1.9 $X2=0
+ $Y2=0
cc_403 N_A_792_48#_M1007_g N_A_634_74#_c_609_n 0.00776468f $X=4.035 $Y=0.58
+ $X2=0 $Y2=0
cc_404 N_A_792_48#_c_484_n N_A_634_74#_c_609_n 9.09382e-19 $X=4.88 $Y=1.82 $X2=0
+ $Y2=0
cc_405 N_A_792_48#_c_490_n N_A_634_74#_c_609_n 0.00178976f $X=5.045 $Y=1.9 $X2=0
+ $Y2=0
cc_406 N_A_792_48#_M1007_g N_A_634_74#_c_610_n 0.0093121f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_407 N_A_792_48#_c_476_n N_A_634_74#_c_610_n 0.0122125f $X=5.185 $Y=1.735
+ $X2=0 $Y2=0
cc_408 N_A_792_48#_c_479_n N_A_634_74#_c_610_n 0.00758287f $X=5.11 $Y=0.83 $X2=0
+ $Y2=0
cc_409 N_A_792_48#_c_485_n N_CLK_M1002_g 0.00334108f $X=5.075 $Y=2.24 $X2=0
+ $Y2=0
cc_410 N_A_792_48#_c_486_n N_CLK_M1002_g 0.0111906f $X=5.045 $Y=2.73 $X2=0 $Y2=0
cc_411 N_A_792_48#_c_488_n N_CLK_M1002_g 0.0237889f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_412 N_A_792_48#_c_507_n N_CLK_M1002_g 0.00287335f $X=6.37 $Y=2.24 $X2=0 $Y2=0
cc_413 N_A_792_48#_c_509_n N_CLK_M1002_g 3.21982e-19 $X=6.455 $Y=1.465 $X2=0
+ $Y2=0
cc_414 N_A_792_48#_c_490_n N_CLK_M1002_g 9.86298e-19 $X=5.045 $Y=1.9 $X2=0 $Y2=0
cc_415 N_A_792_48#_c_479_n N_CLK_c_681_n 5.87016e-19 $X=5.11 $Y=0.83 $X2=0 $Y2=0
cc_416 N_A_792_48#_M1019_g N_CLK_M1020_g 0.0186052f $X=7.015 $Y=2.4 $X2=0 $Y2=0
cc_417 N_A_792_48#_c_488_n N_CLK_M1020_g 0.0139224f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_418 N_A_792_48#_c_507_n N_CLK_M1020_g 0.0221652f $X=6.37 $Y=2.24 $X2=0 $Y2=0
cc_419 N_A_792_48#_c_509_n N_CLK_M1020_g 0.00239304f $X=6.455 $Y=1.465 $X2=0
+ $Y2=0
cc_420 N_A_792_48#_c_477_n N_CLK_M1020_g 8.25641e-19 $X=6.865 $Y=1.465 $X2=0
+ $Y2=0
cc_421 N_A_792_48#_M1012_g N_CLK_c_683_n 0.0363224f $X=6.775 $Y=0.74 $X2=0 $Y2=0
cc_422 N_A_792_48#_M1012_g CLK 2.68908e-19 $X=6.775 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A_792_48#_c_509_n CLK 0.0199562f $X=6.455 $Y=1.465 $X2=0 $Y2=0
cc_424 N_A_792_48#_c_488_n N_CLK_c_685_n 0.0028431f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_425 N_A_792_48#_c_509_n N_CLK_c_685_n 0.0148558f $X=6.455 $Y=1.465 $X2=0
+ $Y2=0
cc_426 N_A_792_48#_c_477_n N_CLK_c_685_n 0.00269108f $X=6.865 $Y=1.465 $X2=0
+ $Y2=0
cc_427 N_A_792_48#_c_481_n N_CLK_c_685_n 0.0363224f $X=7.015 $Y=1.465 $X2=0
+ $Y2=0
cc_428 N_A_792_48#_M1019_g N_A_1292_368#_M1009_g 0.0191816f $X=7.015 $Y=2.4
+ $X2=0 $Y2=0
cc_429 N_A_792_48#_M1019_g N_A_1292_368#_c_754_n 0.0140742f $X=7.015 $Y=2.4
+ $X2=0 $Y2=0
cc_430 N_A_792_48#_c_488_n N_A_1292_368#_c_754_n 0.0140087f $X=6.285 $Y=2.325
+ $X2=0 $Y2=0
cc_431 N_A_792_48#_c_507_n N_A_1292_368#_c_754_n 0.0199043f $X=6.37 $Y=2.24
+ $X2=0 $Y2=0
cc_432 N_A_792_48#_M1012_g N_A_1292_368#_c_743_n 0.0119354f $X=6.775 $Y=0.74
+ $X2=0 $Y2=0
cc_433 N_A_792_48#_M1019_g N_A_1292_368#_c_755_n 0.0140935f $X=7.015 $Y=2.4
+ $X2=0 $Y2=0
cc_434 N_A_792_48#_c_477_n N_A_1292_368#_c_755_n 0.00532205f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_435 N_A_792_48#_M1019_g N_A_1292_368#_c_756_n 0.00144884f $X=7.015 $Y=2.4
+ $X2=0 $Y2=0
cc_436 N_A_792_48#_c_507_n N_A_1292_368#_c_756_n 0.0134884f $X=6.37 $Y=2.24
+ $X2=0 $Y2=0
cc_437 N_A_792_48#_c_477_n N_A_1292_368#_c_756_n 0.0280044f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_438 N_A_792_48#_c_481_n N_A_1292_368#_c_756_n 0.00583315f $X=7.015 $Y=1.465
+ $X2=0 $Y2=0
cc_439 N_A_792_48#_M1012_g N_A_1292_368#_c_745_n 0.00395531f $X=6.775 $Y=0.74
+ $X2=0 $Y2=0
cc_440 N_A_792_48#_c_477_n N_A_1292_368#_c_745_n 0.0171756f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_441 N_A_792_48#_c_481_n N_A_1292_368#_c_745_n 0.00716639f $X=7.015 $Y=1.465
+ $X2=0 $Y2=0
cc_442 N_A_792_48#_M1012_g N_A_1292_368#_c_746_n 0.00401978f $X=6.775 $Y=0.74
+ $X2=0 $Y2=0
cc_443 N_A_792_48#_M1019_g N_A_1292_368#_c_747_n 0.00320332f $X=7.015 $Y=2.4
+ $X2=0 $Y2=0
cc_444 N_A_792_48#_c_477_n N_A_1292_368#_c_748_n 0.0175799f $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_445 N_A_792_48#_c_481_n N_A_1292_368#_c_748_n 0.00290882f $X=7.015 $Y=1.465
+ $X2=0 $Y2=0
cc_446 N_A_792_48#_c_477_n N_A_1292_368#_c_749_n 3.3999e-19 $X=6.865 $Y=1.465
+ $X2=0 $Y2=0
cc_447 N_A_792_48#_c_481_n N_A_1292_368#_c_749_n 0.0191816f $X=7.015 $Y=1.465
+ $X2=0 $Y2=0
cc_448 N_A_792_48#_c_484_n N_VPWR_M1014_d 0.002453f $X=4.88 $Y=1.82 $X2=0 $Y2=0
cc_449 N_A_792_48#_c_488_n N_VPWR_M1002_d 0.00822737f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_450 N_A_792_48#_M1014_g N_VPWR_c_865_n 0.0199098f $X=4.27 $Y=2.485 $X2=0
+ $Y2=0
cc_451 N_A_792_48#_c_484_n N_VPWR_c_865_n 0.0197477f $X=4.88 $Y=1.82 $X2=0 $Y2=0
cc_452 N_A_792_48#_c_486_n N_VPWR_c_865_n 0.0170345f $X=5.045 $Y=2.73 $X2=0
+ $Y2=0
cc_453 N_A_792_48#_M1019_g N_VPWR_c_866_n 6.28181e-19 $X=7.015 $Y=2.4 $X2=0
+ $Y2=0
cc_454 N_A_792_48#_c_488_n N_VPWR_c_866_n 0.0219437f $X=6.285 $Y=2.325 $X2=0
+ $Y2=0
cc_455 N_A_792_48#_M1019_g N_VPWR_c_867_n 0.00398325f $X=7.015 $Y=2.4 $X2=0
+ $Y2=0
cc_456 N_A_792_48#_M1019_g N_VPWR_c_871_n 0.005209f $X=7.015 $Y=2.4 $X2=0 $Y2=0
cc_457 N_A_792_48#_M1014_g N_VPWR_c_874_n 0.00492111f $X=4.27 $Y=2.485 $X2=0
+ $Y2=0
cc_458 N_A_792_48#_c_486_n N_VPWR_c_875_n 0.0128035f $X=5.045 $Y=2.73 $X2=0
+ $Y2=0
cc_459 N_A_792_48#_M1014_g N_VPWR_c_862_n 0.00560012f $X=4.27 $Y=2.485 $X2=0
+ $Y2=0
cc_460 N_A_792_48#_M1019_g N_VPWR_c_862_n 0.00983837f $X=7.015 $Y=2.4 $X2=0
+ $Y2=0
cc_461 N_A_792_48#_c_486_n N_VPWR_c_862_n 0.0135456f $X=5.045 $Y=2.73 $X2=0
+ $Y2=0
cc_462 N_A_792_48#_M1007_g N_VGND_c_1135_n 0.00667064f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_463 N_A_792_48#_M1012_g N_VGND_c_1136_n 0.00242918f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_792_48#_c_509_n N_VGND_c_1136_n 0.00198064f $X=6.455 $Y=1.465 $X2=0
+ $Y2=0
cc_465 N_A_792_48#_M1012_g N_VGND_c_1137_n 0.00353511f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_466 N_A_792_48#_M1007_g N_VGND_c_1141_n 0.00444681f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_467 N_A_792_48#_M1012_g N_VGND_c_1145_n 0.00434272f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_468 N_A_792_48#_M1007_g N_VGND_c_1151_n 0.00877228f $X=4.035 $Y=0.58 $X2=0
+ $Y2=0
cc_469 N_A_792_48#_M1012_g N_VGND_c_1151_n 0.00825979f $X=6.775 $Y=0.74 $X2=0
+ $Y2=0
cc_470 N_A_634_74#_M1022_g N_VPWR_c_865_n 0.00561788f $X=4.82 $Y=2.315 $X2=0
+ $Y2=0
cc_471 N_A_634_74#_c_604_n N_VPWR_c_874_n 0.00640144f $X=3.54 $Y=2.07 $X2=0
+ $Y2=0
cc_472 N_A_634_74#_M1022_g N_VPWR_c_875_n 0.00593584f $X=4.82 $Y=2.315 $X2=0
+ $Y2=0
cc_473 N_A_634_74#_M1022_g N_VPWR_c_862_n 0.00622839f $X=4.82 $Y=2.315 $X2=0
+ $Y2=0
cc_474 N_A_634_74#_c_604_n N_VPWR_c_862_n 0.00771299f $X=3.54 $Y=2.07 $X2=0
+ $Y2=0
cc_475 N_A_634_74#_c_604_n N_A_119_143#_c_974_n 0.0183126f $X=3.54 $Y=2.07 $X2=0
+ $Y2=0
cc_476 N_A_634_74#_c_610_n N_VGND_c_1135_n 0.00126498f $X=4.785 $Y=1.235 $X2=0
+ $Y2=0
cc_477 N_A_634_74#_c_610_n N_VGND_c_1143_n 0.00278271f $X=4.785 $Y=1.235 $X2=0
+ $Y2=0
cc_478 N_A_634_74#_c_610_n N_VGND_c_1151_n 0.00361311f $X=4.785 $Y=1.235 $X2=0
+ $Y2=0
cc_479 N_CLK_M1020_g N_A_1292_368#_c_754_n 0.0118845f $X=6.37 $Y=2.4 $X2=0 $Y2=0
cc_480 N_CLK_c_683_n N_A_1292_368#_c_743_n 0.00172581f $X=6.385 $Y=1.22 $X2=0
+ $Y2=0
cc_481 N_CLK_M1020_g N_A_1292_368#_c_756_n 0.00145089f $X=6.37 $Y=2.4 $X2=0
+ $Y2=0
cc_482 N_CLK_c_683_n N_A_1292_368#_c_745_n 7.3019e-19 $X=6.385 $Y=1.22 $X2=0
+ $Y2=0
cc_483 N_CLK_M1002_g N_VPWR_c_866_n 0.00419332f $X=5.835 $Y=2.26 $X2=0 $Y2=0
cc_484 N_CLK_M1020_g N_VPWR_c_866_n 0.0123708f $X=6.37 $Y=2.4 $X2=0 $Y2=0
cc_485 N_CLK_M1020_g N_VPWR_c_871_n 0.00460063f $X=6.37 $Y=2.4 $X2=0 $Y2=0
cc_486 N_CLK_M1002_g N_VPWR_c_875_n 0.00482866f $X=5.835 $Y=2.26 $X2=0 $Y2=0
cc_487 N_CLK_M1002_g N_VPWR_c_862_n 0.00555093f $X=5.835 $Y=2.26 $X2=0 $Y2=0
cc_488 N_CLK_M1020_g N_VPWR_c_862_n 0.00910231f $X=6.37 $Y=2.4 $X2=0 $Y2=0
cc_489 N_CLK_c_681_n N_VGND_c_1136_n 0.00470925f $X=5.885 $Y=1.22 $X2=0 $Y2=0
cc_490 N_CLK_c_683_n N_VGND_c_1136_n 0.0156468f $X=6.385 $Y=1.22 $X2=0 $Y2=0
cc_491 CLK N_VGND_c_1136_n 0.00899f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_492 N_CLK_c_685_n N_VGND_c_1136_n 0.00507991f $X=6.385 $Y=1.385 $X2=0 $Y2=0
cc_493 N_CLK_c_681_n N_VGND_c_1143_n 0.00430908f $X=5.885 $Y=1.22 $X2=0 $Y2=0
cc_494 N_CLK_c_683_n N_VGND_c_1145_n 0.00383152f $X=6.385 $Y=1.22 $X2=0 $Y2=0
cc_495 N_CLK_c_681_n N_VGND_c_1151_n 0.00821115f $X=5.885 $Y=1.22 $X2=0 $Y2=0
cc_496 N_CLK_c_683_n N_VGND_c_1151_n 0.0075725f $X=6.385 $Y=1.22 $X2=0 $Y2=0
cc_497 N_A_1292_368#_c_755_n N_VPWR_M1019_d 0.0021473f $X=7.365 $Y=1.885 $X2=0
+ $Y2=0
cc_498 N_A_1292_368#_c_754_n N_VPWR_c_866_n 0.0193839f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_1292_368#_M1009_g N_VPWR_c_867_n 0.0173258f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_500 N_A_1292_368#_M1010_g N_VPWR_c_867_n 7.732e-19 $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_501 N_A_1292_368#_c_754_n N_VPWR_c_867_n 0.0323093f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_502 N_A_1292_368#_c_755_n N_VPWR_c_867_n 0.0191623f $X=7.365 $Y=1.885 $X2=0
+ $Y2=0
cc_503 N_A_1292_368#_M1010_g N_VPWR_c_868_n 0.00366558f $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_504 N_A_1292_368#_M1016_g N_VPWR_c_868_n 0.00250919f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_505 N_A_1292_368#_M1016_g N_VPWR_c_870_n 6.51372e-19 $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_506 N_A_1292_368#_M1018_g N_VPWR_c_870_n 0.0206339f $X=9.09 $Y=2.4 $X2=0
+ $Y2=0
cc_507 N_A_1292_368#_c_754_n N_VPWR_c_871_n 0.014549f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_508 N_A_1292_368#_M1009_g N_VPWR_c_876_n 0.00460063f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_509 N_A_1292_368#_M1010_g N_VPWR_c_876_n 0.005209f $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_510 N_A_1292_368#_M1016_g N_VPWR_c_877_n 0.005209f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_511 N_A_1292_368#_M1018_g N_VPWR_c_877_n 0.00475445f $X=9.09 $Y=2.4 $X2=0
+ $Y2=0
cc_512 N_A_1292_368#_M1009_g N_VPWR_c_862_n 0.00909733f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_513 N_A_1292_368#_M1010_g N_VPWR_c_862_n 0.00983932f $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_514 N_A_1292_368#_M1016_g N_VPWR_c_862_n 0.00982524f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_515 N_A_1292_368#_M1018_g N_VPWR_c_862_n 0.00939102f $X=9.09 $Y=2.4 $X2=0
+ $Y2=0
cc_516 N_A_1292_368#_c_754_n N_VPWR_c_862_n 0.0119743f $X=6.79 $Y=1.985 $X2=0
+ $Y2=0
cc_517 N_A_1292_368#_M1009_g N_GCLK_c_1067_n 0.0126934f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_518 N_A_1292_368#_M1010_g N_GCLK_c_1067_n 0.014651f $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_519 N_A_1292_368#_M1016_g N_GCLK_c_1067_n 6.79538e-19 $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_520 N_A_1292_368#_M1000_g N_GCLK_c_1062_n 4.94129e-19 $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_1292_368#_M1003_g N_GCLK_c_1062_n 4.49298e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_522 N_A_1292_368#_M1010_g N_GCLK_c_1068_n 0.0132272f $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_523 N_A_1292_368#_M1016_g N_GCLK_c_1068_n 0.015411f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_524 N_A_1292_368#_c_809_p N_GCLK_c_1068_n 0.0294689f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_525 N_A_1292_368#_c_749_n N_GCLK_c_1068_n 0.00367077f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_526 N_A_1292_368#_M1009_g N_GCLK_c_1069_n 0.00152174f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_527 N_A_1292_368#_M1010_g N_GCLK_c_1069_n 0.00140601f $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_528 N_A_1292_368#_c_755_n N_GCLK_c_1069_n 0.0149283f $X=7.365 $Y=1.885 $X2=0
+ $Y2=0
cc_529 N_A_1292_368#_c_809_p N_GCLK_c_1069_n 0.0276965f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_530 N_A_1292_368#_c_749_n N_GCLK_c_1069_n 0.00572037f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_531 N_A_1292_368#_M1003_g N_GCLK_c_1063_n 0.0124838f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_532 N_A_1292_368#_M1015_g N_GCLK_c_1063_n 0.0140403f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_533 N_A_1292_368#_c_809_p N_GCLK_c_1063_n 0.0234532f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_534 N_A_1292_368#_c_749_n N_GCLK_c_1063_n 0.00298567f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_535 N_A_1292_368#_M1000_g N_GCLK_c_1064_n 2.44239e-19 $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_536 N_A_1292_368#_c_744_n N_GCLK_c_1064_n 0.0053088f $X=7.365 $Y=1.045 $X2=0
+ $Y2=0
cc_537 N_A_1292_368#_c_809_p N_GCLK_c_1064_n 0.0210853f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_538 N_A_1292_368#_c_749_n N_GCLK_c_1064_n 0.00408598f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_539 N_A_1292_368#_M1010_g N_GCLK_c_1070_n 6.46654e-19 $X=8.095 $Y=2.4 $X2=0
+ $Y2=0
cc_540 N_A_1292_368#_M1016_g N_GCLK_c_1070_n 0.013943f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_541 N_A_1292_368#_M1018_g N_GCLK_c_1070_n 4.36913e-19 $X=9.09 $Y=2.4 $X2=0
+ $Y2=0
cc_542 N_A_1292_368#_M1003_g N_GCLK_c_1065_n 6.74842e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_543 N_A_1292_368#_M1015_g N_GCLK_c_1065_n 0.00889459f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_A_1292_368#_M1027_g N_GCLK_c_1065_n 0.00783249f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_545 N_A_1292_368#_M1016_g N_GCLK_c_1066_n 0.00457227f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_546 N_A_1292_368#_M1018_g N_GCLK_c_1066_n 0.00472196f $X=9.09 $Y=2.4 $X2=0
+ $Y2=0
cc_547 N_A_1292_368#_c_749_n N_GCLK_c_1066_n 0.0216837f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_548 N_A_1292_368#_M1016_g N_GCLK_c_1072_n 0.00175698f $X=8.595 $Y=2.4 $X2=0
+ $Y2=0
cc_549 N_A_1292_368#_M1018_g N_GCLK_c_1072_n 8.65021e-19 $X=9.09 $Y=2.4 $X2=0
+ $Y2=0
cc_550 N_A_1292_368#_M1003_g N_GCLK_c_1106_n 9.05544e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_551 N_A_1292_368#_M1015_g N_GCLK_c_1106_n 0.00624222f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_552 N_A_1292_368#_M1027_g N_GCLK_c_1106_n 0.0114427f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_553 N_A_1292_368#_c_809_p N_GCLK_c_1106_n 0.0168342f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_554 N_A_1292_368#_c_749_n N_GCLK_c_1106_n 0.0160322f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_555 N_A_1292_368#_c_744_n N_VGND_M1000_d 0.00421825f $X=7.365 $Y=1.045 $X2=0
+ $Y2=0
cc_556 N_A_1292_368#_c_743_n N_VGND_c_1136_n 0.0193094f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_557 N_A_1292_368#_c_745_n N_VGND_c_1136_n 0.00168579f $X=7.155 $Y=1.045 $X2=0
+ $Y2=0
cc_558 N_A_1292_368#_M1000_g N_VGND_c_1137_n 0.00416717f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_A_1292_368#_c_743_n N_VGND_c_1137_n 0.0290535f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_560 N_A_1292_368#_c_744_n N_VGND_c_1137_n 0.0135013f $X=7.365 $Y=1.045 $X2=0
+ $Y2=0
cc_561 N_A_1292_368#_c_809_p N_VGND_c_1137_n 0.00344427f $X=8.27 $Y=1.465 $X2=0
+ $Y2=0
cc_562 N_A_1292_368#_c_749_n N_VGND_c_1137_n 0.00252623f $X=9.105 $Y=1.465 $X2=0
+ $Y2=0
cc_563 N_A_1292_368#_M1000_g N_VGND_c_1138_n 4.61576e-19 $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_564 N_A_1292_368#_M1003_g N_VGND_c_1138_n 0.00903345f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_565 N_A_1292_368#_M1015_g N_VGND_c_1138_n 0.00307459f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_566 N_A_1292_368#_M1027_g N_VGND_c_1140_n 0.00647412f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_567 N_A_1292_368#_c_743_n N_VGND_c_1145_n 0.0145639f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_568 N_A_1292_368#_M1000_g N_VGND_c_1146_n 0.00461464f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_569 N_A_1292_368#_M1003_g N_VGND_c_1146_n 0.00383152f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_570 N_A_1292_368#_M1015_g N_VGND_c_1147_n 0.00434272f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_571 N_A_1292_368#_M1027_g N_VGND_c_1147_n 0.00434272f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_572 N_A_1292_368#_M1000_g N_VGND_c_1151_n 0.0091381f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_573 N_A_1292_368#_M1003_g N_VGND_c_1151_n 0.00758019f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_574 N_A_1292_368#_M1015_g N_VGND_c_1151_n 0.00820284f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_575 N_A_1292_368#_M1027_g N_VGND_c_1151_n 0.00823942f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_576 N_A_1292_368#_c_743_n N_VGND_c_1151_n 0.0119984f $X=6.99 $Y=0.515 $X2=0
+ $Y2=0
cc_577 N_VPWR_M1004_s N_A_119_143#_c_974_n 0.0183801f $X=1.565 $Y=2.12 $X2=0
+ $Y2=0
cc_578 N_VPWR_c_874_n N_A_119_143#_c_974_n 0.00751736f $X=4.43 $Y=3.33 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_862_n N_A_119_143#_c_974_n 0.0319205f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_580 N_VPWR_c_864_n N_A_119_143#_c_976_n 0.0103229f $X=0.28 $Y=2.12 $X2=0
+ $Y2=0
cc_581 N_VPWR_c_873_n N_A_119_143#_c_976_n 0.00870779f $X=1.545 $Y=3.33 $X2=0
+ $Y2=0
cc_582 N_VPWR_c_878_n N_A_119_143#_c_976_n 0.0130874f $X=1.99 $Y=2.775 $X2=0
+ $Y2=0
cc_583 N_VPWR_c_862_n N_A_119_143#_c_976_n 0.0106996f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_584 N_VPWR_M1004_s N_A_119_143#_c_977_n 0.00614178f $X=1.565 $Y=2.12 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_864_n N_A_119_143#_c_977_n 0.016114f $X=0.28 $Y=2.12 $X2=0 $Y2=0
cc_586 N_VPWR_c_878_n N_A_119_143#_c_977_n 0.0448167f $X=1.99 $Y=2.775 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_862_n N_A_119_143#_c_977_n 0.0108289f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_867_n N_GCLK_c_1067_n 0.0485389f $X=7.29 $Y=2.305 $X2=0 $Y2=0
cc_589 N_VPWR_c_868_n N_GCLK_c_1067_n 0.0283501f $X=8.32 $Y=2.305 $X2=0 $Y2=0
cc_590 N_VPWR_c_876_n N_GCLK_c_1067_n 0.014549f $X=8.235 $Y=3.33 $X2=0 $Y2=0
cc_591 N_VPWR_c_862_n N_GCLK_c_1067_n 0.0119743f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_M1010_s N_GCLK_c_1068_n 0.00218982f $X=8.185 $Y=1.84 $X2=0 $Y2=0
cc_593 N_VPWR_c_868_n N_GCLK_c_1068_n 0.0167599f $X=8.32 $Y=2.305 $X2=0 $Y2=0
cc_594 N_VPWR_c_868_n N_GCLK_c_1070_n 0.0322767f $X=8.32 $Y=2.305 $X2=0 $Y2=0
cc_595 N_VPWR_c_870_n N_GCLK_c_1070_n 0.0386881f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_596 N_VPWR_c_877_n N_GCLK_c_1070_n 0.014549f $X=9.155 $Y=3.33 $X2=0 $Y2=0
cc_597 N_VPWR_c_862_n N_GCLK_c_1070_n 0.0119743f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_598 N_VPWR_c_870_n N_GCLK_c_1072_n 0.00654083f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_599 N_VPWR_c_864_n N_VGND_c_1133_n 3.21545e-19 $X=0.28 $Y=2.12 $X2=0 $Y2=0
cc_600 N_A_119_143#_c_968_n N_VGND_M1026_d 0.0155317f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_601 N_A_119_143#_c_970_n N_VGND_M1026_d 0.00677158f $X=1.57 $Y=1.955 $X2=0
+ $Y2=0
cc_602 N_A_119_143#_c_1021_n N_VGND_M1026_d 8.26265e-19 $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_603 N_A_119_143#_c_967_n N_VGND_c_1133_n 0.0178065f $X=0.78 $Y=0.99 $X2=0
+ $Y2=0
cc_604 N_A_119_143#_c_969_n N_VGND_c_1133_n 0.00875128f $X=0.945 $Y=0.7 $X2=0
+ $Y2=0
cc_605 N_A_119_143#_c_968_n N_VGND_c_1134_n 0.00317977f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_606 N_A_119_143#_c_969_n N_VGND_c_1134_n 0.00690349f $X=0.945 $Y=0.7 $X2=0
+ $Y2=0
cc_607 N_A_119_143#_c_1021_n N_VGND_c_1141_n 0.0012259f $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_608 N_A_119_143#_c_971_n N_VGND_c_1141_n 0.0144289f $X=2.525 $Y=0.62 $X2=0
+ $Y2=0
cc_609 N_A_119_143#_c_972_n N_VGND_c_1141_n 0.011464f $X=2.305 $Y=0.622 $X2=0
+ $Y2=0
cc_610 N_A_119_143#_c_968_n N_VGND_c_1148_n 0.027214f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_611 N_A_119_143#_c_1021_n N_VGND_c_1148_n 0.00659988f $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_612 N_A_119_143#_c_968_n N_VGND_c_1151_n 0.00679534f $X=1.485 $Y=0.7 $X2=0
+ $Y2=0
cc_613 N_A_119_143#_c_969_n N_VGND_c_1151_n 0.0101259f $X=0.945 $Y=0.7 $X2=0
+ $Y2=0
cc_614 N_A_119_143#_c_1021_n N_VGND_c_1151_n 0.00319493f $X=1.57 $Y=0.7 $X2=0
+ $Y2=0
cc_615 N_A_119_143#_c_971_n N_VGND_c_1151_n 0.0120887f $X=2.525 $Y=0.62 $X2=0
+ $Y2=0
cc_616 N_A_119_143#_c_972_n N_VGND_c_1151_n 0.0187306f $X=2.305 $Y=0.622 $X2=0
+ $Y2=0
cc_617 N_GCLK_c_1063_n N_VGND_M1003_d 0.00176461f $X=8.725 $Y=1.045 $X2=0 $Y2=0
cc_618 N_GCLK_c_1062_n N_VGND_c_1137_n 0.00122648f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_619 N_GCLK_c_1062_n N_VGND_c_1138_n 0.0158413f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_620 N_GCLK_c_1063_n N_VGND_c_1138_n 0.0153337f $X=8.725 $Y=1.045 $X2=0 $Y2=0
cc_621 N_GCLK_c_1065_n N_VGND_c_1138_n 0.0164981f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_622 N_GCLK_c_1065_n N_VGND_c_1140_n 0.0293763f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_623 N_GCLK_c_1062_n N_VGND_c_1146_n 0.011066f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_624 N_GCLK_c_1065_n N_VGND_c_1147_n 0.0144922f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_625 N_GCLK_c_1062_n N_VGND_c_1151_n 0.00915947f $X=8.03 $Y=0.515 $X2=0 $Y2=0
cc_626 N_GCLK_c_1065_n N_VGND_c_1151_n 0.0118826f $X=8.89 $Y=0.515 $X2=0 $Y2=0

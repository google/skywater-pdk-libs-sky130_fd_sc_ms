* File: sky130_fd_sc_ms__einvn_1.pex.spice
* Created: Wed Sep  2 12:08:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EINVN_1%TE_B 3 5 7 8 10 12 18 24 26
c47 5 0 7.54751e-20 $X=0.82 $Y=1.43
r48 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.82 $Y=1.595
+ $X2=0.895 $Y2=1.595
r49 22 23 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.78 $Y=1.595 $X2=0.82
+ $Y2=1.595
r50 18 26 3.83775 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=1.085 $Y2=1.605
r51 16 22 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.62 $Y=1.595
+ $X2=0.78 $Y2=1.595
r52 15 26 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.62 $Y=1.595
+ $X2=1.085 $Y2=1.595
r53 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.595 $X2=0.62 $Y2=1.595
r54 10 12 171.378 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=1.315 $Y=1.76
+ $X2=1.315 $Y2=2.4
r55 8 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.225 $Y=1.685
+ $X2=1.315 $Y2=1.76
r56 8 24 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.225 $Y=1.685
+ $X2=0.895 $Y2=1.685
r57 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.82 $Y=1.43
+ $X2=0.82 $Y2=1.595
r58 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.82 $Y=1.43 $X2=0.82
+ $Y2=1.11
r59 1 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.78 $Y=1.76
+ $X2=0.78 $Y2=1.595
r60 1 3 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=0.78 $Y=1.76 $X2=0.78
+ $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_1%A_22_46# 1 2 9 11 13 15 17 21 22 26 31 34
c45 21 0 1.65003e-19 $X=0.615 $Y=0.395
r46 28 31 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.195 $Y=2.015
+ $X2=0.555 $Y2=2.015
r47 26 27 10.5469 $w=6.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=1.085
+ $X2=0.44 $Y2=1.25
r48 22 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.615 $Y=0.395
+ $X2=0.78 $Y2=0.395
r49 21 24 2.94557 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.395
+ $X2=0.445 $Y2=0.56
r50 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=0.395 $X2=0.615 $Y2=0.395
r51 17 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.195 $Y=1.93
+ $X2=0.195 $Y2=2.015
r52 17 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.195 $Y=1.93
+ $X2=0.195 $Y2=1.25
r53 15 26 2.9902 $w=6.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=0.92
+ $X2=0.44 $Y2=1.085
r54 15 24 6.52406 $w=6.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.44 $Y=0.92
+ $X2=0.44 $Y2=0.56
r55 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.33 $Y=0.425
+ $X2=1.33 $Y2=0.87
r56 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.255 $Y=0.35
+ $X2=1.33 $Y2=0.425
r57 9 34 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.255 $Y=0.35
+ $X2=0.78 $Y2=0.35
r58 2 31 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.41
+ $Y=1.92 $X2=0.555 $Y2=2.075
r59 1 26 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=0.455
+ $Y=0.9 $X2=0.605 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_1%A 3 6 8 11 12 13
r33 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.515
+ $X2=1.81 $Y2=1.68
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.515
+ $X2=1.81 $Y2=1.35
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.515 $X2=1.81 $Y2=1.515
r36 8 12 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=1.77 $Y=1.665
+ $X2=1.77 $Y2=1.515
r37 6 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.735 $Y=2.4
+ $X2=1.735 $Y2=1.68
r38 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.72 $Y=0.87 $X2=1.72
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_1%VPWR 1 6 10 12 19 20 23
r24 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r25 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.09 $Y2=3.33
r26 17 19 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.09 $Y2=3.33
r29 12 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 10 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 6 9 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=2.115 $X2=1.09
+ $Y2=2.815
r34 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=3.245 $X2=1.09
+ $Y2=3.33
r35 4 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.09 $Y=3.245 $X2=1.09
+ $Y2=2.815
r36 1 9 600 $w=1.7e-07 $l=9.98962e-07 $layer=licon1_PDIFF $count=1 $X=0.87
+ $Y=1.92 $X2=1.09 $Y2=2.815
r37 1 6 300 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_PDIFF $count=2 $X=0.87
+ $Y=1.92 $X2=1.09 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_1%Z 1 2 11 12 14 17 18
r24 18 26 0.869875 $w=5.48e-07 $l=4e-08 $layer=LI1_cond $X=2.04 $Y=2.775
+ $X2=2.04 $Y2=2.815
r25 17 18 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.04 $Y=2.405
+ $X2=2.04 $Y2=2.775
r26 14 16 17.9201 $w=5.43e-07 $l=5.35e-07 $layer=LI1_cond $X=2.042 $Y=0.645
+ $X2=2.042 $Y2=1.18
r27 12 16 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.23 $Y=1.95
+ $X2=2.23 $Y2=1.18
r28 11 12 8.09223 $w=5.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.035
+ $X2=2.04 $Y2=1.95
r29 9 17 3.91444 $w=5.48e-07 $l=1.8e-07 $layer=LI1_cond $X=2.04 $Y=2.225
+ $X2=2.04 $Y2=2.405
r30 9 11 4.13191 $w=5.48e-07 $l=1.9e-07 $layer=LI1_cond $X=2.04 $Y=2.225
+ $X2=2.04 $Y2=2.035
r31 2 26 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.84 $X2=1.96 $Y2=2.815
r32 2 11 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.84 $X2=1.96 $Y2=2.035
r33 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.795
+ $Y=0.5 $X2=1.935 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_1%VGND 1 6 10 12 19 20 23
c27 20 0 6.02012e-21 $X=2.16 $Y=0
r28 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r29 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.115
+ $Y2=0
r30 17 19 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=2.16
+ $Y2=0
r31 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r32 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.115
+ $Y2=0
r33 12 14 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.72
+ $Y2=0
r34 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r35 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r36 10 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r37 6 8 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.115 $Y=0.645
+ $X2=1.115 $Y2=1.095
r38 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r39 4 6 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.645
r40 1 8 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=0.895
+ $Y=0.9 $X2=1.115 $Y2=1.095
r41 1 6 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=0.895
+ $Y=0.9 $X2=1.115 $Y2=0.645
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
X0 VPWR a_27_120# a_588_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 Q a_842_405# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_672_392# a_369_392# a_875_139# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_588_392# a_369_392# a_672_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_794_503# a_842_405# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X5 a_369_392# a_232_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 VPWR a_672_392# a_842_405# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VGND GATE_N a_232_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_672_392# a_842_405# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND a_842_405# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Q a_842_405# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_27_120# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X12 a_369_392# a_232_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_672_392# a_232_82# a_794_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X14 a_658_79# a_232_82# a_672_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VPWR GATE_N a_232_82# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X16 a_875_139# a_842_405# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 VPWR a_842_405# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 VGND a_27_120# a_658_79# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_27_120# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
.ends

* File: sky130_fd_sc_ms__a222o_1.spice
* Created: Wed Sep  2 11:52:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a222o_1.pex.spice"
.subckt sky130_fd_sc_ms__a222o_1  VNB VPB C1 C2 B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1005 A_119_74# N_C1_M1005_g N_A_32_74#_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_C2_M1000_g A_119_74# VNB NLOWVT L=0.15 W=0.64 AD=0.2544
+ AS=0.0768 PD=1.435 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75000.6 SB=75003.6
+ A=0.096 P=1.58 MULT=1
MM1006 A_386_74# N_B2_M1006_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.2544 PD=0.88 PS=1.435 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75001.5 SB=75002.7
+ A=0.096 P=1.58 MULT=1
MM1007 N_A_32_74#_M1007_d N_B1_M1007_g A_386_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.2512 AS=0.0768 PD=1.425 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.9
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1004 A_651_74# N_A1_M1004_g N_A_32_74#_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.2512 PD=0.88 PS=1.425 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75002.9
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g A_651_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.185229 AS=0.0768 PD=1.22899 PS=0.88 NRD=21.552 NRS=12.18 M=1 R=4.26667
+ SA=75003.3 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1002 N_X_M1002_d N_A_32_74#_M1002_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.214171 PD=2.05 PS=1.42101 NRD=0 NRS=30.804 M=1 R=4.93333
+ SA=75003.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_32_74#_M1001_d N_C1_M1001_g N_A_27_390#_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.2125 AS=0.28 PD=1.425 PS=2.56 NRD=29.55 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_390#_M1009_d N_C2_M1009_g N_A_32_74#_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.2125 PD=1.32 PS=1.425 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.8
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1008 N_A_340_390#_M1008_d N_B2_M1008_g N_A_27_390#_M1009_d VPB PSHORT L=0.18
+ W=1 AD=0.205 AS=0.16 PD=1.41 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90001.3
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1010 N_A_27_390#_M1010_d N_B1_M1010_g N_A_340_390#_M1008_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.205 PD=2.56 PS=1.41 NRD=0 NRS=16.7253 M=1 R=5.55556
+ SA=90001.9 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_A_340_390#_M1011_d N_A1_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.33 PD=1.27 PS=2.66 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.2
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A2_M1012_g N_A_340_390#_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.206887 AS=0.135 PD=1.43868 PS=1.27 NRD=15.7403 NRS=0 M=1 R=5.55556
+ SA=90000.7 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1013 N_X_M1013_d N_A_32_74#_M1013_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.231713 PD=2.8 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__a222o_1.pxi.spice"
*
.ends
*
*

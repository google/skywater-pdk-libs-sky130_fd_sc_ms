* File: sky130_fd_sc_ms__and4_4.pex.spice
* Created: Fri Aug 28 17:13:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4_4%A 1 3 6 10 14 16 23
c51 16 0 5.84547e-20 $X=1.2 $Y=1.665
r52 21 23 21.3457 $w=3.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.225 $Y=1.66
+ $X2=1.38 $Y2=1.66
r53 19 21 37.1829 $w=3.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.955 $Y=1.66
+ $X2=1.225 $Y2=1.66
r54 18 19 0.688571 $w=3.5e-07 $l=5e-09 $layer=POLY_cond $X=0.95 $Y=1.66
+ $X2=0.955 $Y2=1.66
r55 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.615 $X2=1.225 $Y2=1.615
r56 12 23 3.44286 $w=3.5e-07 $l=2.5e-08 $layer=POLY_cond $X=1.405 $Y=1.66
+ $X2=1.38 $Y2=1.66
r57 12 14 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.405 $Y=1.78
+ $X2=1.405 $Y2=2.46
r58 8 23 22.6286 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.38 $Y=1.45 $X2=1.38
+ $Y2=1.66
r59 8 10 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.38 $Y=1.45 $X2=1.38
+ $Y2=0.915
r60 4 18 22.6286 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.95 $Y=1.45 $X2=0.95
+ $Y2=1.66
r61 4 6 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.95 $Y=1.45 $X2=0.95
+ $Y2=0.915
r62 1 19 18.307 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.955 $Y=1.87
+ $X2=0.955 $Y2=1.66
r63 1 3 157.989 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=0.955 $Y=1.87
+ $X2=0.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%B 3 8 9 10 14 17 19 22 23 24 27 28
c65 22 0 5.28639e-20 $X=1.832 $Y=1.46
c66 19 0 2.53319e-19 $X=1.87 $Y=2.46
c67 17 0 1.26182e-19 $X=1.87 $Y=1.79
r68 27 30 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.78
r69 27 29 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.615
+ $X2=0.407 $Y2=1.45
r70 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r71 24 28 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r72 22 23 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.855 $Y=1.46
+ $X2=1.855 $Y2=1.7
r73 21 22 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=1.832 $Y=1.31
+ $X2=1.832 $Y2=1.46
r74 17 23 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.87 $Y=1.79 $X2=1.87
+ $Y2=1.7
r75 17 19 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=1.87 $Y=1.79
+ $X2=1.87 $Y2=2.46
r76 14 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.81 $Y=0.915
+ $X2=1.81 $Y2=1.31
r77 11 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.81 $Y=0.255
+ $X2=1.81 $Y2=0.915
r78 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.735 $Y=0.18
+ $X2=1.81 $Y2=0.255
r79 9 10 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=1.735 $Y=0.18
+ $X2=0.595 $Y2=0.18
r80 8 29 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.52 $Y=0.915
+ $X2=0.52 $Y2=1.45
r81 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.52 $Y=0.255
+ $X2=0.595 $Y2=0.18
r82 5 8 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.52 $Y=0.255 $X2=0.52
+ $Y2=0.915
r83 3 30 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.505 $Y=2.46
+ $X2=0.505 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%D 1 3 6 8 10 11 12 15 17
c57 17 0 4.10416e-20 $X=3.12 $Y=1.665
c58 15 0 1.72297e-19 $X=3.705 $Y=2.46
r59 22 24 19.9323 $w=3.99e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.572
+ $X2=3.26 $Y2=1.572
r60 20 22 33.2206 $w=3.99e-07 $l=2.75e-07 $layer=POLY_cond $X=2.82 $Y=1.572
+ $X2=3.095 $Y2=1.572
r61 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=1.635 $X2=3.095 $Y2=1.635
r62 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.705 $Y=1.8
+ $X2=3.705 $Y2=2.46
r63 12 24 28.6936 $w=3.99e-07 $l=1.86773e-07 $layer=POLY_cond $X=3.335 $Y=1.725
+ $X2=3.26 $Y2=1.572
r64 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.615 $Y=1.725
+ $X2=3.705 $Y2=1.8
r65 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.615 $Y=1.725
+ $X2=3.335 $Y2=1.725
r66 8 24 25.8008 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=3.26 $Y=1.345
+ $X2=3.26 $Y2=1.572
r67 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.26 $Y=1.345
+ $X2=3.26 $Y2=0.915
r68 4 20 21.4026 $w=1.8e-07 $l=2.28e-07 $layer=POLY_cond $X=2.82 $Y=1.8 $X2=2.82
+ $Y2=1.572
r69 4 6 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.82 $Y=1.8 $X2=2.82
+ $Y2=2.46
r70 1 20 18.1203 $w=3.99e-07 $l=2.92539e-07 $layer=POLY_cond $X=2.67 $Y=1.345
+ $X2=2.82 $Y2=1.572
r71 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.67 $Y=1.345 $X2=2.67
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%C 4 9 10 11 14 16 20 23 25 26 27 28 29 32 33
c97 27 0 4.10416e-20 $X=2.347 $Y=1.885
r98 32 34 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.2 $Y=1.51 $X2=4.2
+ $Y2=1.675
r99 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.2
+ $Y=1.51 $X2=4.2 $Y2=1.51
r100 29 33 4.63971 $w=3.83e-07 $l=1.55e-07 $layer=LI1_cond $X=4.172 $Y=1.665
+ $X2=4.172 $Y2=1.51
r101 26 27 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.347 $Y=1.735
+ $X2=2.347 $Y2=1.885
r102 25 26 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.31 $Y=1.46
+ $X2=2.31 $Y2=1.735
r103 24 25 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.275 $Y=1.31
+ $X2=2.275 $Y2=1.46
r104 23 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.2 $Y=1.345
+ $X2=4.2 $Y2=1.51
r105 22 23 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=4.2 $Y=0.255
+ $X2=4.2 $Y2=1.345
r106 20 34 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=4.205 $Y=2.46
+ $X2=4.205 $Y2=1.675
r107 17 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=0.18
+ $X2=3.69 $Y2=0.18
r108 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.125 $Y=0.18
+ $X2=4.2 $Y2=0.255
r109 16 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.125 $Y=0.18
+ $X2=3.765 $Y2=0.18
r110 12 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=0.255
+ $X2=3.69 $Y2=0.18
r111 12 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.69 $Y=0.255
+ $X2=3.69 $Y2=0.915
r112 10 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.615 $Y=0.18
+ $X2=3.69 $Y2=0.18
r113 10 11 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=3.615 $Y=0.18
+ $X2=2.315 $Y2=0.18
r114 9 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.37 $Y=2.46
+ $X2=2.37 $Y2=1.885
r115 4 24 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.24 $Y=0.915
+ $X2=2.24 $Y2=1.31
r116 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.24 $Y=0.255
+ $X2=2.315 $Y2=0.18
r117 1 4 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.24 $Y=0.255
+ $X2=2.24 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%A_119_392# 1 2 3 4 5 18 22 26 30 34 38 42 46
+ 49 50 52 54 57 60 62 63 65 68 70 74 76 79 80 85 91 93 95 106
c199 91 0 1.61898e-19 $X=1.645 $Y=2.105
c200 79 0 1.74227e-19 $X=4.62 $Y=1.95
c201 74 0 1.72297e-19 $X=3.98 $Y=2.815
c202 65 0 1.55561e-20 $X=2.595 $Y=1.97
c203 60 0 1.51907e-19 $X=1.645 $Y=2.46
c204 50 0 1.43623e-19 $X=0.89 $Y=1.13
c205 18 0 1.8401e-19 $X=4.75 $Y=0.74
r206 105 106 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.14 $Y=1.465
+ $X2=6.165 $Y2=1.465
r207 104 105 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=5.715 $Y=1.465
+ $X2=6.14 $Y2=1.465
r208 103 104 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=5.71 $Y=1.465
+ $X2=5.715 $Y2=1.465
r209 100 101 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=5.21 $Y=1.465
+ $X2=5.265 $Y2=1.465
r210 96 98 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.75 $Y=1.465
+ $X2=4.765 $Y2=1.465
r211 86 103 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=5.52 $Y=1.465
+ $X2=5.71 $Y2=1.465
r212 86 101 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=5.52 $Y=1.465
+ $X2=5.265 $Y2=1.465
r213 85 86 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.465 $X2=5.52 $Y2=1.465
r214 83 100 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=4.84 $Y=1.465
+ $X2=5.21 $Y2=1.465
r215 83 98 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.84 $Y=1.465
+ $X2=4.765 $Y2=1.465
r216 82 85 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.84 $Y=1.465
+ $X2=5.52 $Y2=1.465
r217 82 83 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.84
+ $Y=1.465 $X2=4.84 $Y2=1.465
r218 80 82 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.705 $Y=1.465
+ $X2=4.84 $Y2=1.465
r219 78 80 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.62 $Y=1.63
+ $X2=4.705 $Y2=1.465
r220 78 79 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.62 $Y=1.63
+ $X2=4.62 $Y2=1.95
r221 77 95 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=4.145 $Y=2.035
+ $X2=3.98 $Y2=2.045
r222 76 79 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.535 $Y=2.035
+ $X2=4.62 $Y2=1.95
r223 76 77 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.535 $Y=2.035
+ $X2=4.145 $Y2=2.035
r224 72 95 0.89609 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.98 $Y=2.14
+ $X2=3.98 $Y2=2.045
r225 72 74 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.98 $Y=2.14
+ $X2=3.98 $Y2=2.815
r226 71 93 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=2.055
+ $X2=2.595 $Y2=2.055
r227 70 95 8.61065 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=3.815 $Y=2.055
+ $X2=3.98 $Y2=2.045
r228 70 71 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=3.815 $Y=2.055
+ $X2=2.76 $Y2=2.055
r229 66 93 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=2.14
+ $X2=2.595 $Y2=2.055
r230 66 68 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.595 $Y=2.14
+ $X2=2.595 $Y2=2.815
r231 65 93 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.97
+ $X2=2.595 $Y2=2.055
r232 64 65 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.595 $Y=1.77
+ $X2=2.595 $Y2=1.97
r233 62 64 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.43 $Y=1.685
+ $X2=2.595 $Y2=1.77
r234 62 63 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.43 $Y=1.685
+ $X2=1.73 $Y2=1.685
r235 58 91 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.645 $Y=2.24
+ $X2=1.645 $Y2=2.095
r236 58 60 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.645 $Y=2.24
+ $X2=1.645 $Y2=2.46
r237 57 91 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.645 $Y=1.95
+ $X2=1.645 $Y2=2.095
r238 56 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=1.77
+ $X2=1.73 $Y2=1.685
r239 56 57 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.645 $Y=1.77
+ $X2=1.645 $Y2=1.95
r240 55 89 3.14085 $w=2.9e-07 $l=1.63e-07 $layer=LI1_cond $X=0.89 $Y=2.095
+ $X2=0.727 $Y2=2.095
r241 54 91 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=2.095
+ $X2=1.645 $Y2=2.095
r242 54 55 26.6254 $w=2.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.56 $Y=2.095
+ $X2=0.89 $Y2=2.095
r243 50 52 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.89 $Y=1.13
+ $X2=1.165 $Y2=1.13
r244 49 89 4.29699 $w=1.7e-07 $l=1.79819e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.727 $Y2=2.095
r245 48 50 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.805 $Y=1.255
+ $X2=0.89 $Y2=1.13
r246 48 49 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.805 $Y=1.255
+ $X2=0.805 $Y2=1.95
r247 44 106 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.63
+ $X2=6.165 $Y2=1.465
r248 44 46 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.165 $Y=1.63
+ $X2=6.165 $Y2=2.4
r249 40 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.3
+ $X2=6.14 $Y2=1.465
r250 40 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.14 $Y=1.3
+ $X2=6.14 $Y2=0.74
r251 36 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.71 $Y=1.3
+ $X2=5.71 $Y2=1.465
r252 36 38 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.71 $Y=1.3
+ $X2=5.71 $Y2=0.74
r253 32 104 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.63
+ $X2=5.715 $Y2=1.465
r254 32 34 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.715 $Y=1.63
+ $X2=5.715 $Y2=2.4
r255 28 101 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.63
+ $X2=5.265 $Y2=1.465
r256 28 30 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.265 $Y=1.63
+ $X2=5.265 $Y2=2.4
r257 24 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.3
+ $X2=5.21 $Y2=1.465
r258 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.21 $Y=1.3
+ $X2=5.21 $Y2=0.74
r259 20 98 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.63
+ $X2=4.765 $Y2=1.465
r260 20 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.765 $Y=1.63
+ $X2=4.765 $Y2=2.4
r261 16 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=1.3
+ $X2=4.75 $Y2=1.465
r262 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.75 $Y=1.3
+ $X2=4.75 $Y2=0.74
r263 5 95 400 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.96 $X2=3.98 $Y2=2.115
r264 5 74 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.96 $X2=3.98 $Y2=2.815
r265 4 93 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.96 $X2=2.595 $Y2=2.105
r266 4 68 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.96 $X2=2.595 $Y2=2.815
r267 3 91 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.96 $X2=1.645 $Y2=2.105
r268 3 60 300 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.96 $X2=1.645 $Y2=2.46
r269 2 89 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.115
r270 1 52 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.595 $X2=1.165 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 40 44 48 50 52
+ 56 58 63 68 73 78 83 92 95 98 101 104 108
r101 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r102 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r105 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r107 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r108 87 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 87 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r111 84 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.655 $Y=3.33
+ $X2=5.53 $Y2=3.33
r112 84 86 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.655 $Y=3.33 $X2=6
+ $Y2=3.33
r113 83 107 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r114 83 86 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r115 82 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r116 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 79 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.48 $Y2=3.33
r119 79 81 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 78 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.53 $Y2=3.33
r121 78 81 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r123 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 74 98 13.8148 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.287 $Y2=3.33
r125 74 76 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 73 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.48 $Y2=3.33
r127 73 76 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.08 $Y2=3.33
r128 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r129 72 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r131 69 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.095 $Y2=3.33
r132 69 71 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 68 98 13.8148 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=3.287 $Y2=3.33
r134 68 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 67 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r136 67 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r137 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r138 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r139 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 63 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=2.095 $Y2=3.33
r141 63 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 62 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r143 62 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 59 89 4.27358 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r146 59 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 58 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r148 58 61 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r149 56 77 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 56 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r151 52 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.44 $Y=1.985
+ $X2=6.44 $Y2=2.815
r152 50 107 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r153 50 55 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.815
r154 46 104 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=3.33
r155 46 48 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.305
r156 42 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r157 42 44 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.455
r158 38 98 2.90666 $w=7.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.287 $Y=3.245
+ $X2=3.287 $Y2=3.33
r159 38 40 12.8808 $w=7.13e-07 $l=7.7e-07 $layer=LI1_cond $X=3.287 $Y=3.245
+ $X2=3.287 $Y2=2.475
r160 34 37 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.095 $Y=2.105
+ $X2=2.095 $Y2=2.815
r161 32 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=3.33
r162 32 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=2.815
r163 28 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r164 28 30 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.495
r165 24 27 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=0.255 $Y=2.115
+ $X2=0.255 $Y2=2.815
r166 22 89 3.08647 $w=2.8e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.197 $Y2=3.33
r167 22 27 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r168 7 55 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.84 $X2=6.44 $Y2=2.815
r169 7 52 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.84 $X2=6.44 $Y2=1.985
r170 6 48 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.84 $X2=5.49 $Y2=2.305
r171 5 44 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=4.295
+ $Y=1.96 $X2=4.48 $Y2=2.455
r172 4 40 150 $w=1.7e-07 $l=7.86416e-07 $layer=licon1_PDIFF $count=4 $X=2.91
+ $Y=1.96 $X2=3.48 $Y2=2.475
r173 3 37 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.96 $X2=2.095 $Y2=2.815
r174 3 34 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.96 $X2=2.095 $Y2=2.105
r175 2 30 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.96 $X2=1.18 $Y2=2.495
r176 1 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r177 1 24 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%X 1 2 3 4 15 19 23 24 25 26 29 32 35 39 41 42
+ 43 44 47
c80 32 0 8.56004e-20 $X=5.98 $Y=1.8
c81 24 0 1.8401e-19 $X=5.08 $Y=1.045
r82 46 47 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=6.48 $Y=1.48
+ $X2=6.48 $Y2=1.295
r83 45 47 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=1.13
+ $X2=6.48 $Y2=1.295
r84 41 46 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.365 $Y=1.565
+ $X2=6.48 $Y2=1.48
r85 41 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.365 $Y=1.565
+ $X2=6.105 $Y2=1.565
r86 40 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.09 $Y=1.045
+ $X2=5.925 $Y2=1.045
r87 39 45 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.365 $Y=1.045
+ $X2=6.48 $Y2=1.13
r88 39 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.365 $Y=1.045
+ $X2=6.09 $Y2=1.045
r89 35 37 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.98 $Y=1.985
+ $X2=5.98 $Y2=2.815
r90 33 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=1.97 $X2=5.98
+ $Y2=1.885
r91 33 35 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=5.98 $Y=1.97
+ $X2=5.98 $Y2=1.985
r92 32 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=1.8 $X2=5.98
+ $Y2=1.885
r93 31 42 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.98 $Y=1.65
+ $X2=6.105 $Y2=1.565
r94 31 32 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.98 $Y=1.65
+ $X2=5.98 $Y2=1.8
r95 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=0.96
+ $X2=5.925 $Y2=1.045
r96 27 29 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.925 $Y=0.96
+ $X2=5.925 $Y2=0.515
r97 25 44 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.855 $Y=1.885
+ $X2=5.98 $Y2=1.885
r98 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.855 $Y=1.885
+ $X2=5.205 $Y2=1.885
r99 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=1.045
+ $X2=5.925 $Y2=1.045
r100 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.76 $Y=1.045
+ $X2=5.08 $Y2=1.045
r101 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.04 $Y=1.985
+ $X2=5.04 $Y2=2.815
r102 17 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.04 $Y=1.97
+ $X2=5.205 $Y2=1.885
r103 17 19 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.04 $Y=1.97
+ $X2=5.04 $Y2=1.985
r104 13 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.955 $Y=0.96
+ $X2=5.08 $Y2=1.045
r105 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.955 $Y=0.96
+ $X2=4.955 $Y2=0.515
r106 4 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.94 $Y2=2.815
r107 4 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.94 $Y2=1.985
r108 3 21 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.84 $X2=5.04 $Y2=2.815
r109 3 19 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.84 $X2=5.04 $Y2=1.985
r110 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.785
+ $Y=0.37 $X2=5.925 $Y2=0.515
r111 1 15 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.37 $X2=4.995 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%A_32_119# 1 2 3 12 14 15 19 20 21
c48 21 0 1.20592e-19 $X=2.11 $Y=1.215
r49 20 23 14.9533 $w=2.29e-07 $l=2.97061e-07 $layer=LI1_cond $X=3.64 $Y=1.215
+ $X2=3.905 $Y2=1.147
r50 20 21 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=3.64 $Y=1.215
+ $X2=2.11 $Y2=1.215
r51 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.025 $Y=1.13
+ $X2=2.11 $Y2=1.215
r52 17 19 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.025 $Y=1.13
+ $X2=2.025 $Y2=0.74
r53 16 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.025 $Y=0.485
+ $X2=2.025 $Y2=0.74
r54 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.94 $Y=0.4
+ $X2=2.025 $Y2=0.485
r55 14 15 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=1.94 $Y=0.4
+ $X2=0.39 $Y2=0.4
r56 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.265 $Y=0.485
+ $X2=0.39 $Y2=0.4
r57 10 12 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.265 $Y=0.485
+ $X2=0.265 $Y2=0.74
r58 3 23 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.595 $X2=3.905 $Y2=1.085
r59 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.885
+ $Y=0.595 $X2=2.025 $Y2=0.74
r60 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%A_119_119# 1 2 11
r10 8 11 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=0.735 $Y=0.745
+ $X2=1.595 $Y2=0.745
r11 2 11 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.455
+ $Y=0.595 $X2=1.595 $Y2=0.745
r12 1 8 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.595 $X2=0.735 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%A_463_119# 1 2 7 10 15
r29 15 16 5.88214 $w=2.8e-07 $l=1.35e-07 $layer=LI1_cond $X=3.47 $Y=0.74
+ $X2=3.47 $Y2=0.875
r30 10 12 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.455 $Y=0.765
+ $X2=2.455 $Y2=0.875
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=0.875
+ $X2=2.455 $Y2=0.875
r32 7 16 3.65648 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.3 $Y=0.875 $X2=3.47
+ $Y2=0.875
r33 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.3 $Y=0.875 $X2=2.62
+ $Y2=0.875
r34 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.335
+ $Y=0.595 $X2=3.475 $Y2=0.74
r35 1 10 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.595 $X2=2.455 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_4%VGND 1 2 3 4 15 19 23 25 27 30 31 32 34 42 51
+ 56 59 63
r74 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r75 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r76 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r77 54 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r78 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r79 51 62 3.99713 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6.49
+ $Y2=0
r80 51 53 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.26 $Y=0 $X2=6
+ $Y2=0
r81 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r82 50 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r83 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r84 47 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.495
+ $Y2=0
r85 47 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=5.04
+ $Y2=0
r86 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r87 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r88 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=2.965
+ $Y2=0
r89 43 45 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=4.08
+ $Y2=0
r90 42 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.495
+ $Y2=0
r91 42 45 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=0 $X2=4.08
+ $Y2=0
r92 41 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r93 40 41 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 37 41 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r95 36 40 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r96 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.965
+ $Y2=0
r98 34 40 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r99 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r100 32 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r101 30 49 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r102 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.425
+ $Y2=0
r103 29 53 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=6
+ $Y2=0
r104 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.425
+ $Y2=0
r105 25 62 3.21509 $w=2.6e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.49 $Y2=0
r106 25 27 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0.515
r107 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0
r108 21 23 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0.625
r109 17 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0
r110 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.495 $Y=0.085
+ $X2=4.495 $Y2=0.515
r111 13 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=2.965 $Y2=0
r112 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.965 $Y=0.085
+ $X2=2.965 $Y2=0.535
r113 4 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.215
+ $Y=0.37 $X2=6.355 $Y2=0.515
r114 3 23 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.37 $X2=5.425 $Y2=0.625
r115 2 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.35
+ $Y=0.37 $X2=4.495 $Y2=0.515
r116 1 15 182 $w=1.7e-07 $l=2.48193e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.595 $X2=2.965 $Y2=0.535
.ends


* File: sky130_fd_sc_ms__a21oi_2.pex.spice
* Created: Wed Sep  2 11:51:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21OI_2%B1 3 5 7 9 10 12 14 15 16 23
r44 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.48 $Y=1.6 $X2=0.555
+ $Y2=1.6
r45 19 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.27 $Y=1.6 $X2=0.48
+ $Y2=1.6
r46 16 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.6 $X2=0.27 $Y2=1.6
r47 12 14 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r48 11 15 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.095 $Y=1.69
+ $X2=1.005 $Y2=1.69
r49 10 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.365 $Y=1.69
+ $X2=1.455 $Y2=1.765
r50 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.365 $Y=1.69
+ $X2=1.095 $Y2=1.69
r51 7 15 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.69
r52 7 9 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r53 5 15 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.915 $Y=1.69 $X2=1.005
+ $Y2=1.69
r54 5 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.915 $Y=1.69
+ $X2=0.555 $Y2=1.69
r55 1 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.435
+ $X2=0.48 $Y2=1.6
r56 1 3 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.48 $Y=1.435
+ $X2=0.48 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%A2 1 3 6 10 14 16 18 29
c55 14 0 6.65152e-20 $X=2.45 $Y=0.74
r56 29 30 5.44194 $w=3.1e-07 $l=3.5e-08 $layer=POLY_cond $X=2.415 $Y=1.515
+ $X2=2.45 $Y2=1.515
r57 27 29 2.33226 $w=3.1e-07 $l=1.5e-08 $layer=POLY_cond $X=2.4 $Y=1.515
+ $X2=2.415 $Y2=1.515
r58 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.515 $X2=2.4 $Y2=1.515
r59 25 27 76.9645 $w=3.1e-07 $l=4.95e-07 $layer=POLY_cond $X=1.905 $Y=1.515
+ $X2=2.4 $Y2=1.515
r60 18 28 4.78431 $w=5.98e-07 $l=2.4e-07 $layer=LI1_cond $X=2.64 $Y=1.48 $X2=2.4
+ $Y2=1.48
r61 16 28 4.78431 $w=5.98e-07 $l=2.4e-07 $layer=LI1_cond $X=2.16 $Y=1.48 $X2=2.4
+ $Y2=1.48
r62 12 30 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.35
+ $X2=2.45 $Y2=1.515
r63 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.45 $Y=1.35
+ $X2=2.45 $Y2=0.74
r64 8 29 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.68
+ $X2=2.415 $Y2=1.515
r65 8 10 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.415 $Y=1.68
+ $X2=2.415 $Y2=2.4
r66 4 25 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=1.515
r67 4 6 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.905 $Y=1.68
+ $X2=1.905 $Y2=2.4
r68 1 25 16.3258 $w=3.1e-07 $l=2.11069e-07 $layer=POLY_cond $X=1.8 $Y=1.35
+ $X2=1.905 $Y2=1.515
r69 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.8 $Y=1.35 $X2=1.8
+ $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%A1 3 7 11 15 17 24 26
c49 15 0 1.44963e-19 $X=3.31 $Y=0.74
r50 25 26 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=3.31 $Y=1.515
+ $X2=3.315 $Y2=1.515
r51 23 25 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.185 $Y=1.515
+ $X2=3.31 $Y2=1.515
r52 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.515 $X2=3.185 $Y2=1.515
r53 21 23 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.88 $Y=1.515
+ $X2=3.185 $Y2=1.515
r54 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=2.88 $Y2=1.515
r55 17 24 5.01062 $w=3.43e-07 $l=1.5e-07 $layer=LI1_cond $X=3.177 $Y=1.665
+ $X2=3.177 $Y2=1.515
r56 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.35
+ $X2=3.31 $Y2=1.515
r57 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.31 $Y=1.35
+ $X2=3.31 $Y2=0.74
r58 9 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.68
+ $X2=3.315 $Y2=1.515
r59 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.315 $Y=1.68
+ $X2=3.315 $Y2=2.4
r60 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.35
+ $X2=2.88 $Y2=1.515
r61 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.88 $Y=1.35 $X2=2.88
+ $Y2=0.74
r62 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.68
+ $X2=2.865 $Y2=1.515
r63 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.865 $Y=1.68
+ $X2=2.865 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%A_131_368# 1 2 3 4 15 19 20 21 22 23 27 34
+ 36
c51 2 0 1.99095e-19 $X=1.545 $Y=1.84
r52 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.375
+ $X2=2.64 $Y2=2.375
r53 27 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=2.375
+ $X2=3.54 $Y2=2.375
r54 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.375 $Y=2.375
+ $X2=2.805 $Y2=2.375
r55 24 32 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.845 $Y=2.375
+ $X2=1.705 $Y2=2.375
r56 23 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=2.375
+ $X2=2.64 $Y2=2.375
r57 23 24 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.475 $Y=2.375
+ $X2=1.845 $Y2=2.375
r58 21 32 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.46
+ $X2=1.705 $Y2=2.375
r59 21 22 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=1.705 $Y=2.46
+ $X2=1.705 $Y2=2.905
r60 19 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=1.705 $Y2=2.905
r61 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=2.99
+ $X2=0.895 $Y2=2.99
r62 15 18 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=0.755 $Y=2.115
+ $X2=0.755 $Y2=2.815
r63 13 20 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.755 $Y=2.905
+ $X2=0.895 $Y2=2.99
r64 13 18 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=0.755 $Y=2.905
+ $X2=0.755 $Y2=2.815
r65 4 36 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.84 $X2=3.54 $Y2=2.455
r66 3 34 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.505
+ $Y=1.84 $X2=2.64 $Y2=2.455
r67 2 32 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.455
r68 1 18 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.84 $X2=0.78 $Y2=2.815
r69 1 15 400 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.84 $X2=0.78 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%Y 1 2 3 12 15 16 18 20 24 25 30 31
c56 25 0 1.44963e-19 $X=3.055 $Y=0.835
r57 31 37 23.4497 $w=2.28e-07 $l=4.68e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=0.732 $Y2=1.665
r58 30 37 0.601275 $w=2.28e-07 $l=1.2e-08 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.732 $Y2=1.665
r59 25 28 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=3.055 $Y=0.835
+ $X2=3.055 $Y2=0.94
r60 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.23 $Y=1.97
+ $X2=1.23 $Y2=2.65
r61 18 31 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=1.23 $Y=1.665 $X2=1.2
+ $Y2=1.665
r62 18 20 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.23 $Y=1.78
+ $X2=1.23 $Y2=1.97
r63 17 24 2.83584 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.86 $Y=0.835
+ $X2=0.732 $Y2=0.835
r64 16 25 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.93 $Y=0.835
+ $X2=3.055 $Y2=0.835
r65 16 17 135.048 $w=1.68e-07 $l=2.07e-06 $layer=LI1_cond $X=2.93 $Y=0.835
+ $X2=0.86 $Y2=0.835
r66 15 37 0.103554 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=0.732 $Y=1.55
+ $X2=0.732 $Y2=1.665
r67 14 24 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=0.92
+ $X2=0.732 $Y2=0.835
r68 14 15 28.4721 $w=2.53e-07 $l=6.3e-07 $layer=LI1_cond $X=0.732 $Y=0.92
+ $X2=0.732 $Y2=1.55
r69 10 24 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=0.75
+ $X2=0.732 $Y2=0.835
r70 10 12 10.6206 $w=2.53e-07 $l=2.35e-07 $layer=LI1_cond $X=0.732 $Y=0.75
+ $X2=0.732 $Y2=0.515
r71 3 22 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.65
r72 3 20 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=1.97
r73 2 28 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.37 $X2=3.095 $Y2=0.94
r74 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.37 $X2=0.695 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 31 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 28 37 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.175 $Y2=3.33
r49 28 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 23 27 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 22 26 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 20 37 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.175 $Y2=3.33
r55 20 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 18 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 16 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=3.09 $Y2=3.33
r60 15 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.09 $Y2=3.33
r62 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=3.33
r63 11 13 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=2.805
r64 7 37 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=3.245
+ $X2=2.175 $Y2=3.33
r65 7 9 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=2.175 $Y=3.245
+ $X2=2.175 $Y2=2.805
r66 2 13 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.84 $X2=3.09 $Y2=2.805
r67 1 9 600 $w=1.7e-07 $l=1.03263e-06 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.84 $X2=2.135 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%VGND 1 2 7 9 13 15 17 30 31 37
r37 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r40 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r41 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r42 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r43 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.165
+ $Y2=0
r45 25 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.64
+ $Y2=0
r46 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r48 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r49 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r50 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 18 34 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r52 18 20 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r53 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.165
+ $Y2=0
r54 17 23 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.68 $Y2=0
r55 15 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r56 15 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r57 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r58 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.495
r59 7 34 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.215 $Y2=0
r60 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.515
r61 2 13 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.535 $X2=2.165 $Y2=0.495
r62 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_2%A_280_107# 1 2 3 10 11 12 13 14 18 19 21 29
c65 11 0 2.6561e-19 $X=1.67 $Y=1.95
r66 21 29 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.605 $Y=1.95
+ $X2=3.605 $Y2=1.13
r67 19 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=0.965
+ $X2=3.525 $Y2=1.13
r68 18 28 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.525 $Y=0.58
+ $X2=3.525 $Y2=0.455
r69 18 19 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.525 $Y=0.58
+ $X2=3.525 $Y2=0.965
r70 14 28 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=0.455
+ $X2=3.525 $Y2=0.455
r71 14 16 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.36 $Y=0.455
+ $X2=2.665 $Y2=0.455
r72 12 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.52 $Y=2.035
+ $X2=3.605 $Y2=1.95
r73 12 13 113.845 $w=1.68e-07 $l=1.745e-06 $layer=LI1_cond $X=3.52 $Y=2.035
+ $X2=1.775 $Y2=2.035
r74 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.67 $Y=1.95
+ $X2=1.775 $Y2=2.035
r75 10 23 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.67 $Y=1.175
+ $X2=1.525 $Y2=1.175
r76 10 11 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.67 $Y=1.26
+ $X2=1.67 $Y2=1.95
r77 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.37 $X2=3.525 $Y2=0.515
r78 2 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.37 $X2=2.665 $Y2=0.495
r79 1 23 182 $w=1.7e-07 $l=6.99714e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.535 $X2=1.525 $Y2=1.175
.ends


* File: sky130_fd_sc_ms__and2b_2.spice
* Created: Wed Sep  2 11:57:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and2b_2.pex.spice"
.subckt sky130_fd_sc_ms__and2b_2  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_N_M1007_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.11874 AS=0.15675 PD=0.989147 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.6 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1007_d N_A_198_48#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15976 AS=0.1036 PD=1.33085 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_198_48#_M1009_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.29785 AS=0.1036 PD=1.545 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1000 A_505_74# N_B_M1000_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.29785 PD=0.98 PS=1.545 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75002 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_198_48#_M1001_d N_A_27_74#_M1001_g A_505_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.18 W=0.84
+ AD=0.203443 AS=0.2352 PD=1.34571 PS=2.24 NRD=43.8916 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1002 N_VPWR_M1003_d N_A_198_48#_M1002_g N_X_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.271257 AS=0.1512 PD=1.79429 PS=1.39 NRD=14.0658 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A_198_48#_M1008_g N_X_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.371264 AS=0.1512 PD=1.87019 PS=1.39 NRD=24.625 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1005 N_A_198_48#_M1005_d N_B_M1005_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.331486 PD=1.27 PS=1.66981 NRD=0 NRS=45.2903 M=1 R=5.55556
+ SA=90002 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_74#_M1006_g N_A_198_48#_M1005_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__and2b_2.pxi.spice"
*
.ends
*
*

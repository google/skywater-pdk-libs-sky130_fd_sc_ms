* File: sky130_fd_sc_ms__xor3_2.pxi.spice
* Created: Fri Aug 28 18:19:48 2020
* 
x_PM_SKY130_FD_SC_MS__XOR3_2%A_83_289# N_A_83_289#_M1000_d N_A_83_289#_M1021_d
+ N_A_83_289#_M1008_d N_A_83_289#_M1013_d N_A_83_289#_M1018_g
+ N_A_83_289#_M1006_g N_A_83_289#_c_196_n N_A_83_289#_c_197_n
+ N_A_83_289#_c_204_n N_A_83_289#_c_261_p N_A_83_289#_c_215_p
+ N_A_83_289#_c_198_n N_A_83_289#_c_206_n N_A_83_289#_c_207_n
+ N_A_83_289#_c_208_n N_A_83_289#_c_209_n N_A_83_289#_c_210_n
+ N_A_83_289#_c_199_n N_A_83_289#_c_200_n PM_SKY130_FD_SC_MS__XOR3_2%A_83_289#
x_PM_SKY130_FD_SC_MS__XOR3_2%A N_A_M1008_g N_A_c_309_n N_A_M1000_g A N_A_c_311_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A
x_PM_SKY130_FD_SC_MS__XOR3_2%A_440_315# N_A_440_315#_M1011_s
+ N_A_440_315#_M1022_s N_A_440_315#_M1001_g N_A_440_315#_M1010_g
+ N_A_440_315#_c_348_n N_A_440_315#_c_349_n N_A_440_315#_M1013_g
+ N_A_440_315#_c_350_n N_A_440_315#_M1021_g N_A_440_315#_c_352_n
+ N_A_440_315#_c_353_n N_A_440_315#_c_354_n N_A_440_315#_c_355_n
+ N_A_440_315#_c_356_n N_A_440_315#_c_357_n N_A_440_315#_c_358_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A_440_315#
x_PM_SKY130_FD_SC_MS__XOR3_2%B N_B_M1023_g N_B_c_467_n N_B_c_468_n N_B_M1020_g
+ N_B_c_453_n N_B_c_454_n N_B_M1003_g N_B_c_470_n N_B_M1017_g N_B_c_456_n
+ N_B_c_457_n N_B_c_458_n N_B_c_459_n N_B_M1022_g N_B_c_461_n N_B_M1011_g
+ N_B_c_473_n N_B_c_462_n B N_B_c_464_n N_B_c_465_n PM_SKY130_FD_SC_MS__XOR3_2%B
x_PM_SKY130_FD_SC_MS__XOR3_2%A_1162_379# N_A_1162_379#_M1019_s
+ N_A_1162_379#_M1016_s N_A_1162_379#_c_586_n N_A_1162_379#_M1015_g
+ N_A_1162_379#_M1005_g N_A_1162_379#_c_587_n N_A_1162_379#_c_588_n
+ N_A_1162_379#_c_589_n N_A_1162_379#_c_590_n N_A_1162_379#_c_591_n
+ N_A_1162_379#_c_592_n N_A_1162_379#_c_581_n N_A_1162_379#_c_582_n
+ N_A_1162_379#_c_583_n N_A_1162_379#_c_584_n N_A_1162_379#_c_585_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A_1162_379#
x_PM_SKY130_FD_SC_MS__XOR3_2%C N_C_M1012_g N_C_c_687_n N_C_M1009_g N_C_c_688_n
+ N_C_c_689_n N_C_c_690_n N_C_M1016_g N_C_c_692_n N_C_c_693_n N_C_c_694_n
+ N_C_M1019_g N_C_c_695_n C PM_SKY130_FD_SC_MS__XOR3_2%C
x_PM_SKY130_FD_SC_MS__XOR3_2%A_1198_424# N_A_1198_424#_M1005_d
+ N_A_1198_424#_M1015_d N_A_1198_424#_M1004_g N_A_1198_424#_M1002_g
+ N_A_1198_424#_c_783_n N_A_1198_424#_M1007_g N_A_1198_424#_M1014_g
+ N_A_1198_424#_c_786_n N_A_1198_424#_c_787_n N_A_1198_424#_c_788_n
+ N_A_1198_424#_c_789_n N_A_1198_424#_c_790_n N_A_1198_424#_c_791_n
+ N_A_1198_424#_c_795_n N_A_1198_424#_c_796_n N_A_1198_424#_c_792_n
+ N_A_1198_424#_c_838_p N_A_1198_424#_c_798_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A_1198_424#
x_PM_SKY130_FD_SC_MS__XOR3_2%A_27_134# N_A_27_134#_M1018_s N_A_27_134#_M1010_d
+ N_A_27_134#_M1006_s N_A_27_134#_M1001_d N_A_27_134#_c_888_n
+ N_A_27_134#_c_889_n N_A_27_134#_c_890_n N_A_27_134#_c_891_n
+ N_A_27_134#_c_892_n N_A_27_134#_c_893_n N_A_27_134#_c_894_n
+ N_A_27_134#_c_895_n N_A_27_134#_c_896_n N_A_27_134#_c_901_n
+ N_A_27_134#_c_897_n N_A_27_134#_c_898_n N_A_27_134#_c_899_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A_27_134#
x_PM_SKY130_FD_SC_MS__XOR3_2%VPWR N_VPWR_M1006_d N_VPWR_M1022_d N_VPWR_M1016_d
+ N_VPWR_M1007_s N_VPWR_c_976_n N_VPWR_c_977_n N_VPWR_c_978_n N_VPWR_c_979_n
+ N_VPWR_c_980_n N_VPWR_c_981_n N_VPWR_c_982_n N_VPWR_c_983_n N_VPWR_c_1027_n
+ VPWR N_VPWR_c_984_n N_VPWR_c_985_n N_VPWR_c_986_n N_VPWR_c_987_n
+ N_VPWR_c_988_n N_VPWR_c_975_n PM_SKY130_FD_SC_MS__XOR3_2%VPWR
x_PM_SKY130_FD_SC_MS__XOR3_2%A_375_419# N_A_375_419#_M1017_d
+ N_A_375_419#_M1005_s N_A_375_419#_M1023_d N_A_375_419#_M1012_d
+ N_A_375_419#_c_1084_n N_A_375_419#_c_1085_n N_A_375_419#_c_1097_n
+ N_A_375_419#_c_1074_n N_A_375_419#_c_1075_n N_A_375_419#_c_1076_n
+ N_A_375_419#_c_1122_n N_A_375_419#_c_1077_n N_A_375_419#_c_1126_n
+ N_A_375_419#_c_1078_n N_A_375_419#_c_1079_n N_A_375_419#_c_1080_n
+ N_A_375_419#_c_1087_n N_A_375_419#_c_1088_n N_A_375_419#_c_1089_n
+ N_A_375_419#_c_1081_n N_A_375_419#_c_1082_n N_A_375_419#_c_1083_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A_375_419#
x_PM_SKY130_FD_SC_MS__XOR3_2%A_416_113# N_A_416_113#_M1020_d
+ N_A_416_113#_M1009_d N_A_416_113#_M1003_d N_A_416_113#_M1015_s
+ N_A_416_113#_c_1219_n N_A_416_113#_c_1220_n N_A_416_113#_c_1221_n
+ N_A_416_113#_c_1228_n N_A_416_113#_c_1229_n N_A_416_113#_c_1222_n
+ N_A_416_113#_c_1223_n N_A_416_113#_c_1278_n N_A_416_113#_c_1279_n
+ N_A_416_113#_c_1224_n N_A_416_113#_c_1225_n N_A_416_113#_c_1230_n
+ N_A_416_113#_c_1247_n N_A_416_113#_c_1231_n N_A_416_113#_c_1232_n
+ N_A_416_113#_c_1233_n N_A_416_113#_c_1226_n N_A_416_113#_c_1227_n
+ PM_SKY130_FD_SC_MS__XOR3_2%A_416_113#
x_PM_SKY130_FD_SC_MS__XOR3_2%X N_X_M1002_s N_X_M1004_d X X X X X X X
+ PM_SKY130_FD_SC_MS__XOR3_2%X
x_PM_SKY130_FD_SC_MS__XOR3_2%VGND N_VGND_M1018_d N_VGND_M1011_d N_VGND_M1019_d
+ N_VGND_M1014_d N_VGND_c_1364_n N_VGND_c_1365_n N_VGND_c_1366_n N_VGND_c_1367_n
+ VGND N_VGND_c_1368_n N_VGND_c_1369_n N_VGND_c_1370_n N_VGND_c_1371_n
+ N_VGND_c_1372_n N_VGND_c_1373_n N_VGND_c_1374_n N_VGND_c_1375_n
+ PM_SKY130_FD_SC_MS__XOR3_2%VGND
cc_1 VNB N_A_83_289#_M1018_g 0.025899f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_2 VNB N_A_83_289#_c_196_n 0.00288335f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_3 VNB N_A_83_289#_c_197_n 0.0213525f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_4 VNB N_A_83_289#_c_198_n 0.00787075f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_5 VNB N_A_83_289#_c_199_n 0.00297214f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.905
cc_6 VNB N_A_83_289#_c_200_n 8.48484e-19 $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.1
cc_7 VNB N_A_c_309_n 0.0210019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A 0.00137659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_311_n 0.0296322f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_10 VNB N_A_440_315#_M1010_g 0.0365935f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.445
cc_11 VNB N_A_440_315#_c_348_n 0.0212212f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_12 VNB N_A_440_315#_c_349_n 0.0123703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_440_315#_c_350_n 0.0108329f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.92
cc_14 VNB N_A_440_315#_M1021_g 0.0193825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_440_315#_c_352_n 0.00897801f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.24
cc_16 VNB N_A_440_315#_c_353_n 0.00122356f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_17 VNB N_A_440_315#_c_354_n 0.00935992f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_18 VNB N_A_440_315#_c_355_n 3.26207e-19 $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_19 VNB N_A_440_315#_c_356_n 0.0065592f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=2.99
cc_20 VNB N_A_440_315#_c_357_n 0.00140635f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.07
cc_21 VNB N_A_440_315#_c_358_n 0.024011f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.905
cc_22 VNB N_B_M1020_g 0.0412954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_453_n 0.0694559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_454_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_M1017_g 0.0335493f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.92
cc_26 VNB N_B_c_456_n 0.089017f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_27 VNB N_B_c_457_n 0.0180259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_458_n 0.00660556f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_29 VNB N_B_c_459_n 0.0579081f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.09
cc_30 VNB N_B_M1022_g 0.00745313f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_31 VNB N_B_c_461_n 0.0199242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_c_462_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_33 VNB B 0.0062914f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.905
cc_34 VNB N_B_c_464_n 0.0190806f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.07
cc_35 VNB N_B_c_465_n 0.0429467f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_36 VNB N_A_1162_379#_M1005_g 0.0259339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1162_379#_c_581_n 4.38491e-19 $X=-0.19 $Y=-0.245 $X2=0.745
+ $Y2=2.005
cc_38 VNB N_A_1162_379#_c_582_n 0.00454486f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.09
cc_39 VNB N_A_1162_379#_c_583_n 0.00752181f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.24
cc_40 VNB N_A_1162_379#_c_584_n 0.00213207f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.165
cc_41 VNB N_A_1162_379#_c_585_n 0.034674f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_42 VNB N_C_c_687_n 0.0206136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_C_c_688_n 0.0352899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_C_c_689_n 0.0359645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_C_c_690_n 0.0206211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_C_M1016_g 0.00397265f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_47 VNB N_C_c_692_n 0.027196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_C_c_693_n 0.011937f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.775
cc_49 VNB N_C_c_694_n 0.0174959f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.435
cc_50 VNB N_C_c_695_n 0.0105498f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.92
cc_51 VNB C 7.99339e-19 $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.61
cc_52 VNB N_A_1198_424#_M1004_g 5.55144e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1198_424#_M1002_g 0.0221192f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.445
cc_54 VNB N_A_1198_424#_c_783_n 0.00970685f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.99
cc_55 VNB N_A_1198_424#_M1007_g 0.0151082f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=2.435
cc_56 VNB N_A_1198_424#_M1014_g 0.0248256f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_57 VNB N_A_1198_424#_c_786_n 0.0413116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1198_424#_c_787_n 0.0100011f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=2.005
cc_59 VNB N_A_1198_424#_c_788_n 0.012538f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.005
cc_60 VNB N_A_1198_424#_c_789_n 0.00243198f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.24
cc_61 VNB N_A_1198_424#_c_790_n 0.00555163f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.165
cc_62 VNB N_A_1198_424#_c_791_n 0.00493017f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=2.99
cc_63 VNB N_A_1198_424#_c_792_n 0.0010115f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.905
cc_64 VNB N_A_27_134#_c_888_n 0.0122262f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.445
cc_65 VNB N_A_27_134#_c_889_n 0.0103833f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_66 VNB N_A_27_134#_c_890_n 0.00553396f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.775
cc_67 VNB N_A_27_134#_c_891_n 0.00184736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_134#_c_892_n 0.011717f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.92
cc_69 VNB N_A_27_134#_c_893_n 0.0038752f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.61
cc_70 VNB N_A_27_134#_c_894_n 4.4909e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_134#_c_895_n 0.00200956f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.09
cc_72 VNB N_A_27_134#_c_896_n 0.00710642f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.24
cc_73 VNB N_A_27_134#_c_897_n 0.0180441f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_74 VNB N_A_27_134#_c_898_n 0.0054336f $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=2.99
cc_75 VNB N_A_27_134#_c_899_n 0.00346141f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.265
cc_76 VNB N_VPWR_c_975_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_375_419#_c_1074_n 0.00979392f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.61
cc_78 VNB N_A_375_419#_c_1075_n 0.021596f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_79 VNB N_A_375_419#_c_1076_n 0.00289389f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_80 VNB N_A_375_419#_c_1077_n 0.00673931f $X=-0.19 $Y=-0.245 $X2=0.745
+ $Y2=2.005
cc_81 VNB N_A_375_419#_c_1078_n 0.00540474f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=2.24
cc_82 VNB N_A_375_419#_c_1079_n 0.0332271f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.24
cc_83 VNB N_A_375_419#_c_1080_n 0.00432252f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_84 VNB N_A_375_419#_c_1081_n 0.00361673f $X=-0.19 $Y=-0.245 $X2=4.31
+ $Y2=1.265
cc_85 VNB N_A_375_419#_c_1082_n 0.0166275f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.92
cc_86 VNB N_A_375_419#_c_1083_n 0.00844405f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_87 VNB N_A_416_113#_c_1219_n 0.00163083f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.99
cc_88 VNB N_A_416_113#_c_1220_n 0.0128498f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=1.775
cc_89 VNB N_A_416_113#_c_1221_n 0.00351336f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=2.435
cc_90 VNB N_A_416_113#_c_1222_n 0.0141251f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.24
cc_91 VNB N_A_416_113#_c_1223_n 0.00344537f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_92 VNB N_A_416_113#_c_1224_n 0.00643748f $X=-0.19 $Y=-0.245 $X2=3.81
+ $Y2=2.755
cc_93 VNB N_A_416_113#_c_1225_n 0.00230384f $X=-0.19 $Y=-0.245 $X2=3.81
+ $Y2=2.905
cc_94 VNB N_A_416_113#_c_1226_n 0.00505131f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_95 VNB N_A_416_113#_c_1227_n 0.0107302f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.775
cc_96 VNB X 0.00248472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1364_n 0.00766793f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_98 VNB N_VGND_c_1365_n 0.0157044f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.435
cc_99 VNB N_VGND_c_1366_n 0.011316f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.61
cc_100 VNB N_VGND_c_1367_n 0.0467556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1368_n 0.102977f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_102 VNB N_VGND_c_1369_n 0.0640359f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.92
cc_103 VNB N_VGND_c_1370_n 0.0191116f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_104 VNB N_VGND_c_1371_n 0.0197198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1372_n 0.037346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1373_n 0.00477918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1374_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1375_n 0.506431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VPB N_A_83_289#_M1006_g 0.0272886f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_110 VPB N_A_83_289#_c_196_n 0.00133739f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_111 VPB N_A_83_289#_c_197_n 0.013212f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_112 VPB N_A_83_289#_c_204_n 0.00844789f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=2.005
cc_113 VPB N_A_83_289#_c_198_n 0.00680237f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_114 VPB N_A_83_289#_c_206_n 0.0347134f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_115 VPB N_A_83_289#_c_207_n 0.00250443f $X=-0.19 $Y=1.66 $X2=1.64 $Y2=2.99
cc_116 VPB N_A_83_289#_c_208_n 0.00521917f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.905
cc_117 VPB N_A_83_289#_c_209_n 0.00564279f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.92
cc_118 VPB N_A_83_289#_c_210_n 0.0104086f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.07
cc_119 VPB N_A_83_289#_c_199_n 0.00329913f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.905
cc_120 VPB N_A_M1008_g 0.024288f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.935
cc_121 VPB A 0.00190989f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_c_311_n 0.0152984f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_123 VPB N_A_440_315#_M1001_g 0.0361358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_440_315#_c_348_n 0.0166673f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_125 VPB N_A_440_315#_c_349_n 0.0080272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_440_315#_M1013_g 0.0232978f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_127 VPB N_A_440_315#_c_350_n 0.0127697f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.92
cc_128 VPB N_A_440_315#_c_352_n 0.00124171f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.24
cc_129 VPB N_A_440_315#_c_356_n 0.00562608f $X=-0.19 $Y=1.66 $X2=1.64 $Y2=2.99
cc_130 VPB N_A_440_315#_c_357_n 4.64599e-19 $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.07
cc_131 VPB N_A_440_315#_c_358_n 0.0135441f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.905
cc_132 VPB N_B_M1023_g 0.0247735f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.935
cc_133 VPB N_B_c_467_n 0.0501476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_B_c_468_n 0.0141058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_B_M1003_g 0.0353391f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_136 VPB N_B_c_470_n 0.113778f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.775
cc_137 VPB N_B_c_458_n 0.0886941f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=2.005
cc_138 VPB N_B_M1022_g 0.0269886f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_139 VPB N_B_c_473_n 0.00898883f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.755
cc_140 VPB N_A_1162_379#_c_586_n 0.0216259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1162_379#_c_587_n 0.00869713f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_142 VPB N_A_1162_379#_c_588_n 0.0278891f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_143 VPB N_A_1162_379#_c_589_n 0.00327346f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.92
cc_144 VPB N_A_1162_379#_c_590_n 0.0223653f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.61
cc_145 VPB N_A_1162_379#_c_591_n 0.00304973f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_146 VPB N_A_1162_379#_c_592_n 0.0126724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1162_379#_c_581_n 0.00884912f $X=-0.19 $Y=1.66 $X2=0.745
+ $Y2=2.005
cc_148 VPB N_A_1162_379#_c_584_n 0.00170428f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_149 VPB N_A_1162_379#_c_585_n 0.0044609f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_150 VPB N_C_M1012_g 0.0433896f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.935
cc_151 VPB N_C_c_689_n 0.0137087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_C_M1016_g 0.0299316f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_153 VPB C 0.00197916f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.61
cc_154 VPB N_A_1198_424#_M1004_g 0.0246517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_1198_424#_M1007_g 0.0274207f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_156 VPB N_A_1198_424#_c_795_n 0.010092f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.905
cc_157 VPB N_A_1198_424#_c_796_n 0.00211174f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.92
cc_158 VPB N_A_1198_424#_c_792_n 0.00275279f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.905
cc_159 VPB N_A_1198_424#_c_798_n 0.00298453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_27_134#_c_894_n 0.00207959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_27_134#_c_901_n 0.0380117f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_162 VPB N_A_27_134#_c_897_n 0.028539f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_163 VPB N_VPWR_c_976_n 0.0107599f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_164 VPB N_VPWR_c_977_n 0.00805719f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.435
cc_165 VPB N_VPWR_c_978_n 0.00566306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_979_n 0.013253f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.09
cc_167 VPB N_VPWR_c_980_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.905
cc_168 VPB N_VPWR_c_981_n 0.0592247f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.24
cc_169 VPB N_VPWR_c_982_n 0.0227085f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_170 VPB N_VPWR_c_983_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.64 $Y2=2.99
cc_171 VPB N_VPWR_c_984_n 0.0940373f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=1.1
cc_172 VPB N_VPWR_c_985_n 0.0711732f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.775
cc_173 VPB N_VPWR_c_986_n 0.0198086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_987_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_988_n 0.0106494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_975_n 0.108563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_375_419#_c_1084_n 0.0047726f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_178 VPB N_A_375_419#_c_1085_n 7.88827e-19 $X=-0.19 $Y=1.66 $X2=0.655
+ $Y2=1.775
cc_179 VPB N_A_375_419#_c_1074_n 0.00371464f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.61
cc_180 VPB N_A_375_419#_c_1087_n 0.00791988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_375_419#_c_1088_n 0.00674591f $X=-0.19 $Y=1.66 $X2=1.64 $Y2=2.99
cc_182 VPB N_A_375_419#_c_1089_n 0.00450367f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.755
cc_183 VPB N_A_375_419#_c_1081_n 0.00441721f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.265
cc_184 VPB N_A_416_113#_c_1228_n 3.66705e-19 $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.92
cc_185 VPB N_A_416_113#_c_1229_n 0.0136231f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.005
cc_186 VPB N_A_416_113#_c_1230_n 0.011909f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.905
cc_187 VPB N_A_416_113#_c_1231_n 0.00298204f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.905
cc_188 VPB N_A_416_113#_c_1232_n 0.00684386f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=1.1
cc_189 VPB N_A_416_113#_c_1233_n 0.00925538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_416_113#_c_1226_n 0.00151514f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.61
cc_191 VPB N_A_416_113#_c_1227_n 0.00698548f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.775
cc_192 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 N_A_83_289#_c_196_n N_A_M1008_g 9.79754e-19 $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_194 N_A_83_289#_c_197_n N_A_M1008_g 0.0239165f $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_195 N_A_83_289#_c_204_n N_A_M1008_g 0.0143872f $X=1.31 $Y=2.005 $X2=0 $Y2=0
cc_196 N_A_83_289#_c_215_p N_A_M1008_g 0.0135769f $X=1.475 $Y=2.24 $X2=0 $Y2=0
cc_197 N_A_83_289#_c_198_n N_A_M1008_g 0.00627066f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_198 N_A_83_289#_c_207_n N_A_M1008_g 0.00425757f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_199 N_A_83_289#_c_209_n N_A_M1008_g 0.00387221f $X=1.31 $Y=1.92 $X2=0 $Y2=0
cc_200 N_A_83_289#_M1018_g N_A_c_309_n 0.0147663f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_201 N_A_83_289#_c_198_n N_A_c_309_n 0.0111091f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_202 N_A_83_289#_M1018_g A 0.00405976f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_203 N_A_83_289#_c_196_n A 0.0192835f $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_204 N_A_83_289#_c_197_n A 0.00106229f $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_205 N_A_83_289#_c_204_n A 0.0253825f $X=1.31 $Y=2.005 $X2=0 $Y2=0
cc_206 N_A_83_289#_c_198_n A 0.0378672f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_207 N_A_83_289#_M1018_g N_A_c_311_n 8.70324e-19 $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_208 N_A_83_289#_c_196_n N_A_c_311_n 0.00112373f $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_209 N_A_83_289#_c_197_n N_A_c_311_n 0.0190167f $X=0.58 $Y=1.61 $X2=0 $Y2=0
cc_210 N_A_83_289#_c_204_n N_A_c_311_n 0.00143809f $X=1.31 $Y=2.005 $X2=0 $Y2=0
cc_211 N_A_83_289#_c_209_n N_A_c_311_n 0.00290313f $X=1.31 $Y=1.92 $X2=0 $Y2=0
cc_212 N_A_83_289#_c_206_n N_A_440_315#_M1001_g 0.00138057f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_213 N_A_83_289#_c_209_n N_A_440_315#_M1001_g 0.00144782f $X=1.31 $Y=1.92
+ $X2=0 $Y2=0
cc_214 N_A_83_289#_c_198_n N_A_440_315#_c_349_n 0.00853359f $X=1.54 $Y=1.165
+ $X2=0 $Y2=0
cc_215 N_A_83_289#_c_206_n N_A_440_315#_M1013_g 0.00138057f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_216 N_A_83_289#_c_210_n N_A_440_315#_M1013_g 0.00595695f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_217 N_A_83_289#_c_199_n N_A_440_315#_M1021_g 4.86955e-19 $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_218 N_A_83_289#_c_200_n N_A_440_315#_M1021_g 0.00119421f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_219 N_A_83_289#_c_199_n N_A_440_315#_c_353_n 0.00794453f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_220 N_A_83_289#_M1021_d N_A_440_315#_c_354_n 0.0066978f $X=3.84 $Y=0.625
+ $X2=0 $Y2=0
cc_221 N_A_83_289#_c_200_n N_A_440_315#_c_354_n 0.0483684f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_222 N_A_83_289#_c_199_n N_A_440_315#_c_356_n 0.102962f $X=4.06 $Y=1.905 $X2=0
+ $Y2=0
cc_223 N_A_83_289#_c_210_n N_A_440_315#_c_357_n 0.0250643f $X=3.81 $Y=2.07 $X2=0
+ $Y2=0
cc_224 N_A_83_289#_c_199_n N_A_440_315#_c_357_n 0.0225071f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_225 N_A_83_289#_c_210_n N_A_440_315#_c_358_n 0.00811391f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_226 N_A_83_289#_c_199_n N_A_440_315#_c_358_n 0.00113401f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_227 N_A_83_289#_c_215_p N_B_M1023_g 0.00440392f $X=1.475 $Y=2.24 $X2=0 $Y2=0
cc_228 N_A_83_289#_c_206_n N_B_M1023_g 0.0180969f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_229 N_A_83_289#_c_209_n N_B_M1023_g 0.00369495f $X=1.31 $Y=1.92 $X2=0 $Y2=0
cc_230 N_A_83_289#_c_206_n N_B_c_467_n 0.010967f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_231 N_A_83_289#_c_198_n N_B_M1020_g 9.19484e-19 $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_232 N_A_83_289#_c_206_n N_B_M1003_g 0.0149959f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_233 N_A_83_289#_c_206_n N_B_c_470_n 0.0200985f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_234 N_A_83_289#_c_210_n N_B_c_470_n 0.00629714f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_235 N_A_83_289#_c_199_n N_B_c_457_n 0.0075973f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_236 N_A_83_289#_c_200_n N_B_c_457_n 0.00195237f $X=4.31 $Y=1.1 $X2=0 $Y2=0
cc_237 N_A_83_289#_c_206_n N_B_c_458_n 0.00546456f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_238 N_A_83_289#_c_208_n N_B_c_458_n 0.00399845f $X=3.81 $Y=2.905 $X2=0 $Y2=0
cc_239 N_A_83_289#_c_210_n N_B_c_458_n 0.0344368f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_240 N_A_83_289#_c_199_n N_B_c_458_n 0.00950883f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_241 N_A_83_289#_c_200_n N_B_c_459_n 0.00788621f $X=4.31 $Y=1.1 $X2=0 $Y2=0
cc_242 N_A_83_289#_c_261_p N_A_27_134#_M1006_s 0.00262546f $X=0.745 $Y=2.005
+ $X2=0 $Y2=0
cc_243 N_A_83_289#_M1018_g N_A_27_134#_c_888_n 0.00162247f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_244 N_A_83_289#_M1018_g N_A_27_134#_c_889_n 0.0115093f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_245 N_A_83_289#_M1000_d N_A_27_134#_c_890_n 0.0132999f $X=1.4 $Y=0.67 $X2=0
+ $Y2=0
cc_246 N_A_83_289#_M1018_g N_A_27_134#_c_890_n 0.0109735f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_247 N_A_83_289#_c_196_n N_A_27_134#_c_890_n 0.00736351f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_248 N_A_83_289#_c_197_n N_A_27_134#_c_890_n 6.87726e-19 $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_249 N_A_83_289#_c_198_n N_A_27_134#_c_890_n 0.0135869f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_250 N_A_83_289#_M1000_d N_A_27_134#_c_891_n 0.00424046f $X=1.4 $Y=0.67 $X2=0
+ $Y2=0
cc_251 N_A_83_289#_c_198_n N_A_27_134#_c_891_n 0.0290186f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_252 N_A_83_289#_c_198_n N_A_27_134#_c_893_n 0.0143578f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_253 N_A_83_289#_M1018_g N_A_27_134#_c_896_n 0.00602985f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_254 N_A_83_289#_c_196_n N_A_27_134#_c_896_n 0.0015079f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_255 N_A_83_289#_M1006_g N_A_27_134#_c_901_n 0.00906091f $X=0.655 $Y=2.435
+ $X2=0 $Y2=0
cc_256 N_A_83_289#_c_197_n N_A_27_134#_c_901_n 8.08053e-19 $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_257 N_A_83_289#_c_261_p N_A_27_134#_c_901_n 0.00987335f $X=0.745 $Y=2.005
+ $X2=0 $Y2=0
cc_258 N_A_83_289#_M1018_g N_A_27_134#_c_897_n 0.00411368f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_259 N_A_83_289#_M1006_g N_A_27_134#_c_897_n 0.00520723f $X=0.655 $Y=2.435
+ $X2=0 $Y2=0
cc_260 N_A_83_289#_c_196_n N_A_27_134#_c_897_n 0.0361693f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_261 N_A_83_289#_c_197_n N_A_27_134#_c_897_n 0.00748597f $X=0.58 $Y=1.61 $X2=0
+ $Y2=0
cc_262 N_A_83_289#_c_261_p N_A_27_134#_c_897_n 0.0140829f $X=0.745 $Y=2.005
+ $X2=0 $Y2=0
cc_263 N_A_83_289#_c_204_n N_VPWR_M1006_d 0.00391623f $X=1.31 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_264 N_A_83_289#_M1006_g N_VPWR_c_976_n 0.00354172f $X=0.655 $Y=2.435 $X2=0
+ $Y2=0
cc_265 N_A_83_289#_c_204_n N_VPWR_c_976_n 0.0237567f $X=1.31 $Y=2.005 $X2=0
+ $Y2=0
cc_266 N_A_83_289#_c_215_p N_VPWR_c_976_n 0.0417667f $X=1.475 $Y=2.24 $X2=0
+ $Y2=0
cc_267 N_A_83_289#_c_207_n N_VPWR_c_976_n 0.0119461f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_268 N_A_83_289#_M1006_g N_VPWR_c_982_n 0.00640648f $X=0.655 $Y=2.435 $X2=0
+ $Y2=0
cc_269 N_A_83_289#_c_206_n N_VPWR_c_984_n 0.144765f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_270 N_A_83_289#_c_207_n N_VPWR_c_984_n 0.0236566f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_271 N_A_83_289#_c_210_n N_VPWR_c_984_n 0.0112583f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_272 N_A_83_289#_M1006_g N_VPWR_c_975_n 0.00645424f $X=0.655 $Y=2.435 $X2=0
+ $Y2=0
cc_273 N_A_83_289#_c_206_n N_VPWR_c_975_n 0.0758332f $X=3.725 $Y=2.99 $X2=0
+ $Y2=0
cc_274 N_A_83_289#_c_207_n N_VPWR_c_975_n 0.0128296f $X=1.64 $Y=2.99 $X2=0 $Y2=0
cc_275 N_A_83_289#_c_210_n N_VPWR_c_975_n 0.01371f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_276 N_A_83_289#_c_206_n N_A_375_419#_M1023_d 0.00213299f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_277 N_A_83_289#_c_215_p N_A_375_419#_c_1084_n 0.0151273f $X=1.475 $Y=2.24
+ $X2=0 $Y2=0
cc_278 N_A_83_289#_c_209_n N_A_375_419#_c_1084_n 0.00107941f $X=1.31 $Y=1.92
+ $X2=0 $Y2=0
cc_279 N_A_83_289#_M1013_d N_A_375_419#_c_1085_n 0.00315924f $X=3.365 $Y=1.895
+ $X2=0 $Y2=0
cc_280 N_A_83_289#_c_206_n N_A_375_419#_c_1085_n 0.0852097f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_281 N_A_83_289#_c_210_n N_A_375_419#_c_1085_n 0.0152397f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_282 N_A_83_289#_c_206_n N_A_375_419#_c_1097_n 0.0191859f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_283 N_A_83_289#_M1013_d N_A_375_419#_c_1074_n 0.0100038f $X=3.365 $Y=1.895
+ $X2=0 $Y2=0
cc_284 N_A_83_289#_c_210_n N_A_375_419#_c_1074_n 0.0514618f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_285 N_A_83_289#_c_199_n N_A_375_419#_c_1074_n 0.00493854f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_286 N_A_83_289#_M1013_d N_A_416_113#_c_1230_n 0.00983478f $X=3.365 $Y=1.895
+ $X2=0 $Y2=0
cc_287 N_A_83_289#_c_210_n N_A_416_113#_c_1230_n 0.0691818f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_288 N_A_83_289#_M1018_g N_VGND_c_1371_n 0.00305419f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_289 N_A_83_289#_M1018_g N_VGND_c_1375_n 0.00457172f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_290 N_A_M1008_g N_B_M1023_g 0.0206361f $X=1.25 $Y=2.435 $X2=0 $Y2=0
cc_291 N_A_c_309_n N_B_M1020_g 0.0120059f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_292 N_A_c_309_n N_A_27_134#_c_890_n 0.0172797f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_293 A N_A_27_134#_c_890_n 0.01258f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_294 N_A_c_311_n N_A_27_134#_c_890_n 0.00104475f $X=1.325 $Y=1.585 $X2=0 $Y2=0
cc_295 N_A_c_309_n N_A_27_134#_c_891_n 0.00341356f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_296 A N_A_27_134#_c_896_n 0.0031593f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_297 N_A_M1008_g N_VPWR_c_976_n 0.00800247f $X=1.25 $Y=2.435 $X2=0 $Y2=0
cc_298 N_A_M1008_g N_VPWR_c_984_n 0.00578564f $X=1.25 $Y=2.435 $X2=0 $Y2=0
cc_299 N_A_M1008_g N_VPWR_c_975_n 0.00537853f $X=1.25 $Y=2.435 $X2=0 $Y2=0
cc_300 A N_VGND_M1018_d 0.00601105f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_301 N_A_c_309_n N_VGND_c_1368_n 0.00305517f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_302 N_A_c_309_n N_VGND_c_1375_n 0.00457172f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_303 N_A_440_315#_M1001_g N_B_M1023_g 0.00905957f $X=2.29 $Y=2.415 $X2=0 $Y2=0
cc_304 N_A_440_315#_M1001_g N_B_c_467_n 0.0105864f $X=2.29 $Y=2.415 $X2=0 $Y2=0
cc_305 N_A_440_315#_M1010_g N_B_M1020_g 0.0109333f $X=2.505 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_440_315#_M1010_g N_B_c_453_n 0.00355453f $X=2.505 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_440_315#_M1001_g N_B_M1003_g 0.0258878f $X=2.29 $Y=2.415 $X2=0 $Y2=0
cc_308 N_A_440_315#_c_348_n N_B_M1003_g 0.0116044f $X=3.185 $Y=1.65 $X2=0 $Y2=0
cc_309 N_A_440_315#_M1013_g N_B_M1003_g 0.0239677f $X=3.275 $Y=2.315 $X2=0 $Y2=0
cc_310 N_A_440_315#_M1013_g N_B_c_470_n 0.0105864f $X=3.275 $Y=2.315 $X2=0 $Y2=0
cc_311 N_A_440_315#_M1010_g N_B_M1017_g 0.0121494f $X=2.505 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_440_315#_c_348_n N_B_M1017_g 0.00890903f $X=3.185 $Y=1.65 $X2=0 $Y2=0
cc_313 N_A_440_315#_M1021_g N_B_M1017_g 0.0152172f $X=3.765 $Y=0.945 $X2=0 $Y2=0
cc_314 N_A_440_315#_M1021_g N_B_c_456_n 0.00737859f $X=3.765 $Y=0.945 $X2=0
+ $Y2=0
cc_315 N_A_440_315#_M1021_g N_B_c_457_n 7.80508e-19 $X=3.765 $Y=0.945 $X2=0
+ $Y2=0
cc_316 N_A_440_315#_c_353_n N_B_c_457_n 4.54349e-19 $X=3.81 $Y=1.435 $X2=0 $Y2=0
cc_317 N_A_440_315#_c_356_n N_B_c_457_n 0.00112154f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_440_315#_c_357_n N_B_c_457_n 3.32909e-19 $X=3.89 $Y=1.57 $X2=0 $Y2=0
cc_319 N_A_440_315#_c_358_n N_B_c_457_n 0.0180459f $X=3.89 $Y=1.57 $X2=0 $Y2=0
cc_320 N_A_440_315#_c_356_n N_B_c_458_n 0.0134394f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A_440_315#_M1021_g N_B_c_459_n 0.0167537f $X=3.765 $Y=0.945 $X2=0 $Y2=0
cc_322 N_A_440_315#_c_354_n N_B_c_459_n 0.0210838f $X=4.58 $Y=0.68 $X2=0 $Y2=0
cc_323 N_A_440_315#_c_356_n N_B_c_461_n 0.00418241f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_440_315#_c_356_n B 0.0272067f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A_440_315#_c_354_n N_B_c_464_n 7.32755e-19 $X=4.58 $Y=0.68 $X2=0 $Y2=0
cc_326 N_A_440_315#_c_356_n N_B_c_464_n 0.0141116f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A_440_315#_c_356_n N_B_c_465_n 0.0091612f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_440_315#_M1010_g N_A_27_134#_c_891_n 0.00139233f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_329 N_A_440_315#_c_349_n N_A_27_134#_c_892_n 0.00739683f $X=2.58 $Y=1.65
+ $X2=0 $Y2=0
cc_330 N_A_440_315#_M1001_g N_A_27_134#_c_894_n 0.023046f $X=2.29 $Y=2.415 $X2=0
+ $Y2=0
cc_331 N_A_440_315#_M1010_g N_A_27_134#_c_894_n 3.68706e-19 $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_332 N_A_440_315#_c_348_n N_A_27_134#_c_894_n 0.0067172f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_333 N_A_440_315#_c_349_n N_A_27_134#_c_894_n 0.013482f $X=2.58 $Y=1.65 $X2=0
+ $Y2=0
cc_334 N_A_440_315#_M1013_g N_A_27_134#_c_894_n 0.00120588f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_335 N_A_440_315#_M1010_g N_A_27_134#_c_895_n 0.00622153f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_336 N_A_440_315#_M1010_g N_A_27_134#_c_898_n 0.0133067f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_337 N_A_440_315#_M1010_g N_A_27_134#_c_899_n 0.0140064f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_338 N_A_440_315#_c_348_n N_A_27_134#_c_899_n 0.00629061f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_339 N_A_440_315#_c_356_n N_VPWR_c_977_n 0.0393878f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_440_315#_c_356_n N_VPWR_c_984_n 0.00749631f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_440_315#_c_356_n N_VPWR_c_975_n 0.0062048f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_440_315#_M1001_g N_A_375_419#_c_1085_n 0.0131663f $X=2.29 $Y=2.415
+ $X2=0 $Y2=0
cc_343 N_A_440_315#_M1013_g N_A_375_419#_c_1085_n 0.0132347f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_344 N_A_440_315#_M1013_g N_A_375_419#_c_1074_n 0.017567f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_345 N_A_440_315#_c_350_n N_A_375_419#_c_1074_n 0.0145675f $X=3.69 $Y=1.65
+ $X2=0 $Y2=0
cc_346 N_A_440_315#_M1021_g N_A_375_419#_c_1074_n 0.013414f $X=3.765 $Y=0.945
+ $X2=0 $Y2=0
cc_347 N_A_440_315#_c_353_n N_A_375_419#_c_1074_n 0.0471932f $X=3.81 $Y=1.435
+ $X2=0 $Y2=0
cc_348 N_A_440_315#_c_355_n N_A_375_419#_c_1074_n 0.0133618f $X=3.895 $Y=0.68
+ $X2=0 $Y2=0
cc_349 N_A_440_315#_c_357_n N_A_375_419#_c_1074_n 0.0219455f $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_350 N_A_440_315#_M1011_s N_A_375_419#_c_1075_n 0.00231738f $X=4.585 $Y=0.37
+ $X2=0 $Y2=0
cc_351 N_A_440_315#_M1021_g N_A_375_419#_c_1075_n 0.00174767f $X=3.765 $Y=0.945
+ $X2=0 $Y2=0
cc_352 N_A_440_315#_c_354_n N_A_375_419#_c_1075_n 0.0642029f $X=4.58 $Y=0.68
+ $X2=0 $Y2=0
cc_353 N_A_440_315#_c_355_n N_A_375_419#_c_1075_n 0.0129683f $X=3.895 $Y=0.68
+ $X2=0 $Y2=0
cc_354 N_A_440_315#_M1010_g N_A_416_113#_c_1219_n 0.00586918f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_355 N_A_440_315#_M1010_g N_A_416_113#_c_1220_n 0.0029704f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_356 N_A_440_315#_M1013_g N_A_416_113#_c_1228_n 0.00496375f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_357 N_A_440_315#_M1022_s N_A_416_113#_c_1230_n 0.00611506f $X=4.52 $Y=1.84
+ $X2=0 $Y2=0
cc_358 N_A_440_315#_M1013_g N_A_416_113#_c_1230_n 0.0071737f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_359 N_A_440_315#_c_350_n N_A_416_113#_c_1230_n 0.00372063f $X=3.69 $Y=1.65
+ $X2=0 $Y2=0
cc_360 N_A_440_315#_c_356_n N_A_416_113#_c_1230_n 0.0196075f $X=4.665 $Y=1.985
+ $X2=0 $Y2=0
cc_361 N_A_440_315#_c_357_n N_A_416_113#_c_1230_n 0.00212633f $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_362 N_A_440_315#_c_358_n N_A_416_113#_c_1230_n 9.6797e-19 $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_363 N_A_440_315#_M1013_g N_A_416_113#_c_1247_n 0.00259711f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_364 N_A_440_315#_M1001_g N_A_416_113#_c_1231_n 3.98213e-19 $X=2.29 $Y=2.415
+ $X2=0 $Y2=0
cc_365 N_A_440_315#_c_348_n N_A_416_113#_c_1231_n 0.006398f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_366 N_A_440_315#_M1013_g N_A_416_113#_c_1231_n 0.00282008f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_367 N_A_440_315#_M1001_g N_A_416_113#_c_1226_n 5.37562e-19 $X=2.29 $Y=2.415
+ $X2=0 $Y2=0
cc_368 N_A_440_315#_M1010_g N_A_416_113#_c_1226_n 0.00190803f $X=2.505 $Y=0.995
+ $X2=0 $Y2=0
cc_369 N_A_440_315#_c_348_n N_A_416_113#_c_1226_n 0.00840933f $X=3.185 $Y=1.65
+ $X2=0 $Y2=0
cc_370 N_A_440_315#_M1013_g N_A_416_113#_c_1226_n 0.00427356f $X=3.275 $Y=2.315
+ $X2=0 $Y2=0
cc_371 N_A_440_315#_c_352_n N_A_416_113#_c_1226_n 0.00276536f $X=3.275 $Y=1.65
+ $X2=0 $Y2=0
cc_372 N_B_c_465_n N_A_1162_379#_c_585_n 0.00261039f $X=5.085 $Y=1.385 $X2=0
+ $Y2=0
cc_373 N_B_M1020_g N_A_27_134#_c_890_n 0.00578498f $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_374 N_B_M1020_g N_A_27_134#_c_891_n 0.0128816f $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_375 N_B_M1020_g N_A_27_134#_c_892_n 0.00536183f $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_376 N_B_M1023_g N_A_27_134#_c_893_n 0.00270621f $X=1.785 $Y=2.515 $X2=0 $Y2=0
cc_377 N_B_M1023_g N_A_27_134#_c_894_n 5.97507e-19 $X=1.785 $Y=2.515 $X2=0 $Y2=0
cc_378 N_B_M1003_g N_A_27_134#_c_894_n 0.00736636f $X=2.74 $Y=2.415 $X2=0 $Y2=0
cc_379 N_B_M1020_g N_A_27_134#_c_895_n 3.62456e-19 $X=2.005 $Y=0.885 $X2=0 $Y2=0
cc_380 N_B_M1017_g N_A_27_134#_c_895_n 3.86096e-19 $X=3.175 $Y=0.885 $X2=0 $Y2=0
cc_381 N_B_M1017_g N_A_27_134#_c_899_n 0.00169191f $X=3.175 $Y=0.885 $X2=0 $Y2=0
cc_382 N_B_c_468_n N_VPWR_c_976_n 0.00232846f $X=1.875 $Y=3.15 $X2=0 $Y2=0
cc_383 N_B_c_470_n N_VPWR_c_977_n 0.00229165f $X=4.295 $Y=3.15 $X2=0 $Y2=0
cc_384 N_B_c_458_n N_VPWR_c_977_n 8.59752e-19 $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_385 N_B_M1022_g N_VPWR_c_977_n 0.0205358f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_386 B N_VPWR_c_977_n 0.0133645f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_387 N_B_c_465_n N_VPWR_c_977_n 0.00163639f $X=5.085 $Y=1.385 $X2=0 $Y2=0
cc_388 N_B_c_468_n N_VPWR_c_984_n 0.0612182f $X=1.875 $Y=3.15 $X2=0 $Y2=0
cc_389 N_B_M1022_g N_VPWR_c_984_n 0.00460063f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_390 N_B_c_467_n N_VPWR_c_975_n 0.0182655f $X=2.65 $Y=3.15 $X2=0 $Y2=0
cc_391 N_B_c_468_n N_VPWR_c_975_n 0.00678686f $X=1.875 $Y=3.15 $X2=0 $Y2=0
cc_392 N_B_c_470_n N_VPWR_c_975_n 0.0436088f $X=4.295 $Y=3.15 $X2=0 $Y2=0
cc_393 N_B_M1022_g N_VPWR_c_975_n 0.00909358f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_394 N_B_c_473_n N_VPWR_c_975_n 0.00445015f $X=2.74 $Y=3.15 $X2=0 $Y2=0
cc_395 N_B_M1023_g N_A_375_419#_c_1084_n 0.00644408f $X=1.785 $Y=2.515 $X2=0
+ $Y2=0
cc_396 N_B_M1003_g N_A_375_419#_c_1085_n 0.0163577f $X=2.74 $Y=2.415 $X2=0 $Y2=0
cc_397 N_B_M1023_g N_A_375_419#_c_1097_n 0.0023625f $X=1.785 $Y=2.515 $X2=0
+ $Y2=0
cc_398 N_B_M1017_g N_A_375_419#_c_1074_n 0.00780549f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_399 N_B_c_456_n N_A_375_419#_c_1075_n 0.0143527f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_400 N_B_c_459_n N_A_375_419#_c_1075_n 0.0121042f $X=4.435 $Y=1.22 $X2=0 $Y2=0
cc_401 N_B_c_461_n N_A_375_419#_c_1075_n 0.0134432f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_402 N_B_M1017_g N_A_375_419#_c_1076_n 0.00724099f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_403 N_B_c_456_n N_A_375_419#_c_1076_n 0.00420304f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_404 N_B_c_459_n N_A_375_419#_c_1122_n 8.24696e-19 $X=4.435 $Y=1.22 $X2=0
+ $Y2=0
cc_405 N_B_c_461_n N_A_375_419#_c_1122_n 0.00826933f $X=4.935 $Y=1.22 $X2=0
+ $Y2=0
cc_406 B N_A_375_419#_c_1077_n 0.0050401f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_407 N_B_c_465_n N_A_375_419#_c_1077_n 5.83726e-19 $X=5.085 $Y=1.385 $X2=0
+ $Y2=0
cc_408 N_B_c_461_n N_A_375_419#_c_1126_n 0.00670237f $X=4.935 $Y=1.22 $X2=0
+ $Y2=0
cc_409 B N_A_375_419#_c_1126_n 0.00729471f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_410 N_B_c_465_n N_A_375_419#_c_1126_n 6.76062e-19 $X=5.085 $Y=1.385 $X2=0
+ $Y2=0
cc_411 N_B_c_453_n N_A_416_113#_c_1220_n 0.0129409f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_412 N_B_M1017_g N_A_416_113#_c_1220_n 0.00870892f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_413 N_B_M1020_g N_A_416_113#_c_1221_n 0.0064969f $X=2.005 $Y=0.885 $X2=0
+ $Y2=0
cc_414 N_B_c_453_n N_A_416_113#_c_1221_n 0.00305251f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_415 N_B_c_461_n N_A_416_113#_c_1223_n 0.00482248f $X=4.935 $Y=1.22 $X2=0
+ $Y2=0
cc_416 B N_A_416_113#_c_1223_n 3.28587e-19 $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_417 N_B_c_457_n N_A_416_113#_c_1230_n 0.00154074f $X=4.37 $Y=1.52 $X2=0 $Y2=0
cc_418 N_B_c_458_n N_A_416_113#_c_1230_n 0.00524423f $X=4.37 $Y=3.075 $X2=0
+ $Y2=0
cc_419 N_B_M1022_g N_A_416_113#_c_1230_n 0.0114668f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_420 B N_A_416_113#_c_1230_n 0.00403396f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_421 N_B_c_464_n N_A_416_113#_c_1230_n 0.00248958f $X=4.8 $Y=1.385 $X2=0 $Y2=0
cc_422 N_B_M1003_g N_A_416_113#_c_1231_n 0.00280848f $X=2.74 $Y=2.415 $X2=0
+ $Y2=0
cc_423 N_B_M1022_g N_A_416_113#_c_1233_n 0.00212654f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_424 N_B_M1017_g N_A_416_113#_c_1226_n 0.0203921f $X=3.175 $Y=0.885 $X2=0
+ $Y2=0
cc_425 N_B_M1022_g N_A_416_113#_c_1227_n 0.00670504f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_426 B N_A_416_113#_c_1227_n 0.020093f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_427 N_B_c_465_n N_A_416_113#_c_1227_n 0.0052234f $X=5.085 $Y=1.385 $X2=0
+ $Y2=0
cc_428 N_B_c_461_n N_VGND_c_1364_n 0.00174649f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_429 N_B_c_454_n N_VGND_c_1368_n 0.0625641f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_430 N_B_c_461_n N_VGND_c_1368_n 0.00278237f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_431 N_B_c_453_n N_VGND_c_1375_n 0.0268561f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_432 N_B_c_454_n N_VGND_c_1375_n 0.0104612f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_433 N_B_c_456_n N_VGND_c_1375_n 0.0367758f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_434 N_B_c_461_n N_VGND_c_1375_n 0.00359083f $X=4.935 $Y=1.22 $X2=0 $Y2=0
cc_435 N_B_c_462_n N_VGND_c_1375_n 0.00512617f $X=3.175 $Y=0.18 $X2=0 $Y2=0
cc_436 N_A_1162_379#_c_586_n N_C_M1012_g 0.0108913f $X=5.9 $Y=2.045 $X2=0 $Y2=0
cc_437 N_A_1162_379#_c_587_n N_C_M1012_g 0.00850299f $X=6.155 $Y=1.895 $X2=0
+ $Y2=0
cc_438 N_A_1162_379#_c_589_n N_C_M1012_g 0.00509764f $X=6.095 $Y=2.905 $X2=0
+ $Y2=0
cc_439 N_A_1162_379#_c_590_n N_C_M1012_g 0.0179723f $X=7.28 $Y=2.99 $X2=0 $Y2=0
cc_440 N_A_1162_379#_c_592_n N_C_M1012_g 0.00543171f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_441 N_A_1162_379#_M1005_g N_C_c_687_n 0.00796138f $X=6.155 $Y=0.855 $X2=0
+ $Y2=0
cc_442 N_A_1162_379#_c_581_n N_C_c_688_n 0.00405392f $X=7.72 $Y=2.195 $X2=0
+ $Y2=0
cc_443 N_A_1162_379#_c_582_n N_C_c_688_n 0.002567f $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_444 N_A_1162_379#_c_584_n N_C_c_689_n 2.17322e-19 $X=6.015 $Y=1.52 $X2=0
+ $Y2=0
cc_445 N_A_1162_379#_c_585_n N_C_c_689_n 0.0164644f $X=6.015 $Y=1.52 $X2=0 $Y2=0
cc_446 N_A_1162_379#_c_583_n N_C_c_690_n 0.00961036f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_447 N_A_1162_379#_c_592_n N_C_M1016_g 0.00245686f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_448 N_A_1162_379#_c_581_n N_C_M1016_g 0.0378294f $X=7.72 $Y=2.195 $X2=0 $Y2=0
cc_449 N_A_1162_379#_c_582_n N_C_M1016_g 0.00140204f $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_450 N_A_1162_379#_c_582_n N_C_c_692_n 5.32204e-19 $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_451 N_A_1162_379#_c_583_n N_C_c_692_n 0.0128944f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_452 N_A_1162_379#_c_583_n N_C_c_693_n 0.00248458f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_453 N_A_1162_379#_c_583_n N_C_c_694_n 0.00802643f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_454 N_A_1162_379#_c_582_n N_C_c_695_n 0.0101509f $X=7.9 $Y=1.435 $X2=0 $Y2=0
cc_455 N_A_1162_379#_c_583_n N_C_c_695_n 0.00286998f $X=7.86 $Y=0.6 $X2=0 $Y2=0
cc_456 N_A_1162_379#_c_589_n N_A_1198_424#_M1015_d 0.0130668f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_457 N_A_1162_379#_c_590_n N_A_1198_424#_M1015_d 0.00897796f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_458 N_A_1162_379#_c_591_n N_A_1198_424#_M1015_d 4.04887e-19 $X=6.18 $Y=2.99
+ $X2=0 $Y2=0
cc_459 N_A_1162_379#_c_583_n N_A_1198_424#_M1002_g 0.00421174f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_460 N_A_1162_379#_c_582_n N_A_1198_424#_c_786_n 0.00141437f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_461 N_A_1162_379#_c_583_n N_A_1198_424#_c_786_n 0.00100179f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_462 N_A_1162_379#_M1005_g N_A_1198_424#_c_789_n 0.00398659f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_463 N_A_1162_379#_c_584_n N_A_1198_424#_c_790_n 0.0495155f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_464 N_A_1162_379#_c_585_n N_A_1198_424#_c_790_n 0.00304279f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_465 N_A_1162_379#_c_581_n N_A_1198_424#_c_791_n 0.00164698f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_466 N_A_1162_379#_c_582_n N_A_1198_424#_c_791_n 0.0135398f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_467 N_A_1162_379#_c_583_n N_A_1198_424#_c_791_n 0.00890402f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_468 N_A_1162_379#_M1016_s N_A_1198_424#_c_795_n 0.00536549f $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_469 N_A_1162_379#_c_581_n N_A_1198_424#_c_795_n 0.0259303f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_470 N_A_1162_379#_c_582_n N_A_1198_424#_c_795_n 0.00698104f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_471 N_A_1162_379#_c_588_n N_A_1198_424#_c_796_n 0.00253348f $X=6.155 $Y=1.97
+ $X2=0 $Y2=0
cc_472 N_A_1162_379#_c_589_n N_A_1198_424#_c_796_n 0.00729123f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_473 N_A_1162_379#_c_587_n N_A_1198_424#_c_792_n 0.00304279f $X=6.155 $Y=1.895
+ $X2=0 $Y2=0
cc_474 N_A_1162_379#_c_589_n N_A_1198_424#_c_792_n 0.0495155f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_475 N_A_1162_379#_c_590_n N_A_1198_424#_c_792_n 0.0122348f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_476 N_A_1162_379#_c_581_n N_A_1198_424#_c_798_n 0.00541743f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_477 N_A_1162_379#_c_586_n N_VPWR_c_977_n 0.00249745f $X=5.9 $Y=2.045 $X2=0
+ $Y2=0
cc_478 N_A_1162_379#_c_588_n N_VPWR_c_977_n 0.00201311f $X=6.155 $Y=1.97 $X2=0
+ $Y2=0
cc_479 N_A_1162_379#_c_581_n N_VPWR_c_978_n 0.05018f $X=7.72 $Y=2.195 $X2=0
+ $Y2=0
cc_480 N_A_1162_379#_c_582_n N_VPWR_c_978_n 0.00322867f $X=7.9 $Y=1.435 $X2=0
+ $Y2=0
cc_481 N_A_1162_379#_c_590_n N_VPWR_c_979_n 0.00703128f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_482 N_A_1162_379#_c_592_n N_VPWR_c_1027_n 0.0145254f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_483 N_A_1162_379#_c_586_n N_VPWR_c_985_n 0.005209f $X=5.9 $Y=2.045 $X2=0
+ $Y2=0
cc_484 N_A_1162_379#_c_590_n N_VPWR_c_985_n 0.0823131f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_485 N_A_1162_379#_c_591_n N_VPWR_c_985_n 0.0121867f $X=6.18 $Y=2.99 $X2=0
+ $Y2=0
cc_486 N_A_1162_379#_c_586_n N_VPWR_c_975_n 0.00990867f $X=5.9 $Y=2.045 $X2=0
+ $Y2=0
cc_487 N_A_1162_379#_c_590_n N_VPWR_c_975_n 0.0471112f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_488 N_A_1162_379#_c_591_n N_VPWR_c_975_n 0.00660921f $X=6.18 $Y=2.99 $X2=0
+ $Y2=0
cc_489 N_A_1162_379#_c_581_n N_VPWR_c_975_n 0.0125625f $X=7.72 $Y=2.195 $X2=0
+ $Y2=0
cc_490 N_A_1162_379#_c_590_n N_A_375_419#_M1012_d 0.00292446f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_491 N_A_1162_379#_M1005_g N_A_375_419#_c_1078_n 0.00442722f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_492 N_A_1162_379#_M1005_g N_A_375_419#_c_1079_n 0.00730004f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_493 N_A_1162_379#_c_583_n N_A_375_419#_c_1079_n 0.00472011f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_494 N_A_1162_379#_c_590_n N_A_375_419#_c_1087_n 0.0151051f $X=7.28 $Y=2.99
+ $X2=0 $Y2=0
cc_495 N_A_1162_379#_c_592_n N_A_375_419#_c_1087_n 0.0119875f $X=7.365 $Y=2.905
+ $X2=0 $Y2=0
cc_496 N_A_1162_379#_c_581_n N_A_375_419#_c_1087_n 0.0235137f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_497 N_A_1162_379#_M1016_s N_A_375_419#_c_1088_n 0.00357637f $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_498 N_A_1162_379#_c_581_n N_A_375_419#_c_1088_n 0.0204983f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_499 N_A_1162_379#_M1016_s N_A_375_419#_c_1081_n 2.42181e-19 $X=7.3 $Y=1.84
+ $X2=0 $Y2=0
cc_500 N_A_1162_379#_c_581_n N_A_375_419#_c_1081_n 0.0181632f $X=7.72 $Y=2.195
+ $X2=0 $Y2=0
cc_501 N_A_1162_379#_c_582_n N_A_375_419#_c_1081_n 0.0130101f $X=7.9 $Y=1.435
+ $X2=0 $Y2=0
cc_502 N_A_1162_379#_c_583_n N_A_375_419#_c_1081_n 0.0076654f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_503 N_A_1162_379#_c_583_n N_A_375_419#_c_1082_n 0.0505046f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_504 N_A_1162_379#_c_583_n N_A_375_419#_c_1083_n 0.0130296f $X=7.86 $Y=0.6
+ $X2=0 $Y2=0
cc_505 N_A_1162_379#_c_586_n N_A_416_113#_c_1229_n 0.0140432f $X=5.9 $Y=2.045
+ $X2=0 $Y2=0
cc_506 N_A_1162_379#_c_591_n N_A_416_113#_c_1229_n 0.00383535f $X=6.18 $Y=2.99
+ $X2=0 $Y2=0
cc_507 N_A_1162_379#_M1005_g N_A_416_113#_c_1222_n 0.0150552f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_508 N_A_1162_379#_c_584_n N_A_416_113#_c_1222_n 0.0251443f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_509 N_A_1162_379#_c_585_n N_A_416_113#_c_1222_n 0.00161433f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_510 N_A_1162_379#_M1005_g N_A_416_113#_c_1278_n 0.0107362f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_511 N_A_1162_379#_M1005_g N_A_416_113#_c_1279_n 0.00552867f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_512 N_A_1162_379#_c_589_n N_A_416_113#_c_1232_n 0.00107267f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_513 N_A_1162_379#_c_586_n N_A_416_113#_c_1233_n 0.00264311f $X=5.9 $Y=2.045
+ $X2=0 $Y2=0
cc_514 N_A_1162_379#_c_588_n N_A_416_113#_c_1233_n 0.0060626f $X=6.155 $Y=1.97
+ $X2=0 $Y2=0
cc_515 N_A_1162_379#_c_589_n N_A_416_113#_c_1233_n 0.0440126f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_516 N_A_1162_379#_M1005_g N_A_416_113#_c_1227_n 0.00453554f $X=6.155 $Y=0.855
+ $X2=0 $Y2=0
cc_517 N_A_1162_379#_c_588_n N_A_416_113#_c_1227_n 6.6135e-19 $X=6.155 $Y=1.97
+ $X2=0 $Y2=0
cc_518 N_A_1162_379#_c_589_n N_A_416_113#_c_1227_n 0.0110355f $X=6.095 $Y=2.905
+ $X2=0 $Y2=0
cc_519 N_A_1162_379#_c_584_n N_A_416_113#_c_1227_n 0.0248017f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_520 N_A_1162_379#_c_585_n N_A_416_113#_c_1227_n 0.00507613f $X=6.015 $Y=1.52
+ $X2=0 $Y2=0
cc_521 N_A_1162_379#_M1005_g N_VGND_c_1364_n 2.09474e-19 $X=6.155 $Y=0.855 $X2=0
+ $Y2=0
cc_522 N_A_1162_379#_c_583_n N_VGND_c_1365_n 0.0415257f $X=7.86 $Y=0.6 $X2=0
+ $Y2=0
cc_523 N_A_1162_379#_M1005_g N_VGND_c_1369_n 6.51701e-19 $X=6.155 $Y=0.855 $X2=0
+ $Y2=0
cc_524 N_A_1162_379#_c_583_n N_VGND_c_1369_n 0.0101731f $X=7.86 $Y=0.6 $X2=0
+ $Y2=0
cc_525 N_A_1162_379#_c_583_n N_VGND_c_1375_n 0.00902782f $X=7.86 $Y=0.6 $X2=0
+ $Y2=0
cc_526 N_C_M1016_g N_A_1198_424#_M1004_g 0.00729948f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_527 N_C_c_694_n N_A_1198_424#_M1002_g 0.0144313f $X=8.075 $Y=0.885 $X2=0
+ $Y2=0
cc_528 N_C_c_690_n N_A_1198_424#_c_786_n 0.00538345f $X=7.735 $Y=1.355 $X2=0
+ $Y2=0
cc_529 N_C_c_695_n N_A_1198_424#_c_786_n 0.00464217f $X=7.66 $Y=1.355 $X2=0
+ $Y2=0
cc_530 N_C_c_687_n N_A_1198_424#_c_789_n 0.00167979f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_531 C N_A_1198_424#_c_789_n 0.023585f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_532 N_C_c_689_n N_A_1198_424#_c_790_n 0.00754199f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_533 N_C_M1012_g N_A_1198_424#_c_795_n 0.00993509f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_534 N_C_c_688_n N_A_1198_424#_c_795_n 0.00341283f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_535 N_C_c_689_n N_A_1198_424#_c_795_n 8.5126e-19 $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_536 N_C_M1016_g N_A_1198_424#_c_795_n 0.00320669f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_537 C N_A_1198_424#_c_795_n 0.00148248f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_538 N_C_M1012_g N_A_1198_424#_c_796_n 0.00212698f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_539 N_C_M1012_g N_A_1198_424#_c_792_n 0.0248884f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_540 N_C_c_689_n N_A_1198_424#_c_792_n 0.0054384f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_541 C N_A_1198_424#_c_792_n 0.00784722f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_542 N_C_M1016_g N_A_1198_424#_c_798_n 0.0016766f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_543 N_C_M1016_g N_VPWR_c_978_n 0.0087502f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_544 N_C_M1012_g N_VPWR_c_985_n 0.00333926f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_545 N_C_M1016_g N_VPWR_c_985_n 0.00377165f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_546 N_C_M1012_g N_VPWR_c_975_n 0.00430191f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_547 N_C_M1016_g N_VPWR_c_975_n 0.00493777f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_548 N_C_c_687_n N_A_375_419#_c_1079_n 0.00455332f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_549 N_C_c_694_n N_A_375_419#_c_1079_n 0.00234865f $X=8.075 $Y=0.885 $X2=0
+ $Y2=0
cc_550 N_C_M1012_g N_A_375_419#_c_1087_n 0.00565088f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_551 N_C_M1016_g N_A_375_419#_c_1087_n 0.00198175f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_552 N_C_c_688_n N_A_375_419#_c_1088_n 0.00435379f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_553 N_C_c_689_n N_A_375_419#_c_1088_n 0.00112054f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_554 N_C_M1016_g N_A_375_419#_c_1088_n 0.0012064f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_555 C N_A_375_419#_c_1088_n 0.00530888f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_556 N_C_M1012_g N_A_375_419#_c_1089_n 0.00396157f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_557 N_C_c_689_n N_A_375_419#_c_1089_n 0.00576853f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_558 C N_A_375_419#_c_1089_n 0.0141845f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_559 N_C_M1012_g N_A_375_419#_c_1081_n 0.00399377f $X=6.66 $Y=2.54 $X2=0 $Y2=0
cc_560 N_C_c_687_n N_A_375_419#_c_1081_n 3.87848e-19 $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_561 N_C_c_688_n N_A_375_419#_c_1081_n 0.0133863f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_562 N_C_c_689_n N_A_375_419#_c_1081_n 0.00180986f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_563 N_C_c_690_n N_A_375_419#_c_1081_n 0.00178741f $X=7.735 $Y=1.355 $X2=0
+ $Y2=0
cc_564 N_C_M1016_g N_A_375_419#_c_1081_n 0.00141422f $X=7.75 $Y=2.16 $X2=0 $Y2=0
cc_565 N_C_c_695_n N_A_375_419#_c_1081_n 3.52513e-19 $X=7.66 $Y=1.355 $X2=0
+ $Y2=0
cc_566 C N_A_375_419#_c_1081_n 0.0307052f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_567 N_C_c_687_n N_A_375_419#_c_1082_n 0.00692779f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_568 N_C_c_693_n N_A_375_419#_c_1082_n 0.00547767f $X=7.81 $Y=0.96 $X2=0 $Y2=0
cc_569 N_C_c_694_n N_A_375_419#_c_1082_n 9.09628e-19 $X=8.075 $Y=0.885 $X2=0
+ $Y2=0
cc_570 N_C_c_687_n N_A_375_419#_c_1083_n 0.00194033f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_571 N_C_c_688_n N_A_375_419#_c_1083_n 0.00513991f $X=7.66 $Y=1.43 $X2=0 $Y2=0
cc_572 N_C_c_690_n N_A_375_419#_c_1083_n 0.00375665f $X=7.735 $Y=1.355 $X2=0
+ $Y2=0
cc_573 C N_A_375_419#_c_1083_n 0.00675568f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_574 C N_A_416_113#_M1009_d 0.00270076f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_575 N_C_c_687_n N_A_416_113#_c_1278_n 0.00141899f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_576 N_C_c_687_n N_A_416_113#_c_1224_n 0.00409002f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_577 N_C_c_689_n N_A_416_113#_c_1224_n 0.00460589f $X=7.14 $Y=1.43 $X2=0 $Y2=0
cc_578 C N_A_416_113#_c_1224_n 0.0110577f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_579 N_C_c_687_n N_A_416_113#_c_1225_n 0.0113393f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_580 C N_A_416_113#_c_1225_n 3.08063e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_581 N_C_c_690_n N_VGND_c_1365_n 5.24626e-19 $X=7.735 $Y=1.355 $X2=0 $Y2=0
cc_582 N_C_c_694_n N_VGND_c_1365_n 0.00684806f $X=8.075 $Y=0.885 $X2=0 $Y2=0
cc_583 N_C_c_694_n N_VGND_c_1369_n 0.00537471f $X=8.075 $Y=0.885 $X2=0 $Y2=0
cc_584 N_C_c_693_n N_VGND_c_1375_n 0.00289176f $X=7.81 $Y=0.96 $X2=0 $Y2=0
cc_585 N_C_c_694_n N_VGND_c_1375_n 0.00539454f $X=8.075 $Y=0.885 $X2=0 $Y2=0
cc_586 N_A_1198_424#_c_795_n N_VPWR_M1016_d 0.00991372f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_587 N_A_1198_424#_c_838_p N_VPWR_M1016_d 0.00624964f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_588 N_A_1198_424#_c_798_n N_VPWR_M1016_d 0.00582584f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_A_1198_424#_M1004_g N_VPWR_c_978_n 0.00177932f $X=8.645 $Y=2.4 $X2=0
+ $Y2=0
cc_590 N_A_1198_424#_c_795_n N_VPWR_c_978_n 0.0202422f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_591 N_A_1198_424#_c_838_p N_VPWR_c_978_n 0.00275409f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_592 N_A_1198_424#_c_798_n N_VPWR_c_978_n 0.0227956f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_593 N_A_1198_424#_M1004_g N_VPWR_c_979_n 0.00564635f $X=8.645 $Y=2.4 $X2=0
+ $Y2=0
cc_594 N_A_1198_424#_M1007_g N_VPWR_c_981_n 0.00649215f $X=9.095 $Y=2.4 $X2=0
+ $Y2=0
cc_595 N_A_1198_424#_c_786_n N_VPWR_c_1027_n 0.00132101f $X=8.555 $Y=1.485 $X2=0
+ $Y2=0
cc_596 N_A_1198_424#_c_791_n N_VPWR_c_1027_n 0.00123758f $X=8.36 $Y=1.485 $X2=0
+ $Y2=0
cc_597 N_A_1198_424#_c_795_n N_VPWR_c_1027_n 0.00448577f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_598 N_A_1198_424#_c_838_p N_VPWR_c_1027_n 0.00428557f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_599 N_A_1198_424#_c_798_n N_VPWR_c_1027_n 0.0136724f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_600 N_A_1198_424#_M1004_g N_VPWR_c_986_n 0.005209f $X=8.645 $Y=2.4 $X2=0
+ $Y2=0
cc_601 N_A_1198_424#_M1007_g N_VPWR_c_986_n 0.005209f $X=9.095 $Y=2.4 $X2=0
+ $Y2=0
cc_602 N_A_1198_424#_M1004_g N_VPWR_c_975_n 0.00986839f $X=8.645 $Y=2.4 $X2=0
+ $Y2=0
cc_603 N_A_1198_424#_M1007_g N_VPWR_c_975_n 0.00986008f $X=9.095 $Y=2.4 $X2=0
+ $Y2=0
cc_604 N_A_1198_424#_c_795_n N_A_375_419#_c_1087_n 0.0191656f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_605 N_A_1198_424#_c_796_n N_A_375_419#_c_1087_n 0.0011513f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_606 N_A_1198_424#_c_792_n N_A_375_419#_c_1087_n 0.0248614f $X=6.48 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_A_1198_424#_c_795_n N_A_375_419#_c_1088_n 0.0189311f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_A_1198_424#_c_795_n N_A_375_419#_c_1089_n 0.00661589f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_609 N_A_1198_424#_c_796_n N_A_375_419#_c_1089_n 0.00118398f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_A_1198_424#_c_792_n N_A_375_419#_c_1089_n 0.0117642f $X=6.48 $Y=2.035
+ $X2=0 $Y2=0
cc_611 N_A_1198_424#_M1005_d N_A_416_113#_c_1222_n 0.00152064f $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_612 N_A_1198_424#_c_789_n N_A_416_113#_c_1222_n 0.0138486f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_613 N_A_1198_424#_c_790_n N_A_416_113#_c_1222_n 0.00129791f $X=6.527 $Y=1.525
+ $X2=0 $Y2=0
cc_614 N_A_1198_424#_M1005_d N_A_416_113#_c_1278_n 0.00304149f $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_615 N_A_1198_424#_c_789_n N_A_416_113#_c_1278_n 0.00577431f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_616 N_A_1198_424#_M1005_d N_A_416_113#_c_1279_n 8.211e-19 $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_617 N_A_1198_424#_M1005_d N_A_416_113#_c_1225_n 0.00779558f $X=6.23 $Y=0.535
+ $X2=0 $Y2=0
cc_618 N_A_1198_424#_c_789_n N_A_416_113#_c_1225_n 0.0134906f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_619 N_A_1198_424#_c_790_n N_A_416_113#_c_1225_n 0.00575786f $X=6.527 $Y=1.525
+ $X2=0 $Y2=0
cc_620 N_A_1198_424#_M1004_g X 0.0206202f $X=8.645 $Y=2.4 $X2=0 $Y2=0
cc_621 N_A_1198_424#_M1002_g X 0.0188787f $X=8.655 $Y=0.76 $X2=0 $Y2=0
cc_622 N_A_1198_424#_c_783_n X 0.008373f $X=9.005 $Y=1.395 $X2=0 $Y2=0
cc_623 N_A_1198_424#_M1007_g X 0.0353121f $X=9.095 $Y=2.4 $X2=0 $Y2=0
cc_624 N_A_1198_424#_M1014_g X 0.0192976f $X=9.085 $Y=0.76 $X2=0 $Y2=0
cc_625 N_A_1198_424#_c_787_n X 0.00777273f $X=8.645 $Y=1.485 $X2=0 $Y2=0
cc_626 N_A_1198_424#_c_788_n X 0.00663376f $X=9.095 $Y=1.395 $X2=0 $Y2=0
cc_627 N_A_1198_424#_c_791_n X 0.050671f $X=8.36 $Y=1.485 $X2=0 $Y2=0
cc_628 N_A_1198_424#_c_838_p X 0.00732723f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_629 N_A_1198_424#_M1002_g N_VGND_c_1365_n 0.00969831f $X=8.655 $Y=0.76 $X2=0
+ $Y2=0
cc_630 N_A_1198_424#_c_786_n N_VGND_c_1365_n 0.0029613f $X=8.555 $Y=1.485 $X2=0
+ $Y2=0
cc_631 N_A_1198_424#_c_791_n N_VGND_c_1365_n 0.0278705f $X=8.36 $Y=1.485 $X2=0
+ $Y2=0
cc_632 N_A_1198_424#_M1014_g N_VGND_c_1367_n 0.00650727f $X=9.085 $Y=0.76 $X2=0
+ $Y2=0
cc_633 N_A_1198_424#_M1002_g N_VGND_c_1370_n 0.00537471f $X=8.655 $Y=0.76 $X2=0
+ $Y2=0
cc_634 N_A_1198_424#_M1014_g N_VGND_c_1370_n 0.00537471f $X=9.085 $Y=0.76 $X2=0
+ $Y2=0
cc_635 N_A_1198_424#_M1002_g N_VGND_c_1375_n 0.00539454f $X=8.655 $Y=0.76 $X2=0
+ $Y2=0
cc_636 N_A_1198_424#_M1014_g N_VGND_c_1375_n 0.00539454f $X=9.085 $Y=0.76 $X2=0
+ $Y2=0
cc_637 N_A_27_134#_c_901_n N_VPWR_c_976_n 0.0286637f $X=0.43 $Y=2.425 $X2=0
+ $Y2=0
cc_638 N_A_27_134#_c_901_n N_VPWR_c_982_n 0.0205351f $X=0.43 $Y=2.425 $X2=0
+ $Y2=0
cc_639 N_A_27_134#_c_901_n N_VPWR_c_975_n 0.0184615f $X=0.43 $Y=2.425 $X2=0
+ $Y2=0
cc_640 N_A_27_134#_c_892_n N_A_375_419#_c_1084_n 0.00838799f $X=2.35 $Y=1.48
+ $X2=0 $Y2=0
cc_641 N_A_27_134#_c_893_n N_A_375_419#_c_1084_n 0.00484309f $X=1.965 $Y=1.48
+ $X2=0 $Y2=0
cc_642 N_A_27_134#_c_894_n N_A_375_419#_c_1084_n 0.0127976f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_643 N_A_27_134#_M1001_d N_A_375_419#_c_1085_n 0.00304139f $X=2.38 $Y=2.095
+ $X2=0 $Y2=0
cc_644 N_A_27_134#_c_894_n N_A_375_419#_c_1085_n 0.0170259f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_645 N_A_27_134#_c_891_n N_A_416_113#_c_1219_n 0.0140676f $X=1.88 $Y=1.395
+ $X2=0 $Y2=0
cc_646 N_A_27_134#_c_892_n N_A_416_113#_c_1219_n 0.0141889f $X=2.35 $Y=1.48
+ $X2=0 $Y2=0
cc_647 N_A_27_134#_c_899_n N_A_416_113#_c_1219_n 0.0296524f $X=2.79 $Y=0.995
+ $X2=0 $Y2=0
cc_648 N_A_27_134#_M1010_d N_A_416_113#_c_1220_n 0.00913335f $X=2.58 $Y=0.785
+ $X2=0 $Y2=0
cc_649 N_A_27_134#_c_899_n N_A_416_113#_c_1220_n 0.0277569f $X=2.79 $Y=0.995
+ $X2=0 $Y2=0
cc_650 N_A_27_134#_c_894_n N_A_416_113#_c_1247_n 0.00133559f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_651 N_A_27_134#_c_894_n N_A_416_113#_c_1231_n 0.0236501f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_652 N_A_27_134#_c_894_n N_A_416_113#_c_1226_n 0.0132322f $X=2.515 $Y=2.275
+ $X2=0 $Y2=0
cc_653 N_A_27_134#_c_895_n N_A_416_113#_c_1226_n 0.00752401f $X=2.595 $Y=1.395
+ $X2=0 $Y2=0
cc_654 N_A_27_134#_c_898_n N_A_416_113#_c_1226_n 0.00844652f $X=2.515 $Y=1.48
+ $X2=0 $Y2=0
cc_655 N_A_27_134#_c_899_n N_A_416_113#_c_1226_n 0.0194534f $X=2.79 $Y=0.995
+ $X2=0 $Y2=0
cc_656 N_A_27_134#_c_890_n N_VGND_M1018_d 0.02171f $X=1.795 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_657 N_A_27_134#_c_890_n N_VGND_c_1368_n 0.0125374f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_658 N_A_27_134#_c_888_n N_VGND_c_1371_n 0.00698834f $X=0.265 $Y=0.83 $X2=0
+ $Y2=0
cc_659 N_A_27_134#_c_890_n N_VGND_c_1371_n 0.00286374f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_660 N_A_27_134#_c_890_n N_VGND_c_1372_n 0.0436747f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_661 N_A_27_134#_c_888_n N_VGND_c_1375_n 0.0107515f $X=0.265 $Y=0.83 $X2=0
+ $Y2=0
cc_662 N_A_27_134#_c_890_n N_VGND_c_1375_n 0.0288798f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_985_n N_A_416_113#_c_1229_n 0.0192342f $X=7.975 $Y=3.33 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_975_n N_A_416_113#_c_1229_n 0.0158523f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_665 N_VPWR_M1022_d N_A_416_113#_c_1230_n 0.00323229f $X=4.98 $Y=1.84 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_977_n N_A_416_113#_c_1230_n 0.0239351f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_977_n N_A_416_113#_c_1232_n 0.00263503f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_977_n N_A_416_113#_c_1233_n 0.0726098f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_977_n N_A_416_113#_c_1227_n 0.00496383f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_670 N_VPWR_c_978_n X 0.0049173f $X=8.06 $Y=1.985 $X2=0 $Y2=0
cc_671 N_VPWR_c_979_n X 0.0250331f $X=8.252 $Y=3.245 $X2=0 $Y2=0
cc_672 N_VPWR_c_981_n X 0.0395687f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_673 N_VPWR_c_986_n X 0.0144623f $X=9.235 $Y=3.33 $X2=0 $Y2=0
cc_674 N_VPWR_c_975_n X 0.0118344f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_675 N_VPWR_c_981_n N_VGND_c_1367_n 0.00814581f $X=9.32 $Y=1.985 $X2=0 $Y2=0
cc_676 N_A_375_419#_c_1085_n N_A_416_113#_M1003_d 0.00461307f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_677 N_A_375_419#_c_1074_n N_A_416_113#_c_1220_n 0.0135079f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_678 N_A_375_419#_c_1085_n N_A_416_113#_c_1228_n 0.0209219f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_679 N_A_375_419#_M1005_s N_A_416_113#_c_1222_n 0.00315345f $X=5.805 $Y=0.535
+ $X2=0 $Y2=0
cc_680 N_A_375_419#_c_1077_n N_A_416_113#_c_1222_n 0.00707829f $X=5.775 $Y=0.76
+ $X2=0 $Y2=0
cc_681 N_A_375_419#_c_1078_n N_A_416_113#_c_1222_n 0.0200365f $X=5.9 $Y=0.675
+ $X2=0 $Y2=0
cc_682 N_A_375_419#_c_1079_n N_A_416_113#_c_1222_n 0.00363379f $X=7.435 $Y=0.34
+ $X2=0 $Y2=0
cc_683 N_A_375_419#_c_1077_n N_A_416_113#_c_1223_n 0.0142807f $X=5.775 $Y=0.76
+ $X2=0 $Y2=0
cc_684 N_A_375_419#_c_1079_n N_A_416_113#_c_1279_n 0.0105973f $X=7.435 $Y=0.34
+ $X2=0 $Y2=0
cc_685 N_A_375_419#_c_1082_n N_A_416_113#_c_1224_n 0.0270814f $X=7.52 $Y=1.095
+ $X2=0 $Y2=0
cc_686 N_A_375_419#_c_1079_n N_A_416_113#_c_1225_n 0.0644024f $X=7.435 $Y=0.34
+ $X2=0 $Y2=0
cc_687 N_A_375_419#_c_1085_n N_A_416_113#_c_1230_n 0.00337922f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_688 N_A_375_419#_c_1074_n N_A_416_113#_c_1230_n 0.0188093f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_689 N_A_375_419#_c_1085_n N_A_416_113#_c_1247_n 0.00259371f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_690 N_A_375_419#_c_1074_n N_A_416_113#_c_1247_n 0.00237204f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_691 N_A_375_419#_c_1074_n N_A_416_113#_c_1226_n 0.112445f $X=3.47 $Y=0.71
+ $X2=0 $Y2=0
cc_692 N_A_375_419#_c_1075_n N_VGND_M1011_d 0.00247003f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_693 N_A_375_419#_c_1122_n N_VGND_M1011_d 0.00410163f $X=5.06 $Y=0.675 $X2=0
+ $Y2=0
cc_694 N_A_375_419#_c_1077_n N_VGND_M1011_d 0.0200041f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_695 N_A_375_419#_c_1126_n N_VGND_M1011_d 9.76702e-19 $X=5.145 $Y=0.76 $X2=0
+ $Y2=0
cc_696 N_A_375_419#_c_1075_n N_VGND_c_1364_n 0.0141996f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_697 N_A_375_419#_c_1122_n N_VGND_c_1364_n 0.00594708f $X=5.06 $Y=0.675 $X2=0
+ $Y2=0
cc_698 N_A_375_419#_c_1077_n N_VGND_c_1364_n 0.0192217f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_699 N_A_375_419#_c_1078_n N_VGND_c_1364_n 0.00547381f $X=5.9 $Y=0.675 $X2=0
+ $Y2=0
cc_700 N_A_375_419#_c_1080_n N_VGND_c_1364_n 0.0127057f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_701 N_A_375_419#_c_1079_n N_VGND_c_1365_n 0.00418126f $X=7.435 $Y=0.34 $X2=0
+ $Y2=0
cc_702 N_A_375_419#_c_1075_n N_VGND_c_1368_n 0.102488f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_703 N_A_375_419#_c_1076_n N_VGND_c_1368_n 0.0115893f $X=3.555 $Y=0.34 $X2=0
+ $Y2=0
cc_704 N_A_375_419#_c_1077_n N_VGND_c_1368_n 0.00270711f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_705 N_A_375_419#_c_1077_n N_VGND_c_1369_n 0.00350729f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_706 N_A_375_419#_c_1079_n N_VGND_c_1369_n 0.102958f $X=7.435 $Y=0.34 $X2=0
+ $Y2=0
cc_707 N_A_375_419#_c_1080_n N_VGND_c_1369_n 0.0177305f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_708 N_A_375_419#_c_1075_n N_VGND_c_1375_n 0.0553628f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_709 N_A_375_419#_c_1076_n N_VGND_c_1375_n 0.00583135f $X=3.555 $Y=0.34 $X2=0
+ $Y2=0
cc_710 N_A_375_419#_c_1077_n N_VGND_c_1375_n 0.0116289f $X=5.775 $Y=0.76 $X2=0
+ $Y2=0
cc_711 N_A_375_419#_c_1079_n N_VGND_c_1375_n 0.0596141f $X=7.435 $Y=0.34 $X2=0
+ $Y2=0
cc_712 N_A_375_419#_c_1080_n N_VGND_c_1375_n 0.00968346f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_713 N_A_416_113#_c_1223_n N_VGND_M1011_d 0.00213745f $X=5.68 $Y=1.1 $X2=0
+ $Y2=0
cc_714 N_A_416_113#_c_1220_n N_VGND_c_1368_n 0.0284116f $X=3.045 $Y=0.51 $X2=0
+ $Y2=0
cc_715 N_A_416_113#_c_1221_n N_VGND_c_1368_n 0.00581481f $X=2.305 $Y=0.51 $X2=0
+ $Y2=0
cc_716 N_A_416_113#_c_1220_n N_VGND_c_1375_n 0.0270015f $X=3.045 $Y=0.51 $X2=0
+ $Y2=0
cc_717 N_A_416_113#_c_1221_n N_VGND_c_1375_n 0.00530552f $X=2.305 $Y=0.51 $X2=0
+ $Y2=0
cc_718 X N_VGND_c_1365_n 0.0308484f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_719 X N_VGND_c_1367_n 0.0294122f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_720 X N_VGND_c_1370_n 0.0134077f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_721 X N_VGND_c_1375_n 0.0119261f $X=8.795 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o311ai_1.pxi.spice
* Created: Fri Aug 28 18:01:12 2020
* 
x_PM_SKY130_FD_SC_MS__O311AI_1%A1 N_A1_M1003_g N_A1_M1002_g A1 N_A1_c_55_n
+ N_A1_c_56_n PM_SKY130_FD_SC_MS__O311AI_1%A1
x_PM_SKY130_FD_SC_MS__O311AI_1%A2 N_A2_M1008_g N_A2_M1004_g A2 A2 A2 A2
+ N_A2_c_82_n N_A2_c_83_n PM_SKY130_FD_SC_MS__O311AI_1%A2
x_PM_SKY130_FD_SC_MS__O311AI_1%A3 N_A3_M1007_g N_A3_M1009_g A3 N_A3_c_121_n
+ N_A3_c_122_n PM_SKY130_FD_SC_MS__O311AI_1%A3
x_PM_SKY130_FD_SC_MS__O311AI_1%B1 N_B1_M1005_g N_B1_M1006_g B1 N_B1_c_153_n
+ N_B1_c_154_n PM_SKY130_FD_SC_MS__O311AI_1%B1
x_PM_SKY130_FD_SC_MS__O311AI_1%C1 N_C1_c_186_n N_C1_M1001_g N_C1_M1000_g C1
+ N_C1_c_189_n PM_SKY130_FD_SC_MS__O311AI_1%C1
x_PM_SKY130_FD_SC_MS__O311AI_1%VPWR N_VPWR_M1002_s N_VPWR_M1005_d N_VPWR_c_214_n
+ N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_218_n VPWR
+ N_VPWR_c_219_n N_VPWR_c_213_n PM_SKY130_FD_SC_MS__O311AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O311AI_1%Y N_Y_M1001_d N_Y_M1007_d N_Y_M1000_d N_Y_c_252_n
+ N_Y_c_253_n N_Y_c_254_n N_Y_c_250_n N_Y_c_251_n N_Y_c_256_n Y Y Y N_Y_c_257_n
+ PM_SKY130_FD_SC_MS__O311AI_1%Y
x_PM_SKY130_FD_SC_MS__O311AI_1%VGND N_VGND_M1003_s N_VGND_M1008_d N_VGND_c_302_n
+ N_VGND_c_303_n N_VGND_c_304_n VGND N_VGND_c_305_n N_VGND_c_306_n
+ N_VGND_c_307_n N_VGND_c_308_n PM_SKY130_FD_SC_MS__O311AI_1%VGND
x_PM_SKY130_FD_SC_MS__O311AI_1%A_128_74# N_A_128_74#_M1003_d N_A_128_74#_M1009_d
+ N_A_128_74#_c_337_n N_A_128_74#_c_345_n N_A_128_74#_c_338_n
+ N_A_128_74#_c_353_n N_A_128_74#_c_339_n PM_SKY130_FD_SC_MS__O311AI_1%A_128_74#
cc_1 VNB N_A1_M1003_g 0.0316595f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_2 VNB N_A1_c_55_n 0.0290951f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_3 VNB N_A1_c_56_n 0.0178902f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_4 VNB N_A2_M1008_g 0.0280323f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_5 VNB N_A2_c_82_n 0.0251117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A2_c_83_n 0.00519747f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.565
cc_7 VNB N_A3_M1007_g 0.00652164f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_8 VNB A3 0.00613168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_c_121_n 0.0335647f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_10 VNB N_A3_c_122_n 0.020506f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_11 VNB N_B1_M1005_g 0.0071114f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_12 VNB B1 0.00839315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_153_n 0.0306255f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_14 VNB N_B1_c_154_n 0.0181734f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_15 VNB N_C1_c_186_n 0.0227334f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.35
cc_16 VNB N_C1_M1000_g 0.00919457f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_17 VNB C1 0.0124946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C1_c_189_n 0.0667459f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_19 VNB N_VPWR_c_213_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_250_n 0.00413443f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.565
cc_21 VNB N_Y_c_251_n 0.030059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_302_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_23 VNB N_VGND_c_303_n 0.0451868f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_VGND_c_304_n 0.0115377f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_25 VNB N_VGND_c_305_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_306_n 0.049013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_307_n 0.214603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_308_n 0.0107715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_128_74#_c_337_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_30 VNB N_A_128_74#_c_338_n 0.0102186f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.515
cc_31 VNB N_A_128_74#_c_339_n 0.00294871f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.68
cc_32 VPB N_A1_M1002_g 0.0253535f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_33 VPB N_A1_c_55_n 0.00579078f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_34 VPB N_A1_c_56_n 0.0125724f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_35 VPB N_A2_M1004_g 0.0223898f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_36 VPB N_A2_c_82_n 0.00557768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A2_c_83_n 0.00171527f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.565
cc_38 VPB N_A3_M1007_g 0.0260971f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_39 VPB N_B1_M1005_g 0.0246456f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_40 VPB N_C1_M1000_g 0.0300392f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_41 VPB N_VPWR_c_214_n 0.0155055f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_42 VPB N_VPWR_c_215_n 0.0484671f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_43 VPB N_VPWR_c_216_n 0.00976275f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.68
cc_44 VPB N_VPWR_c_217_n 0.0498463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_218_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_219_n 0.0225072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_213_n 0.0810881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_Y_c_252_n 0.00285226f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.515
cc_49 VPB N_Y_c_253_n 0.00685577f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_50 VPB N_Y_c_254_n 0.0104749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_Y_c_250_n 7.3943e-19 $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.565
cc_52 VPB N_Y_c_256_n 0.0109693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_Y_c_257_n 0.0502116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 N_A1_M1003_g N_A2_M1008_g 0.0181074f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_55 N_A1_M1002_g N_A2_M1004_g 0.0443527f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_56 N_A1_c_55_n N_A2_c_82_n 0.0443527f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_57 N_A1_c_56_n N_A2_c_82_n 0.00153198f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_58 N_A1_M1002_g N_A2_c_83_n 0.00453772f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_59 N_A1_c_55_n N_A2_c_83_n 5.46266e-19 $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_60 N_A1_c_56_n N_A2_c_83_n 0.0257291f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_61 N_A1_M1002_g N_VPWR_c_215_n 0.0222746f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A1_c_55_n N_VPWR_c_215_n 7.79182e-19 $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_63 N_A1_c_56_n N_VPWR_c_215_n 0.0262242f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_64 N_A1_M1002_g N_VPWR_c_217_n 0.00460063f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_65 N_A1_M1002_g N_VPWR_c_213_n 0.00908371f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A1_M1003_g N_VGND_c_303_n 0.0184904f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_67 N_A1_c_55_n N_VGND_c_303_n 0.00156574f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_68 N_A1_c_56_n N_VGND_c_303_n 0.0236882f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A1_M1003_g N_VGND_c_305_n 0.00434272f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A1_M1003_g N_VGND_c_307_n 0.0082426f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A1_M1003_g N_A_128_74#_c_337_n 0.00632535f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A1_M1003_g N_A_128_74#_c_338_n 0.00375706f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A1_c_55_n N_A_128_74#_c_338_n 0.00171791f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A1_c_56_n N_A_128_74#_c_338_n 0.00625586f $X=0.54 $Y=1.515 $X2=0 $Y2=0
cc_75 N_A2_M1004_g N_A3_M1007_g 0.0387697f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A2_M1008_g A3 0.00151734f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A2_c_82_n A3 2.36557e-19 $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A2_c_83_n A3 0.0141439f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A2_M1008_g N_A3_c_121_n 0.00407278f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A2_c_82_n N_A3_c_121_n 0.0171673f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A2_c_83_n N_A3_c_121_n 0.0174397f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A2_M1008_g N_A3_c_122_n 0.0162896f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A2_M1004_g N_VPWR_c_215_n 0.00345211f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A2_c_83_n N_VPWR_c_215_n 0.0364692f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A2_M1004_g N_VPWR_c_217_n 0.00365007f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A2_c_83_n N_VPWR_c_217_n 0.0105186f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A2_M1004_g N_VPWR_c_213_n 0.00444515f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A2_c_83_n N_VPWR_c_213_n 0.011939f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A2_c_83_n A_225_368# 0.0163138f $X=1.11 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_90 N_A2_c_83_n N_Y_c_252_n 0.0380302f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A2_c_83_n N_Y_c_254_n 0.00726162f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_92 N_A2_M1008_g N_VGND_c_304_n 0.00488678f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A2_M1008_g N_VGND_c_305_n 0.00461464f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A2_M1008_g N_VGND_c_307_n 0.00465508f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A2_M1008_g N_A_128_74#_c_337_n 4.71232e-19 $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A2_M1008_g N_A_128_74#_c_345_n 0.0120154f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A2_c_82_n N_A_128_74#_c_345_n 9.22244e-19 $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A2_c_83_n N_A_128_74#_c_345_n 0.0155033f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A2_M1008_g N_A_128_74#_c_338_n 0.00106811f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A3_M1007_g N_B1_M1005_g 0.0269438f $X=1.605 $Y=2.4 $X2=0 $Y2=0
cc_101 A3 B1 0.0261333f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_102 N_A3_c_122_n B1 0.00229487f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_103 A3 N_B1_c_153_n 3.90318e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A3_c_121_n N_B1_c_153_n 0.0174805f $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_105 N_A3_c_122_n N_B1_c_154_n 0.0200745f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A3_M1007_g N_VPWR_c_217_n 0.00553757f $X=1.605 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A3_M1007_g N_VPWR_c_213_n 0.0109203f $X=1.605 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A3_M1007_g N_Y_c_252_n 0.0152086f $X=1.605 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A3_M1007_g N_Y_c_254_n 0.00241247f $X=1.605 $Y=2.4 $X2=0 $Y2=0
cc_110 A3 N_Y_c_254_n 0.00503923f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A3_c_121_n N_Y_c_254_n 4.61395e-19 $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_112 N_A3_c_122_n N_VGND_c_304_n 0.00603858f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A3_c_122_n N_VGND_c_306_n 0.00461464f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A3_c_122_n N_VGND_c_307_n 0.00465894f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_115 A3 N_A_128_74#_c_345_n 0.0228656f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A3_c_121_n N_A_128_74#_c_345_n 9.98643e-19 $X=1.68 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A3_c_122_n N_A_128_74#_c_345_n 0.0134555f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_118 N_A3_c_122_n N_A_128_74#_c_339_n 0.00281817f $X=1.68 $Y=1.22 $X2=0 $Y2=0
cc_119 N_B1_c_154_n N_C1_c_186_n 0.0363339f $X=2.25 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_120 N_B1_M1005_g N_C1_M1000_g 0.0254685f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_121 B1 N_C1_c_189_n 3.61714e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_c_153_n N_C1_c_189_n 0.0174432f $X=2.25 $Y=1.385 $X2=0 $Y2=0
cc_123 N_B1_M1005_g N_VPWR_c_216_n 0.00347203f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B1_M1005_g N_VPWR_c_217_n 0.005209f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B1_M1005_g N_VPWR_c_213_n 0.00983871f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_126 N_B1_M1005_g N_Y_c_252_n 0.0151624f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B1_M1005_g N_Y_c_253_n 0.0135147f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_128 B1 N_Y_c_253_n 0.0221856f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_c_153_n N_Y_c_253_n 0.00104284f $X=2.25 $Y=1.385 $X2=0 $Y2=0
cc_130 N_B1_M1005_g N_Y_c_254_n 0.00242245f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_131 B1 N_Y_c_254_n 0.00592165f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_M1005_g N_Y_c_250_n 0.00337768f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_133 B1 N_Y_c_250_n 0.0282201f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B1_c_153_n N_Y_c_250_n 0.00187211f $X=2.25 $Y=1.385 $X2=0 $Y2=0
cc_135 N_B1_c_154_n N_Y_c_251_n 0.00893686f $X=2.25 $Y=1.22 $X2=0 $Y2=0
cc_136 N_B1_M1005_g N_Y_c_257_n 7.06246e-19 $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_137 N_B1_c_154_n N_VGND_c_306_n 0.00433834f $X=2.25 $Y=1.22 $X2=0 $Y2=0
cc_138 N_B1_c_154_n N_VGND_c_307_n 0.00822046f $X=2.25 $Y=1.22 $X2=0 $Y2=0
cc_139 B1 N_A_128_74#_c_353_n 0.0124978f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_c_153_n N_A_128_74#_c_353_n 6.10381e-19 $X=2.25 $Y=1.385 $X2=0 $Y2=0
cc_141 N_B1_c_154_n N_A_128_74#_c_353_n 0.00280745f $X=2.25 $Y=1.22 $X2=0 $Y2=0
cc_142 N_B1_c_154_n N_A_128_74#_c_339_n 0.00863906f $X=2.25 $Y=1.22 $X2=0 $Y2=0
cc_143 N_C1_M1000_g N_VPWR_c_216_n 0.00879843f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_144 N_C1_M1000_g N_VPWR_c_219_n 0.005209f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_145 N_C1_M1000_g N_VPWR_c_213_n 0.00987248f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_146 N_C1_M1000_g N_Y_c_252_n 9.55194e-19 $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_147 N_C1_c_186_n N_Y_c_250_n 0.00786229f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_148 N_C1_M1000_g N_Y_c_250_n 0.00728919f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_149 C1 N_Y_c_250_n 0.0265523f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_150 N_C1_c_189_n N_Y_c_250_n 0.00898252f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_151 N_C1_c_186_n N_Y_c_251_n 0.0179308f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_152 C1 N_Y_c_251_n 0.0160699f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_153 N_C1_c_189_n N_Y_c_251_n 0.00520334f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_154 N_C1_M1000_g N_Y_c_256_n 0.0190313f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_155 C1 N_Y_c_256_n 0.0263919f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_156 N_C1_c_189_n N_Y_c_256_n 0.00648981f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_157 N_C1_M1000_g N_Y_c_257_n 0.0163047f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_158 N_C1_c_186_n N_VGND_c_306_n 0.00291513f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_159 N_C1_c_186_n N_VGND_c_307_n 0.00363424f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_160 N_C1_c_186_n N_A_128_74#_c_339_n 5.78724e-19 $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_161 N_VPWR_c_216_n N_Y_c_252_n 0.0353111f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_162 N_VPWR_c_217_n N_Y_c_252_n 0.014549f $X=2.285 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_c_213_n N_Y_c_252_n 0.0119743f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_M1005_d N_Y_c_253_n 0.00286648f $X=2.265 $Y=1.84 $X2=0 $Y2=0
cc_165 N_VPWR_c_216_n N_Y_c_253_n 0.0213608f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_166 N_VPWR_c_216_n N_Y_c_256_n 0.0011721f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_167 N_VPWR_c_216_n N_Y_c_257_n 0.0336136f $X=2.45 $Y=2.145 $X2=0 $Y2=0
cc_168 N_VPWR_c_219_n N_Y_c_257_n 0.0190111f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VPWR_c_213_n N_Y_c_257_n 0.0156676f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_170 N_Y_c_251_n N_VGND_c_306_n 0.0228546f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_171 N_Y_c_251_n N_VGND_c_307_n 0.0185794f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_172 N_Y_c_251_n N_A_128_74#_c_353_n 0.00803923f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_173 N_Y_c_251_n N_A_128_74#_c_339_n 0.0219699f $X=2.945 $Y=0.515 $X2=0 $Y2=0
cc_174 N_Y_c_250_n A_469_74# 0.0013188f $X=2.67 $Y=1.72 $X2=-0.19 $Y2=-0.245
cc_175 N_Y_c_251_n A_469_74# 0.00783876f $X=2.945 $Y=0.515 $X2=-0.19 $Y2=-0.245
cc_176 N_VGND_c_303_n N_A_128_74#_c_337_n 0.0191389f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_177 N_VGND_c_304_n N_A_128_74#_c_337_n 0.0132958f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_178 N_VGND_c_305_n N_A_128_74#_c_337_n 0.0145639f $X=1.115 $Y=0 $X2=0 $Y2=0
cc_179 N_VGND_c_307_n N_A_128_74#_c_337_n 0.0119984f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_180 N_VGND_M1008_d N_A_128_74#_c_345_n 0.0183532f $X=1.095 $Y=0.37 $X2=0
+ $Y2=0
cc_181 N_VGND_c_304_n N_A_128_74#_c_345_n 0.0352958f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_182 N_VGND_c_307_n N_A_128_74#_c_345_n 0.0130717f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_c_303_n N_A_128_74#_c_338_n 0.0124832f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_184 N_VGND_c_304_n N_A_128_74#_c_339_n 0.00286618f $X=1.405 $Y=0.515 $X2=0
+ $Y2=0
cc_185 N_VGND_c_306_n N_A_128_74#_c_339_n 0.0158357f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_307_n N_A_128_74#_c_339_n 0.0121432f $X=3.12 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o31a_1.spice
* Created: Fri Aug 28 18:02:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o31a_1.pex.spice"
.subckt sky130_fd_sc_ms__o31a_1  VNB VPB A1 A2 A3 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_84_48#_M1008_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.2109 PD=1.25478 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1007 N_A_230_94#_M1007_d N_A1_M1007_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1136 AS=0.144093 PD=0.995 PS=1.08522 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75000.8 SB=75002 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_230_94#_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1136 PD=1.21 PS=0.995 NRD=28.116 NRS=14.052 M=1 R=4.26667
+ SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_230_94#_M1000_d N_A3_M1000_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1104 AS=0.1824 PD=0.985 PS=1.21 NRD=12.18 NRS=26.244 M=1 R=4.26667
+ SA=75002 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1001 N_A_84_48#_M1001_d N_B1_M1001_g N_A_230_94#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2272 AS=0.1104 PD=1.99 PS=0.985 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75002.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A_84_48#_M1006_g N_X_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.290355 AS=0.3136 PD=1.72226 PS=2.8 NRD=19.7788 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1004 A_259_368# N_A1_M1004_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.259245 PD=1.24 PS=1.53774 NRD=12.7853 NRS=23.64 M=1 R=5.55556 SA=90000.9
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1009 A_343_368# N_A2_M1009_g A_259_368# VPB PSHORT L=0.18 W=1 AD=0.165 AS=0.12
+ PD=1.33 PS=1.24 NRD=21.6503 NRS=12.7853 M=1 R=5.55556 SA=90001.3 SB=90001.3
+ A=0.18 P=2.36 MULT=1
MM1002 N_A_84_48#_M1002_d N_A3_M1002_g A_343_368# VPB PSHORT L=0.18 W=1
+ AD=0.188696 AS=0.165 PD=1.47826 PS=1.33 NRD=0 NRS=21.6503 M=1 R=5.55556
+ SA=90001.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g N_A_84_48#_M1002_d VPB PSHORT L=0.18 W=0.84
+ AD=0.3864 AS=0.158504 PD=2.6 PS=1.24174 NRD=0 NRS=20.3107 M=1 R=4.66667
+ SA=90002.3 SB=90000.4 A=0.1512 P=2.04 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__o31a_1.pxi.spice"
*
.ends
*
*

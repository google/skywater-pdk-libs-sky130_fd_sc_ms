# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__and4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.450000 1.390000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.980000 1.345000 4.365000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.930000 1.470000 3.260000 1.800000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.097400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.830000 0.350000 5.080000 0.960000 ;
        RECT 4.830000 0.960000 6.595000 1.130000 ;
        RECT 4.875000 1.800000 6.105000 1.970000 ;
        RECT 4.875000 1.970000 5.205000 2.980000 ;
        RECT 5.760000 0.350000 6.090000 0.960000 ;
        RECT 5.855000 1.480000 6.595000 1.650000 ;
        RECT 5.855000 1.650000 6.105000 1.800000 ;
        RECT 5.855000 1.970000 6.105000 2.980000 ;
        RECT 6.365000 1.130000 6.595000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  1.950000 0.395000 3.245000 ;
      RECT 0.140000  0.315000 2.110000 0.485000 ;
      RECT 0.140000  0.485000 0.390000 1.255000 ;
      RECT 0.565000  1.950000 1.730000 2.240000 ;
      RECT 0.570000  0.655000 1.760000 0.835000 ;
      RECT 0.720000  1.005000 1.330000 1.255000 ;
      RECT 0.720000  1.255000 0.890000 1.950000 ;
      RECT 1.015000  2.410000 1.345000 3.245000 ;
      RECT 1.560000  1.600000 2.760000 1.770000 ;
      RECT 1.560000  1.770000 1.730000 1.950000 ;
      RECT 1.560000  2.240000 1.730000 2.980000 ;
      RECT 1.930000  1.940000 2.260000 3.245000 ;
      RECT 1.940000  0.485000 2.110000 1.130000 ;
      RECT 1.940000  1.130000 4.070000 1.175000 ;
      RECT 1.940000  1.175000 3.810000 1.300000 ;
      RECT 2.290000  0.575000 2.620000 0.790000 ;
      RECT 2.290000  0.790000 3.640000 0.825000 ;
      RECT 2.290000  0.825000 3.470000 0.960000 ;
      RECT 2.430000  1.770000 2.760000 1.970000 ;
      RECT 2.430000  1.970000 4.705000 2.120000 ;
      RECT 2.430000  2.120000 4.145000 2.140000 ;
      RECT 2.430000  2.140000 2.760000 2.980000 ;
      RECT 2.800000  0.085000 3.130000 0.620000 ;
      RECT 2.930000  2.310000 3.645000 3.245000 ;
      RECT 3.300000  0.575000 3.640000 0.790000 ;
      RECT 3.640000  0.995000 4.070000 1.130000 ;
      RECT 3.815000  1.950000 4.705000 1.970000 ;
      RECT 3.815000  2.140000 4.145000 2.980000 ;
      RECT 4.315000  2.290000 4.645000 3.245000 ;
      RECT 4.330000  0.085000 4.660000 1.130000 ;
      RECT 4.535000  1.300000 5.685000 1.630000 ;
      RECT 4.535000  1.630000 4.705000 1.950000 ;
      RECT 5.260000  0.085000 5.590000 0.790000 ;
      RECT 5.405000  2.140000 5.655000 3.245000 ;
      RECT 6.260000  0.085000 6.520000 0.680000 ;
      RECT 6.275000  1.820000 6.605000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ms__and4_4
END LIBRARY

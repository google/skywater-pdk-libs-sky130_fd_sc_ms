# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sedfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sedfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.28000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.835000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.485000 0.350000 15.825000 2.150000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.355000 0.350000 16.685000 0.960000 ;
        RECT 16.355000 0.960000 17.165000 1.130000 ;
        RECT 16.435000 1.805000 17.165000 1.975000 ;
        RECT 16.435000 1.975000 16.665000 3.010000 ;
        RECT 16.700000 1.130000 17.165000 1.805000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.125000 1.180000 5.635000 1.510000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.180000 4.915000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.705000 1.180000 7.045000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 17.280000 0.085000 ;
        RECT  1.070000  0.085000  1.400000 0.810000 ;
        RECT  2.180000  0.085000  2.510000 1.005000 ;
        RECT  4.960000  0.085000  5.290000 1.010000 ;
        RECT  6.415000  0.085000  6.745000 0.920000 ;
        RECT  7.555000  0.085000  7.725000 1.130000 ;
        RECT 10.270000  0.085000 10.520000 0.680000 ;
        RECT 11.710000  0.085000 11.960000 0.680000 ;
        RECT 13.320000  0.085000 14.335000 0.600000 ;
        RECT 14.065000  0.600000 14.335000 1.120000 ;
        RECT 15.065000  0.085000 15.315000 1.130000 ;
        RECT 16.005000  0.085000 16.175000 1.130000 ;
        RECT 16.855000  0.085000 17.115000 0.790000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
        RECT 16.955000 -0.085000 17.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 17.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 17.280000 3.415000 ;
        RECT  1.065000 2.630000  1.315000 3.245000 ;
        RECT  2.505000 2.630000  2.755000 3.245000 ;
        RECT  5.035000 2.595000  5.305000 3.245000 ;
        RECT  6.485000 2.650000  6.735000 3.245000 ;
        RECT  7.795000 2.650000  8.125000 3.245000 ;
        RECT 10.225000 2.730000 10.555000 3.245000 ;
        RECT 11.320000 2.730000 11.650000 3.245000 ;
        RECT 13.765000 2.650000 14.305000 3.245000 ;
        RECT 15.035000 2.660000 15.365000 3.245000 ;
        RECT 15.935000 2.660000 16.265000 3.245000 ;
        RECT 16.835000 2.145000 17.165000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
        RECT 16.475000 3.245000 16.645000 3.415000 ;
        RECT 16.955000 3.245000 17.125000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 17.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.420000  0.580000 0.730000 ;
      RECT  0.085000 0.730000  0.255000 2.290000 ;
      RECT  0.085000 2.290000  1.655000 2.460000 ;
      RECT  0.085000 2.460000  0.525000 2.980000 ;
      RECT  1.005000 1.110000  2.010000 1.280000 ;
      RECT  1.005000 1.280000  1.335000 1.950000 ;
      RECT  1.005000 1.950000  2.635000 2.120000 ;
      RECT  1.485000 2.460000  1.655000 2.905000 ;
      RECT  1.485000 2.905000  2.335000 3.075000 ;
      RECT  1.680000 0.545000  2.010000 1.110000 ;
      RECT  1.825000 2.120000  1.995000 2.735000 ;
      RECT  2.165000 2.290000  3.545000 2.460000 ;
      RECT  2.165000 2.460000  2.335000 2.905000 ;
      RECT  2.305000 1.515000  2.635000 1.950000 ;
      RECT  2.875000 1.515000  3.205000 1.845000 ;
      RECT  3.000000 0.545000  3.330000 1.175000 ;
      RECT  3.000000 1.175000  3.545000 1.345000 ;
      RECT  3.265000 2.460000  3.545000 2.970000 ;
      RECT  3.375000 1.345000  3.545000 2.290000 ;
      RECT  3.500000 0.545000  3.885000 1.005000 ;
      RECT  3.715000 1.005000  3.885000 2.290000 ;
      RECT  3.715000 2.290000  3.965000 2.905000 ;
      RECT  3.715000 2.905000  4.865000 3.075000 ;
      RECT  4.055000 0.365000  4.305000 0.605000 ;
      RECT  4.055000 0.605000  4.790000 1.010000 ;
      RECT  4.055000 1.010000  4.305000 1.680000 ;
      RECT  4.055000 1.680000  6.135000 1.850000 ;
      RECT  4.055000 1.850000  4.305000 2.055000 ;
      RECT  4.135000 2.055000  4.305000 2.245000 ;
      RECT  4.135000 2.245000  4.525000 2.735000 ;
      RECT  4.695000 2.255000  6.475000 2.310000 ;
      RECT  4.695000 2.310000  8.465000 2.425000 ;
      RECT  4.695000 2.425000  4.865000 2.905000 ;
      RECT  5.805000 1.430000  6.135000 1.680000 ;
      RECT  5.805000 1.850000  6.135000 2.085000 ;
      RECT  5.820000 0.605000  6.150000 1.090000 ;
      RECT  5.820000 1.090000  6.475000 1.260000 ;
      RECT  5.845000 2.425000  8.465000 2.480000 ;
      RECT  5.845000 2.480000  6.305000 2.925000 ;
      RECT  6.305000 1.260000  6.475000 2.255000 ;
      RECT  6.855000 1.820000  7.655000 2.140000 ;
      RECT  6.915000 0.350000  7.385000 1.010000 ;
      RECT  7.215000 1.010000  7.385000 1.470000 ;
      RECT  7.215000 1.470000  7.655000 1.820000 ;
      RECT  7.905000 0.255000  9.735000 0.425000 ;
      RECT  7.905000 0.425000  8.235000 1.130000 ;
      RECT  7.905000 1.480000  8.715000 1.650000 ;
      RECT  7.905000 1.650000  8.075000 2.310000 ;
      RECT  8.245000 1.820000  9.055000 2.140000 ;
      RECT  8.295000 2.480000  9.055000 2.650000 ;
      RECT  8.465000 0.595000  8.715000 1.480000 ;
      RECT  8.725000 2.140000  9.055000 2.305000 ;
      RECT  8.805000 2.650000  9.055000 2.980000 ;
      RECT  8.885000 0.425000  9.055000 1.820000 ;
      RECT  9.225000 0.595000  9.395000 1.690000 ;
      RECT  9.225000 1.690000 10.940000 1.860000 ;
      RECT  9.225000 1.860000  9.395000 2.530000 ;
      RECT  9.225000 2.530000  9.585000 2.980000 ;
      RECT  9.565000 0.425000  9.735000 0.850000 ;
      RECT  9.565000 0.850000 10.860000 1.020000 ;
      RECT  9.565000 1.020000  9.855000 1.345000 ;
      RECT  9.565000 2.030000  9.925000 2.360000 ;
      RECT  9.755000 2.360000  9.925000 2.390000 ;
      RECT  9.755000 2.390000 12.720000 2.560000 ;
      RECT 10.065000 1.190000 11.885000 1.360000 ;
      RECT 10.065000 1.360000 10.395000 1.520000 ;
      RECT 10.610000 1.530000 10.940000 1.690000 ;
      RECT 10.690000 0.255000 11.540000 0.425000 ;
      RECT 10.690000 0.425000 10.860000 0.850000 ;
      RECT 10.760000 2.050000 11.385000 2.220000 ;
      RECT 11.030000 0.595000 11.200000 1.190000 ;
      RECT 11.215000 1.360000 11.885000 1.520000 ;
      RECT 11.215000 1.520000 11.385000 2.050000 ;
      RECT 11.370000 0.425000 11.540000 0.850000 ;
      RECT 11.370000 0.850000 12.250000 1.020000 ;
      RECT 12.080000 1.020000 12.250000 1.130000 ;
      RECT 12.080000 1.130000 13.525000 1.300000 ;
      RECT 12.080000 1.300000 12.380000 1.800000 ;
      RECT 12.420000 0.350000 12.750000 0.770000 ;
      RECT 12.420000 0.770000 13.865000 0.940000 ;
      RECT 12.550000 1.470000 12.985000 1.800000 ;
      RECT 12.550000 1.800000 12.720000 2.390000 ;
      RECT 12.890000 2.520000 13.325000 2.980000 ;
      RECT 13.155000 1.715000 13.865000 1.885000 ;
      RECT 13.155000 1.885000 13.325000 2.520000 ;
      RECT 13.195000 1.300000 13.525000 1.545000 ;
      RECT 13.585000 2.055000 15.235000 2.320000 ;
      RECT 13.585000 2.320000 16.185000 2.380000 ;
      RECT 13.695000 0.940000 13.865000 1.300000 ;
      RECT 13.695000 1.300000 14.495000 1.630000 ;
      RECT 13.695000 1.630000 13.865000 1.715000 ;
      RECT 14.475000 1.800000 15.235000 2.055000 ;
      RECT 14.475000 2.380000 16.185000 2.490000 ;
      RECT 14.475000 2.490000 14.835000 2.980000 ;
      RECT 14.505000 0.350000 14.835000 1.130000 ;
      RECT 14.665000 1.130000 14.835000 1.550000 ;
      RECT 14.665000 1.550000 15.235000 1.800000 ;
      RECT 15.995000 1.300000 16.510000 1.635000 ;
      RECT 15.995000 1.635000 16.185000 2.320000 ;
    LAYER mcon ;
      RECT  3.035000 1.580000  3.205000 1.750000 ;
      RECT 15.035000 1.580000 15.205000 1.750000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000 15.265000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT 14.975000 1.550000 15.265000 1.595000 ;
      RECT 14.975000 1.735000 15.265000 1.780000 ;
  END
END sky130_fd_sc_ms__sedfxbp_2

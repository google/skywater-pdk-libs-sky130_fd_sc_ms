* File: sky130_fd_sc_ms__dfxbp_1.pex.spice
* Created: Fri Aug 28 17:24:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFXBP_1%CLK 3 5 7 8 12 15
c33 12 0 2.6712e-20 $X=0.335 $Y=1.385
c34 3 0 1.76233e-19 $X=0.5 $Y=2.4
r35 14 15 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.5 $Y2=1.385
r36 11 14 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.335 $Y=1.385
+ $X2=0.495 $Y2=1.385
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.335
+ $Y=1.385 $X2=0.335 $Y2=1.385
r38 8 12 2.95898 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.335 $Y2=1.365
r39 5 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r40 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
r41 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.55 $X2=0.5
+ $Y2=1.385
r42 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.5 $Y=1.55 $X2=0.5
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_27_74# 1 2 9 11 13 16 20 22 24 26 30 33 37
+ 41 45 48 49 50 51 53 55 56 59 60 61 62 65 68 70 75 76 78 80 83 84 85 89
c241 89 0 2.50478e-20 $X=1.135 $Y=1.385
c242 80 0 4.89519e-20 $X=0.965 $Y=1.385
c243 75 0 6.57199e-20 $X=5.55 $Y=0.455
c244 65 0 1.87448e-19 $X=3.285 $Y=1.91
c245 37 0 6.7972e-20 $X=5.64 $Y=1.3
c246 30 0 1.76992e-19 $X=5.64 $Y=0.94
c247 26 0 3.57825e-20 $X=5.34 $Y=1.895
c248 20 0 1.32495e-19 $X=3.175 $Y=2.75
c249 16 0 4.57052e-20 $X=3.015 $Y=0.805
c250 11 0 2.6712e-20 $X=1.135 $Y=1.22
c251 9 0 9.05393e-20 $X=0.95 $Y=2.4
r252 91 93 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.015 $Y=1.91
+ $X2=3.175 $Y2=1.91
r253 84 85 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.48 $Y=0.52
+ $X2=4.65 $Y2=0.52
r254 81 89 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.965 $Y=1.385
+ $X2=1.135 $Y2=1.385
r255 81 86 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.965 $Y=1.385
+ $X2=0.95 $Y2=1.385
r256 80 82 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=1.385
+ $X2=0.88 $Y2=1.55
r257 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.385 $X2=0.965 $Y2=1.385
r258 76 98 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.55 $Y=0.455
+ $X2=5.55 $Y2=0.62
r259 75 85 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=5.55 $Y=0.455
+ $X2=4.65 $Y2=0.455
r260 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=0.455 $X2=5.55 $Y2=0.455
r261 72 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.665
+ $X2=3.57 $Y2=0.665
r262 72 84 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.655 $Y=0.665
+ $X2=4.48 $Y2=0.665
r263 69 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.75
+ $X2=3.57 $Y2=0.665
r264 69 70 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.57 $Y=0.75 $X2=3.57
+ $Y2=1.75
r265 68 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.58
+ $X2=3.57 $Y2=0.665
r266 67 68 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.57 $Y=0.425
+ $X2=3.57 $Y2=0.58
r267 65 93 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.285 $Y=1.91
+ $X2=3.175 $Y2=1.91
r268 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.285
+ $Y=1.91 $X2=3.285 $Y2=1.91
r269 62 70 7.72402 $w=3.25e-07 $l=2.00035e-07 $layer=LI1_cond $X=3.485 $Y=1.912
+ $X2=3.57 $Y2=1.75
r270 62 64 7.09196 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=3.485 $Y=1.912
+ $X2=3.285 $Y2=1.912
r271 60 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.485 $Y=0.34
+ $X2=3.57 $Y2=0.425
r272 60 61 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.485 $Y=0.34
+ $X2=2.545 $Y2=0.34
r273 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=0.425
+ $X2=2.545 $Y2=0.34
r274 58 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.46 $Y=0.425
+ $X2=2.46 $Y2=0.73
r275 57 78 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.09 $Y=0.815
+ $X2=0.88 $Y2=0.815
r276 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=0.815
+ $X2=2.46 $Y2=0.73
r277 56 57 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=2.375 $Y=0.815
+ $X2=1.09 $Y2=0.815
r278 55 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.755 $Y=1.72
+ $X2=0.755 $Y2=1.55
r279 53 80 1.23476 $w=4.18e-07 $l=4.5e-08 $layer=LI1_cond $X=0.88 $Y=1.34
+ $X2=0.88 $Y2=1.385
r280 52 78 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0.9 $X2=0.88
+ $Y2=0.815
r281 52 53 12.0732 $w=4.18e-07 $l=4.4e-07 $layer=LI1_cond $X=0.88 $Y=0.9
+ $X2=0.88 $Y2=1.34
r282 50 78 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.67 $Y=0.815
+ $X2=0.88 $Y2=0.815
r283 50 51 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.67 $Y=0.815
+ $X2=0.445 $Y2=0.815
r284 48 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.67 $Y=1.805
+ $X2=0.755 $Y2=1.72
r285 48 49 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.67 $Y=1.805
+ $X2=0.36 $Y2=1.805
r286 45 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.73
+ $X2=0.445 $Y2=0.815
r287 45 47 1.84848 $w=3.3e-07 $l=5e-08 $layer=LI1_cond $X=0.28 $Y=0.73 $X2=0.28
+ $Y2=0.68
r288 41 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.235 $Y=1.985
+ $X2=0.235 $Y2=2.815
r289 39 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.235 $Y=1.89
+ $X2=0.36 $Y2=1.805
r290 39 41 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.235 $Y=1.89
+ $X2=0.235 $Y2=1.985
r291 35 37 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.34 $Y=1.3 $X2=5.64
+ $Y2=1.3
r292 30 98 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.64 $Y=0.94
+ $X2=5.64 $Y2=0.62
r293 28 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.64 $Y=1.225
+ $X2=5.64 $Y2=1.3
r294 28 30 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.64 $Y=1.225
+ $X2=5.64 $Y2=0.94
r295 26 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.34 $Y=1.895
+ $X2=5.34 $Y2=1.97
r296 25 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.34 $Y=1.375
+ $X2=5.34 $Y2=1.3
r297 25 26 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.34 $Y=1.375
+ $X2=5.34 $Y2=1.895
r298 22 33 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=5.18 $Y=1.97
+ $X2=5.34 $Y2=1.97
r299 22 24 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.18 $Y=2.045
+ $X2=5.18 $Y2=2.54
r300 18 93 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=2.075
+ $X2=3.175 $Y2=1.91
r301 18 20 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.175 $Y=2.075
+ $X2=3.175 $Y2=2.75
r302 14 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.015 $Y=1.745
+ $X2=3.015 $Y2=1.91
r303 14 16 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.015 $Y=1.745
+ $X2=3.015 $Y2=0.805
r304 11 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.22
+ $X2=1.135 $Y2=1.385
r305 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.135 $Y=1.22
+ $X2=1.135 $Y2=0.74
r306 7 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.55
+ $X2=0.95 $Y2=1.385
r307 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.95 $Y=1.55 $X2=0.95
+ $Y2=2.4
r308 2 43 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=2.815
r309 2 41 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=1.985
r310 1 47 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%D 3 5 7 9 11 16 18 19 25 27 39
c62 39 0 8.5492e-20 $X=2.16 $Y=1.665
c63 25 0 3.08123e-19 $X=2.025 $Y=2.19
c64 18 0 4.57052e-20 $X=2.16 $Y=1.295
c65 16 0 1.99054e-19 $X=1.995 $Y=2.19
c66 5 0 1.35673e-19 $X=2.51 $Y=1.2
r67 33 39 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=2.09 $Y=1.6 $X2=2.09
+ $Y2=1.665
r68 27 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.175 $Y=1.2 $X2=2.175
+ $Y2=1.29
r69 19 41 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.09 $Y2=1.78
r70 19 39 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=2.09 $Y=1.675
+ $X2=2.09 $Y2=1.665
r71 19 33 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=2.09 $Y=1.59 $X2=2.09
+ $Y2=1.6
r72 18 19 9.60369 $w=3.58e-07 $l=3e-07 $layer=LI1_cond $X=2.09 $Y=1.29 $X2=2.09
+ $Y2=1.59
r73 18 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.175
+ $Y=1.29 $X2=2.175 $Y2=1.29
r74 14 25 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.865 $Y=2.19
+ $X2=2.025 $Y2=2.19
r75 13 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.865 $Y=2.19
+ $X2=1.995 $Y2=2.19
r76 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=2.19 $X2=1.865 $Y2=2.19
r77 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=2.025
+ $X2=1.995 $Y2=2.19
r78 11 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.995 $Y=2.025
+ $X2=1.995 $Y2=1.78
r79 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.585 $Y=1.125
+ $X2=2.585 $Y2=0.805
r80 6 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.2
+ $X2=2.175 $Y2=1.2
r81 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.51 $Y=1.2
+ $X2=2.585 $Y2=1.125
r82 5 6 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.51 $Y=1.2 $X2=2.34
+ $Y2=1.2
r83 1 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=2.355
+ $X2=2.025 $Y2=2.19
r84 1 3 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.025 $Y=2.355
+ $X2=2.025 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_208_368# 1 2 9 10 11 15 19 23 27 30 33 35
+ 37 39 41 44 45 48 51 54 55 58 62 66 72 74 76 78 79 83
c228 78 0 1.10354e-19 $X=5.825 $Y=1.78
c229 72 0 1.49219e-19 $X=4.89 $Y=1.52
c230 55 0 1.76233e-19 $X=1.222 $Y=2.63
c231 54 0 4.89519e-20 $X=1.635 $Y=1.65
c232 51 0 1.3952e-19 $X=1.43 $Y=1.756
c233 37 0 1.65203e-19 $X=3.12 $Y=2.8
c234 19 0 4.21193e-20 $X=3.49 $Y=0.72
c235 11 0 1.08514e-19 $X=2.55 $Y=1.74
r236 79 89 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.825 $Y=1.78
+ $X2=5.715 $Y2=1.78
r237 78 81 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=1.78
+ $X2=5.825 $Y2=1.945
r238 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.825
+ $Y=1.78 $X2=5.825 $Y2=1.78
r239 72 87 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.52
+ $X2=4.89 $Y2=1.355
r240 71 74 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.89 $Y=1.52
+ $X2=5.065 $Y2=1.52
r241 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.89
+ $Y=1.52 $X2=4.89 $Y2=1.52
r242 62 64 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.205 $Y=2.67
+ $X2=3.205 $Y2=2.8
r243 58 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.14 $Y=2.63
+ $X2=2.14 $Y2=2.8
r244 55 57 6.14986 $w=3.67e-07 $l=1.85e-07 $layer=LI1_cond $X=1.222 $Y=2.63
+ $X2=1.222 $Y2=2.815
r245 54 84 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.635 $Y=1.65
+ $X2=1.635 $Y2=1.74
r246 54 83 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.65
+ $X2=1.635 $Y2=1.485
r247 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.65 $X2=1.635 $Y2=1.65
r248 51 53 7.39941 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=1.43 $Y=1.756
+ $X2=1.635 $Y2=1.756
r249 50 51 9.20414 $w=3.38e-07 $l=3.51312e-07 $layer=LI1_cond $X=1.175 $Y=1.985
+ $X2=1.43 $Y2=1.756
r250 48 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.905 $Y=2.905
+ $X2=5.905 $Y2=1.945
r251 46 76 4.10697 $w=2.22e-07 $l=1.08305e-07 $layer=LI1_cond $X=5.15 $Y=2.99
+ $X2=5.065 $Y2=2.937
r252 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.82 $Y=2.99
+ $X2=5.905 $Y2=2.905
r253 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.82 $Y=2.99
+ $X2=5.15 $Y2=2.99
r254 44 76 2.32734 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=5.065 $Y=2.8
+ $X2=5.065 $Y2=2.937
r255 43 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=1.685
+ $X2=5.065 $Y2=1.52
r256 43 44 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.065 $Y=1.685
+ $X2=5.065 $Y2=2.8
r257 42 66 17.4193 $w=1.68e-07 $l=2.67e-07 $layer=LI1_cond $X=4.385 $Y=2.937
+ $X2=4.385 $Y2=2.67
r258 41 76 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.937
+ $X2=5.065 $Y2=2.937
r259 41 42 21.3726 $w=2.73e-07 $l=5.1e-07 $layer=LI1_cond $X=4.98 $Y=2.937
+ $X2=4.47 $Y2=2.937
r260 40 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=2.67
+ $X2=3.205 $Y2=2.67
r261 39 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=2.67
+ $X2=4.385 $Y2=2.67
r262 39 40 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.3 $Y=2.67
+ $X2=3.29 $Y2=2.67
r263 38 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.8
+ $X2=2.14 $Y2=2.8
r264 37 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.8
+ $X2=3.205 $Y2=2.8
r265 37 38 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.12 $Y=2.8
+ $X2=2.225 $Y2=2.8
r266 36 55 5.25812 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=1.435 $Y=2.63
+ $X2=1.222 $Y2=2.63
r267 35 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.63
+ $X2=2.14 $Y2=2.63
r268 35 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.055 $Y=2.63
+ $X2=1.435 $Y2=2.63
r269 31 51 0.862142 $w=3.3e-07 $l=2.71e-07 $layer=LI1_cond $X=1.43 $Y=1.485
+ $X2=1.43 $Y2=1.756
r270 31 33 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.43 $Y=1.485
+ $X2=1.43 $Y2=1.155
r271 30 55 2.70071 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.222 $Y=2.545
+ $X2=1.222 $Y2=2.63
r272 30 50 14.0462 $w=4.23e-07 $l=5.18e-07 $layer=LI1_cond $X=1.222 $Y=2.545
+ $X2=1.222 $Y2=2.027
r273 25 89 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.945
+ $X2=5.715 $Y2=1.78
r274 25 27 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.715 $Y=1.945
+ $X2=5.715 $Y2=2.62
r275 23 87 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.95 $Y=0.875
+ $X2=4.95 $Y2=1.355
r276 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.49 $Y=0.255
+ $X2=3.49 $Y2=0.72
r277 13 15 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.64 $Y=1.815
+ $X2=2.64 $Y2=2.445
r278 12 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.74
+ $X2=1.635 $Y2=1.74
r279 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.55 $Y=1.74
+ $X2=2.64 $Y2=1.815
r280 11 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.55 $Y=1.74
+ $X2=1.8 $Y2=1.74
r281 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.415 $Y=0.18
+ $X2=3.49 $Y2=0.255
r282 9 10 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=3.415 $Y=0.18
+ $X2=1.8 $Y2=0.18
r283 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.725 $Y=0.255
+ $X2=1.8 $Y2=0.18
r284 7 83 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.725 $Y=0.255
+ $X2=1.725 $Y2=1.485
r285 2 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.84 $X2=1.175 $Y2=2.815
r286 2 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.84 $X2=1.175 $Y2=1.985
r287 1 33 182 $w=1.7e-07 $l=8.88214e-07 $layer=licon1_NDIFF $count=1 $X=1.21
+ $Y=0.37 $X2=1.43 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_701_463# 1 2 7 9 11 12 14 17 19 25 28 32
+ 34 37 40
c89 34 0 1.27123e-19 $X=4.45 $Y=1.015
c90 28 0 1.76992e-19 $X=4.735 $Y=1.005
c91 19 0 4.21193e-20 $X=4.45 $Y=1.192
r92 35 37 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.535 $Y=1.94
+ $X2=4.725 $Y2=1.94
r93 30 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.725 $Y=2.025
+ $X2=4.725 $Y2=1.94
r94 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.725 $Y=2.025
+ $X2=4.725 $Y2=2.42
r95 26 34 3.05675 $w=3.1e-07 $l=1.8759e-07 $layer=LI1_cond $X=4.62 $Y=1.052
+ $X2=4.45 $Y2=1.015
r96 26 28 5.00117 $w=2.63e-07 $l=1.15e-07 $layer=LI1_cond $X=4.62 $Y=1.052
+ $X2=4.735 $Y2=1.052
r97 25 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=1.855
+ $X2=4.535 $Y2=1.94
r98 24 34 3.57226 $w=1.7e-07 $l=3.95221e-07 $layer=LI1_cond $X=4.535 $Y=1.37
+ $X2=4.45 $Y2=1.015
r99 24 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.535 $Y=1.37
+ $X2=4.535 $Y2=1.855
r100 22 40 20.6994 $w=3.26e-07 $l=1.4e-07 $layer=POLY_cond $X=3.99 $Y=1.23
+ $X2=3.85 $Y2=1.23
r101 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.99
+ $Y=1.205 $X2=3.99 $Y2=1.205
r102 19 34 3.05675 $w=3.1e-07 $l=1.77e-07 $layer=LI1_cond $X=4.45 $Y=1.192
+ $X2=4.45 $Y2=1.015
r103 19 21 14.9331 $w=3.53e-07 $l=4.6e-07 $layer=LI1_cond $X=4.45 $Y=1.192
+ $X2=3.99 $Y2=1.192
r104 12 40 20.933 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.85 $Y=1.04
+ $X2=3.85 $Y2=1.23
r105 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.85 $Y=1.04
+ $X2=3.85 $Y2=0.72
r106 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.735 $Y=2.315
+ $X2=3.735 $Y2=2.39
r107 10 40 17.0031 $w=3.26e-07 $l=2.40728e-07 $layer=POLY_cond $X=3.735 $Y=1.42
+ $X2=3.85 $Y2=1.23
r108 10 11 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=3.735 $Y=1.42
+ $X2=3.735 $Y2=2.315
r109 7 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.595 $Y=2.39
+ $X2=3.735 $Y2=2.39
r110 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.595 $Y=2.465
+ $X2=3.595 $Y2=2.75
r111 2 32 600 $w=1.7e-07 $l=3.91152e-07 $layer=licon1_PDIFF $count=1 $X=4.515
+ $Y=2.12 $X2=4.725 $Y2=2.42
r112 1 28 182 $w=1.7e-07 $l=7.26722e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.38 $X2=4.735 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_546_447# 1 2 9 13 16 17 19 21 25 37
c88 21 0 1.35673e-19 $X=3.23 $Y=0.77
r89 36 37 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.425 $Y=1.795
+ $X2=4.44 $Y2=1.795
r90 26 36 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=4.185 $Y=1.795
+ $X2=4.425 $Y2=1.795
r91 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.795 $X2=4.185 $Y2=1.795
r92 23 25 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=4.15 $Y=2.245
+ $X2=4.15 $Y2=1.795
r93 19 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.19 $Y=1.495
+ $X2=2.865 $Y2=1.495
r94 19 21 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=3.19 $Y=1.41
+ $X2=3.19 $Y2=0.77
r95 18 33 3.40825 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.95 $Y=2.33
+ $X2=2.865 $Y2=2.395
r96 17 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.02 $Y=2.33
+ $X2=4.15 $Y2=2.245
r97 17 18 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.02 $Y=2.33
+ $X2=2.95 $Y2=2.33
r98 16 33 3.40825 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.865 $Y=2.245
+ $X2=2.865 $Y2=2.395
r99 15 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.58
+ $X2=2.865 $Y2=1.495
r100 15 16 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.865 $Y=1.58
+ $X2=2.865 $Y2=2.245
r101 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.44 $Y=1.63
+ $X2=4.44 $Y2=1.795
r102 11 13 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=4.44 $Y=1.63
+ $X2=4.44 $Y2=0.655
r103 7 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.96
+ $X2=4.425 $Y2=1.795
r104 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.425 $Y=1.96
+ $X2=4.425 $Y2=2.54
r105 2 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.235 $X2=2.865 $Y2=2.38
r106 1 21 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.09
+ $Y=0.595 $X2=3.23 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_1191_120# 1 2 7 9 10 12 17 21 23 27 31 35
+ 40 43 44 47 51 53 54 55 56 61 65 66 67
c142 66 0 3.58297e-19 $X=7.565 $Y=1.515
c143 35 0 4.23824e-20 $X=6.305 $Y=1.3
c144 7 0 1.54211e-19 $X=6.03 $Y=1.225
r145 65 68 6.96826 $w=4.28e-07 $l=2.6e-07 $layer=LI1_cond $X=7.515 $Y=1.515
+ $X2=7.515 $Y2=1.775
r146 65 67 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.515 $Y=1.515
+ $X2=7.515 $Y2=1.35
r147 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.565
+ $Y=1.515 $X2=7.565 $Y2=1.515
r148 60 63 9.97615 $w=5.87e-07 $l=4.8e-07 $layer=LI1_cond $X=6.395 $Y=1.885
+ $X2=6.875 $Y2=1.885
r149 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.395
+ $Y=1.715 $X2=6.395 $Y2=1.715
r150 57 67 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.385 $Y=1.02
+ $X2=7.385 $Y2=1.35
r151 56 63 10.2728 $w=5.87e-07 $l=2.13014e-07 $layer=LI1_cond $X=7.04 $Y=1.775
+ $X2=6.875 $Y2=1.885
r152 55 68 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=7.3 $Y=1.775
+ $X2=7.515 $Y2=1.775
r153 55 56 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.3 $Y=1.775
+ $X2=7.04 $Y2=1.775
r154 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=0.935
+ $X2=7.385 $Y2=1.02
r155 53 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.3 $Y=0.935
+ $X2=6.97 $Y2=0.935
r156 49 63 4.10774 $w=3.3e-07 $l=3.35e-07 $layer=LI1_cond $X=6.875 $Y=2.22
+ $X2=6.875 $Y2=1.885
r157 49 51 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=6.875 $Y=2.22
+ $X2=6.875 $Y2=2.695
r158 45 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.805 $Y=0.85
+ $X2=6.97 $Y2=0.935
r159 45 47 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.805 $Y=0.85
+ $X2=6.805 $Y2=0.645
r160 43 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.395 $Y=1.55
+ $X2=6.395 $Y2=1.715
r161 40 61 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=6.395 $Y=2.185
+ $X2=6.395 $Y2=1.715
r162 33 35 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=6.03 $Y=1.3
+ $X2=6.305 $Y2=1.3
r163 29 44 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=8.595 $Y=1.68
+ $X2=8.505 $Y2=1.35
r164 29 31 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=8.595 $Y=1.68
+ $X2=8.595 $Y2=2.26
r165 25 44 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.58 $Y=1.35
+ $X2=8.505 $Y2=1.35
r166 25 27 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=8.58 $Y=1.35
+ $X2=8.58 $Y2=0.835
r167 24 66 3.90195 $w=3.3e-07 $l=1.48e-07 $layer=POLY_cond $X=7.695 $Y=1.515
+ $X2=7.547 $Y2=1.515
r168 23 44 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.505 $Y=1.515
+ $X2=8.505 $Y2=1.35
r169 23 24 141.638 $w=3.3e-07 $l=8.1e-07 $layer=POLY_cond $X=8.505 $Y=1.515
+ $X2=7.695 $Y2=1.515
r170 19 66 34.7346 $w=1.65e-07 $l=1.9182e-07 $layer=POLY_cond $X=7.605 $Y=1.68
+ $X2=7.547 $Y2=1.515
r171 19 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.605 $Y=1.68
+ $X2=7.605 $Y2=2.4
r172 15 66 34.7346 $w=1.65e-07 $l=1.85257e-07 $layer=POLY_cond $X=7.59 $Y=1.35
+ $X2=7.547 $Y2=1.515
r173 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.59 $Y=1.35
+ $X2=7.59 $Y2=0.74
r174 13 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.305 $Y=1.375
+ $X2=6.305 $Y2=1.3
r175 13 43 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.305 $Y=1.375
+ $X2=6.305 $Y2=1.55
r176 10 40 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.105 $Y=2.26
+ $X2=6.395 $Y2=2.26
r177 10 12 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.105 $Y=2.335
+ $X2=6.105 $Y2=2.62
r178 7 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.03 $Y=1.225
+ $X2=6.03 $Y2=1.3
r179 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.03 $Y=1.225 $X2=6.03
+ $Y2=0.94
r180 2 63 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.875 $Y2=1.985
r181 2 51 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.875 $Y2=2.695
r182 1 47 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.66
+ $Y=0.37 $X2=6.805 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_1005_120# 1 2 9 11 13 15 17 19 26 28 30
c83 28 0 2.55347e-19 $X=6.965 $Y=1.355
c84 15 0 5.7879e-20 $X=5.405 $Y=1.38
c85 9 0 2.43826e-20 $X=7.02 $Y=0.645
r86 28 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.965 $Y=1.355
+ $X2=6.8 $Y2=1.355
r87 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.965
+ $Y=1.355 $X2=6.965 $Y2=1.355
r88 24 25 10.9446 $w=3.79e-07 $l=3.4e-07 $layer=LI1_cond $X=5.357 $Y=0.955
+ $X2=5.357 $Y2=1.295
r89 22 25 5.45184 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=5.357 $Y2=1.295
r90 22 30 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=6.8 $Y2=1.295
r91 17 26 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.445 $Y=2.24
+ $X2=5.445 $Y2=2.115
r92 17 19 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.445 $Y=2.24
+ $X2=5.445 $Y2=2.545
r93 15 25 6.49482 $w=3.79e-07 $l=1.06325e-07 $layer=LI1_cond $X=5.405 $Y=1.38
+ $X2=5.357 $Y2=1.295
r94 15 26 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.405 $Y=1.38
+ $X2=5.405 $Y2=2.115
r95 11 29 47.5149 $w=3.21e-07 $l=3.02985e-07 $layer=POLY_cond $X=7.1 $Y=1.61
+ $X2=6.995 $Y2=1.355
r96 11 13 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=7.1 $Y=1.61 $X2=7.1
+ $Y2=2.34
r97 7 29 38.5532 $w=3.21e-07 $l=1.77059e-07 $layer=POLY_cond $X=7.02 $Y=1.19
+ $X2=6.995 $Y2=1.355
r98 7 9 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.02 $Y=1.19 $X2=7.02
+ $Y2=0.645
r99 2 19 600 $w=1.7e-07 $l=4.87852e-07 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=2.12 $X2=5.405 $Y2=2.545
r100 1 24 182 $w=1.7e-07 $l=4.69148e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.6 $X2=5.29 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_1644_112# 1 2 9 13 17 21 25 26 28
r53 26 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.465
+ $X2=9.06 $Y2=1.63
r54 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.465
+ $X2=9.06 $Y2=1.3
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.06
+ $Y=1.465 $X2=9.06 $Y2=1.465
r56 23 28 0.182887 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=8.53 $Y=1.465
+ $X2=8.405 $Y2=1.465
r57 23 25 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.53 $Y=1.465
+ $X2=9.06 $Y2=1.465
r58 19 28 7.32358 $w=2.12e-07 $l=1.83016e-07 $layer=LI1_cond $X=8.367 $Y=1.63
+ $X2=8.405 $Y2=1.465
r59 19 21 22.4987 $w=1.73e-07 $l=3.55e-07 $layer=LI1_cond $X=8.367 $Y=1.63
+ $X2=8.367 $Y2=1.985
r60 15 28 7.32358 $w=2.12e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=1.3
+ $X2=8.405 $Y2=1.465
r61 15 17 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.405 $Y=1.3
+ $X2=8.405 $Y2=0.835
r62 13 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.09 $Y=0.74
+ $X2=9.09 $Y2=1.3
r63 9 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=9.1 $Y=2.4 $X2=9.1
+ $Y2=1.63
r64 2 21 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.235
+ $Y=1.84 $X2=8.37 $Y2=1.985
r65 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.56 $X2=8.365 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 40 41 42 44
+ 49 54 66 70 77 78 81 84 87 94 97
c120 21 0 2.50478e-20 $X=0.725 $Y=2.225
r121 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 87 90 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=3.935 $Y=3.01
+ $X2=3.935 $Y2=3.33
r125 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r126 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 78 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r129 75 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=8.82 $Y2=3.33
r130 75 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=9.36 $Y2=3.33
r131 74 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 74 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r134 71 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.49 $Y=3.33
+ $X2=7.365 $Y2=3.33
r135 71 73 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=7.49 $Y=3.33 $X2=8.4
+ $Y2=3.33
r136 70 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.655 $Y=3.33
+ $X2=8.82 $Y2=3.33
r137 70 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.655 $Y=3.33
+ $X2=8.4 $Y2=3.33
r138 69 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r139 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r140 66 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=7.365 $Y2=3.33
r141 66 68 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r142 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r143 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r144 62 90 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=3.935 $Y2=3.33
r145 62 64 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=4.13 $Y=3.33 $X2=6
+ $Y2=3.33
r146 61 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r147 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 58 61 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 57 60 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r151 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 55 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.72 $Y2=3.33
r153 55 57 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.16 $Y2=3.33
r154 54 90 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.74 $Y=3.33
+ $X2=3.935 $Y2=3.33
r155 54 60 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.74 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 53 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r157 53 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r158 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r159 50 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=0.685 $Y2=3.33
r160 50 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=1.2 $Y2=3.33
r161 49 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.72 $Y2=3.33
r162 49 52 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 47 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r165 44 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.685 $Y2=3.33
r166 44 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r167 42 65 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=3.33 $X2=6
+ $Y2=3.33
r168 42 91 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 40 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6 $Y2=3.33
r170 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.33 $Y2=3.33
r171 39 68 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.96 $Y2=3.33
r172 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.33 $Y2=3.33
r173 35 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=3.33
r174 35 37 44.0024 $w=3.28e-07 $l=1.26e-06 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=1.985
r175 31 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.365 $Y=3.245
+ $X2=7.365 $Y2=3.33
r176 31 33 48.4026 $w=2.48e-07 $l=1.05e-06 $layer=LI1_cond $X=7.365 $Y=3.245
+ $X2=7.365 $Y2=2.195
r177 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=3.33
r178 27 29 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=2.62
r179 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.33
r180 23 25 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.05
r181 19 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=3.245
+ $X2=0.685 $Y2=3.33
r182 19 21 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.685 $Y=3.245
+ $X2=0.685 $Y2=2.225
r183 6 37 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.685
+ $Y=1.84 $X2=8.82 $Y2=1.985
r184 5 33 300 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_PDIFF $count=2 $X=7.19
+ $Y=1.84 $X2=7.325 $Y2=2.195
r185 4 29 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=6.195
+ $Y=2.41 $X2=6.33 $Y2=2.62
r186 3 87 600 $w=1.7e-07 $l=5.81722e-07 $layer=licon1_PDIFF $count=1 $X=3.685
+ $Y=2.54 $X2=3.935 $Y2=3.01
r187 2 25 600 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=2.515 $X2=1.72 $Y2=3.05
r188 1 21 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.84 $X2=0.725 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%A_423_503# 1 2 8 11 16 20
c39 16 0 1.54739e-19 $X=2.525 $Y=2.21
c40 8 0 1.68603e-19 $X=2.525 $Y=2.045
r41 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.525 $Y=1.155
+ $X2=2.8 $Y2=1.155
r42 14 16 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.335 $Y=2.21
+ $X2=2.525 $Y2=2.21
r43 9 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=1.07 $X2=2.8
+ $Y2=1.155
r44 9 11 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.8 $Y=1.07 $X2=2.8
+ $Y2=0.815
r45 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.045
+ $X2=2.525 $Y2=2.21
r46 7 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.24
+ $X2=2.525 $Y2=1.155
r47 7 8 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.525 $Y=1.24
+ $X2=2.525 $Y2=2.045
r48 2 14 600 $w=1.7e-07 $l=4.00156e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=2.515 $X2=2.335 $Y2=2.21
r49 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.595 $X2=2.8 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%Q 1 2 9 13 16 17 18 19
c35 13 0 2.43826e-20 $X=7.855 $Y=1.13
r36 18 19 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=7.867 $Y=2.405
+ $X2=7.867 $Y2=2.775
r37 16 17 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.867 $Y=2.195
+ $X2=7.867 $Y2=2.03
r38 14 18 4.92278 $w=4.03e-07 $l=1.73e-07 $layer=LI1_cond $X=7.867 $Y=2.232
+ $X2=7.867 $Y2=2.405
r39 14 16 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=7.867 $Y=2.232
+ $X2=7.867 $Y2=2.195
r40 13 17 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.985 $Y=1.13
+ $X2=7.985 $Y2=2.03
r41 7 13 10.1249 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.855 $Y=0.915
+ $X2=7.855 $Y2=1.13
r42 7 9 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=7.855 $Y=0.915 $X2=7.855
+ $Y2=0.515
r43 2 16 300 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_PDIFF $count=2 $X=7.695
+ $Y=1.84 $X2=7.83 $Y2=2.195
r44 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.665
+ $Y=0.37 $X2=7.805 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%Q_N 1 2 9 13 14 15 16 23 32
r25 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=9.337 $Y=1.997
+ $X2=9.337 $Y2=2.035
r26 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=9.337 $Y=2.405
+ $X2=9.337 $Y2=2.775
r27 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=9.337 $Y=1.973
+ $X2=9.337 $Y2=1.997
r28 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=9.337 $Y=1.973
+ $X2=9.337 $Y2=1.82
r29 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=9.337 $Y=2.058
+ $X2=9.337 $Y2=2.405
r30 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=9.337 $Y=2.058
+ $X2=9.337 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.43 $Y=1.13 $X2=9.43
+ $Y2=1.82
r32 7 13 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=9.327 $Y=0.943
+ $X2=9.327 $Y2=1.13
r33 7 9 13.1532 $w=3.73e-07 $l=4.28e-07 $layer=LI1_cond $X=9.327 $Y=0.943
+ $X2=9.327 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.84 $X2=9.325 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.84 $X2=9.325 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.165
+ $Y=0.37 $X2=9.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 42 43 45 46
+ 47 49 54 59 71 80 81 84 87 91 97
c120 33 0 1.91441e-19 $X=7.305 $Y=0.515
r121 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r122 91 94 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.145 $Y=0
+ $X2=4.145 $Y2=0.325
r123 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r124 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r125 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r127 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r128 78 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r129 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r130 75 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=7.305
+ $Y2=0
r131 75 77 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=8.4
+ $Y2=0
r132 74 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r133 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r134 71 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=7.305
+ $Y2=0
r135 71 73 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.14 $Y=0 $X2=6.96
+ $Y2=0
r136 70 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r137 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r138 67 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r139 66 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r140 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r141 64 91 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.145
+ $Y2=0
r142 64 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.56
+ $Y2=0
r143 63 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r144 63 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r145 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 60 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.03
+ $Y2=0
r147 60 62 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=3.6 $Y2=0
r148 59 91 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=4.145
+ $Y2=0
r149 59 62 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=3.6
+ $Y2=0
r150 58 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r151 58 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r152 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r153 55 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.815
+ $Y2=0
r154 55 57 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=1.68 $Y2=0
r155 54 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.03
+ $Y2=0
r156 54 57 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.68 $Y2=0
r157 52 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r158 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r159 49 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.815
+ $Y2=0
r160 49 51 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r161 47 70 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6
+ $Y2=0
r162 47 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r163 45 77 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.71 $Y=0 $X2=8.4
+ $Y2=0
r164 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.71 $Y=0 $X2=8.835
+ $Y2=0
r165 44 80 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.96 $Y=0 $X2=9.36
+ $Y2=0
r166 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.96 $Y=0 $X2=8.835
+ $Y2=0
r167 42 69 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.08 $Y=0 $X2=6 $Y2=0
r168 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=6.245
+ $Y2=0
r169 41 73 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.96
+ $Y2=0
r170 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.41 $Y=0 $X2=6.245
+ $Y2=0
r171 37 39 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=8.835 $Y=0.515
+ $X2=8.835 $Y2=0.965
r172 35 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=0.085
+ $X2=8.835 $Y2=0
r173 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.835 $Y=0.085
+ $X2=8.835 $Y2=0.515
r174 31 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0
r175 31 33 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0.515
r176 27 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0
r177 27 29 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0.875
r178 23 87 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r179 23 25 12.8415 $w=3.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.475
r180 19 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r181 19 21 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.395
r182 6 39 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=8.655
+ $Y=0.56 $X2=8.875 $Y2=0.965
r183 6 37 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=8.655
+ $Y=0.56 $X2=8.875 $Y2=0.515
r184 5 33 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.095
+ $Y=0.37 $X2=7.305 $Y2=0.515
r185 4 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.73 $X2=6.245 $Y2=0.875
r186 3 94 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=3.925
+ $Y=0.51 $X2=4.145 $Y2=0.325
r187 2 25 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.33 $X2=2.03 $Y2=0.475
r188 1 21 182 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.815 $Y2=0.395
.ends


* NGSPICE file created from sky130_fd_sc_ms__dlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_83_244# a_315_338# a_267_392# VPB pshort w=1e+06u l=180000u
+  ad=4.054e+11p pd=3.24e+06u as=2.4e+11p ps=2.48e+06u
M1001 a_1044_387# CLK VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=2.5157e+12p ps=1.567e+07u
M1002 a_511_508# a_315_48# a_83_244# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1003 GCLK a_1044_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.45355e+12p ps=1.19e+07u
M1004 VPWR a_83_244# a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1005 VPWR a_27_74# a_1044_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_27_74# a_511_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_494_118# a_315_338# a_83_244# VNB nlowvt w=420000u l=150000u
+  ad=1.54875e+11p pd=1.7e+06u as=3.049e+11p ps=2.47e+06u
M1008 a_315_338# a_315_48# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1009 VGND a_1044_387# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_74# a_494_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_315_338# a_315_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 VPWR CLK a_315_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.52e+11p ps=2.28e+06u
M1013 a_83_244# a_315_48# a_267_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1014 a_267_74# GATE VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND CLK a_315_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 GCLK a_1044_387# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1017 a_1044_387# a_27_74# a_1044_119# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.554e+11p ps=1.9e+06u
M1018 VPWR a_1044_387# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1044_119# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_267_392# GATE VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_83_244# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends


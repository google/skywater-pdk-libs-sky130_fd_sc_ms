* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and2b_4 A_N B VGND VNB VPB VPWR X
X0 VPWR a_221_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_233_74# a_27_392# a_221_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VPWR a_221_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 X a_221_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_27_392# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VGND B a_233_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR a_27_392# a_221_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X7 VPWR B a_221_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 a_233_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_27_392# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 X a_221_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 X a_221_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 VGND a_221_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 X a_221_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_221_424# a_27_392# a_233_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_221_424# a_27_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X16 a_221_424# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X17 VGND a_221_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

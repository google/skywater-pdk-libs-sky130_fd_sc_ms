* File: sky130_fd_sc_ms__o221a_1.pxi.spice
* Created: Wed Sep  2 12:22:50 2020
* 
x_PM_SKY130_FD_SC_MS__O221A_1%A_83_264# N_A_83_264#_M1006_d N_A_83_264#_M1002_d
+ N_A_83_264#_M1009_d N_A_83_264#_M1007_g N_A_83_264#_M1004_g N_A_83_264#_c_85_n
+ N_A_83_264#_c_86_n N_A_83_264#_c_145_p N_A_83_264#_c_87_n N_A_83_264#_c_114_p
+ N_A_83_264#_c_88_n N_A_83_264#_c_80_n N_A_83_264#_c_81_n N_A_83_264#_c_82_n
+ N_A_83_264#_c_90_n N_A_83_264#_c_83_n N_A_83_264#_c_91_n
+ PM_SKY130_FD_SC_MS__O221A_1%A_83_264#
x_PM_SKY130_FD_SC_MS__O221A_1%A1 N_A1_M1003_g N_A1_M1010_g A1 N_A1_c_176_n
+ PM_SKY130_FD_SC_MS__O221A_1%A1
x_PM_SKY130_FD_SC_MS__O221A_1%A2 N_A2_M1000_g N_A2_M1002_g A2 N_A2_c_215_n
+ PM_SKY130_FD_SC_MS__O221A_1%A2
x_PM_SKY130_FD_SC_MS__O221A_1%B2 N_B2_M1011_g N_B2_c_248_n N_B2_c_249_n
+ N_B2_c_250_n N_B2_M1001_g B2 N_B2_c_252_n N_B2_c_253_n
+ PM_SKY130_FD_SC_MS__O221A_1%B2
x_PM_SKY130_FD_SC_MS__O221A_1%B1 N_B1_M1005_g N_B1_M1008_g B1 N_B1_c_294_n
+ PM_SKY130_FD_SC_MS__O221A_1%B1
x_PM_SKY130_FD_SC_MS__O221A_1%C1 N_C1_c_328_n N_C1_M1006_g N_C1_M1009_g
+ N_C1_c_329_n C1 C1 N_C1_c_331_n N_C1_c_332_n PM_SKY130_FD_SC_MS__O221A_1%C1
x_PM_SKY130_FD_SC_MS__O221A_1%X N_X_M1004_s N_X_M1007_s N_X_c_368_n N_X_c_369_n
+ N_X_c_365_n X X N_X_c_367_n X PM_SKY130_FD_SC_MS__O221A_1%X
x_PM_SKY130_FD_SC_MS__O221A_1%VPWR N_VPWR_M1007_d N_VPWR_M1005_d N_VPWR_c_389_n
+ N_VPWR_c_390_n VPWR N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_388_n
+ N_VPWR_c_394_n N_VPWR_c_395_n PM_SKY130_FD_SC_MS__O221A_1%VPWR
x_PM_SKY130_FD_SC_MS__O221A_1%VGND N_VGND_M1004_d N_VGND_M1000_d N_VGND_c_432_n
+ N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n VGND N_VGND_c_436_n
+ N_VGND_c_437_n N_VGND_c_438_n PM_SKY130_FD_SC_MS__O221A_1%VGND
x_PM_SKY130_FD_SC_MS__O221A_1%A_245_94# N_A_245_94#_M1003_d N_A_245_94#_M1001_d
+ N_A_245_94#_c_476_n N_A_245_94#_c_477_n N_A_245_94#_c_478_n
+ N_A_245_94#_c_495_n PM_SKY130_FD_SC_MS__O221A_1%A_245_94#
x_PM_SKY130_FD_SC_MS__O221A_1%A_456_74# N_A_456_74#_M1001_s N_A_456_74#_M1008_d
+ N_A_456_74#_c_512_n N_A_456_74#_c_513_n N_A_456_74#_c_514_n
+ N_A_456_74#_c_522_n PM_SKY130_FD_SC_MS__O221A_1%A_456_74#
cc_1 VNB N_A_83_264#_M1007_g 5.80156e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_264#_M1004_g 0.0301825f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_3 VNB N_A_83_264#_c_80_n 0.0333404f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.96
cc_4 VNB N_A_83_264#_c_81_n 0.00390048f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.485
cc_5 VNB N_A_83_264#_c_82_n 0.0384287f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.485
cc_6 VNB N_A_83_264#_c_83_n 0.0271336f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=0.525
cc_7 VNB N_A1_M1003_g 0.0313341f $X=-0.19 $Y=-0.245 $X2=3.905 $Y2=1.96
cc_8 VNB A1 0.00325184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_c_176_n 0.0198088f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_10 VNB N_A2_M1000_g 0.0316315f $X=-0.19 $Y=-0.245 $X2=3.905 $Y2=1.96
cc_11 VNB A2 0.00299813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_215_n 0.0166132f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_13 VNB N_B2_c_248_n 0.0194238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B2_c_249_n 0.0199768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_250_n 0.0194669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B2 0.00444804f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_17 VNB N_B2_c_252_n 0.0282098f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_18 VNB N_B2_c_253_n 0.00280391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_M1008_g 0.0359828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.00248798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_294_n 0.0262171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C1_c_328_n 0.0206367f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=1.96
cc_23 VNB N_C1_c_329_n 0.00594779f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_24 VNB C1 0.00795525f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_25 VNB N_C1_c_331_n 0.0237545f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_26 VNB N_C1_c_332_n 0.0218548f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.65
cc_27 VNB N_X_c_365_n 0.0249958f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.74
cc_28 VNB X 0.0145164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_367_n 0.0273847f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.815
cc_30 VNB N_VPWR_c_388_n 0.183584f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.815
cc_31 VNB N_VGND_c_432_n 0.0236354f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_32 VNB N_VGND_c_433_n 0.016373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_434_n 0.01947f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.035
cc_34 VNB N_VGND_c_435_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_35 VNB N_VGND_c_436_n 0.0587016f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=0.95
cc_36 VNB N_VGND_c_437_n 0.267882f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.96
cc_37 VNB N_VGND_c_438_n 0.0272997f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.485
cc_38 VNB N_A_245_94#_c_476_n 0.00327588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_245_94#_c_477_n 0.0216121f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_40 VNB N_A_245_94#_c_478_n 0.00406832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_41 VNB N_A_456_74#_c_512_n 0.00465728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_456_74#_c_513_n 0.00490525f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_43 VNB N_A_456_74#_c_514_n 0.00489174f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_44 VPB N_A_83_264#_M1007_g 0.0310437f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_45 VPB N_A_83_264#_c_85_n 0.00289574f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_46 VPB N_A_83_264#_c_86_n 0.010377f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=2.035
cc_47 VPB N_A_83_264#_c_87_n 0.00285226f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=2.815
cc_48 VPB N_A_83_264#_c_88_n 0.0348765f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.815
cc_49 VPB N_A_83_264#_c_80_n 0.0140682f $X=-0.19 $Y=1.66 $X2=4.12 $Y2=1.96
cc_50 VPB N_A_83_264#_c_90_n 0.00363208f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=2.115
cc_51 VPB N_A_83_264#_c_91_n 0.0100225f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.125
cc_52 VPB N_A1_M1010_g 0.0257216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB A1 0.00138199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A1_c_176_n 0.0134373f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_55 VPB N_A2_M1002_g 0.0243062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB A2 0.00174709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A2_c_215_n 0.0105862f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_58 VPB N_B2_M1011_g 0.0262234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB B2 0.00311741f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_60 VPB N_B2_c_253_n 0.0108889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_B1_M1005_g 0.0302616f $X=-0.19 $Y=1.66 $X2=3.905 $Y2=1.96
cc_62 VPB B1 0.00304223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B1_c_294_n 0.0214588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_C1_M1009_g 0.0334843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_C1_c_329_n 0.0168738f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_66 VPB C1 0.00314059f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_67 VPB N_X_c_368_n 0.0116338f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_68 VPB N_X_c_369_n 0.0403824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_X_c_365_n 0.00728828f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.74
cc_70 VPB N_VPWR_c_389_n 0.0105243f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_71 VPB N_VPWR_c_390_n 0.0118351f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=0.74
cc_72 VPB N_VPWR_c_391_n 0.0546548f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_73 VPB N_VPWR_c_392_n 0.0191515f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.815
cc_74 VPB N_VPWR_c_388_n 0.0895845f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.815
cc_75 VPB N_VPWR_c_394_n 0.0285033f $X=-0.19 $Y=1.66 $X2=4.12 $Y2=1.96
cc_76 VPB N_VPWR_c_395_n 0.0159371f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.485
cc_77 N_A_83_264#_M1004_g N_A1_M1003_g 0.0202137f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A_83_264#_c_81_n N_A1_M1003_g 8.05667e-19 $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_79 N_A_83_264#_c_82_n N_A1_M1003_g 0.00601582f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_80 N_A_83_264#_M1007_g N_A1_M1010_g 0.0192758f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A_83_264#_c_85_n N_A1_M1010_g 0.0031117f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_82 N_A_83_264#_c_86_n N_A1_M1010_g 0.018003f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_83 N_A_83_264#_c_87_n N_A1_M1010_g 0.0028279f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_84 N_A_83_264#_c_86_n A1 0.0241033f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_83_264#_c_81_n A1 0.0202352f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_86 N_A_83_264#_c_82_n A1 7.26157e-19 $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_87 N_A_83_264#_M1007_g N_A1_c_176_n 0.00285059f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_83_264#_c_85_n N_A1_c_176_n 9.8453e-19 $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_89 N_A_83_264#_c_86_n N_A1_c_176_n 0.00104284f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A_83_264#_c_81_n N_A1_c_176_n 7.10742e-19 $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_82_n N_A1_c_176_n 0.011617f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_86_n N_A2_M1002_g 0.0127019f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_83_264#_c_87_n N_A2_M1002_g 0.0175268f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_94 N_A_83_264#_c_90_n N_A2_M1002_g 0.0012159f $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_95 N_A_83_264#_c_86_n A2 0.0114708f $X=1.725 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_83_264#_c_90_n A2 0.0150447f $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_97 N_A_83_264#_c_90_n N_A2_c_215_n 0.00349435f $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_98 N_A_83_264#_c_87_n N_B2_M1011_g 0.0233307f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_114_p N_B2_M1011_g 0.0184144f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_90_n N_B2_M1011_g 3.18422e-19 $X=1.89 $Y=2.115 $X2=0 $Y2=0
cc_101 N_A_83_264#_c_114_p B2 0.0395872f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_114_p N_B2_c_253_n 0.00375045f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_103 N_A_83_264#_c_114_p N_B1_M1005_g 0.0227208f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_104 N_A_83_264#_c_114_p B1 0.0233927f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_114_p N_B1_c_294_n 0.00224137f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_106 N_A_83_264#_c_114_p N_C1_M1009_g 0.016577f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_107 N_A_83_264#_c_88_n N_C1_M1009_g 0.0161131f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_91_n N_C1_M1009_g 0.00196977f $X=4.04 $Y=2.125 $X2=0 $Y2=0
cc_109 N_A_83_264#_c_114_p N_C1_c_329_n 0.00147604f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_110 N_A_83_264#_c_114_p C1 0.0242561f $X=3.875 $Y=2.045 $X2=0 $Y2=0
cc_111 N_A_83_264#_c_80_n C1 0.0429988f $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_112 N_A_83_264#_c_83_n C1 0.00409207f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_80_n N_C1_c_331_n 0.0211211f $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_83_n N_C1_c_331_n 0.00420768f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_80_n N_C1_c_332_n 0.00352354f $X=4.12 $Y=1.96 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_83_n N_C1_c_332_n 0.0114582f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_117 N_A_83_264#_M1007_g N_X_c_368_n 0.00373617f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_85_n N_X_c_368_n 0.00559274f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_119 N_A_83_264#_M1007_g N_X_c_369_n 0.0200238f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_83_264#_M1004_g N_X_c_365_n 0.00457487f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_83_264#_c_85_n N_X_c_365_n 0.0056675f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_122 N_A_83_264#_c_81_n N_X_c_365_n 0.0248004f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_123 N_A_83_264#_c_82_n N_X_c_365_n 0.0106457f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_124 N_A_83_264#_M1004_g X 0.00285885f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_83_264#_c_81_n X 0.00479823f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_126 N_A_83_264#_c_82_n X 0.00224231f $X=0.62 $Y=1.485 $X2=0 $Y2=0
cc_127 N_A_83_264#_M1004_g N_X_c_367_n 0.00787957f $X=0.57 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_85_n N_VPWR_M1007_d 0.00228953f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_83_264#_c_86_n N_VPWR_M1007_d 0.00832454f $X=1.725 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_83_264#_c_145_p N_VPWR_M1007_d 0.0036995f $X=0.785 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_83_264#_c_114_p N_VPWR_M1005_d 0.0246619f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_132 N_A_83_264#_M1007_g N_VPWR_c_389_n 0.0112844f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_83_264#_c_86_n N_VPWR_c_389_n 0.0222558f $X=1.725 $Y=2.035 $X2=0
+ $Y2=0
cc_134 N_A_83_264#_c_145_p N_VPWR_c_389_n 0.00933174f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_135 N_A_83_264#_c_87_n N_VPWR_c_389_n 0.0183098f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_136 N_A_83_264#_c_82_n N_VPWR_c_389_n 3.20969e-19 $X=0.62 $Y=1.485 $X2=0
+ $Y2=0
cc_137 N_A_83_264#_c_114_p N_VPWR_c_390_n 0.0604197f $X=3.875 $Y=2.045 $X2=0
+ $Y2=0
cc_138 N_A_83_264#_c_88_n N_VPWR_c_390_n 0.0263973f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_139 N_A_83_264#_c_87_n N_VPWR_c_391_n 0.014549f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_140 N_A_83_264#_c_88_n N_VPWR_c_392_n 0.014549f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_141 N_A_83_264#_M1007_g N_VPWR_c_388_n 0.00989052f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_83_264#_c_87_n N_VPWR_c_388_n 0.0119743f $X=1.89 $Y=2.815 $X2=0 $Y2=0
cc_143 N_A_83_264#_c_88_n N_VPWR_c_388_n 0.0119743f $X=4.04 $Y=2.815 $X2=0 $Y2=0
cc_144 N_A_83_264#_M1007_g N_VPWR_c_394_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_83_264#_c_86_n A_267_392# 0.0048076f $X=1.725 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_83_264#_c_114_p A_465_392# 0.0136052f $X=3.875 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_83_264#_M1004_g N_VGND_c_432_n 0.00946427f $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_83_264#_c_81_n N_VGND_c_432_n 0.00762027f $X=0.62 $Y=1.485 $X2=0
+ $Y2=0
cc_149 N_A_83_264#_c_82_n N_VGND_c_432_n 7.25643e-19 $X=0.62 $Y=1.485 $X2=0
+ $Y2=0
cc_150 N_A_83_264#_c_83_n N_VGND_c_436_n 0.018459f $X=3.935 $Y=0.525 $X2=0 $Y2=0
cc_151 N_A_83_264#_M1004_g N_VGND_c_437_n 0.00828947f $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_83_264#_c_83_n N_VGND_c_437_n 0.0158482f $X=3.935 $Y=0.525 $X2=0
+ $Y2=0
cc_153 N_A_83_264#_M1004_g N_VGND_c_438_n 0.00434272f $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_83_264#_c_86_n N_A_245_94#_c_477_n 9.96677e-19 $X=1.725 $Y=2.035
+ $X2=0 $Y2=0
cc_155 N_A_83_264#_c_90_n N_A_245_94#_c_477_n 0.00484566f $X=1.89 $Y=2.115 $X2=0
+ $Y2=0
cc_156 N_A_83_264#_M1004_g N_A_245_94#_c_478_n 6.79941e-19 $X=0.57 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A_83_264#_c_86_n N_A_245_94#_c_478_n 0.00632799f $X=1.725 $Y=2.035
+ $X2=0 $Y2=0
cc_158 N_A_83_264#_c_83_n N_A_456_74#_c_513_n 0.00313012f $X=3.935 $Y=0.525
+ $X2=0 $Y2=0
cc_159 N_A1_M1003_g N_A2_M1000_g 0.0248377f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_160 N_A1_M1010_g N_A2_M1002_g 0.0441054f $X=1.245 $Y=2.46 $X2=0 $Y2=0
cc_161 A1 A2 0.020843f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A1_c_176_n A2 0.00200717f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_163 A1 N_A2_c_215_n 4.11485e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A1_c_176_n N_A2_c_215_n 0.0441054f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_165 N_A1_M1010_g N_VPWR_c_389_n 0.0149908f $X=1.245 $Y=2.46 $X2=0 $Y2=0
cc_166 N_A1_M1010_g N_VPWR_c_391_n 0.00553757f $X=1.245 $Y=2.46 $X2=0 $Y2=0
cc_167 N_A1_M1010_g N_VPWR_c_388_n 0.0109174f $X=1.245 $Y=2.46 $X2=0 $Y2=0
cc_168 N_A1_M1003_g N_VGND_c_432_n 0.00744236f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_169 A1 N_VGND_c_432_n 6.86881e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_M1003_g N_VGND_c_433_n 6.44645e-19 $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_171 N_A1_M1003_g N_VGND_c_434_n 0.00485498f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_172 N_A1_M1003_g N_VGND_c_437_n 0.00514438f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_173 N_A1_M1003_g N_A_245_94#_c_476_n 0.00748716f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_174 N_A1_M1003_g N_A_245_94#_c_478_n 0.0062738f $X=1.15 $Y=0.79 $X2=0 $Y2=0
cc_175 A1 N_A_245_94#_c_478_n 0.0112432f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A1_c_176_n N_A_245_94#_c_478_n 8.52409e-19 $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_177 N_A2_M1002_g N_B2_M1011_g 0.0231714f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_178 N_A2_M1000_g N_B2_c_249_n 0.011086f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_179 A2 B2 0.0197629f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A2_c_215_n B2 4.16298e-19 $X=1.74 $Y=1.615 $X2=0 $Y2=0
cc_181 A2 N_B2_c_252_n 4.19338e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_182 N_A2_c_215_n N_B2_c_252_n 0.0181454f $X=1.74 $Y=1.615 $X2=0 $Y2=0
cc_183 N_A2_M1002_g N_VPWR_c_391_n 0.005209f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_184 N_A2_M1002_g N_VPWR_c_388_n 0.00984319f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_185 N_A2_M1000_g N_VGND_c_433_n 0.0122599f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_186 N_A2_M1000_g N_VGND_c_434_n 0.00421418f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_187 N_A2_M1000_g N_VGND_c_437_n 0.00432128f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_188 N_A2_M1000_g N_A_245_94#_c_476_n 0.00350341f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_189 N_A2_M1000_g N_A_245_94#_c_477_n 0.0153207f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_190 A2 N_A_245_94#_c_477_n 0.0250329f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A2_c_215_n N_A_245_94#_c_477_n 0.0041539f $X=1.74 $Y=1.615 $X2=0 $Y2=0
cc_192 N_A2_M1000_g N_A_456_74#_c_512_n 0.00116577f $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_193 N_A2_M1000_g N_A_456_74#_c_514_n 3.62451e-19 $X=1.65 $Y=0.79 $X2=0 $Y2=0
cc_194 N_B2_c_250_n N_B1_M1008_g 0.0275047f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_195 B2 N_B1_M1008_g 2.17586e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_196 N_B2_c_252_n N_B1_M1008_g 0.00510377f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_197 B2 B1 0.0260436f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_198 N_B2_c_252_n B1 2.35705e-19 $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_199 N_B2_M1011_g N_B1_c_294_n 0.0413135f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_200 N_B2_c_248_n N_B1_c_294_n 0.00239154f $X=2.645 $Y=1.175 $X2=0 $Y2=0
cc_201 B2 N_B1_c_294_n 0.00659348f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_202 N_B2_c_252_n N_B1_c_294_n 0.00387701f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_203 N_B2_c_253_n N_B1_c_294_n 0.00773329f $X=2.31 $Y=1.78 $X2=0 $Y2=0
cc_204 N_B2_M1011_g N_VPWR_c_390_n 0.00356673f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_205 N_B2_M1011_g N_VPWR_c_391_n 0.00553757f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_206 N_B2_M1011_g N_VPWR_c_388_n 0.0109203f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_207 N_B2_c_250_n N_VGND_c_433_n 7.83914e-19 $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_208 N_B2_c_250_n N_VGND_c_436_n 0.00278271f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_209 N_B2_c_250_n N_VGND_c_437_n 0.00358525f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_210 N_B2_c_248_n N_A_245_94#_c_477_n 0.0178297f $X=2.645 $Y=1.175 $X2=0 $Y2=0
cc_211 N_B2_c_249_n N_A_245_94#_c_477_n 0.0118983f $X=2.475 $Y=1.175 $X2=0 $Y2=0
cc_212 B2 N_A_245_94#_c_477_n 0.0457618f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B2_c_252_n N_A_245_94#_c_477_n 0.0063832f $X=2.31 $Y=1.615 $X2=0 $Y2=0
cc_214 N_B2_c_248_n N_A_245_94#_c_495_n 5.20128e-19 $X=2.645 $Y=1.175 $X2=0
+ $Y2=0
cc_215 N_B2_c_250_n N_A_245_94#_c_495_n 0.0123389f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_216 N_B2_c_249_n N_A_456_74#_c_512_n 0.00812328f $X=2.475 $Y=1.175 $X2=0
+ $Y2=0
cc_217 N_B2_c_250_n N_A_456_74#_c_513_n 0.0133401f $X=2.72 $Y=1.1 $X2=0 $Y2=0
cc_218 B1 N_C1_c_328_n 4.13026e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B1_c_294_n N_C1_c_328_n 0.0178735f $X=3.09 $Y=1.625 $X2=0 $Y2=0
cc_220 N_B1_M1008_g C1 0.00496568f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_221 B1 C1 0.0208926f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B1_c_294_n C1 0.00207338f $X=3.09 $Y=1.625 $X2=0 $Y2=0
cc_223 N_B1_M1008_g N_C1_c_331_n 0.0147786f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_224 N_B1_M1008_g N_C1_c_332_n 0.017212f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_225 N_B1_M1005_g N_VPWR_c_390_n 0.0228889f $X=2.805 $Y=2.46 $X2=0 $Y2=0
cc_226 N_B1_M1005_g N_VPWR_c_391_n 0.00460063f $X=2.805 $Y=2.46 $X2=0 $Y2=0
cc_227 N_B1_M1005_g N_VPWR_c_388_n 0.00909693f $X=2.805 $Y=2.46 $X2=0 $Y2=0
cc_228 N_B1_M1008_g N_VGND_c_436_n 0.00278271f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_229 N_B1_M1008_g N_VGND_c_437_n 0.00354237f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_230 N_B1_M1008_g N_A_245_94#_c_477_n 0.00516704f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_231 B1 N_A_245_94#_c_477_n 0.0140154f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B1_c_294_n N_A_245_94#_c_477_n 0.00705294f $X=3.09 $Y=1.625 $X2=0 $Y2=0
cc_233 N_B1_M1008_g N_A_245_94#_c_495_n 0.0084974f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_234 N_B1_M1008_g N_A_456_74#_c_513_n 0.0133206f $X=3.15 $Y=0.69 $X2=0 $Y2=0
cc_235 N_C1_M1009_g N_VPWR_c_390_n 0.00668958f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_236 N_C1_M1009_g N_VPWR_c_392_n 0.005209f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_237 N_C1_M1009_g N_VPWR_c_388_n 0.00990469f $X=3.815 $Y=2.46 $X2=0 $Y2=0
cc_238 N_C1_c_332_n N_VGND_c_436_n 0.00430908f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_239 N_C1_c_332_n N_VGND_c_437_n 0.00821503f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_240 C1 N_A_245_94#_c_477_n 0.00728498f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_241 N_C1_c_332_n N_A_245_94#_c_495_n 6.13134e-19 $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_242 N_C1_c_332_n N_A_456_74#_c_513_n 0.00735461f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_243 C1 N_A_456_74#_c_522_n 0.00723658f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_244 N_C1_c_331_n N_A_456_74#_c_522_n 4.53017e-19 $X=3.66 $Y=1.285 $X2=0 $Y2=0
cc_245 N_C1_c_332_n N_A_456_74#_c_522_n 0.0059147f $X=3.7 $Y=1.12 $X2=0 $Y2=0
cc_246 N_X_c_369_n N_VPWR_c_389_n 0.0422698f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_247 N_X_c_369_n N_VPWR_c_388_n 0.0119743f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_248 N_X_c_369_n N_VPWR_c_394_n 0.014549f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_249 N_X_c_367_n N_VGND_c_432_n 0.0317414f $X=0.355 $Y=0.515 $X2=0 $Y2=0
cc_250 N_X_c_367_n N_VGND_c_437_n 0.0147684f $X=0.355 $Y=0.515 $X2=0 $Y2=0
cc_251 N_X_c_367_n N_VGND_c_438_n 0.0179105f $X=0.355 $Y=0.515 $X2=0 $Y2=0
cc_252 N_VGND_c_432_n N_A_245_94#_c_476_n 0.0243787f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_253 N_VGND_c_433_n N_A_245_94#_c_476_n 0.0191765f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_254 N_VGND_c_434_n N_A_245_94#_c_476_n 0.0103491f $X=1.7 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_437_n N_A_245_94#_c_476_n 0.0113354f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_433_n N_A_245_94#_c_477_n 0.0244412f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_257 N_VGND_c_432_n N_A_245_94#_c_478_n 0.00156673f $X=0.855 $Y=0.515 $X2=0
+ $Y2=0
cc_258 N_VGND_c_433_n N_A_456_74#_c_512_n 0.0346871f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_259 N_VGND_c_436_n N_A_456_74#_c_513_n 0.0664804f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_437_n N_A_456_74#_c_513_n 0.0369159f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_433_n N_A_456_74#_c_514_n 0.0121618f $X=1.865 $Y=0.735 $X2=0
+ $Y2=0
cc_262 N_VGND_c_436_n N_A_456_74#_c_514_n 0.0236697f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_437_n N_A_456_74#_c_514_n 0.0128321f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_264 N_A_245_94#_c_477_n N_A_456_74#_c_512_n 0.0258597f $X=2.77 $Y=1.195 $X2=0
+ $Y2=0
cc_265 N_A_245_94#_M1001_d N_A_456_74#_c_513_n 0.00176461f $X=2.795 $Y=0.37
+ $X2=0 $Y2=0
cc_266 N_A_245_94#_c_495_n N_A_456_74#_c_513_n 0.016064f $X=2.935 $Y=0.81 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__dlrtn_2.pxi.spice
* Created: Wed Sep  2 12:05:30 2020
* 
x_PM_SKY130_FD_SC_MS__DLRTN_2%D N_D_M1017_g N_D_M1015_g D N_D_c_145_n
+ PM_SKY130_FD_SC_MS__DLRTN_2%D
x_PM_SKY130_FD_SC_MS__DLRTN_2%GATE_N N_GATE_N_M1001_g N_GATE_N_M1011_g GATE_N
+ N_GATE_N_c_175_n PM_SKY130_FD_SC_MS__DLRTN_2%GATE_N
x_PM_SKY130_FD_SC_MS__DLRTN_2%A_232_98# N_A_232_98#_M1001_d N_A_232_98#_M1011_d
+ N_A_232_98#_c_212_n N_A_232_98#_M1021_g N_A_232_98#_M1007_g
+ N_A_232_98#_M1014_g N_A_232_98#_M1012_g N_A_232_98#_c_216_n
+ N_A_232_98#_c_217_n N_A_232_98#_c_223_n N_A_232_98#_c_218_n
+ N_A_232_98#_c_225_n N_A_232_98#_c_226_n N_A_232_98#_c_227_n
+ N_A_232_98#_c_228_n N_A_232_98#_c_229_n N_A_232_98#_c_230_n
+ N_A_232_98#_c_219_n PM_SKY130_FD_SC_MS__DLRTN_2%A_232_98#
x_PM_SKY130_FD_SC_MS__DLRTN_2%A_27_136# N_A_27_136#_M1017_s N_A_27_136#_M1015_s
+ N_A_27_136#_c_331_n N_A_27_136#_M1003_g N_A_27_136#_c_333_n
+ N_A_27_136#_c_334_n N_A_27_136#_M1016_g N_A_27_136#_c_335_n
+ N_A_27_136#_c_336_n N_A_27_136#_c_337_n N_A_27_136#_c_338_n
+ N_A_27_136#_c_339_n N_A_27_136#_c_342_n N_A_27_136#_c_340_n
+ PM_SKY130_FD_SC_MS__DLRTN_2%A_27_136#
x_PM_SKY130_FD_SC_MS__DLRTN_2%A_373_82# N_A_373_82#_M1007_s N_A_373_82#_M1021_s
+ N_A_373_82#_M1010_g N_A_373_82#_M1020_g N_A_373_82#_c_416_n
+ N_A_373_82#_c_417_n N_A_373_82#_c_409_n N_A_373_82#_c_410_n
+ N_A_373_82#_c_411_n N_A_373_82#_c_412_n N_A_373_82#_c_413_n
+ N_A_373_82#_c_419_n N_A_373_82#_c_414_n PM_SKY130_FD_SC_MS__DLRTN_2%A_373_82#
x_PM_SKY130_FD_SC_MS__DLRTN_2%A_913_406# N_A_913_406#_M1002_s
+ N_A_913_406#_M1008_d N_A_913_406#_M1005_g N_A_913_406#_M1018_g
+ N_A_913_406#_c_519_n N_A_913_406#_c_504_n N_A_913_406#_M1006_g
+ N_A_913_406#_M1004_g N_A_913_406#_c_507_n N_A_913_406#_M1009_g
+ N_A_913_406#_M1013_g N_A_913_406#_c_510_n N_A_913_406#_c_511_n
+ N_A_913_406#_c_522_n N_A_913_406#_c_523_n N_A_913_406#_c_512_n
+ N_A_913_406#_c_524_n N_A_913_406#_c_525_n N_A_913_406#_c_513_n
+ N_A_913_406#_c_526_n N_A_913_406#_c_514_n N_A_913_406#_c_515_n
+ N_A_913_406#_c_529_n N_A_913_406#_c_516_n
+ PM_SKY130_FD_SC_MS__DLRTN_2%A_913_406#
x_PM_SKY130_FD_SC_MS__DLRTN_2%A_673_392# N_A_673_392#_M1014_d
+ N_A_673_392#_M1010_d N_A_673_392#_M1008_g N_A_673_392#_M1002_g
+ N_A_673_392#_c_641_n N_A_673_392#_c_642_n N_A_673_392#_c_651_n
+ N_A_673_392#_c_652_n N_A_673_392#_c_653_n N_A_673_392#_c_654_n
+ N_A_673_392#_c_643_n N_A_673_392#_c_644_n N_A_673_392#_c_645_n
+ N_A_673_392#_c_646_n N_A_673_392#_c_647_n
+ PM_SKY130_FD_SC_MS__DLRTN_2%A_673_392#
x_PM_SKY130_FD_SC_MS__DLRTN_2%RESET_B N_RESET_B_M1000_g N_RESET_B_M1019_g
+ RESET_B N_RESET_B_c_741_n N_RESET_B_c_742_n N_RESET_B_c_743_n
+ PM_SKY130_FD_SC_MS__DLRTN_2%RESET_B
x_PM_SKY130_FD_SC_MS__DLRTN_2%VPWR N_VPWR_M1015_d N_VPWR_M1021_d N_VPWR_M1005_d
+ N_VPWR_M1019_d N_VPWR_M1009_s N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n
+ N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n N_VPWR_c_784_n VPWR
+ N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n N_VPWR_c_788_n N_VPWR_c_789_n
+ N_VPWR_c_790_n N_VPWR_c_791_n N_VPWR_c_777_n PM_SKY130_FD_SC_MS__DLRTN_2%VPWR
x_PM_SKY130_FD_SC_MS__DLRTN_2%Q N_Q_M1004_d N_Q_M1006_d N_Q_c_863_n N_Q_c_864_n
+ Q Q Q N_Q_c_867_n N_Q_c_865_n PM_SKY130_FD_SC_MS__DLRTN_2%Q
x_PM_SKY130_FD_SC_MS__DLRTN_2%VGND N_VGND_M1017_d N_VGND_M1007_d N_VGND_M1018_d
+ N_VGND_M1000_d N_VGND_M1013_s N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n
+ N_VGND_c_901_n VGND N_VGND_c_902_n N_VGND_c_903_n N_VGND_c_904_n
+ N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n N_VGND_c_908_n N_VGND_c_909_n
+ N_VGND_c_910_n N_VGND_c_911_n PM_SKY130_FD_SC_MS__DLRTN_2%VGND
cc_1 VNB N_D_M1017_g 0.028834f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_2 VNB D 0.00388042f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_c_145_n 0.0258834f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.615
cc_4 VNB N_GATE_N_M1001_g 0.0314722f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_5 VNB GATE_N 0.0017082f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_GATE_N_c_175_n 0.0197779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_232_98#_c_212_n 0.0157424f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.39
cc_8 VNB N_A_232_98#_M1021_g 0.00884119f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_9 VNB N_A_232_98#_M1007_g 0.0275675f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_10 VNB N_A_232_98#_M1014_g 0.049147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_232_98#_c_216_n 0.00676283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_232_98#_c_217_n 0.00820746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_232_98#_c_218_n 0.0145513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_232_98#_c_219_n 0.0270096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_136#_c_331_n 0.0442213f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.39
cc_16 VNB N_A_27_136#_M1003_g 0.00414833f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A_27_136#_c_333_n 0.0386914f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_18 VNB N_A_27_136#_c_334_n 0.0181563f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_19 VNB N_A_27_136#_c_335_n 0.0125907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_136#_c_336_n 0.0120287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_136#_c_337_n 0.0115633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_136#_c_338_n 0.00498838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_136#_c_339_n 0.0132007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_136#_c_340_n 0.0193493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_373_82#_M1020_g 0.0320396f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_26 VNB N_A_373_82#_c_409_n 0.0159493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_373_82#_c_410_n 0.00173945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_373_82#_c_411_n 0.0196327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_373_82#_c_412_n 0.0312102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_373_82#_c_413_n 0.00442376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_373_82#_c_414_n 0.00351115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_913_406#_M1018_g 0.0652905f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_33 VNB N_A_913_406#_c_504_n 0.0141135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_913_406#_M1006_g 0.00962424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_913_406#_M1004_g 0.0280574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_913_406#_c_507_n 0.00970685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_913_406#_M1009_g 0.0151082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_913_406#_M1013_g 0.0275403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_913_406#_c_510_n 0.00424728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_913_406#_c_511_n 0.012538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_913_406#_c_512_n 0.00885266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_913_406#_c_513_n 0.00415206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_913_406#_c_514_n 0.00286577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_913_406#_c_515_n 0.014959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_913_406#_c_516_n 0.0360511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_673_392#_M1002_g 0.0277598f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_47 VNB N_A_673_392#_c_641_n 0.0345938f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_48 VNB N_A_673_392#_c_642_n 0.0145515f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.615
cc_49 VNB N_A_673_392#_c_643_n 0.0028741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_673_392#_c_644_n 0.0175228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_673_392#_c_645_n 0.00257655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_673_392#_c_646_n 0.010508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_673_392#_c_647_n 0.00694351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_RESET_B_M1019_g 0.00645307f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.39
cc_55 VNB N_RESET_B_c_741_n 0.0289522f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_56 VNB N_RESET_B_c_742_n 0.0157968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_c_743_n 0.0208067f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_58 VNB N_VPWR_c_777_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Q_c_863_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_60 VNB N_Q_c_864_n 3.99771e-19 $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_61 VNB N_Q_c_865_n 0.00123966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_898_n 0.00989418f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.615
cc_63 VNB N_VGND_c_899_n 0.011769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_900_n 0.0125358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_901_n 0.0551324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_902_n 0.0194325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_903_n 0.0439944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_904_n 0.0300433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_905_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_906_n 0.023189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_907_n 0.0382579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_908_n 0.0291695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_909_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_910_n 0.0172179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_911_n 0.453507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VPB N_D_M1015_g 0.0301058f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.39
cc_77 VPB D 0.00196111f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_78 VPB N_D_c_145_n 0.0129489f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.615
cc_79 VPB N_GATE_N_M1011_g 0.0285961f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.39
cc_80 VPB GATE_N 0.00195884f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_81 VPB N_GATE_N_c_175_n 0.0132673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_232_98#_M1021_g 0.0372685f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.615
cc_83 VPB N_A_232_98#_M1014_g 0.0256747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_232_98#_M1012_g 0.0251921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_232_98#_c_223_n 0.00488677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_232_98#_c_218_n 0.00704763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_232_98#_c_225_n 0.00963284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_232_98#_c_226_n 0.00686999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_232_98#_c_227_n 0.00592361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_232_98#_c_228_n 0.054335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_232_98#_c_229_n 0.00911394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_232_98#_c_230_n 0.00526719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_232_98#_c_219_n 0.0100157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_136#_M1003_g 0.030505f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_95 VPB N_A_27_136#_c_342_n 0.0542876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_136#_c_340_n 0.0139522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_373_82#_M1010_g 0.0216089f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_98 VPB N_A_373_82#_c_416_n 0.0150426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_373_82#_c_417_n 6.63005e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_373_82#_c_409_n 0.0139743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_373_82#_c_419_n 0.00675226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_373_82#_c_414_n 0.0022585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_913_406#_M1005_g 0.0303207f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_104 VPB N_A_913_406#_M1018_g 0.00154973f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_105 VPB N_A_913_406#_c_519_n 0.00811541f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_106 VPB N_A_913_406#_M1006_g 0.0253341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_913_406#_M1009_g 0.0273989f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_913_406#_c_522_n 0.0127768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_913_406#_c_523_n 0.0307097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_913_406#_c_524_n 0.00240191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_913_406#_c_525_n 0.00754493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_913_406#_c_526_n 0.00744566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_913_406#_c_514_n 3.58276e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_913_406#_c_515_n 0.00286928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_913_406#_c_529_n 0.0262775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_673_392#_M1008_g 0.0236506f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_117 VPB N_A_673_392#_c_641_n 0.0156573f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_118 VPB N_A_673_392#_c_642_n 7.8261e-19 $X=-0.19 $Y=1.66 $X2=0.675 $Y2=1.615
cc_119 VPB N_A_673_392#_c_651_n 6.56999e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_673_392#_c_652_n 0.00273707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_673_392#_c_653_n 0.0252082f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_673_392#_c_654_n 0.00172416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_673_392#_c_646_n 0.00476225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_RESET_B_M1019_g 0.0249194f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=2.39
cc_125 VPB N_VPWR_c_778_n 0.0308367f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_126 VPB N_VPWR_c_779_n 0.013216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_780_n 0.0102253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_781_n 0.0123832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_782_n 0.0709516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_783_n 0.0241107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_784_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_785_n 0.0348259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_786_n 0.0220361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_787_n 0.028134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_788_n 0.00631473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_789_n 0.0566101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_790_n 0.0286325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_791_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_777_n 0.115523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB Q 0.00429432f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.615
cc_141 VPB N_Q_c_867_n 0.00410866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_Q_c_865_n 0.00103009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 N_D_M1017_g N_GATE_N_M1001_g 0.0245058f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_144 N_D_M1015_g N_GATE_N_M1011_g 0.0141966f $X=0.675 $Y=2.39 $X2=0 $Y2=0
cc_145 D GATE_N 0.0264884f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_146 N_D_c_145_n GATE_N 3.62002e-19 $X=0.675 $Y=1.615 $X2=0 $Y2=0
cc_147 D N_GATE_N_c_175_n 0.00201746f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_148 N_D_c_145_n N_GATE_N_c_175_n 0.0174151f $X=0.675 $Y=1.615 $X2=0 $Y2=0
cc_149 N_D_M1017_g N_A_232_98#_c_217_n 0.00147505f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_150 N_D_M1017_g N_A_27_136#_c_335_n 0.00689961f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_151 N_D_M1017_g N_A_27_136#_c_336_n 0.0118249f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_152 N_D_M1017_g N_A_27_136#_c_337_n 0.00420241f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_153 N_D_M1017_g N_A_27_136#_c_339_n 0.00657237f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_154 D N_A_27_136#_c_339_n 6.29576e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_155 N_D_M1015_g N_A_27_136#_c_342_n 0.0152415f $X=0.675 $Y=2.39 $X2=0 $Y2=0
cc_156 D N_A_27_136#_c_342_n 0.0149649f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_157 N_D_c_145_n N_A_27_136#_c_342_n 0.00475259f $X=0.675 $Y=1.615 $X2=0 $Y2=0
cc_158 N_D_M1017_g N_A_27_136#_c_340_n 0.0128282f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_159 N_D_M1015_g N_A_27_136#_c_340_n 0.0035594f $X=0.675 $Y=2.39 $X2=0 $Y2=0
cc_160 D N_A_27_136#_c_340_n 0.0251401f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_161 N_D_M1015_g N_VPWR_c_778_n 0.00460946f $X=0.675 $Y=2.39 $X2=0 $Y2=0
cc_162 D N_VPWR_c_778_n 0.00433462f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_163 N_D_M1015_g N_VPWR_c_783_n 0.00546844f $X=0.675 $Y=2.39 $X2=0 $Y2=0
cc_164 N_D_M1015_g N_VPWR_c_777_n 0.00599321f $X=0.675 $Y=2.39 $X2=0 $Y2=0
cc_165 N_D_M1017_g N_VGND_c_902_n 0.00297615f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_166 N_D_M1017_g N_VGND_c_911_n 0.00454494f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_167 N_GATE_N_M1001_g N_A_232_98#_c_217_n 0.00829292f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_168 GATE_N N_A_232_98#_c_217_n 0.0138981f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_169 N_GATE_N_c_175_n N_A_232_98#_c_217_n 0.00123995f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_170 N_GATE_N_M1011_g N_A_232_98#_c_223_n 0.0076028f $X=1.225 $Y=2.39 $X2=0
+ $Y2=0
cc_171 N_GATE_N_M1001_g N_A_232_98#_c_218_n 0.00486829f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_172 GATE_N N_A_232_98#_c_218_n 0.0177666f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_173 N_GATE_N_c_175_n N_A_232_98#_c_218_n 0.00135318f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_174 N_GATE_N_M1011_g N_A_232_98#_c_226_n 0.00433562f $X=1.225 $Y=2.39 $X2=0
+ $Y2=0
cc_175 N_GATE_N_M1011_g N_A_232_98#_c_229_n 0.0030318f $X=1.225 $Y=2.39 $X2=0
+ $Y2=0
cc_176 GATE_N N_A_232_98#_c_229_n 0.00393715f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_177 N_GATE_N_M1011_g N_A_232_98#_c_230_n 0.00578119f $X=1.225 $Y=2.39 $X2=0
+ $Y2=0
cc_178 GATE_N N_A_232_98#_c_230_n 0.0082296f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_179 N_GATE_N_c_175_n N_A_232_98#_c_230_n 0.00246407f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_180 N_GATE_N_M1001_g N_A_232_98#_c_219_n 0.00268628f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_181 GATE_N N_A_232_98#_c_219_n 2.42469e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_182 N_GATE_N_c_175_n N_A_232_98#_c_219_n 0.0115984f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_183 N_GATE_N_M1001_g N_A_27_136#_c_335_n 0.00225195f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_184 N_GATE_N_M1001_g N_A_27_136#_c_336_n 0.0176812f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_185 N_GATE_N_M1011_g N_A_373_82#_c_419_n 6.83713e-19 $X=1.225 $Y=2.39 $X2=0
+ $Y2=0
cc_186 N_GATE_N_M1011_g N_VPWR_c_778_n 0.0046091f $X=1.225 $Y=2.39 $X2=0 $Y2=0
cc_187 GATE_N N_VPWR_c_778_n 0.00915244f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_188 N_GATE_N_c_175_n N_VPWR_c_778_n 8.44966e-19 $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_189 N_GATE_N_M1011_g N_VPWR_c_785_n 0.00546038f $X=1.225 $Y=2.39 $X2=0 $Y2=0
cc_190 N_GATE_N_M1011_g N_VPWR_c_777_n 0.00599321f $X=1.225 $Y=2.39 $X2=0 $Y2=0
cc_191 N_GATE_N_M1001_g N_VGND_c_906_n 0.00210264f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_192 N_GATE_N_M1001_g N_VGND_c_907_n 0.00374721f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_193 N_GATE_N_M1001_g N_VGND_c_911_n 0.00508379f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_194 N_A_232_98#_M1007_g N_A_27_136#_c_331_n 0.0167777f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_195 N_A_232_98#_M1021_g N_A_27_136#_M1003_g 0.0384185f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_196 N_A_232_98#_c_225_n N_A_27_136#_M1003_g 0.0157162f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_197 N_A_232_98#_M1014_g N_A_27_136#_c_334_n 0.056201f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_198 N_A_232_98#_M1001_d N_A_27_136#_c_336_n 0.00784312f $X=1.16 $Y=0.49 $X2=0
+ $Y2=0
cc_199 N_A_232_98#_M1007_g N_A_27_136#_c_336_n 0.0176894f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_200 N_A_232_98#_c_217_n N_A_27_136#_c_336_n 0.0238302f $X=1.505 $Y=1.085
+ $X2=0 $Y2=0
cc_201 N_A_232_98#_c_218_n N_A_27_136#_c_336_n 0.0193437f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_202 N_A_232_98#_c_219_n N_A_27_136#_c_336_n 0.00122731f $X=1.74 $Y=1.415
+ $X2=0 $Y2=0
cc_203 N_A_232_98#_M1007_g N_A_27_136#_c_338_n 0.0117503f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_204 N_A_232_98#_c_225_n N_A_373_82#_M1021_s 0.00720588f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_205 N_A_232_98#_M1014_g N_A_373_82#_M1010_g 0.039003f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_206 N_A_232_98#_c_225_n N_A_373_82#_M1010_g 0.0150236f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_207 N_A_232_98#_M1014_g N_A_373_82#_M1020_g 0.0215197f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_208 N_A_232_98#_M1021_g N_A_373_82#_c_416_n 0.0100792f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_209 N_A_232_98#_M1014_g N_A_373_82#_c_416_n 6.13645e-19 $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_210 N_A_232_98#_c_225_n N_A_373_82#_c_416_n 0.0263744f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_211 N_A_232_98#_M1014_g N_A_373_82#_c_417_n 0.00134433f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_212 N_A_232_98#_M1014_g N_A_373_82#_c_409_n 0.0180105f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_213 N_A_232_98#_M1014_g N_A_373_82#_c_411_n 0.0228893f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_214 N_A_232_98#_M1014_g N_A_373_82#_c_412_n 0.021337f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_215 N_A_232_98#_c_228_n N_A_373_82#_c_412_n 0.00434555f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_216 N_A_232_98#_c_212_n N_A_373_82#_c_413_n 0.00469476f $X=2.145 $Y=1.415
+ $X2=0 $Y2=0
cc_217 N_A_232_98#_M1007_g N_A_373_82#_c_413_n 0.00618595f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_218 N_A_232_98#_c_218_n N_A_373_82#_c_413_n 0.0266185f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_219 N_A_232_98#_c_219_n N_A_373_82#_c_413_n 4.35132e-19 $X=1.74 $Y=1.415
+ $X2=0 $Y2=0
cc_220 N_A_232_98#_c_212_n N_A_373_82#_c_419_n 0.00349637f $X=2.145 $Y=1.415
+ $X2=0 $Y2=0
cc_221 N_A_232_98#_M1021_g N_A_373_82#_c_419_n 0.0153854f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_222 N_A_232_98#_c_218_n N_A_373_82#_c_419_n 0.00488298f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_223 N_A_232_98#_c_225_n N_A_373_82#_c_419_n 0.0268578f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_224 N_A_232_98#_c_230_n N_A_373_82#_c_419_n 0.043001f $X=1.48 $Y=1.95 $X2=0
+ $Y2=0
cc_225 N_A_232_98#_c_219_n N_A_373_82#_c_419_n 4.53443e-19 $X=1.74 $Y=1.415
+ $X2=0 $Y2=0
cc_226 N_A_232_98#_c_212_n N_A_373_82#_c_414_n 0.00585489f $X=2.145 $Y=1.415
+ $X2=0 $Y2=0
cc_227 N_A_232_98#_M1021_g N_A_373_82#_c_414_n 0.0117641f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_228 N_A_232_98#_M1007_g N_A_373_82#_c_414_n 0.00598842f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_229 N_A_232_98#_c_216_n N_A_373_82#_c_414_n 0.00360478f $X=2.235 $Y=1.415
+ $X2=0 $Y2=0
cc_230 N_A_232_98#_c_218_n N_A_373_82#_c_414_n 0.0321568f $X=1.59 $Y=1.67 $X2=0
+ $Y2=0
cc_231 N_A_232_98#_c_230_n N_A_373_82#_c_414_n 0.00704491f $X=1.48 $Y=1.95 $X2=0
+ $Y2=0
cc_232 N_A_232_98#_c_219_n N_A_373_82#_c_414_n 5.43459e-19 $X=1.74 $Y=1.415
+ $X2=0 $Y2=0
cc_233 N_A_232_98#_M1012_g N_A_913_406#_M1005_g 0.0123422f $X=3.815 $Y=2.73
+ $X2=0 $Y2=0
cc_234 N_A_232_98#_c_225_n N_A_913_406#_M1005_g 0.0038923f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_235 N_A_232_98#_c_227_n N_A_913_406#_M1005_g 0.00397869f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_236 N_A_232_98#_c_227_n N_A_913_406#_c_522_n 0.0198487f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_237 N_A_232_98#_c_228_n N_A_913_406#_c_522_n 0.00135115f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_238 N_A_232_98#_c_227_n N_A_913_406#_c_523_n 4.19484e-19 $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_239 N_A_232_98#_c_228_n N_A_913_406#_c_523_n 0.0184475f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_240 N_A_232_98#_c_225_n N_A_673_392#_M1010_d 0.00692933f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_241 N_A_232_98#_c_225_n N_A_673_392#_c_651_n 0.0301739f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_242 N_A_232_98#_c_227_n N_A_673_392#_c_651_n 0.013226f $X=4.16 $Y=2.195 $X2=0
+ $Y2=0
cc_243 N_A_232_98#_c_228_n N_A_673_392#_c_651_n 0.00790539f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_244 N_A_232_98#_M1014_g N_A_673_392#_c_652_n 0.0089637f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_245 N_A_232_98#_c_227_n N_A_673_392#_c_652_n 0.010678f $X=4.16 $Y=2.195 $X2=0
+ $Y2=0
cc_246 N_A_232_98#_c_228_n N_A_673_392#_c_652_n 0.00445706f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_247 N_A_232_98#_M1014_g N_A_673_392#_c_653_n 0.00689739f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_248 N_A_232_98#_c_225_n N_A_673_392#_c_653_n 0.00354902f $X=3.995 $Y=2.605
+ $X2=0 $Y2=0
cc_249 N_A_232_98#_c_227_n N_A_673_392#_c_653_n 0.0261498f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_250 N_A_232_98#_c_228_n N_A_673_392#_c_653_n 0.00496075f $X=4.16 $Y=2.195
+ $X2=0 $Y2=0
cc_251 N_A_232_98#_M1014_g N_A_673_392#_c_654_n 0.00393099f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_252 N_A_232_98#_M1014_g N_A_673_392#_c_643_n 7.62689e-19 $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_253 N_A_232_98#_M1014_g N_A_673_392#_c_645_n 0.00113438f $X=3.8 $Y=0.69 $X2=0
+ $Y2=0
cc_254 N_A_232_98#_c_225_n N_VPWR_M1021_d 0.0100288f $X=3.995 $Y=2.605 $X2=0
+ $Y2=0
cc_255 N_A_232_98#_c_226_n N_VPWR_c_778_n 0.0133739f $X=1.675 $Y=2.605 $X2=0
+ $Y2=0
cc_256 N_A_232_98#_c_229_n N_VPWR_c_778_n 0.022655f $X=1.45 $Y=2.115 $X2=0 $Y2=0
cc_257 N_A_232_98#_M1021_g N_VPWR_c_779_n 0.00205413f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_258 N_A_232_98#_c_225_n N_VPWR_c_779_n 0.0249677f $X=3.995 $Y=2.605 $X2=0
+ $Y2=0
cc_259 N_A_232_98#_M1021_g N_VPWR_c_785_n 0.00433266f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_260 N_A_232_98#_c_225_n N_VPWR_c_785_n 0.0112491f $X=3.995 $Y=2.605 $X2=0
+ $Y2=0
cc_261 N_A_232_98#_c_226_n N_VPWR_c_785_n 0.0107106f $X=1.675 $Y=2.605 $X2=0
+ $Y2=0
cc_262 N_A_232_98#_M1012_g N_VPWR_c_789_n 0.00518677f $X=3.815 $Y=2.73 $X2=0
+ $Y2=0
cc_263 N_A_232_98#_c_225_n N_VPWR_c_789_n 0.0252583f $X=3.995 $Y=2.605 $X2=0
+ $Y2=0
cc_264 N_A_232_98#_c_225_n N_VPWR_c_790_n 0.00270878f $X=3.995 $Y=2.605 $X2=0
+ $Y2=0
cc_265 N_A_232_98#_M1021_g N_VPWR_c_777_n 0.00595788f $X=2.235 $Y=2.38 $X2=0
+ $Y2=0
cc_266 N_A_232_98#_M1012_g N_VPWR_c_777_n 0.00647345f $X=3.815 $Y=2.73 $X2=0
+ $Y2=0
cc_267 N_A_232_98#_c_225_n N_VPWR_c_777_n 0.0659417f $X=3.995 $Y=2.605 $X2=0
+ $Y2=0
cc_268 N_A_232_98#_c_226_n N_VPWR_c_777_n 0.0130158f $X=1.675 $Y=2.605 $X2=0
+ $Y2=0
cc_269 N_A_232_98#_c_225_n A_589_392# 0.00450673f $X=3.995 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_270 N_A_232_98#_c_225_n A_781_504# 0.0113875f $X=3.995 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_271 N_A_232_98#_M1014_g N_VGND_c_903_n 0.00461464f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_272 N_A_232_98#_M1007_g N_VGND_c_907_n 0.00414982f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_273 N_A_232_98#_M1007_g N_VGND_c_908_n 0.0060117f $X=2.25 $Y=0.78 $X2=0 $Y2=0
cc_274 N_A_232_98#_M1007_g N_VGND_c_911_n 0.00533081f $X=2.25 $Y=0.78 $X2=0
+ $Y2=0
cc_275 N_A_232_98#_M1014_g N_VGND_c_911_n 0.00909529f $X=3.8 $Y=0.69 $X2=0 $Y2=0
cc_276 N_A_27_136#_c_336_n N_A_373_82#_M1007_s 0.00778716f $X=2.615 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_277 N_A_27_136#_M1003_g N_A_373_82#_M1010_g 0.0735195f $X=2.855 $Y=2.46 $X2=0
+ $Y2=0
cc_278 N_A_27_136#_c_331_n N_A_373_82#_c_416_n 9.68515e-19 $X=2.855 $Y=1.59
+ $X2=0 $Y2=0
cc_279 N_A_27_136#_M1003_g N_A_373_82#_c_416_n 0.014815f $X=2.855 $Y=2.46 $X2=0
+ $Y2=0
cc_280 N_A_27_136#_c_333_n N_A_373_82#_c_416_n 0.00467116f $X=3.335 $Y=1.185
+ $X2=0 $Y2=0
cc_281 N_A_27_136#_c_338_n N_A_373_82#_c_416_n 0.0189066f $X=2.78 $Y=1.425 $X2=0
+ $Y2=0
cc_282 N_A_27_136#_c_331_n N_A_373_82#_c_417_n 0.00166193f $X=2.855 $Y=1.59
+ $X2=0 $Y2=0
cc_283 N_A_27_136#_M1003_g N_A_373_82#_c_417_n 8.66641e-19 $X=2.855 $Y=2.46
+ $X2=0 $Y2=0
cc_284 N_A_27_136#_c_338_n N_A_373_82#_c_417_n 0.00440446f $X=2.78 $Y=1.425
+ $X2=0 $Y2=0
cc_285 N_A_27_136#_c_331_n N_A_373_82#_c_409_n 0.0210237f $X=2.855 $Y=1.59 $X2=0
+ $Y2=0
cc_286 N_A_27_136#_c_333_n N_A_373_82#_c_409_n 0.0214194f $X=3.335 $Y=1.185
+ $X2=0 $Y2=0
cc_287 N_A_27_136#_c_338_n N_A_373_82#_c_409_n 3.06958e-19 $X=2.78 $Y=1.425
+ $X2=0 $Y2=0
cc_288 N_A_27_136#_c_331_n N_A_373_82#_c_410_n 0.00496558f $X=2.855 $Y=1.59
+ $X2=0 $Y2=0
cc_289 N_A_27_136#_c_333_n N_A_373_82#_c_410_n 0.0227079f $X=3.335 $Y=1.185
+ $X2=0 $Y2=0
cc_290 N_A_27_136#_c_338_n N_A_373_82#_c_410_n 0.0231983f $X=2.78 $Y=1.425 $X2=0
+ $Y2=0
cc_291 N_A_27_136#_c_336_n N_A_373_82#_c_413_n 0.0253275f $X=2.615 $Y=0.665
+ $X2=0 $Y2=0
cc_292 N_A_27_136#_c_338_n N_A_373_82#_c_413_n 0.0110325f $X=2.78 $Y=1.425 $X2=0
+ $Y2=0
cc_293 N_A_27_136#_M1003_g N_A_373_82#_c_419_n 0.00177924f $X=2.855 $Y=2.46
+ $X2=0 $Y2=0
cc_294 N_A_27_136#_c_331_n N_A_373_82#_c_414_n 0.00122897f $X=2.855 $Y=1.59
+ $X2=0 $Y2=0
cc_295 N_A_27_136#_M1003_g N_A_373_82#_c_414_n 0.00125361f $X=2.855 $Y=2.46
+ $X2=0 $Y2=0
cc_296 N_A_27_136#_c_338_n N_A_373_82#_c_414_n 0.0163973f $X=2.78 $Y=1.425 $X2=0
+ $Y2=0
cc_297 N_A_27_136#_M1003_g N_A_673_392#_c_651_n 8.04035e-19 $X=2.855 $Y=2.46
+ $X2=0 $Y2=0
cc_298 N_A_27_136#_c_342_n N_VPWR_c_778_n 0.0369382f $X=0.45 $Y=2.115 $X2=0
+ $Y2=0
cc_299 N_A_27_136#_M1003_g N_VPWR_c_779_n 0.00656069f $X=2.855 $Y=2.46 $X2=0
+ $Y2=0
cc_300 N_A_27_136#_c_342_n N_VPWR_c_783_n 0.014253f $X=0.45 $Y=2.115 $X2=0 $Y2=0
cc_301 N_A_27_136#_M1003_g N_VPWR_c_789_n 0.00392086f $X=2.855 $Y=2.46 $X2=0
+ $Y2=0
cc_302 N_A_27_136#_M1003_g N_VPWR_c_777_n 0.00500427f $X=2.855 $Y=2.46 $X2=0
+ $Y2=0
cc_303 N_A_27_136#_c_342_n N_VPWR_c_777_n 0.0172992f $X=0.45 $Y=2.115 $X2=0
+ $Y2=0
cc_304 N_A_27_136#_c_336_n N_VGND_M1017_d 0.0162931f $X=2.615 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_305 N_A_27_136#_c_336_n N_VGND_M1007_d 0.0215978f $X=2.615 $Y=0.665 $X2=0
+ $Y2=0
cc_306 N_A_27_136#_c_338_n N_VGND_M1007_d 0.0106158f $X=2.78 $Y=1.425 $X2=0
+ $Y2=0
cc_307 N_A_27_136#_c_336_n N_VGND_c_902_n 0.00345394f $X=2.615 $Y=0.665 $X2=0
+ $Y2=0
cc_308 N_A_27_136#_c_337_n N_VGND_c_902_n 0.00791634f $X=0.445 $Y=0.665 $X2=0
+ $Y2=0
cc_309 N_A_27_136#_c_334_n N_VGND_c_903_n 0.00461464f $X=3.41 $Y=1.11 $X2=0
+ $Y2=0
cc_310 N_A_27_136#_c_336_n N_VGND_c_906_n 0.0246008f $X=2.615 $Y=0.665 $X2=0
+ $Y2=0
cc_311 N_A_27_136#_c_336_n N_VGND_c_907_n 0.0262718f $X=2.615 $Y=0.665 $X2=0
+ $Y2=0
cc_312 N_A_27_136#_c_334_n N_VGND_c_908_n 0.00642663f $X=3.41 $Y=1.11 $X2=0
+ $Y2=0
cc_313 N_A_27_136#_c_336_n N_VGND_c_908_n 0.0445474f $X=2.615 $Y=0.665 $X2=0
+ $Y2=0
cc_314 N_A_27_136#_c_334_n N_VGND_c_911_n 0.00913019f $X=3.41 $Y=1.11 $X2=0
+ $Y2=0
cc_315 N_A_27_136#_c_336_n N_VGND_c_911_n 0.0521649f $X=2.615 $Y=0.665 $X2=0
+ $Y2=0
cc_316 N_A_27_136#_c_337_n N_VGND_c_911_n 0.011025f $X=0.445 $Y=0.665 $X2=0
+ $Y2=0
cc_317 N_A_373_82#_M1020_g N_A_913_406#_M1018_g 0.0427029f $X=4.275 $Y=0.58
+ $X2=0 $Y2=0
cc_318 N_A_373_82#_c_411_n N_A_913_406#_M1018_g 0.00125716f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_319 N_A_373_82#_c_412_n N_A_913_406#_M1018_g 0.0196496f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_320 N_A_373_82#_c_416_n N_A_673_392#_M1010_d 0.00114581f $X=3.155 $Y=1.925
+ $X2=0 $Y2=0
cc_321 N_A_373_82#_M1010_g N_A_673_392#_c_651_n 0.00406642f $X=3.275 $Y=2.46
+ $X2=0 $Y2=0
cc_322 N_A_373_82#_c_416_n N_A_673_392#_c_651_n 0.00737679f $X=3.155 $Y=1.925
+ $X2=0 $Y2=0
cc_323 N_A_373_82#_c_409_n N_A_673_392#_c_651_n 4.30426e-19 $X=3.32 $Y=1.635
+ $X2=0 $Y2=0
cc_324 N_A_373_82#_c_411_n N_A_673_392#_c_651_n 0.00494788f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_325 N_A_373_82#_M1010_g N_A_673_392#_c_652_n 0.00316171f $X=3.275 $Y=2.46
+ $X2=0 $Y2=0
cc_326 N_A_373_82#_c_416_n N_A_673_392#_c_652_n 0.0125405f $X=3.155 $Y=1.925
+ $X2=0 $Y2=0
cc_327 N_A_373_82#_c_411_n N_A_673_392#_c_653_n 0.0449883f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_328 N_A_373_82#_c_412_n N_A_673_392#_c_653_n 0.00440959f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_329 N_A_373_82#_c_416_n N_A_673_392#_c_654_n 0.00187356f $X=3.155 $Y=1.925
+ $X2=0 $Y2=0
cc_330 N_A_373_82#_c_417_n N_A_673_392#_c_654_n 0.0127726f $X=3.32 $Y=1.635
+ $X2=0 $Y2=0
cc_331 N_A_373_82#_c_409_n N_A_673_392#_c_654_n 7.18648e-19 $X=3.32 $Y=1.635
+ $X2=0 $Y2=0
cc_332 N_A_373_82#_c_411_n N_A_673_392#_c_654_n 0.0141411f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_333 N_A_373_82#_M1020_g N_A_673_392#_c_643_n 0.0102957f $X=4.275 $Y=0.58
+ $X2=0 $Y2=0
cc_334 N_A_373_82#_M1020_g N_A_673_392#_c_644_n 0.00848162f $X=4.275 $Y=0.58
+ $X2=0 $Y2=0
cc_335 N_A_373_82#_c_411_n N_A_673_392#_c_644_n 0.0137779f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_336 N_A_373_82#_c_412_n N_A_673_392#_c_644_n 0.00145734f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_337 N_A_373_82#_M1020_g N_A_673_392#_c_645_n 0.00270231f $X=4.275 $Y=0.58
+ $X2=0 $Y2=0
cc_338 N_A_373_82#_c_411_n N_A_673_392#_c_645_n 0.0284678f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_339 N_A_373_82#_c_412_n N_A_673_392#_c_645_n 0.00267329f $X=4.25 $Y=1.355
+ $X2=0 $Y2=0
cc_340 N_A_373_82#_c_411_n N_A_673_392#_c_647_n 0.010967f $X=4.25 $Y=1.355 $X2=0
+ $Y2=0
cc_341 N_A_373_82#_c_416_n N_VPWR_M1021_d 0.00616791f $X=3.155 $Y=1.925 $X2=0
+ $Y2=0
cc_342 N_A_373_82#_M1010_g N_VPWR_c_789_n 0.00392086f $X=3.275 $Y=2.46 $X2=0
+ $Y2=0
cc_343 N_A_373_82#_M1010_g N_VPWR_c_777_n 0.00501413f $X=3.275 $Y=2.46 $X2=0
+ $Y2=0
cc_344 N_A_373_82#_c_416_n A_589_392# 0.00230006f $X=3.155 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_345 N_A_373_82#_M1020_g N_VGND_c_898_n 0.00151928f $X=4.275 $Y=0.58 $X2=0
+ $Y2=0
cc_346 N_A_373_82#_M1020_g N_VGND_c_903_n 0.00434272f $X=4.275 $Y=0.58 $X2=0
+ $Y2=0
cc_347 N_A_373_82#_M1020_g N_VGND_c_911_n 0.00448673f $X=4.275 $Y=0.58 $X2=0
+ $Y2=0
cc_348 N_A_913_406#_c_523_n N_A_673_392#_M1008_g 0.00367488f $X=4.73 $Y=2.195
+ $X2=0 $Y2=0
cc_349 N_A_913_406#_c_524_n N_A_673_392#_M1008_g 0.0162447f $X=5.88 $Y=2.815
+ $X2=0 $Y2=0
cc_350 N_A_913_406#_c_526_n N_A_673_392#_M1008_g 0.0291822f $X=5.795 $Y=1.805
+ $X2=0 $Y2=0
cc_351 N_A_913_406#_c_514_n N_A_673_392#_M1008_g 0.00159644f $X=5.795 $Y=1.72
+ $X2=0 $Y2=0
cc_352 N_A_913_406#_c_512_n N_A_673_392#_M1002_g 0.0142421f $X=5.475 $Y=0.515
+ $X2=0 $Y2=0
cc_353 N_A_913_406#_c_513_n N_A_673_392#_M1002_g 0.00489327f $X=5.512 $Y=1.13
+ $X2=0 $Y2=0
cc_354 N_A_913_406#_c_514_n N_A_673_392#_M1002_g 0.0070337f $X=5.795 $Y=1.72
+ $X2=0 $Y2=0
cc_355 N_A_913_406#_M1018_g N_A_673_392#_c_641_n 0.0142218f $X=4.7 $Y=0.58 $X2=0
+ $Y2=0
cc_356 N_A_913_406#_c_522_n N_A_673_392#_c_641_n 0.00651642f $X=5.545 $Y=2.195
+ $X2=0 $Y2=0
cc_357 N_A_913_406#_c_513_n N_A_673_392#_c_641_n 0.00768436f $X=5.512 $Y=1.13
+ $X2=0 $Y2=0
cc_358 N_A_913_406#_c_514_n N_A_673_392#_c_641_n 0.0051522f $X=5.795 $Y=1.72
+ $X2=0 $Y2=0
cc_359 N_A_913_406#_c_526_n N_A_673_392#_c_642_n 0.00137552f $X=5.795 $Y=1.805
+ $X2=0 $Y2=0
cc_360 N_A_913_406#_c_514_n N_A_673_392#_c_642_n 0.00925024f $X=5.795 $Y=1.72
+ $X2=0 $Y2=0
cc_361 N_A_913_406#_c_519_n N_A_673_392#_c_653_n 0.00942519f $X=4.715 $Y=1.77
+ $X2=0 $Y2=0
cc_362 N_A_913_406#_c_522_n N_A_673_392#_c_653_n 0.0300742f $X=5.545 $Y=2.195
+ $X2=0 $Y2=0
cc_363 N_A_913_406#_c_523_n N_A_673_392#_c_653_n 0.00359948f $X=4.73 $Y=2.195
+ $X2=0 $Y2=0
cc_364 N_A_913_406#_c_529_n N_A_673_392#_c_653_n 0.00764166f $X=4.73 $Y=2.03
+ $X2=0 $Y2=0
cc_365 N_A_913_406#_M1018_g N_A_673_392#_c_643_n 0.00179535f $X=4.7 $Y=0.58
+ $X2=0 $Y2=0
cc_366 N_A_913_406#_M1018_g N_A_673_392#_c_644_n 0.0153705f $X=4.7 $Y=0.58 $X2=0
+ $Y2=0
cc_367 N_A_913_406#_c_519_n N_A_673_392#_c_644_n 5.25968e-19 $X=4.715 $Y=1.77
+ $X2=0 $Y2=0
cc_368 N_A_913_406#_c_512_n N_A_673_392#_c_644_n 0.0152186f $X=5.475 $Y=0.515
+ $X2=0 $Y2=0
cc_369 N_A_913_406#_c_519_n N_A_673_392#_c_646_n 0.00127151f $X=4.715 $Y=1.77
+ $X2=0 $Y2=0
cc_370 N_A_913_406#_c_522_n N_A_673_392#_c_646_n 0.0349663f $X=5.545 $Y=2.195
+ $X2=0 $Y2=0
cc_371 N_A_913_406#_c_513_n N_A_673_392#_c_646_n 0.00453021f $X=5.512 $Y=1.13
+ $X2=0 $Y2=0
cc_372 N_A_913_406#_c_514_n N_A_673_392#_c_646_n 0.0383995f $X=5.795 $Y=1.72
+ $X2=0 $Y2=0
cc_373 N_A_913_406#_M1018_g N_A_673_392#_c_647_n 0.0147644f $X=4.7 $Y=0.58 $X2=0
+ $Y2=0
cc_374 N_A_913_406#_c_513_n N_A_673_392#_c_647_n 0.00882763f $X=5.512 $Y=1.13
+ $X2=0 $Y2=0
cc_375 N_A_913_406#_c_514_n N_A_673_392#_c_647_n 0.00905133f $X=5.795 $Y=1.72
+ $X2=0 $Y2=0
cc_376 N_A_913_406#_c_524_n N_RESET_B_M1019_g 0.00976453f $X=5.88 $Y=2.815 $X2=0
+ $Y2=0
cc_377 N_A_913_406#_c_525_n N_RESET_B_M1019_g 0.0153121f $X=6.505 $Y=1.805 $X2=0
+ $Y2=0
cc_378 N_A_913_406#_c_526_n N_RESET_B_M1019_g 0.0153355f $X=5.795 $Y=1.805 $X2=0
+ $Y2=0
cc_379 N_A_913_406#_c_514_n N_RESET_B_M1019_g 0.00103957f $X=5.795 $Y=1.72 $X2=0
+ $Y2=0
cc_380 N_A_913_406#_c_515_n N_RESET_B_M1019_g 0.00416663f $X=6.68 $Y=1.485 $X2=0
+ $Y2=0
cc_381 N_A_913_406#_c_516_n N_RESET_B_M1019_g 0.00354122f $X=6.68 $Y=1.395 $X2=0
+ $Y2=0
cc_382 N_A_913_406#_c_525_n N_RESET_B_c_741_n 0.00246626f $X=6.505 $Y=1.805
+ $X2=0 $Y2=0
cc_383 N_A_913_406#_c_526_n N_RESET_B_c_741_n 9.71268e-19 $X=5.795 $Y=1.805
+ $X2=0 $Y2=0
cc_384 N_A_913_406#_c_514_n N_RESET_B_c_741_n 3.21747e-19 $X=5.795 $Y=1.72 $X2=0
+ $Y2=0
cc_385 N_A_913_406#_c_515_n N_RESET_B_c_741_n 7.91684e-19 $X=6.68 $Y=1.485 $X2=0
+ $Y2=0
cc_386 N_A_913_406#_c_516_n N_RESET_B_c_741_n 0.0149678f $X=6.68 $Y=1.395 $X2=0
+ $Y2=0
cc_387 N_A_913_406#_c_525_n N_RESET_B_c_742_n 0.0191514f $X=6.505 $Y=1.805 $X2=0
+ $Y2=0
cc_388 N_A_913_406#_c_526_n N_RESET_B_c_742_n 0.0137614f $X=5.795 $Y=1.805 $X2=0
+ $Y2=0
cc_389 N_A_913_406#_c_514_n N_RESET_B_c_742_n 0.0284564f $X=5.795 $Y=1.72 $X2=0
+ $Y2=0
cc_390 N_A_913_406#_c_515_n N_RESET_B_c_742_n 0.0165051f $X=6.68 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_A_913_406#_c_516_n N_RESET_B_c_742_n 2.8064e-19 $X=6.68 $Y=1.395 $X2=0
+ $Y2=0
cc_392 N_A_913_406#_c_512_n N_RESET_B_c_743_n 0.00309061f $X=5.475 $Y=0.515
+ $X2=0 $Y2=0
cc_393 N_A_913_406#_c_522_n N_VPWR_M1005_d 0.00629756f $X=5.545 $Y=2.195 $X2=0
+ $Y2=0
cc_394 N_A_913_406#_c_525_n N_VPWR_M1019_d 0.00492793f $X=6.505 $Y=1.805 $X2=0
+ $Y2=0
cc_395 N_A_913_406#_c_515_n N_VPWR_M1019_d 0.00366578f $X=6.68 $Y=1.485 $X2=0
+ $Y2=0
cc_396 N_A_913_406#_M1006_g N_VPWR_c_780_n 0.0074535f $X=7.145 $Y=2.4 $X2=0
+ $Y2=0
cc_397 N_A_913_406#_c_525_n N_VPWR_c_780_n 0.0149335f $X=6.505 $Y=1.805 $X2=0
+ $Y2=0
cc_398 N_A_913_406#_c_526_n N_VPWR_c_780_n 0.0499033f $X=5.795 $Y=1.805 $X2=0
+ $Y2=0
cc_399 N_A_913_406#_c_515_n N_VPWR_c_780_n 0.0128156f $X=6.68 $Y=1.485 $X2=0
+ $Y2=0
cc_400 N_A_913_406#_c_516_n N_VPWR_c_780_n 6.19355e-19 $X=6.68 $Y=1.395 $X2=0
+ $Y2=0
cc_401 N_A_913_406#_M1009_g N_VPWR_c_782_n 0.00688324f $X=7.595 $Y=2.4 $X2=0
+ $Y2=0
cc_402 N_A_913_406#_c_524_n N_VPWR_c_786_n 0.0144922f $X=5.88 $Y=2.815 $X2=0
+ $Y2=0
cc_403 N_A_913_406#_M1006_g N_VPWR_c_787_n 0.00349816f $X=7.145 $Y=2.4 $X2=0
+ $Y2=0
cc_404 N_A_913_406#_M1009_g N_VPWR_c_787_n 0.005209f $X=7.595 $Y=2.4 $X2=0 $Y2=0
cc_405 N_A_913_406#_M1005_g N_VPWR_c_789_n 0.00562069f $X=4.655 $Y=2.73 $X2=0
+ $Y2=0
cc_406 N_A_913_406#_M1005_g N_VPWR_c_790_n 0.0235206f $X=4.655 $Y=2.73 $X2=0
+ $Y2=0
cc_407 N_A_913_406#_c_522_n N_VPWR_c_790_n 0.0455143f $X=5.545 $Y=2.195 $X2=0
+ $Y2=0
cc_408 N_A_913_406#_c_523_n N_VPWR_c_790_n 0.00328725f $X=4.73 $Y=2.195 $X2=0
+ $Y2=0
cc_409 N_A_913_406#_c_524_n N_VPWR_c_790_n 0.0140432f $X=5.88 $Y=2.815 $X2=0
+ $Y2=0
cc_410 N_A_913_406#_M1005_g N_VPWR_c_777_n 0.00539454f $X=4.655 $Y=2.73 $X2=0
+ $Y2=0
cc_411 N_A_913_406#_M1006_g N_VPWR_c_777_n 0.00434525f $X=7.145 $Y=2.4 $X2=0
+ $Y2=0
cc_412 N_A_913_406#_M1009_g N_VPWR_c_777_n 0.00985527f $X=7.595 $Y=2.4 $X2=0
+ $Y2=0
cc_413 N_A_913_406#_c_524_n N_VPWR_c_777_n 0.0118826f $X=5.88 $Y=2.815 $X2=0
+ $Y2=0
cc_414 N_A_913_406#_M1004_g N_Q_c_863_n 0.0232839f $X=7.155 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A_913_406#_M1013_g N_Q_c_863_n 0.0193613f $X=7.585 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A_913_406#_M1004_g N_Q_c_864_n 7.75299e-19 $X=7.155 $Y=0.74 $X2=0 $Y2=0
cc_417 N_A_913_406#_c_507_n N_Q_c_864_n 0.0092514f $X=7.505 $Y=1.395 $X2=0 $Y2=0
cc_418 N_A_913_406#_M1013_g N_Q_c_864_n 7.75299e-19 $X=7.585 $Y=0.74 $X2=0 $Y2=0
cc_419 N_A_913_406#_c_510_n N_Q_c_864_n 0.0041437f $X=7.145 $Y=1.395 $X2=0 $Y2=0
cc_420 N_A_913_406#_c_511_n N_Q_c_864_n 0.00663376f $X=7.595 $Y=1.395 $X2=0
+ $Y2=0
cc_421 N_A_913_406#_c_515_n N_Q_c_864_n 0.00619468f $X=6.68 $Y=1.485 $X2=0 $Y2=0
cc_422 N_A_913_406#_M1006_g Q 0.031404f $X=7.145 $Y=2.4 $X2=0 $Y2=0
cc_423 N_A_913_406#_M1009_g Q 0.0106338f $X=7.595 $Y=2.4 $X2=0 $Y2=0
cc_424 N_A_913_406#_c_504_n N_Q_c_867_n 0.0070804f $X=7.055 $Y=1.395 $X2=0 $Y2=0
cc_425 N_A_913_406#_M1006_g N_Q_c_867_n 0.0207518f $X=7.145 $Y=2.4 $X2=0 $Y2=0
cc_426 N_A_913_406#_c_507_n N_Q_c_867_n 2.91044e-19 $X=7.505 $Y=1.395 $X2=0
+ $Y2=0
cc_427 N_A_913_406#_M1009_g N_Q_c_867_n 0.00426872f $X=7.595 $Y=2.4 $X2=0 $Y2=0
cc_428 N_A_913_406#_c_515_n N_Q_c_867_n 0.00632434f $X=6.68 $Y=1.485 $X2=0 $Y2=0
cc_429 N_A_913_406#_M1006_g N_Q_c_865_n 0.00390202f $X=7.145 $Y=2.4 $X2=0 $Y2=0
cc_430 N_A_913_406#_M1009_g N_Q_c_865_n 0.0178406f $X=7.595 $Y=2.4 $X2=0 $Y2=0
cc_431 N_A_913_406#_c_515_n N_Q_c_865_n 0.00420462f $X=6.68 $Y=1.485 $X2=0 $Y2=0
cc_432 N_A_913_406#_M1018_g N_VGND_c_898_n 0.0111821f $X=4.7 $Y=0.58 $X2=0 $Y2=0
cc_433 N_A_913_406#_c_512_n N_VGND_c_898_n 0.0225979f $X=5.475 $Y=0.515 $X2=0
+ $Y2=0
cc_434 N_A_913_406#_c_504_n N_VGND_c_899_n 0.006447f $X=7.055 $Y=1.395 $X2=0
+ $Y2=0
cc_435 N_A_913_406#_M1004_g N_VGND_c_899_n 0.0163364f $X=7.155 $Y=0.74 $X2=0
+ $Y2=0
cc_436 N_A_913_406#_c_512_n N_VGND_c_899_n 0.0258773f $X=5.475 $Y=0.515 $X2=0
+ $Y2=0
cc_437 N_A_913_406#_c_515_n N_VGND_c_899_n 0.018142f $X=6.68 $Y=1.485 $X2=0
+ $Y2=0
cc_438 N_A_913_406#_c_516_n N_VGND_c_899_n 0.00242479f $X=6.68 $Y=1.395 $X2=0
+ $Y2=0
cc_439 N_A_913_406#_M1013_g N_VGND_c_901_n 0.0184907f $X=7.585 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A_913_406#_M1018_g N_VGND_c_903_n 0.00383152f $X=4.7 $Y=0.58 $X2=0
+ $Y2=0
cc_441 N_A_913_406#_c_512_n N_VGND_c_904_n 0.0176863f $X=5.475 $Y=0.515 $X2=0
+ $Y2=0
cc_442 N_A_913_406#_M1004_g N_VGND_c_905_n 0.00434272f $X=7.155 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_913_406#_M1013_g N_VGND_c_905_n 0.00434272f $X=7.585 $Y=0.74 $X2=0
+ $Y2=0
cc_444 N_A_913_406#_M1018_g N_VGND_c_911_n 0.00386109f $X=4.7 $Y=0.58 $X2=0
+ $Y2=0
cc_445 N_A_913_406#_M1004_g N_VGND_c_911_n 0.00825059f $X=7.155 $Y=0.74 $X2=0
+ $Y2=0
cc_446 N_A_913_406#_M1013_g N_VGND_c_911_n 0.00823962f $X=7.585 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_913_406#_c_512_n N_VGND_c_911_n 0.0144066f $X=5.475 $Y=0.515 $X2=0
+ $Y2=0
cc_448 N_A_673_392#_c_642_n N_RESET_B_M1019_g 0.0219346f $X=5.555 $Y=1.35 $X2=0
+ $Y2=0
cc_449 N_A_673_392#_M1002_g N_RESET_B_c_741_n 0.0174816f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_450 N_A_673_392#_c_642_n N_RESET_B_c_741_n 0.00278721f $X=5.555 $Y=1.35 $X2=0
+ $Y2=0
cc_451 N_A_673_392#_M1002_g N_RESET_B_c_742_n 0.00205529f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_673_392#_c_642_n N_RESET_B_c_742_n 3.47714e-19 $X=5.555 $Y=1.35 $X2=0
+ $Y2=0
cc_453 N_A_673_392#_M1002_g N_RESET_B_c_743_n 0.0482898f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_454 N_A_673_392#_c_646_n N_VPWR_M1005_d 9.31261e-19 $X=5.21 $Y=1.515 $X2=0
+ $Y2=0
cc_455 N_A_673_392#_M1008_g N_VPWR_c_786_n 0.0053223f $X=5.645 $Y=2.4 $X2=0
+ $Y2=0
cc_456 N_A_673_392#_M1008_g N_VPWR_c_790_n 0.00593313f $X=5.645 $Y=2.4 $X2=0
+ $Y2=0
cc_457 N_A_673_392#_M1008_g N_VPWR_c_777_n 0.0102337f $X=5.645 $Y=2.4 $X2=0
+ $Y2=0
cc_458 N_A_673_392#_M1002_g N_VGND_c_898_n 0.00335086f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_459 N_A_673_392#_c_643_n N_VGND_c_898_n 0.00984031f $X=4.06 $Y=0.58 $X2=0
+ $Y2=0
cc_460 N_A_673_392#_c_644_n N_VGND_c_898_n 0.0247482f $X=4.97 $Y=0.935 $X2=0
+ $Y2=0
cc_461 N_A_673_392#_M1002_g N_VGND_c_899_n 0.00234534f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_462 N_A_673_392#_c_643_n N_VGND_c_903_n 0.0145482f $X=4.06 $Y=0.58 $X2=0
+ $Y2=0
cc_463 N_A_673_392#_M1002_g N_VGND_c_904_n 0.00349296f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_673_392#_c_643_n N_VGND_c_908_n 6.72815e-19 $X=4.06 $Y=0.58 $X2=0
+ $Y2=0
cc_465 N_A_673_392#_M1002_g N_VGND_c_911_n 0.00550827f $X=5.69 $Y=0.74 $X2=0
+ $Y2=0
cc_466 N_A_673_392#_c_643_n N_VGND_c_911_n 0.0119922f $X=4.06 $Y=0.58 $X2=0
+ $Y2=0
cc_467 N_A_673_392#_c_644_n N_VGND_c_911_n 0.019671f $X=4.97 $Y=0.935 $X2=0
+ $Y2=0
cc_468 N_RESET_B_M1019_g N_VPWR_c_780_n 0.0253158f $X=6.105 $Y=2.4 $X2=0 $Y2=0
cc_469 N_RESET_B_M1019_g N_VPWR_c_786_n 0.005209f $X=6.105 $Y=2.4 $X2=0 $Y2=0
cc_470 N_RESET_B_M1019_g N_VPWR_c_777_n 0.00988702f $X=6.105 $Y=2.4 $X2=0 $Y2=0
cc_471 N_RESET_B_M1019_g N_Q_c_867_n 0.00586595f $X=6.105 $Y=2.4 $X2=0 $Y2=0
cc_472 N_RESET_B_c_741_n N_VGND_c_899_n 9.03586e-19 $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_473 N_RESET_B_c_742_n N_VGND_c_899_n 0.0124443f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_474 N_RESET_B_c_743_n N_VGND_c_899_n 0.0161122f $X=6.14 $Y=1.22 $X2=0 $Y2=0
cc_475 N_RESET_B_c_743_n N_VGND_c_904_n 0.00383152f $X=6.14 $Y=1.22 $X2=0 $Y2=0
cc_476 N_RESET_B_c_743_n N_VGND_c_911_n 0.0075725f $X=6.14 $Y=1.22 $X2=0 $Y2=0
cc_477 N_VPWR_M1019_d Q 0.0099171f $X=6.195 $Y=1.84 $X2=0 $Y2=0
cc_478 N_VPWR_c_787_n Q 0.0300745f $X=7.705 $Y=3.33 $X2=0 $Y2=0
cc_479 N_VPWR_c_777_n Q 0.0244021f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_480 N_VPWR_M1019_d N_Q_c_867_n 0.00567897f $X=6.195 $Y=1.84 $X2=0 $Y2=0
cc_481 N_VPWR_c_780_n N_Q_c_867_n 0.0705528f $X=6.485 $Y=2.225 $X2=0 $Y2=0
cc_482 N_VPWR_c_782_n N_Q_c_867_n 0.0502658f $X=7.875 $Y=1.985 $X2=0 $Y2=0
cc_483 N_Q_c_863_n N_VGND_c_899_n 0.0256468f $X=7.37 $Y=0.515 $X2=0 $Y2=0
cc_484 N_Q_c_863_n N_VGND_c_901_n 0.0308485f $X=7.37 $Y=0.515 $X2=0 $Y2=0
cc_485 N_Q_c_863_n N_VGND_c_905_n 0.0144922f $X=7.37 $Y=0.515 $X2=0 $Y2=0
cc_486 N_Q_c_863_n N_VGND_c_911_n 0.0118826f $X=7.37 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__inv_2.pxi.spice
* Created: Wed Sep  2 12:10:57 2020
* 
x_PM_SKY130_FD_SC_MS__INV_2%A N_A_M1000_g N_A_M1002_g N_A_c_31_n N_A_M1001_g
+ N_A_M1003_g N_A_c_34_n A N_A_c_35_n N_A_c_36_n PM_SKY130_FD_SC_MS__INV_2%A
x_PM_SKY130_FD_SC_MS__INV_2%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_c_69_n
+ N_VPWR_c_70_n N_VPWR_c_71_n N_VPWR_c_72_n VPWR N_VPWR_c_73_n N_VPWR_c_68_n
+ PM_SKY130_FD_SC_MS__INV_2%VPWR
x_PM_SKY130_FD_SC_MS__INV_2%Y N_Y_M1002_d N_Y_M1000_d Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_MS__INV_2%Y
x_PM_SKY130_FD_SC_MS__INV_2%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_c_111_n
+ N_VGND_c_112_n N_VGND_c_113_n N_VGND_c_114_n VGND N_VGND_c_115_n
+ N_VGND_c_116_n PM_SKY130_FD_SC_MS__INV_2%VGND
cc_1 VNB N_A_M1000_g 0.00186993f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A_M1002_g 0.0266858f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_3 VNB N_A_c_31_n 0.00970685f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.375
cc_4 VNB N_A_M1001_g 0.0167069f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_5 VNB N_A_M1003_g 0.0260209f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_6 VNB N_A_c_34_n 0.0122617f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.375
cc_7 VNB N_A_c_35_n 0.00655144f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_8 VNB N_A_c_36_n 0.0555854f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.465
cc_9 VNB N_VPWR_c_68_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_10 VNB Y 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_11 VNB Y 8.14549e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB Y 0.00291429f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.375
cc_13 VNB N_VGND_c_111_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_14 VNB N_VGND_c_112_n 0.0419252f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.375
cc_15 VNB N_VGND_c_113_n 0.0108375f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.45
cc_16 VNB N_VGND_c_114_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_17 VNB N_VGND_c_115_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_18 VNB N_VGND_c_116_n 0.116359f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.465
cc_19 VPB N_A_M1000_g 0.0270574f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_20 VPB N_A_M1001_g 0.0274176f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_21 VPB N_A_c_35_n 0.0072578f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_22 VPB N_VPWR_c_69_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_23 VPB N_VPWR_c_70_n 0.0482811f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.375
cc_24 VPB N_VPWR_c_71_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_25 VPB N_VPWR_c_72_n 0.0642732f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.3
cc_26 VPB N_VPWR_c_73_n 0.0182519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_68_n 0.048697f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_28 VPB Y 0.00396093f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.375
cc_29 N_A_M1000_g N_VPWR_c_70_n 0.0173373f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_30 N_A_M1001_g N_VPWR_c_70_n 6.42904e-19 $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_31 N_A_c_35_n N_VPWR_c_70_n 0.0266029f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_32 N_A_c_36_n N_VPWR_c_70_n 0.00152096f $X=0.585 $Y=1.465 $X2=0 $Y2=0
cc_33 N_A_M1001_g N_VPWR_c_72_n 0.00517083f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_34 N_A_M1000_g N_VPWR_c_73_n 0.00460063f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_35 N_A_M1001_g N_VPWR_c_73_n 0.00515235f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_36 N_A_M1000_g N_VPWR_c_68_n 0.00908554f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_37 N_A_M1001_g N_VPWR_c_68_n 0.00967629f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_38 N_A_M1002_g Y 0.00788704f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_39 N_A_M1003_g Y 0.00788704f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_40 N_A_M1002_g Y 0.00327512f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_41 N_A_M1003_g Y 0.00202916f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_42 N_A_M1002_g Y 0.00465421f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_43 N_A_c_31_n Y 0.0101905f $X=0.855 $Y=1.375 $X2=0 $Y2=0
cc_44 N_A_M1001_g Y 0.0355803f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_45 N_A_M1003_g Y 0.00881083f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_46 N_A_c_34_n Y 0.00658953f $X=0.945 $Y=1.375 $X2=0 $Y2=0
cc_47 N_A_c_35_n Y 0.0369047f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_48 N_A_c_36_n Y 0.00483978f $X=0.585 $Y=1.465 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_VGND_c_112_n 0.00647412f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_50 N_A_c_35_n N_VGND_c_112_n 0.0215684f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_51 N_A_c_36_n N_VGND_c_112_n 0.00196285f $X=0.585 $Y=1.465 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_VGND_c_114_n 0.00647412f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_53 N_A_M1002_g N_VGND_c_115_n 0.00434272f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_54 N_A_M1003_g N_VGND_c_115_n 0.00434272f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_55 N_A_M1002_g N_VGND_c_116_n 0.00823992f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_56 N_A_M1003_g N_VGND_c_116_n 0.00823959f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_57 N_VPWR_c_70_n Y 0.0394212f $X=0.27 $Y=2.115 $X2=0 $Y2=0
cc_58 N_VPWR_c_72_n Y 0.0395076f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_59 N_VPWR_c_73_n Y 0.0125261f $X=1.085 $Y=3.33 $X2=0 $Y2=0
cc_60 N_VPWR_c_68_n Y 0.0102881f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_61 Y N_VGND_c_112_n 0.0293763f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_62 Y N_VGND_c_114_n 0.0293763f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_63 Y N_VGND_c_115_n 0.0144922f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_64 Y N_VGND_c_116_n 0.0118826f $X=0.635 $Y=0.47 $X2=0 $Y2=0

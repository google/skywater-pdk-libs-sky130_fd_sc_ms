* File: sky130_fd_sc_ms__einvn_4.pxi.spice
* Created: Wed Sep  2 12:08:25 2020
* 
x_PM_SKY130_FD_SC_MS__EINVN_4%TE_B N_TE_B_M1015_g N_TE_B_c_109_n N_TE_B_M1014_g
+ N_TE_B_c_100_n N_TE_B_c_111_n N_TE_B_M1000_g N_TE_B_c_101_n N_TE_B_c_113_n
+ N_TE_B_M1002_g N_TE_B_c_102_n N_TE_B_c_115_n N_TE_B_M1004_g N_TE_B_c_103_n
+ N_TE_B_c_117_n N_TE_B_M1005_g N_TE_B_c_104_n N_TE_B_c_105_n N_TE_B_c_106_n
+ TE_B N_TE_B_c_107_n N_TE_B_c_108_n PM_SKY130_FD_SC_MS__EINVN_4%TE_B
x_PM_SKY130_FD_SC_MS__EINVN_4%A_114_74# N_A_114_74#_M1015_d N_A_114_74#_M1014_d
+ N_A_114_74#_c_194_n N_A_114_74#_c_195_n N_A_114_74#_c_196_n
+ N_A_114_74#_M1003_g N_A_114_74#_c_197_n N_A_114_74#_c_198_n
+ N_A_114_74#_M1006_g N_A_114_74#_c_199_n N_A_114_74#_c_200_n
+ N_A_114_74#_M1013_g N_A_114_74#_c_201_n N_A_114_74#_c_202_n
+ N_A_114_74#_M1017_g N_A_114_74#_c_203_n N_A_114_74#_c_204_n
+ N_A_114_74#_c_205_n N_A_114_74#_c_206_n N_A_114_74#_c_207_n
+ N_A_114_74#_c_208_n PM_SKY130_FD_SC_MS__EINVN_4%A_114_74#
x_PM_SKY130_FD_SC_MS__EINVN_4%A N_A_c_289_n N_A_M1008_g N_A_c_283_n N_A_M1001_g
+ N_A_c_290_n N_A_M1009_g N_A_c_284_n N_A_M1007_g N_A_c_291_n N_A_M1010_g
+ N_A_c_285_n N_A_M1012_g N_A_c_292_n N_A_M1011_g N_A_c_286_n N_A_M1016_g A A
+ N_A_c_288_n PM_SKY130_FD_SC_MS__EINVN_4%A
x_PM_SKY130_FD_SC_MS__EINVN_4%VPWR N_VPWR_M1014_s N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n VPWR
+ N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_367_n N_VPWR_c_376_n
+ N_VPWR_c_377_n PM_SKY130_FD_SC_MS__EINVN_4%VPWR
x_PM_SKY130_FD_SC_MS__EINVN_4%A_241_368# N_A_241_368#_M1000_s
+ N_A_241_368#_M1002_s N_A_241_368#_M1005_s N_A_241_368#_M1009_s
+ N_A_241_368#_M1011_s N_A_241_368#_c_432_n N_A_241_368#_c_428_n
+ N_A_241_368#_c_429_n N_A_241_368#_c_433_n N_A_241_368#_c_430_n
+ N_A_241_368#_c_434_n N_A_241_368#_c_435_n N_A_241_368#_c_436_n
+ N_A_241_368#_c_475_n N_A_241_368#_c_437_n N_A_241_368#_c_438_n
+ N_A_241_368#_c_431_n N_A_241_368#_c_439_n
+ PM_SKY130_FD_SC_MS__EINVN_4%A_241_368#
x_PM_SKY130_FD_SC_MS__EINVN_4%Z N_Z_M1001_s N_Z_M1012_s N_Z_M1008_d N_Z_M1010_d
+ N_Z_c_518_n N_Z_c_522_n N_Z_c_527_n N_Z_c_531_n N_Z_c_516_n N_Z_c_537_n Z
+ N_Z_c_517_n PM_SKY130_FD_SC_MS__EINVN_4%Z
x_PM_SKY130_FD_SC_MS__EINVN_4%VGND N_VGND_M1015_s N_VGND_M1003_s N_VGND_M1013_s
+ N_VGND_c_565_n N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n
+ N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n VGND N_VGND_c_573_n
+ N_VGND_c_574_n PM_SKY130_FD_SC_MS__EINVN_4%VGND
x_PM_SKY130_FD_SC_MS__EINVN_4%A_281_74# N_A_281_74#_M1003_d N_A_281_74#_M1006_d
+ N_A_281_74#_M1017_d N_A_281_74#_M1007_d N_A_281_74#_M1016_d
+ N_A_281_74#_c_626_n N_A_281_74#_c_627_n N_A_281_74#_c_628_n
+ N_A_281_74#_c_629_n N_A_281_74#_c_630_n N_A_281_74#_c_631_n
+ N_A_281_74#_c_632_n N_A_281_74#_c_633_n N_A_281_74#_c_634_n
+ N_A_281_74#_c_635_n N_A_281_74#_c_660_n N_A_281_74#_c_636_n
+ PM_SKY130_FD_SC_MS__EINVN_4%A_281_74#
cc_1 VNB N_TE_B_M1015_g 0.0294944f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_TE_B_c_100_n 0.0235348f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.65
cc_3 VNB N_TE_B_c_101_n 0.0055238f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.65
cc_4 VNB N_TE_B_c_102_n 0.00546594f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.65
cc_5 VNB N_TE_B_c_103_n 0.0113338f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.65
cc_6 VNB N_TE_B_c_104_n 0.00370683f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.65
cc_7 VNB N_TE_B_c_105_n 0.00369526f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.65
cc_8 VNB N_TE_B_c_106_n 0.00370683f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.65
cc_9 VNB N_TE_B_c_107_n 0.00440334f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_10 VNB N_TE_B_c_108_n 0.0577209f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.512
cc_11 VNB N_A_114_74#_c_194_n 0.0208628f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_12 VNB N_A_114_74#_c_195_n 0.0139628f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.65
cc_13 VNB N_A_114_74#_c_196_n 0.0166447f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.65
cc_14 VNB N_A_114_74#_c_197_n 0.0122635f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=2.4
cc_15 VNB N_A_114_74#_c_198_n 0.0143129f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.65
cc_16 VNB N_A_114_74#_c_199_n 0.0122635f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.4
cc_17 VNB N_A_114_74#_c_200_n 0.0143129f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.65
cc_18 VNB N_A_114_74#_c_201_n 0.0200435f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.4
cc_19 VNB N_A_114_74#_c_202_n 0.0145547f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=1.65
cc_20 VNB N_A_114_74#_c_203_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.65
cc_21 VNB N_A_114_74#_c_204_n 0.00511435f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.65
cc_22 VNB N_A_114_74#_c_205_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.65
cc_23 VNB N_A_114_74#_c_206_n 0.0146868f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_114_74#_c_207_n 0.0066218f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.512
cc_25 VNB N_A_114_74#_c_208_n 0.0711714f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.512
cc_26 VNB N_A_c_283_n 0.0157318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_284_n 0.0161778f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.725
cc_28 VNB N_A_c_285_n 0.0159974f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.4
cc_29 VNB N_A_c_286_n 0.0207336f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.4
cc_30 VNB A 0.0256668f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=2.4
cc_31 VNB N_A_c_288_n 0.122555f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.512
cc_32 VNB N_VPWR_c_367_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_241_368#_c_428_n 0.00395162f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.4
cc_34 VNB N_A_241_368#_c_429_n 0.00301433f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.65
cc_35 VNB N_A_241_368#_c_430_n 0.00757f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.65
cc_36 VNB N_A_241_368#_c_431_n 0.00151865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Z_c_516_n 4.62656e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_Z_c_517_n 0.00122353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_565_n 0.010678f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.725
cc_40 VNB N_VGND_c_566_n 0.0420905f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=2.4
cc_41 VNB N_VGND_c_567_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=2.4
cc_42 VNB N_VGND_c_568_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.725
cc_43 VNB N_VGND_c_569_n 0.0381462f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.65
cc_44 VNB N_VGND_c_570_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=1.65
cc_45 VNB N_VGND_c_571_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=2.4
cc_46 VNB N_VGND_c_572_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=2.4
cc_47 VNB N_VGND_c_573_n 0.0552148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_574_n 0.305559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_281_74#_c_626_n 0.00221876f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.65
cc_50 VNB N_A_281_74#_c_627_n 0.00627739f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.725
cc_51 VNB N_A_281_74#_c_628_n 2.75804e-19 $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=2.4
cc_52 VNB N_A_281_74#_c_629_n 0.00229766f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=1.65
cc_53 VNB N_A_281_74#_c_630_n 0.0106645f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=2.4
cc_54 VNB N_A_281_74#_c_631_n 0.00251555f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.65
cc_55 VNB N_A_281_74#_c_632_n 2.66637e-19 $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.65
cc_56 VNB N_A_281_74#_c_633_n 0.00304162f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.65
cc_57 VNB N_A_281_74#_c_634_n 0.01171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_281_74#_c_635_n 0.0226357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_281_74#_c_636_n 0.00105952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_TE_B_c_109_n 0.0266811f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.725
cc_61 VPB N_TE_B_c_100_n 0.0286071f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=1.65
cc_62 VPB N_TE_B_c_111_n 0.0221933f $X=-0.19 $Y=1.66 $X2=1.575 $Y2=1.725
cc_63 VPB N_TE_B_c_101_n 0.00378507f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=1.65
cc_64 VPB N_TE_B_c_113_n 0.0184192f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=1.725
cc_65 VPB N_TE_B_c_102_n 0.0044263f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.65
cc_66 VPB N_TE_B_c_115_n 0.0186711f $X=-0.19 $Y=1.66 $X2=2.475 $Y2=1.725
cc_67 VPB N_TE_B_c_103_n 0.00728504f $X=-0.19 $Y=1.66 $X2=2.885 $Y2=1.65
cc_68 VPB N_TE_B_c_117_n 0.0185402f $X=-0.19 $Y=1.66 $X2=2.975 $Y2=1.725
cc_69 VPB N_TE_B_c_104_n 0.00124171f $X=-0.19 $Y=1.66 $X2=1.575 $Y2=1.65
cc_70 VPB N_TE_B_c_105_n 0.00124171f $X=-0.19 $Y=1.66 $X2=2.025 $Y2=1.65
cc_71 VPB N_TE_B_c_106_n 0.00124171f $X=-0.19 $Y=1.66 $X2=2.475 $Y2=1.65
cc_72 VPB N_TE_B_c_107_n 0.00780381f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_73 VPB N_TE_B_c_108_n 0.017666f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.512
cc_74 VPB N_A_114_74#_c_207_n 0.0135911f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.512
cc_75 VPB N_A_c_289_n 0.017773f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_76 VPB N_A_c_290_n 0.0170653f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_77 VPB N_A_c_291_n 0.0170653f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=1.65
cc_78 VPB N_A_c_292_n 0.0227957f $X=-0.19 $Y=1.66 $X2=2.115 $Y2=1.65
cc_79 VPB N_A_c_288_n 0.0302139f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.512
cc_80 VPB N_VPWR_c_368_n 0.012566f $X=-0.19 $Y=1.66 $X2=1.575 $Y2=1.725
cc_81 VPB N_VPWR_c_369_n 0.0495179f $X=-0.19 $Y=1.66 $X2=1.575 $Y2=2.4
cc_82 VPB N_VPWR_c_370_n 0.00645399f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.65
cc_83 VPB N_VPWR_c_371_n 0.00751209f $X=-0.19 $Y=1.66 $X2=2.565 $Y2=1.65
cc_84 VPB N_VPWR_c_372_n 0.0337833f $X=-0.19 $Y=1.66 $X2=2.475 $Y2=1.65
cc_85 VPB N_VPWR_c_373_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_86 VPB N_VPWR_c_374_n 0.0583197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_367_n 0.0824929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_376_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_377_n 0.0061237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_241_368#_c_432_n 0.0142346f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.65
cc_91 VPB N_A_241_368#_c_433_n 0.00304337f $X=-0.19 $Y=1.66 $X2=2.975 $Y2=2.4
cc_92 VPB N_A_241_368#_c_434_n 0.00133034f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_93 VPB N_A_241_368#_c_435_n 0.0026202f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.512
cc_94 VPB N_A_241_368#_c_436_n 0.00159425f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.512
cc_95 VPB N_A_241_368#_c_437_n 0.0119149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_241_368#_c_438_n 0.0425896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_241_368#_c_439_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 N_TE_B_c_104_n N_A_114_74#_c_194_n 0.0163574f $X=1.575 $Y=1.65 $X2=0 $Y2=0
cc_99 N_TE_B_c_100_n N_A_114_74#_c_195_n 0.0163574f $X=1.485 $Y=1.65 $X2=0 $Y2=0
cc_100 N_TE_B_c_108_n N_A_114_74#_c_195_n 0.00138455f $X=0.655 $Y=1.512 $X2=0
+ $Y2=0
cc_101 N_TE_B_c_105_n N_A_114_74#_c_197_n 0.0163574f $X=2.025 $Y=1.65 $X2=0
+ $Y2=0
cc_102 N_TE_B_c_106_n N_A_114_74#_c_199_n 0.0163574f $X=2.475 $Y=1.65 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_101_n N_A_114_74#_c_203_n 0.0163574f $X=1.935 $Y=1.65 $X2=0
+ $Y2=0
cc_104 N_TE_B_c_102_n N_A_114_74#_c_204_n 0.0163574f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_105 N_TE_B_c_103_n N_A_114_74#_c_205_n 0.0163574f $X=2.885 $Y=1.65 $X2=0
+ $Y2=0
cc_106 N_TE_B_M1015_g N_A_114_74#_c_206_n 0.0183768f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_107 N_TE_B_c_100_n N_A_114_74#_c_206_n 0.00181554f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_108 N_TE_B_c_107_n N_A_114_74#_c_206_n 7.97299e-19 $X=0.29 $Y=1.465 $X2=0
+ $Y2=0
cc_109 N_TE_B_c_108_n N_A_114_74#_c_206_n 0.00371785f $X=0.655 $Y=1.512 $X2=0
+ $Y2=0
cc_110 N_TE_B_c_109_n N_A_114_74#_c_207_n 0.0249979f $X=0.565 $Y=1.725 $X2=0
+ $Y2=0
cc_111 N_TE_B_c_100_n N_A_114_74#_c_207_n 0.0189941f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_112 N_TE_B_c_107_n N_A_114_74#_c_207_n 0.0354205f $X=0.29 $Y=1.465 $X2=0
+ $Y2=0
cc_113 N_TE_B_c_108_n N_A_114_74#_c_207_n 0.0120559f $X=0.655 $Y=1.512 $X2=0
+ $Y2=0
cc_114 N_TE_B_M1015_g N_A_114_74#_c_208_n 0.0180863f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_115 N_TE_B_c_117_n N_A_c_289_n 0.0101256f $X=2.975 $Y=1.725 $X2=-0.19
+ $Y2=-0.245
cc_116 N_TE_B_c_103_n N_A_c_288_n 0.0101256f $X=2.885 $Y=1.65 $X2=0 $Y2=0
cc_117 N_TE_B_c_109_n N_VPWR_c_369_n 0.00501904f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_118 N_TE_B_c_107_n N_VPWR_c_369_n 0.0219684f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_119 N_TE_B_c_108_n N_VPWR_c_369_n 0.0016728f $X=0.655 $Y=1.512 $X2=0 $Y2=0
cc_120 N_TE_B_c_111_n N_VPWR_c_370_n 0.0218717f $X=1.575 $Y=1.725 $X2=0 $Y2=0
cc_121 N_TE_B_c_101_n N_VPWR_c_370_n 0.00197117f $X=1.935 $Y=1.65 $X2=0 $Y2=0
cc_122 N_TE_B_c_113_n N_VPWR_c_370_n 0.00202886f $X=2.025 $Y=1.725 $X2=0 $Y2=0
cc_123 N_TE_B_c_113_n N_VPWR_c_371_n 7.38193e-19 $X=2.025 $Y=1.725 $X2=0 $Y2=0
cc_124 N_TE_B_c_115_n N_VPWR_c_371_n 0.0192368f $X=2.475 $Y=1.725 $X2=0 $Y2=0
cc_125 N_TE_B_c_103_n N_VPWR_c_371_n 0.00306626f $X=2.885 $Y=1.65 $X2=0 $Y2=0
cc_126 N_TE_B_c_117_n N_VPWR_c_371_n 0.00185284f $X=2.975 $Y=1.725 $X2=0 $Y2=0
cc_127 N_TE_B_c_109_n N_VPWR_c_372_n 0.005209f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_128 N_TE_B_c_111_n N_VPWR_c_372_n 0.00460063f $X=1.575 $Y=1.725 $X2=0 $Y2=0
cc_129 N_TE_B_c_113_n N_VPWR_c_373_n 0.005209f $X=2.025 $Y=1.725 $X2=0 $Y2=0
cc_130 N_TE_B_c_115_n N_VPWR_c_373_n 0.00460063f $X=2.475 $Y=1.725 $X2=0 $Y2=0
cc_131 N_TE_B_c_117_n N_VPWR_c_374_n 0.00517089f $X=2.975 $Y=1.725 $X2=0 $Y2=0
cc_132 N_TE_B_c_109_n N_VPWR_c_367_n 0.00991332f $X=0.565 $Y=1.725 $X2=0 $Y2=0
cc_133 N_TE_B_c_111_n N_VPWR_c_367_n 0.00913687f $X=1.575 $Y=1.725 $X2=0 $Y2=0
cc_134 N_TE_B_c_113_n N_VPWR_c_367_n 0.00982266f $X=2.025 $Y=1.725 $X2=0 $Y2=0
cc_135 N_TE_B_c_115_n N_VPWR_c_367_n 0.00908554f $X=2.475 $Y=1.725 $X2=0 $Y2=0
cc_136 N_TE_B_c_117_n N_VPWR_c_367_n 0.00977404f $X=2.975 $Y=1.725 $X2=0 $Y2=0
cc_137 N_TE_B_c_109_n N_A_241_368#_c_432_n 0.00246536f $X=0.565 $Y=1.725 $X2=0
+ $Y2=0
cc_138 N_TE_B_c_100_n N_A_241_368#_c_432_n 0.0100406f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_111_n N_A_241_368#_c_432_n 0.00473389f $X=1.575 $Y=1.725 $X2=0
+ $Y2=0
cc_140 N_TE_B_c_100_n N_A_241_368#_c_428_n 0.00269544f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_141 N_TE_B_c_101_n N_A_241_368#_c_428_n 0.00779369f $X=1.935 $Y=1.65 $X2=0
+ $Y2=0
cc_142 N_TE_B_c_104_n N_A_241_368#_c_428_n 0.00922102f $X=1.575 $Y=1.65 $X2=0
+ $Y2=0
cc_143 N_TE_B_c_105_n N_A_241_368#_c_428_n 0.0083671f $X=2.025 $Y=1.65 $X2=0
+ $Y2=0
cc_144 N_TE_B_c_100_n N_A_241_368#_c_429_n 0.00428963f $X=1.485 $Y=1.65 $X2=0
+ $Y2=0
cc_145 N_TE_B_c_108_n N_A_241_368#_c_429_n 4.01997e-19 $X=0.655 $Y=1.512 $X2=0
+ $Y2=0
cc_146 N_TE_B_c_111_n N_A_241_368#_c_433_n 6.90987e-19 $X=1.575 $Y=1.725 $X2=0
+ $Y2=0
cc_147 N_TE_B_c_113_n N_A_241_368#_c_433_n 0.017575f $X=2.025 $Y=1.725 $X2=0
+ $Y2=0
cc_148 N_TE_B_c_102_n N_A_241_368#_c_433_n 0.00710954f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_149 N_TE_B_c_115_n N_A_241_368#_c_433_n 0.00297728f $X=2.475 $Y=1.725 $X2=0
+ $Y2=0
cc_150 N_TE_B_c_105_n N_A_241_368#_c_433_n 0.00227061f $X=2.025 $Y=1.65 $X2=0
+ $Y2=0
cc_151 N_TE_B_c_102_n N_A_241_368#_c_430_n 0.00269544f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_152 N_TE_B_c_103_n N_A_241_368#_c_430_n 0.0172115f $X=2.885 $Y=1.65 $X2=0
+ $Y2=0
cc_153 N_TE_B_c_106_n N_A_241_368#_c_430_n 0.00922102f $X=2.475 $Y=1.65 $X2=0
+ $Y2=0
cc_154 N_TE_B_c_115_n N_A_241_368#_c_434_n 7.32019e-19 $X=2.475 $Y=1.725 $X2=0
+ $Y2=0
cc_155 N_TE_B_c_103_n N_A_241_368#_c_434_n 0.00426948f $X=2.885 $Y=1.65 $X2=0
+ $Y2=0
cc_156 N_TE_B_c_117_n N_A_241_368#_c_434_n 0.0154642f $X=2.975 $Y=1.725 $X2=0
+ $Y2=0
cc_157 N_TE_B_c_117_n N_A_241_368#_c_436_n 0.00337043f $X=2.975 $Y=1.725 $X2=0
+ $Y2=0
cc_158 N_TE_B_c_102_n N_A_241_368#_c_431_n 0.00261868f $X=2.385 $Y=1.65 $X2=0
+ $Y2=0
cc_159 N_TE_B_c_105_n N_A_241_368#_c_431_n 3.61456e-19 $X=2.025 $Y=1.65 $X2=0
+ $Y2=0
cc_160 N_TE_B_c_117_n N_Z_c_518_n 2.49165e-19 $X=2.975 $Y=1.725 $X2=0 $Y2=0
cc_161 N_TE_B_c_103_n Z 2.49165e-19 $X=2.885 $Y=1.65 $X2=0 $Y2=0
cc_162 N_TE_B_M1015_g N_VGND_c_566_n 0.00555851f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_163 N_TE_B_c_107_n N_VGND_c_566_n 0.0206988f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_164 N_TE_B_c_108_n N_VGND_c_566_n 0.00187637f $X=0.655 $Y=1.512 $X2=0 $Y2=0
cc_165 N_TE_B_M1015_g N_VGND_c_569_n 0.00431986f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_166 N_TE_B_M1015_g N_VGND_c_574_n 0.00824594f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_167 N_TE_B_c_104_n N_A_281_74#_c_627_n 7.00196e-19 $X=1.575 $Y=1.65 $X2=0
+ $Y2=0
cc_168 N_TE_B_c_106_n N_A_281_74#_c_630_n 5.79814e-19 $X=2.475 $Y=1.65 $X2=0
+ $Y2=0
cc_169 N_A_114_74#_c_202_n N_A_c_283_n 0.00903267f $X=3.055 $Y=1.185 $X2=0 $Y2=0
cc_170 N_A_114_74#_c_201_n N_A_c_288_n 0.00903267f $X=2.98 $Y=1.26 $X2=0 $Y2=0
cc_171 N_A_114_74#_c_207_n N_VPWR_c_369_n 0.0346097f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_114_74#_c_207_n N_VPWR_c_372_n 0.014549f $X=0.79 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_114_74#_c_207_n N_VPWR_c_367_n 0.0119743f $X=0.79 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_114_74#_c_207_n N_A_241_368#_c_432_n 0.0871686f $X=0.79 $Y=1.985
+ $X2=0 $Y2=0
cc_175 N_A_114_74#_c_194_n N_A_241_368#_c_428_n 0.00442459f $X=1.69 $Y=1.26
+ $X2=0 $Y2=0
cc_176 N_A_114_74#_c_195_n N_A_241_368#_c_429_n 0.0048544f $X=1.295 $Y=1.26
+ $X2=0 $Y2=0
cc_177 N_A_114_74#_c_206_n N_A_241_368#_c_429_n 0.00980665f $X=0.79 $Y=1.31
+ $X2=0 $Y2=0
cc_178 N_A_114_74#_c_207_n N_A_241_368#_c_429_n 0.0114923f $X=0.79 $Y=1.985
+ $X2=0 $Y2=0
cc_179 N_A_114_74#_c_199_n N_A_241_368#_c_430_n 0.00438974f $X=2.55 $Y=1.26
+ $X2=0 $Y2=0
cc_180 N_A_114_74#_c_201_n N_A_241_368#_c_430_n 0.00205135f $X=2.98 $Y=1.26
+ $X2=0 $Y2=0
cc_181 N_A_114_74#_c_197_n N_A_241_368#_c_431_n 0.00188621f $X=2.12 $Y=1.26
+ $X2=0 $Y2=0
cc_182 N_A_114_74#_c_206_n N_VGND_c_566_n 0.0367724f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_183 N_A_114_74#_c_196_n N_VGND_c_567_n 0.0122703f $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_184 N_A_114_74#_c_197_n N_VGND_c_567_n 7.11061e-19 $X=2.12 $Y=1.26 $X2=0
+ $Y2=0
cc_185 N_A_114_74#_c_198_n N_VGND_c_567_n 0.0106722f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_186 N_A_114_74#_c_200_n N_VGND_c_567_n 5.10431e-19 $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_187 N_A_114_74#_c_206_n N_VGND_c_567_n 0.00159476f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_188 N_A_114_74#_c_198_n N_VGND_c_568_n 5.10431e-19 $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_189 N_A_114_74#_c_200_n N_VGND_c_568_n 0.0106722f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_190 N_A_114_74#_c_201_n N_VGND_c_568_n 7.11061e-19 $X=2.98 $Y=1.26 $X2=0
+ $Y2=0
cc_191 N_A_114_74#_c_202_n N_VGND_c_568_n 0.010039f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_192 N_A_114_74#_c_196_n N_VGND_c_569_n 0.00383152f $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_193 N_A_114_74#_c_206_n N_VGND_c_569_n 0.0406574f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_194 N_A_114_74#_c_208_n N_VGND_c_569_n 0.00199209f $X=1.13 $Y=0.465 $X2=0
+ $Y2=0
cc_195 N_A_114_74#_c_198_n N_VGND_c_571_n 0.00383152f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_196 N_A_114_74#_c_200_n N_VGND_c_571_n 0.00383152f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_197 N_A_114_74#_c_202_n N_VGND_c_573_n 0.00383152f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_A_114_74#_c_196_n N_VGND_c_574_n 0.00762539f $X=1.765 $Y=1.185 $X2=0
+ $Y2=0
cc_199 N_A_114_74#_c_198_n N_VGND_c_574_n 0.0075754f $X=2.195 $Y=1.185 $X2=0
+ $Y2=0
cc_200 N_A_114_74#_c_200_n N_VGND_c_574_n 0.0075754f $X=2.625 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_A_114_74#_c_202_n N_VGND_c_574_n 0.00757637f $X=3.055 $Y=1.185 $X2=0
+ $Y2=0
cc_202 N_A_114_74#_c_206_n N_VGND_c_574_n 0.0281533f $X=0.79 $Y=1.31 $X2=0 $Y2=0
cc_203 N_A_114_74#_c_196_n N_A_281_74#_c_626_n 0.00122824f $X=1.765 $Y=1.185
+ $X2=0 $Y2=0
cc_204 N_A_114_74#_c_206_n N_A_281_74#_c_626_n 0.0621205f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_205 N_A_114_74#_c_208_n N_A_281_74#_c_626_n 0.00274841f $X=1.13 $Y=0.465
+ $X2=0 $Y2=0
cc_206 N_A_114_74#_c_194_n N_A_281_74#_c_627_n 8.87202e-19 $X=1.69 $Y=1.26 $X2=0
+ $Y2=0
cc_207 N_A_114_74#_c_196_n N_A_281_74#_c_627_n 0.0075146f $X=1.765 $Y=1.185
+ $X2=0 $Y2=0
cc_208 N_A_114_74#_c_197_n N_A_281_74#_c_627_n 0.00614039f $X=2.12 $Y=1.26 $X2=0
+ $Y2=0
cc_209 N_A_114_74#_c_198_n N_A_281_74#_c_627_n 0.00752307f $X=2.195 $Y=1.185
+ $X2=0 $Y2=0
cc_210 N_A_114_74#_c_199_n N_A_281_74#_c_627_n 8.86022e-19 $X=2.55 $Y=1.26 $X2=0
+ $Y2=0
cc_211 N_A_114_74#_c_203_n N_A_281_74#_c_627_n 0.00251095f $X=1.765 $Y=1.26
+ $X2=0 $Y2=0
cc_212 N_A_114_74#_c_204_n N_A_281_74#_c_627_n 0.00250761f $X=2.195 $Y=1.26
+ $X2=0 $Y2=0
cc_213 N_A_114_74#_c_194_n N_A_281_74#_c_628_n 0.00791143f $X=1.69 $Y=1.26 $X2=0
+ $Y2=0
cc_214 N_A_114_74#_c_206_n N_A_281_74#_c_628_n 0.0145349f $X=0.79 $Y=1.31 $X2=0
+ $Y2=0
cc_215 N_A_114_74#_c_198_n N_A_281_74#_c_629_n 0.00106896f $X=2.195 $Y=1.185
+ $X2=0 $Y2=0
cc_216 N_A_114_74#_c_200_n N_A_281_74#_c_629_n 0.00106896f $X=2.625 $Y=1.185
+ $X2=0 $Y2=0
cc_217 N_A_114_74#_c_199_n N_A_281_74#_c_630_n 8.87202e-19 $X=2.55 $Y=1.26 $X2=0
+ $Y2=0
cc_218 N_A_114_74#_c_200_n N_A_281_74#_c_630_n 0.00753499f $X=2.625 $Y=1.185
+ $X2=0 $Y2=0
cc_219 N_A_114_74#_c_201_n N_A_281_74#_c_630_n 0.0101675f $X=2.98 $Y=1.26 $X2=0
+ $Y2=0
cc_220 N_A_114_74#_c_202_n N_A_281_74#_c_630_n 0.00752307f $X=3.055 $Y=1.185
+ $X2=0 $Y2=0
cc_221 N_A_114_74#_c_205_n N_A_281_74#_c_630_n 0.00251095f $X=2.625 $Y=1.26
+ $X2=0 $Y2=0
cc_222 N_A_114_74#_c_202_n N_A_281_74#_c_631_n 9.48753e-19 $X=3.055 $Y=1.185
+ $X2=0 $Y2=0
cc_223 N_A_114_74#_c_202_n N_A_281_74#_c_632_n 9.80302e-19 $X=3.055 $Y=1.185
+ $X2=0 $Y2=0
cc_224 N_A_114_74#_c_199_n N_A_281_74#_c_660_n 0.00526155f $X=2.55 $Y=1.26 $X2=0
+ $Y2=0
cc_225 N_A_c_289_n N_VPWR_c_374_n 0.00333926f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_226 N_A_c_290_n N_VPWR_c_374_n 0.00333926f $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_227 N_A_c_291_n N_VPWR_c_374_n 0.00333926f $X=4.325 $Y=1.725 $X2=0 $Y2=0
cc_228 N_A_c_292_n N_VPWR_c_374_n 0.00333926f $X=4.775 $Y=1.725 $X2=0 $Y2=0
cc_229 N_A_c_289_n N_VPWR_c_367_n 0.00422798f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_230 N_A_c_290_n N_VPWR_c_367_n 0.00422687f $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_231 N_A_c_291_n N_VPWR_c_367_n 0.00422687f $X=4.325 $Y=1.725 $X2=0 $Y2=0
cc_232 N_A_c_292_n N_VPWR_c_367_n 0.00426429f $X=4.775 $Y=1.725 $X2=0 $Y2=0
cc_233 N_A_c_288_n N_A_241_368#_c_430_n 0.00371655f $X=4.785 $Y=1.472 $X2=0
+ $Y2=0
cc_234 N_A_c_288_n N_A_241_368#_c_434_n 0.0018147f $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_235 N_A_c_289_n N_A_241_368#_c_435_n 0.0139961f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_236 N_A_c_290_n N_A_241_368#_c_435_n 0.0139729f $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_237 N_A_c_288_n N_A_241_368#_c_475_n 4.79064e-19 $X=4.785 $Y=1.472 $X2=0
+ $Y2=0
cc_238 N_A_c_291_n N_A_241_368#_c_437_n 0.0140221f $X=4.325 $Y=1.725 $X2=0 $Y2=0
cc_239 N_A_c_292_n N_A_241_368#_c_437_n 0.0149445f $X=4.775 $Y=1.725 $X2=0 $Y2=0
cc_240 N_A_c_292_n N_A_241_368#_c_438_n 0.00147281f $X=4.775 $Y=1.725 $X2=0
+ $Y2=0
cc_241 A N_A_241_368#_c_438_n 0.0148634f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_242 N_A_c_288_n N_A_241_368#_c_438_n 0.00381921f $X=4.785 $Y=1.472 $X2=0
+ $Y2=0
cc_243 N_A_c_289_n N_Z_c_518_n 0.0104219f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_244 N_A_c_290_n N_Z_c_518_n 0.0116523f $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_245 N_A_c_290_n N_Z_c_522_n 0.0117685f $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_246 N_A_c_291_n N_Z_c_522_n 0.0125297f $X=4.325 $Y=1.725 $X2=0 $Y2=0
cc_247 N_A_c_292_n N_Z_c_522_n 0.00669924f $X=4.775 $Y=1.725 $X2=0 $Y2=0
cc_248 A N_Z_c_522_n 0.0517544f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_249 N_A_c_288_n N_Z_c_522_n 0.0228583f $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_250 N_A_c_284_n N_Z_c_527_n 0.013849f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_251 N_A_c_285_n N_Z_c_527_n 0.0112736f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_252 A N_Z_c_527_n 0.030527f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_253 N_A_c_288_n N_Z_c_527_n 7.06413e-19 $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_254 N_A_c_290_n N_Z_c_531_n 6.45773e-19 $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_255 N_A_c_291_n N_Z_c_531_n 0.0116523f $X=4.325 $Y=1.725 $X2=0 $Y2=0
cc_256 N_A_c_292_n N_Z_c_531_n 0.0109688f $X=4.775 $Y=1.725 $X2=0 $Y2=0
cc_257 N_A_c_283_n N_Z_c_516_n 7.88797e-19 $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A_c_284_n N_Z_c_516_n 0.0045177f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_259 N_A_c_285_n N_Z_c_516_n 6.97036e-19 $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_260 A N_Z_c_537_n 0.0140706f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_261 N_A_c_288_n N_Z_c_537_n 6.72853e-19 $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_262 N_A_c_289_n Z 0.00326583f $X=3.425 $Y=1.725 $X2=0 $Y2=0
cc_263 N_A_c_290_n Z 0.00224404f $X=3.875 $Y=1.725 $X2=0 $Y2=0
cc_264 N_A_c_291_n Z 7.19288e-19 $X=4.325 $Y=1.725 $X2=0 $Y2=0
cc_265 N_A_c_288_n Z 0.0241006f $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_266 N_A_c_284_n N_Z_c_517_n 0.00160429f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_267 A N_Z_c_517_n 0.023376f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_268 N_A_c_288_n N_Z_c_517_n 0.0219011f $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_269 N_A_c_283_n N_VGND_c_568_n 3.79623e-19 $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_270 N_A_c_283_n N_VGND_c_573_n 0.00278247f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_271 N_A_c_284_n N_VGND_c_573_n 0.00278271f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_272 N_A_c_285_n N_VGND_c_573_n 0.00278271f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_273 N_A_c_286_n N_VGND_c_573_n 0.00278247f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_274 N_A_c_283_n N_VGND_c_574_n 0.00353524f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_275 N_A_c_284_n N_VGND_c_574_n 0.00352619f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_276 N_A_c_285_n N_VGND_c_574_n 0.00353528f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A_c_286_n N_VGND_c_574_n 0.00357084f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A_c_283_n N_A_281_74#_c_630_n 0.00174914f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_279 N_A_c_288_n N_A_281_74#_c_630_n 0.00720745f $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_280 N_A_c_283_n N_A_281_74#_c_631_n 0.00194824f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_281 N_A_c_283_n N_A_281_74#_c_632_n 0.00761102f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_282 N_A_c_284_n N_A_281_74#_c_632_n 9.14331e-19 $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_283 N_A_c_283_n N_A_281_74#_c_633_n 0.0146721f $X=3.485 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A_c_284_n N_A_281_74#_c_633_n 0.0130518f $X=3.915 $Y=1.22 $X2=0 $Y2=0
cc_285 N_A_c_288_n N_A_281_74#_c_633_n 2.98044e-19 $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_286 N_A_c_285_n N_A_281_74#_c_634_n 0.00708406f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_287 N_A_c_286_n N_A_281_74#_c_634_n 0.0140292f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_288 N_A_c_285_n N_A_281_74#_c_635_n 5.5198e-19 $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_289 N_A_c_286_n N_A_281_74#_c_635_n 0.0114766f $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_290 A N_A_281_74#_c_635_n 0.0251801f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_291 N_A_c_288_n N_A_281_74#_c_635_n 0.00114736f $X=4.785 $Y=1.472 $X2=0 $Y2=0
cc_292 N_A_c_285_n N_A_281_74#_c_636_n 0.00529157f $X=4.355 $Y=1.22 $X2=0 $Y2=0
cc_293 N_A_c_286_n N_A_281_74#_c_636_n 5.01714e-19 $X=4.785 $Y=1.22 $X2=0 $Y2=0
cc_294 N_VPWR_c_370_n N_A_241_368#_c_432_n 0.0379768f $X=1.8 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_372_n N_A_241_368#_c_432_n 0.011066f $X=1.635 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_367_n N_A_241_368#_c_432_n 0.00915947f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_370_n N_A_241_368#_c_428_n 0.0198465f $X=1.8 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_370_n N_A_241_368#_c_433_n 0.0379768f $X=1.8 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_371_n N_A_241_368#_c_433_n 0.0395686f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_373_n N_A_241_368#_c_433_n 0.0109793f $X=2.535 $Y=3.33 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_367_n N_A_241_368#_c_433_n 0.00901959f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_371_n N_A_241_368#_c_430_n 0.0263013f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_371_n N_A_241_368#_c_434_n 0.0397705f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_374_n N_A_241_368#_c_435_n 0.0458929f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_367_n N_A_241_368#_c_435_n 0.0257967f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_371_n N_A_241_368#_c_436_n 0.0119238f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_374_n N_A_241_368#_c_436_n 0.0177474f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_367_n N_A_241_368#_c_436_n 0.00957218f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_374_n N_A_241_368#_c_437_n 0.0638408f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_367_n N_A_241_368#_c_437_n 0.0355196f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_374_n N_A_241_368#_c_439_n 0.0121867f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_367_n N_A_241_368#_c_439_n 0.00660921f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_A_241_368#_c_435_n N_Z_M1008_d 0.00165831f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_314 N_A_241_368#_c_437_n N_Z_M1010_d 0.00165831f $X=4.915 $Y=2.99 $X2=0 $Y2=0
cc_315 N_A_241_368#_c_435_n N_Z_c_518_n 0.0159318f $X=4.015 $Y=2.99 $X2=0 $Y2=0
cc_316 N_A_241_368#_M1009_s N_Z_c_522_n 0.00165831f $X=3.965 $Y=1.84 $X2=0 $Y2=0
cc_317 N_A_241_368#_c_475_n N_Z_c_522_n 0.0126919f $X=4.1 $Y=2.225 $X2=0 $Y2=0
cc_318 N_A_241_368#_c_438_n N_Z_c_522_n 0.00326551f $X=5 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A_241_368#_c_437_n N_Z_c_531_n 0.0159318f $X=4.915 $Y=2.99 $X2=0 $Y2=0
cc_320 N_A_241_368#_c_430_n Z 0.00746325f $X=3.035 $Y=1.565 $X2=0 $Y2=0
cc_321 N_A_241_368#_c_434_n Z 0.0423689f $X=3.2 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_241_368#_c_430_n N_Z_c_517_n 0.00346621f $X=3.035 $Y=1.565 $X2=0
+ $Y2=0
cc_323 N_A_241_368#_c_428_n N_A_281_74#_c_627_n 0.0320456f $X=2.085 $Y=1.565
+ $X2=0 $Y2=0
cc_324 N_A_241_368#_c_431_n N_A_281_74#_c_627_n 0.0192612f $X=2.21 $Y=1.565
+ $X2=0 $Y2=0
cc_325 N_A_241_368#_c_428_n N_A_281_74#_c_628_n 0.0135853f $X=2.085 $Y=1.565
+ $X2=0 $Y2=0
cc_326 N_A_241_368#_c_430_n N_A_281_74#_c_630_n 0.0600906f $X=3.035 $Y=1.565
+ $X2=0 $Y2=0
cc_327 N_A_241_368#_c_430_n N_A_281_74#_c_660_n 0.0127483f $X=3.035 $Y=1.565
+ $X2=0 $Y2=0
cc_328 N_A_241_368#_c_431_n N_A_281_74#_c_660_n 8.91514e-19 $X=2.21 $Y=1.565
+ $X2=0 $Y2=0
cc_329 N_Z_c_527_n N_A_281_74#_M1007_d 0.00351264f $X=4.485 $Y=0.89 $X2=0 $Y2=0
cc_330 N_Z_c_517_n N_A_281_74#_c_630_n 0.0127735f $X=3.65 $Y=1.55 $X2=0 $Y2=0
cc_331 N_Z_c_516_n N_A_281_74#_c_632_n 0.0137359f $X=3.74 $Y=0.89 $X2=0 $Y2=0
cc_332 N_Z_M1001_s N_A_281_74#_c_633_n 0.00171549f $X=3.56 $Y=0.37 $X2=0 $Y2=0
cc_333 N_Z_c_527_n N_A_281_74#_c_633_n 0.023966f $X=4.485 $Y=0.89 $X2=0 $Y2=0
cc_334 N_Z_c_516_n N_A_281_74#_c_633_n 0.0154405f $X=3.74 $Y=0.89 $X2=0 $Y2=0
cc_335 N_Z_M1012_s N_A_281_74#_c_634_n 0.00176461f $X=4.43 $Y=0.37 $X2=0 $Y2=0
cc_336 N_Z_c_527_n N_A_281_74#_c_634_n 0.00424866f $X=4.485 $Y=0.89 $X2=0 $Y2=0
cc_337 N_Z_c_537_n N_A_281_74#_c_634_n 0.0121701f $X=4.57 $Y=0.8 $X2=0 $Y2=0
cc_338 N_VGND_c_567_n N_A_281_74#_c_626_n 0.0229082f $X=1.98 $Y=0.515 $X2=0
+ $Y2=0
cc_339 N_VGND_c_569_n N_A_281_74#_c_626_n 0.00749631f $X=1.815 $Y=0 $X2=0 $Y2=0
cc_340 N_VGND_c_574_n N_A_281_74#_c_626_n 0.0062048f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_567_n N_A_281_74#_c_627_n 0.0216086f $X=1.98 $Y=0.515 $X2=0
+ $Y2=0
cc_342 N_VGND_c_567_n N_A_281_74#_c_629_n 0.0229082f $X=1.98 $Y=0.515 $X2=0
+ $Y2=0
cc_343 N_VGND_c_568_n N_A_281_74#_c_629_n 0.0229082f $X=2.84 $Y=0.515 $X2=0
+ $Y2=0
cc_344 N_VGND_c_571_n N_A_281_74#_c_629_n 0.00749631f $X=2.675 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_c_574_n N_A_281_74#_c_629_n 0.0062048f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_568_n N_A_281_74#_c_630_n 0.0216086f $X=2.84 $Y=0.515 $X2=0
+ $Y2=0
cc_347 N_VGND_c_568_n N_A_281_74#_c_631_n 0.0175237f $X=2.84 $Y=0.515 $X2=0
+ $Y2=0
cc_348 N_VGND_c_573_n N_A_281_74#_c_631_n 0.0178338f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_574_n N_A_281_74#_c_631_n 0.00960503f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_573_n N_A_281_74#_c_633_n 0.0912556f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_574_n N_A_281_74#_c_633_n 0.0506361f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_573_n N_A_281_74#_c_634_n 0.0235688f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_574_n N_A_281_74#_c_634_n 0.0127152f $X=5.04 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__fah_4.pex.spice
* Created: Fri Aug 28 17:35:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FAH_4%A 3 7 11 15 17 23 24
c44 7 0 1.40087e-19 $X=0.495 $Y=0.69
c45 3 0 1.1782e-19 $X=0.505 $Y=2.46
r46 23 25 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=0.93 $Y=1.635
+ $X2=0.955 $Y2=1.635
r47 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.635 $X2=0.93 $Y2=1.635
r48 21 23 0.734756 $w=3.28e-07 $l=5e-09 $layer=POLY_cond $X=0.925 $Y=1.635
+ $X2=0.93 $Y2=1.635
r49 20 21 61.7195 $w=3.28e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.635
+ $X2=0.925 $Y2=1.635
r50 19 20 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.635
+ $X2=0.505 $Y2=1.635
r51 17 24 8.34528 $w=2.88e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=1.655
+ $X2=0.93 $Y2=1.655
r52 13 25 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.8
+ $X2=0.955 $Y2=1.635
r53 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.8
+ $X2=0.955 $Y2=2.46
r54 9 21 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.47
+ $X2=0.925 $Y2=1.635
r55 9 11 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.925 $Y=1.47
+ $X2=0.925 $Y2=0.69
r56 5 19 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=1.635
r57 5 7 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=0.69
r58 1 20 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.8
+ $X2=0.505 $Y2=1.635
r59 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.8 $X2=0.505
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_27_74# 1 2 7 11 13 15 16 19 23 25 29 31 32
+ 33 39
c71 39 0 5.85186e-20 $X=1.5 $Y=1.395
r72 37 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.5 $Y=1.485 $X2=1.5
+ $Y2=1.395
r73 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.5
+ $Y=1.485 $X2=1.5 $Y2=1.485
r74 33 36 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.5 $Y=1.255 $X2=1.5
+ $Y2=1.485
r75 30 31 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.255
+ $X2=0.225 $Y2=1.255
r76 29 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=1.255
+ $X2=1.5 $Y2=1.255
r77 29 30 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.335 $Y=1.255
+ $X2=0.365 $Y2=1.255
r78 25 27 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.225 $Y=2.135
+ $X2=0.225 $Y2=2.815
r79 23 32 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=2.11
+ $X2=0.225 $Y2=1.97
r80 23 25 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.225 $Y=2.11
+ $X2=0.225 $Y2=2.135
r81 21 31 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.17 $Y=1.34
+ $X2=0.225 $Y2=1.255
r82 21 32 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.17 $Y=1.34
+ $X2=0.17 $Y2=1.97
r83 17 31 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=1.17
+ $X2=0.225 $Y2=1.255
r84 17 19 26.9589 $w=2.78e-07 $l=6.55e-07 $layer=LI1_cond $X=0.225 $Y=1.17
+ $X2=0.225 $Y2=0.515
r85 13 16 18.8402 $w=1.65e-07 $l=9.40744e-08 $layer=POLY_cond $X=2.13 $Y=1.32
+ $X2=2.087 $Y2=1.395
r86 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.13 $Y=1.32 $X2=2.13
+ $Y2=0.84
r87 9 16 18.8402 $w=1.65e-07 $l=8.74643e-08 $layer=POLY_cond $X=2.06 $Y=1.47
+ $X2=2.087 $Y2=1.395
r88 9 11 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=2.06 $Y=1.47 $X2=2.06
+ $Y2=2.37
r89 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.395
+ $X2=1.5 $Y2=1.395
r90 7 16 6.66866 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=1.97 $Y=1.395
+ $X2=2.087 $Y2=1.395
r91 7 8 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.97 $Y=1.395
+ $X2=1.665 $Y2=1.395
r92 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r93 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.135
r94 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_586_257# 1 2 3 10 12 17 18 19 23 26 30 33 36
+ 37 41 43 44 45 46 48 50 52 54
c167 52 0 1.99791e-19 $X=5.94 $Y=2.815
c168 50 0 1.35704e-20 $X=5.94 $Y=2.12
c169 37 0 1.58586e-19 $X=4.385 $Y=0.79
c170 26 0 1.73206e-19 $X=4.09 $Y=2.23
c171 23 0 4.11294e-20 $X=4.015 $Y=0.97
c172 12 0 1.11098e-19 $X=3.02 $Y=2.23
r173 50 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.035
r174 50 52 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.815
r175 46 48 171.257 $w=1.68e-07 $l=2.625e-06 $layer=LI1_cond $X=5.405 $Y=0.34
+ $X2=8.03 $Y2=0.34
r176 44 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=5.94 $Y2=2.035
r177 44 45 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.855 $Y=2.035
+ $X2=5.265 $Y2=2.035
r178 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.18 $Y=1.95
+ $X2=5.265 $Y2=2.035
r179 42 54 3.84343 $w=2.4e-07 $l=1.38651e-07 $layer=LI1_cond $X=5.18 $Y=0.92
+ $X2=5.25 $Y2=0.812
r180 42 43 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=5.18 $Y=0.92
+ $X2=5.18 $Y2=1.95
r181 39 54 3.84343 $w=2.4e-07 $l=1.07e-07 $layer=LI1_cond $X=5.25 $Y=0.705
+ $X2=5.25 $Y2=0.812
r182 39 41 7.80687 $w=3.08e-07 $l=2.1e-07 $layer=LI1_cond $X=5.25 $Y=0.705
+ $X2=5.25 $Y2=0.495
r183 38 46 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.25 $Y=0.425
+ $X2=5.405 $Y2=0.34
r184 38 41 2.60229 $w=3.08e-07 $l=7e-08 $layer=LI1_cond $X=5.25 $Y=0.425
+ $X2=5.25 $Y2=0.495
r185 36 54 2.60907 $w=1.7e-07 $l=1.65635e-07 $layer=LI1_cond $X=5.095 $Y=0.79
+ $X2=5.25 $Y2=0.812
r186 36 37 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.095 $Y=0.79
+ $X2=4.385 $Y2=0.79
r187 34 60 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.162 $Y=0.375
+ $X2=4.162 $Y2=0.54
r188 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.22
+ $Y=0.375 $X2=4.22 $Y2=0.375
r189 31 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.22 $Y=0.705
+ $X2=4.385 $Y2=0.79
r190 31 33 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.22 $Y=0.705
+ $X2=4.22 $Y2=0.375
r191 29 30 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.06 $Y=1.365
+ $X2=4.06 $Y2=1.515
r192 26 30 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=4.09 $Y=2.23
+ $X2=4.09 $Y2=1.515
r193 23 29 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.015 $Y=0.97
+ $X2=4.015 $Y2=1.365
r194 23 60 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.015 $Y=0.97
+ $X2=4.015 $Y2=0.54
r195 18 34 21.2463 $w=4.45e-07 $l=1.7e-07 $layer=POLY_cond $X=4.162 $Y=0.205
+ $X2=4.162 $Y2=0.375
r196 18 19 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.94 $Y=0.205
+ $X2=3.11 $Y2=0.205
r197 17 28 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=0.89
+ $X2=3.035 $Y2=1.285
r198 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.035 $Y=0.28
+ $X2=3.11 $Y2=0.205
r199 14 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.035 $Y=0.28
+ $X2=3.035 $Y2=0.89
r200 10 28 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.02 $Y=1.375
+ $X2=3.02 $Y2=1.285
r201 10 12 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=3.02 $Y=1.375
+ $X2=3.02 $Y2=2.23
r202 3 56 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.94 $Y2=2.115
r203 3 52 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.94 $Y2=2.815
r204 2 48 182 $w=1.7e-07 $l=4.92874e-07 $layer=licon1_NDIFF $count=1 $X=7.81
+ $Y=0.735 $X2=8.03 $Y2=0.34
r205 1 41 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.1
+ $Y=0.37 $X2=5.24 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%B 4 7 9 10 13 18 19 23 24 26 28 30 32 33 34 38
+ 39 43 44 45 54
c148 43 0 3.01964e-20 $X=4.8 $Y=2.065
c149 38 0 4.11294e-20 $X=4.8 $Y=1.385
c150 32 0 3.09806e-19 $X=3.6 $Y=1.735
c151 26 0 1.70742e-19 $X=5.715 $Y=1.765
r152 48 55 8.97022 $w=4.65e-07 $l=7.5e-08 $layer=POLY_cond $X=4.867 $Y=1.765
+ $X2=4.867 $Y2=1.69
r153 44 45 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.915 $Y=2.405
+ $X2=4.915 $Y2=2.775
r154 44 57 5.60012 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.915 $Y=2.405
+ $X2=4.915 $Y2=2.29
r155 44 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.8
+ $Y=2.405 $X2=4.8 $Y2=2.405
r156 43 51 40.665 $w=4.65e-07 $l=3.4e-07 $layer=POLY_cond $X=4.867 $Y=2.065
+ $X2=4.867 $Y2=2.405
r157 43 48 35.8809 $w=4.65e-07 $l=3e-07 $layer=POLY_cond $X=4.867 $Y=2.065
+ $X2=4.867 $Y2=1.765
r158 42 57 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=4.8 $Y=2.065
+ $X2=4.8 $Y2=2.29
r159 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=2.065 $X2=4.8 $Y2=2.065
r160 39 55 36.4789 $w=4.65e-07 $l=3.05e-07 $layer=POLY_cond $X=4.867 $Y=1.385
+ $X2=4.867 $Y2=1.69
r161 39 54 47.3569 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.867 $Y=1.385
+ $X2=4.867 $Y2=1.22
r162 38 42 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.8 $Y=1.385
+ $X2=4.8 $Y2=2.065
r163 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=1.385 $X2=4.8 $Y2=1.385
r164 34 51 32.6516 $w=4.65e-07 $l=2.73e-07 $layer=POLY_cond $X=4.867 $Y=2.678
+ $X2=4.867 $Y2=2.405
r165 31 32 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.6 $Y=1.585
+ $X2=3.6 $Y2=1.735
r166 29 30 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.577 $Y=1.45
+ $X2=2.577 $Y2=1.6
r167 26 28 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.715 $Y=1.765
+ $X2=5.715 $Y2=2.4
r168 25 55 29.5843 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.1 $Y=1.69
+ $X2=4.867 $Y2=1.69
r169 24 26 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.625 $Y=1.69
+ $X2=5.715 $Y2=1.765
r170 24 25 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.625 $Y=1.69
+ $X2=5.1 $Y2=1.69
r171 23 54 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.025 $Y=0.74
+ $X2=5.025 $Y2=1.22
r172 20 33 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.73 $Y=3.095
+ $X2=3.64 $Y2=3.095
r173 19 34 49.4222 $w=4.65e-07 $l=5.20224e-07 $layer=POLY_cond $X=4.635 $Y=3.095
+ $X2=4.867 $Y2=2.678
r174 19 20 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=4.635 $Y=3.095
+ $X2=3.73 $Y2=3.095
r175 18 32 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.64 $Y=2.23
+ $X2=3.64 $Y2=1.735
r176 16 33 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.64 $Y=3.02
+ $X2=3.64 $Y2=3.095
r177 16 18 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=3.64 $Y=3.02
+ $X2=3.64 $Y2=2.23
r178 13 31 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.545 $Y=0.97
+ $X2=3.545 $Y2=1.585
r179 9 33 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.55 $Y=3.095 $X2=3.64
+ $Y2=3.095
r180 9 10 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=3.55 $Y=3.095
+ $X2=2.655 $Y2=3.095
r181 7 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.605 $Y=0.89
+ $X2=2.605 $Y2=1.45
r182 4 30 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.565 $Y=2.23
+ $X2=2.565 $Y2=1.6
r183 2 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.565 $Y=3.02
+ $X2=2.655 $Y2=3.095
r184 2 4 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.565 $Y=3.02
+ $X2=2.565 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_531_362# 1 2 7 12 13 15 16 17 18 20 25 26 31
+ 35 37 42 43 45 46 47 48 51 55 57 58
c205 58 0 3.01964e-20 $X=5.52 $Y=1.665
c206 55 0 1.58586e-19 $X=4.08 $Y=1.665
c207 37 0 3.83589e-19 $X=3.885 $Y=1.657
c208 26 0 9.38637e-20 $X=6.275 $Y=1.3
c209 13 0 3.0708e-19 $X=6.315 $Y=1.225
r210 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r211 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r212 51 68 14.4306 $w=2.28e-07 $l=2.88e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=2.832 $Y2=1.665
r213 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r214 48 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r215 47 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=5.52 $Y2=1.665
r216 47 48 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=4.225 $Y2=1.665
r217 46 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r218 45 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r219 45 46 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=3.265 $Y2=1.665
r220 43 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.64 $Y=1.21 $X2=5.64
+ $Y2=1.3
r221 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.21 $X2=5.64 $Y2=1.21
r222 39 58 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=5.535 $Y=1.375
+ $X2=5.535 $Y2=1.665
r223 38 42 4.24584 $w=2.83e-07 $l=1.05e-07 $layer=LI1_cond $X=5.535 $Y=1.232
+ $X2=5.64 $Y2=1.232
r224 38 39 2.81168 $w=2e-07 $l=1.43e-07 $layer=LI1_cond $X=5.535 $Y=1.232
+ $X2=5.535 $Y2=1.375
r225 37 55 10.4524 $w=2.13e-07 $l=1.95e-07 $layer=LI1_cond $X=3.885 $Y=1.657
+ $X2=4.08 $Y2=1.657
r226 33 37 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.8 $Y=1.55
+ $X2=3.885 $Y2=1.657
r227 33 35 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.8 $Y=1.55
+ $X2=3.8 $Y2=0.795
r228 29 68 0.103554 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=2.832 $Y=1.78
+ $X2=2.832 $Y2=1.665
r229 29 31 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=2.832 $Y=1.78
+ $X2=2.832 $Y2=1.955
r230 23 25 209.903 $w=1.8e-07 $l=5.4e-07 $layer=POLY_cond $X=7.485 $Y=3.075
+ $X2=7.485 $Y2=2.535
r231 22 25 211.847 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=7.485 $Y=1.99
+ $X2=7.485 $Y2=2.535
r232 18 22 54.566 $w=2.12e-07 $l=4.2332e-07 $layer=POLY_cond $X=7.245 $Y=1.67
+ $X2=7.485 $Y2=1.99
r233 18 20 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=7.245 $Y=1.67
+ $X2=7.245 $Y2=0.945
r234 16 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.395 $Y=3.15
+ $X2=7.485 $Y2=3.075
r235 16 17 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=7.395 $Y=3.15
+ $X2=6.34 $Y2=3.15
r236 13 26 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=6.315 $Y=1.225
+ $X2=6.275 $Y2=1.3
r237 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.315 $Y=1.225
+ $X2=6.315 $Y2=0.83
r238 10 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.25 $Y=3.075
+ $X2=6.34 $Y2=3.15
r239 10 12 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=6.25 $Y=3.075
+ $X2=6.25 $Y2=2.315
r240 9 26 18.8402 $w=1.65e-07 $l=8.66025e-08 $layer=POLY_cond $X=6.25 $Y=1.375
+ $X2=6.275 $Y2=1.3
r241 9 12 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=6.25 $Y=1.375
+ $X2=6.25 $Y2=2.315
r242 8 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=1.3
+ $X2=5.64 $Y2=1.3
r243 7 26 6.66866 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=6.16 $Y=1.3
+ $X2=6.275 $Y2=1.3
r244 7 8 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.16 $Y=1.3
+ $X2=5.805 $Y2=1.3
r245 2 31 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=1.81 $X2=2.79 $Y2=1.955
r246 1 35 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=3.62
+ $Y=0.65 $X2=3.8 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_536_114# 1 2 10 13 15 16 20 22 23 24 25 27
+ 30 34 36 37 39 40 41 42 48 52 53 58
c196 58 0 1.03543e-19 $X=3.865 $Y=2.025
c197 53 0 4.2619e-20 $X=6.795 $Y=1.57
c198 52 0 8.74051e-20 $X=6.795 $Y=1.57
c199 42 0 3.55926e-19 $X=3.745 $Y=2.035
c200 41 0 1.8874e-19 $X=6.815 $Y=2.035
c201 39 0 1.73206e-19 $X=3.46 $Y=1.935
c202 30 0 1.35123e-19 $X=7.89 $Y=1.525
c203 23 0 5.38428e-20 $X=8.345 $Y=1.965
r204 52 55 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.57
+ $X2=6.795 $Y2=1.735
r205 52 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.57
+ $X2=6.795 $Y2=1.405
r206 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.795
+ $Y=1.57 $X2=6.795 $Y2=1.57
r207 49 53 12.7592 $w=4.18e-07 $l=4.65e-07 $layer=LI1_cond $X=6.865 $Y=2.035
+ $X2=6.865 $Y2=1.57
r208 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r209 45 58 15.887 $w=1.83e-07 $l=2.65e-07 $layer=LI1_cond $X=3.6 $Y=2.027
+ $X2=3.865 $Y2=2.027
r210 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r211 42 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r212 41 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=6.96 $Y2=2.035
r213 41 42 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=3.745 $Y2=2.035
r214 40 45 3.2973 $w=1.83e-07 $l=5.5e-08 $layer=LI1_cond $X=3.545 $Y=2.027
+ $X2=3.6 $Y2=2.027
r215 39 40 6.83233 $w=1.85e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.46 $Y=1.935
+ $X2=3.545 $Y2=2.027
r216 38 39 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.46 $Y=1.38
+ $X2=3.46 $Y2=1.935
r217 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.375 $Y=1.295
+ $X2=3.46 $Y2=1.38
r218 36 37 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.375 $Y=1.295
+ $X2=2.985 $Y2=1.295
r219 32 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.82 $Y=1.21
+ $X2=2.985 $Y2=1.295
r220 32 34 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.82 $Y=1.21
+ $X2=2.82 $Y2=0.745
r221 28 30 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.735 $Y=1.525
+ $X2=7.89 $Y2=1.525
r222 25 27 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.435 $Y=2.04
+ $X2=8.435 $Y2=2.535
r223 23 25 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.345 $Y=1.965
+ $X2=8.435 $Y2=2.04
r224 23 24 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=8.345 $Y=1.965
+ $X2=7.965 $Y2=1.965
r225 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.89 $Y=1.89
+ $X2=7.965 $Y2=1.965
r226 21 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.89 $Y=1.6
+ $X2=7.89 $Y2=1.525
r227 21 22 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.89 $Y=1.6
+ $X2=7.89 $Y2=1.89
r228 18 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.735 $Y=1.45
+ $X2=7.735 $Y2=1.525
r229 18 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.735 $Y=1.45
+ $X2=7.735 $Y2=1.055
r230 17 20 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.735 $Y=0.255
+ $X2=7.735 $Y2=1.055
r231 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.66 $Y=0.18
+ $X2=7.735 $Y2=0.255
r232 15 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.66 $Y=0.18
+ $X2=6.89 $Y2=0.18
r233 13 55 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.845 $Y=2.315
+ $X2=6.845 $Y2=1.735
r234 10 54 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.815 $Y=0.945
+ $X2=6.815 $Y2=1.405
r235 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.815 $Y=0.255
+ $X2=6.89 $Y2=0.18
r236 7 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.815 $Y=0.255
+ $X2=6.815 $Y2=0.945
r237 2 58 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.81 $X2=3.865 $Y2=2.025
r238 1 34 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.68
+ $Y=0.57 $X2=2.82 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_1378_125# 1 2 3 4 15 17 19 21 22 23 25 27 29
+ 31 32 33 37 39 40 42 44 47 52 53 55 59 62 63 65 66 67 68 73 74
c221 62 0 1.37274e-19 $X=7.03 $Y=1.11
c222 59 0 9.38637e-20 $X=6.4 $Y=2.065
c223 42 0 1.35123e-19 $X=8.37 $Y=1.485
c224 39 0 1.70833e-19 $X=7.875 $Y=1.565
c225 27 0 1.69806e-19 $X=6.4 $Y=1.98
c226 22 0 5.40791e-20 $X=8.88 $Y=1.485
r227 73 74 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=12.505 $Y=2.035
+ $X2=12.505 $Y2=1.95
r228 68 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.63 $Y=2.695
+ $X2=8.63 $Y2=2.99
r229 62 63 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.03 $Y=1.115
+ $X2=6.865 $Y2=1.115
r230 57 59 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.28 $Y=2.065
+ $X2=6.4 $Y2=2.065
r231 53 55 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=12.465 $Y=1.095
+ $X2=12.69 $Y2=1.095
r232 52 76 2.84834 $w=4.2e-07 $l=1.25e-07 $layer=LI1_cond $X=12.505 $Y=2.61
+ $X2=12.505 $Y2=2.735
r233 51 73 3.42989 $w=4.18e-07 $l=1.25e-07 $layer=LI1_cond $X=12.505 $Y=2.16
+ $X2=12.505 $Y2=2.035
r234 51 52 12.3476 $w=4.18e-07 $l=4.5e-07 $layer=LI1_cond $X=12.505 $Y=2.16
+ $X2=12.505 $Y2=2.61
r235 49 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.38 $Y=1.18
+ $X2=12.465 $Y2=1.095
r236 49 74 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=12.38 $Y=1.18
+ $X2=12.38 $Y2=1.95
r237 48 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=2.695
+ $X2=8.63 $Y2=2.695
r238 47 76 5.69669 $w=1.7e-07 $l=2.29129e-07 $layer=LI1_cond $X=12.295 $Y=2.695
+ $X2=12.505 $Y2=2.735
r239 47 48 233.561 $w=1.68e-07 $l=3.58e-06 $layer=LI1_cond $X=12.295 $Y=2.695
+ $X2=8.715 $Y2=2.695
r240 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.71
+ $Y=1.485 $X2=8.71 $Y2=1.485
r241 42 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.37 $Y=1.485
+ $X2=8.205 $Y2=1.485
r242 42 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.37 $Y=1.485
+ $X2=8.71 $Y2=1.485
r243 41 66 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.875 $Y=2.99
+ $X2=7.79 $Y2=2.9
r244 40 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=8.63 $Y2=2.99
r245 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=7.875 $Y2=2.99
r246 39 67 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.875 $Y=1.565
+ $X2=8.205 $Y2=1.565
r247 37 66 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.79 $Y=2.725
+ $X2=7.79 $Y2=2.9
r248 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.79 $Y=1.65
+ $X2=7.875 $Y2=1.565
r249 36 37 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=7.79 $Y=1.65
+ $X2=7.79 $Y2=2.725
r250 33 65 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=7.165 $Y=2.9
+ $X2=6.99 $Y2=2.9
r251 33 35 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=7.165 $Y=2.9
+ $X2=7.205 $Y2=2.9
r252 32 66 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.705 $Y=2.9
+ $X2=7.79 $Y2=2.9
r253 32 35 16.4635 $w=3.48e-07 $l=5e-07 $layer=LI1_cond $X=7.705 $Y=2.9
+ $X2=7.205 $Y2=2.9
r254 31 63 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.485 $Y=1.13
+ $X2=6.865 $Y2=1.13
r255 29 65 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.365 $Y=2.99
+ $X2=6.99 $Y2=2.99
r256 27 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=1.98 $X2=6.4
+ $Y2=2.065
r257 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.4 $Y=1.215
+ $X2=6.485 $Y2=1.13
r258 26 27 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.4 $Y=1.215
+ $X2=6.4 $Y2=1.98
r259 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.28 $Y=2.905
+ $X2=6.365 $Y2=2.99
r260 24 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=2.15
+ $X2=6.28 $Y2=2.065
r261 24 25 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.28 $Y=2.15
+ $X2=6.28 $Y2=2.905
r262 22 45 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=8.88 $Y=1.485
+ $X2=8.71 $Y2=1.485
r263 22 23 15.9654 $w=2.4e-07 $l=9e-08 $layer=POLY_cond $X=8.88 $Y=1.485
+ $X2=8.97 $Y2=1.485
r264 19 21 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=9.425 $Y=1.32
+ $X2=9.425 $Y2=0.92
r265 18 23 15.9654 $w=2.4e-07 $l=1.27279e-07 $layer=POLY_cond $X=9.06 $Y=1.395
+ $X2=8.97 $Y2=1.485
r266 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.35 $Y=1.395
+ $X2=9.425 $Y2=1.32
r267 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.35 $Y=1.395
+ $X2=9.06 $Y2=1.395
r268 13 23 9.46703 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.97 $Y=1.65
+ $X2=8.97 $Y2=1.485
r269 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=8.97 $Y=1.65
+ $X2=8.97 $Y2=2.34
r270 4 76 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=12.405
+ $Y=1.84 $X2=12.55 $Y2=2.715
r271 4 73 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=12.405
+ $Y=1.84 $X2=12.55 $Y2=2.035
r272 3 35 600 $w=1.7e-07 $l=1.04129e-06 $layer=licon1_PDIFF $count=1 $X=6.935
+ $Y=1.895 $X2=7.205 $Y2=2.81
r273 2 55 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=12.545
+ $Y=0.6 $X2=12.69 $Y2=1.095
r274 1 62 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=6.89
+ $Y=0.625 $X2=7.03 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_1268_379# 1 2 9 13 15 17 18 20 23 27 29 31
+ 32 34 35 38 39 42 43 44 46 47 48 50 53 56 61 77
c174 38 0 8.74051e-20 $X=7.45 $Y=2.32
c175 35 0 1.8874e-19 $X=7.365 $Y=2.405
r176 77 78 62.6163 $w=3.31e-07 $l=4.3e-07 $layer=POLY_cond $X=11.405 $Y=1.517
+ $X2=11.835 $Y2=1.517
r177 76 77 8.00906 $w=3.31e-07 $l=5.5e-08 $layer=POLY_cond $X=11.35 $Y=1.517
+ $X2=11.405 $Y2=1.517
r178 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.905
+ $Y=1.515 $X2=9.905 $Y2=1.515
r179 64 65 8.82039 $w=3.18e-07 $l=1.75e-07 $layer=LI1_cond $X=7.525 $Y=1.11
+ $X2=7.525 $Y2=1.285
r180 61 64 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=7.525 $Y=1.02
+ $X2=7.525 $Y2=1.11
r181 56 59 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=6.66 $Y=2.405
+ $X2=6.66 $Y2=2.525
r182 54 74 39.3172 $w=3.31e-07 $l=2.7e-07 $layer=POLY_cond $X=10.585 $Y=1.517
+ $X2=10.855 $Y2=1.517
r183 54 72 23.2991 $w=3.31e-07 $l=1.6e-07 $layer=POLY_cond $X=10.585 $Y=1.517
+ $X2=10.425 $Y2=1.517
r184 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.585
+ $Y=1.515 $X2=10.585 $Y2=1.515
r185 51 67 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.515
+ $X2=9.865 $Y2=1.515
r186 51 53 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=9.95 $Y=1.515
+ $X2=10.585 $Y2=1.515
r187 50 67 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.35
+ $X2=9.865 $Y2=1.515
r188 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.865 $Y=1.18
+ $X2=9.865 $Y2=1.35
r189 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.78 $Y=1.095
+ $X2=9.865 $Y2=1.18
r190 47 48 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.78 $Y=1.095
+ $X2=9.555 $Y2=1.095
r191 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.47 $Y=1.01
+ $X2=9.555 $Y2=1.095
r192 45 46 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.47 $Y=0.765
+ $X2=9.47 $Y2=1.01
r193 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.385 $Y=0.68
+ $X2=9.47 $Y2=0.765
r194 43 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.385 $Y=0.68
+ $X2=8.875 $Y2=0.68
r195 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.79 $Y=0.765
+ $X2=8.875 $Y2=0.68
r196 41 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.79 $Y=0.765
+ $X2=8.79 $Y2=0.935
r197 40 61 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.685 $Y=1.02
+ $X2=7.525 $Y2=1.02
r198 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.705 $Y=1.02
+ $X2=8.79 $Y2=0.935
r199 39 40 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.705 $Y=1.02
+ $X2=7.685 $Y2=1.02
r200 38 65 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=7.45 $Y=2.32
+ $X2=7.45 $Y2=1.285
r201 36 56 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=2.405
+ $X2=6.66 $Y2=2.405
r202 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=2.405
+ $X2=7.45 $Y2=2.32
r203 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.365 $Y=2.405
+ $X2=6.785 $Y2=2.405
r204 32 78 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=11.835 $Y=1.35
+ $X2=11.835 $Y2=1.517
r205 32 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.835 $Y=1.35
+ $X2=11.835 $Y2=0.87
r206 29 77 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=11.405 $Y=1.35
+ $X2=11.405 $Y2=1.517
r207 29 31 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.405 $Y=1.35
+ $X2=11.405 $Y2=0.87
r208 25 76 17.0024 $w=1.8e-07 $l=1.68e-07 $layer=POLY_cond $X=11.35 $Y=1.685
+ $X2=11.35 $Y2=1.517
r209 25 27 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=11.35 $Y=1.685
+ $X2=11.35 $Y2=2.4
r210 21 76 65.5287 $w=3.31e-07 $l=4.5e-07 $layer=POLY_cond $X=10.9 $Y=1.517
+ $X2=11.35 $Y2=1.517
r211 21 74 6.55287 $w=3.31e-07 $l=4.5e-08 $layer=POLY_cond $X=10.9 $Y=1.517
+ $X2=10.855 $Y2=1.517
r212 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.9 $Y=1.68
+ $X2=10.9 $Y2=2.4
r213 18 74 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=10.855 $Y=1.35
+ $X2=10.855 $Y2=1.517
r214 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.855 $Y=1.35
+ $X2=10.855 $Y2=0.87
r215 15 72 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=10.425 $Y=1.35
+ $X2=10.425 $Y2=1.517
r216 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.425 $Y=1.35
+ $X2=10.425 $Y2=0.87
r217 11 72 21.1148 $w=3.31e-07 $l=1.45e-07 $layer=POLY_cond $X=10.28 $Y=1.517
+ $X2=10.425 $Y2=1.517
r218 11 68 54.6073 $w=3.31e-07 $l=3.75e-07 $layer=POLY_cond $X=10.28 $Y=1.517
+ $X2=9.905 $Y2=1.517
r219 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.28 $Y=1.68
+ $X2=10.28 $Y2=2.4
r220 7 68 10.9215 $w=3.31e-07 $l=7.5e-08 $layer=POLY_cond $X=9.83 $Y=1.517
+ $X2=9.905 $Y2=1.517
r221 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.83 $Y=1.68 $X2=9.83
+ $Y2=2.4
r222 2 59 600 $w=1.7e-07 $l=7.57166e-07 $layer=licon1_PDIFF $count=1 $X=6.34
+ $Y=1.895 $X2=6.62 $Y2=2.525
r223 1 64 182 $w=1.7e-07 $l=5.7639e-07 $layer=licon1_NDIFF $count=1 $X=7.32
+ $Y=0.625 $X2=7.52 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%CI 3 7 8 11 12 13
r38 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.815 $Y=1.515
+ $X2=12.815 $Y2=1.68
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.815 $Y=1.515
+ $X2=12.815 $Y2=1.35
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.815
+ $Y=1.515 $X2=12.815 $Y2=1.515
r41 8 12 5.01062 $w=3.43e-07 $l=1.5e-07 $layer=LI1_cond $X=12.807 $Y=1.665
+ $X2=12.807 $Y2=1.515
r42 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.905 $Y=0.92
+ $X2=12.905 $Y2=1.35
r43 3 14 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=12.775 $Y=2.34
+ $X2=12.775 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_1278_102# 1 2 9 11 13 16 18 20 23 25 27 28
+ 30 33 35 38 39 41 42 44 45 46 48 49 52 53 58 64 66 70 79
c216 66 0 5.40791e-20 $X=8.21 $Y=2.26
c217 18 0 1.44963e-19 $X=13.935 $Y=1.35
r218 79 80 2.19757 $w=3.29e-07 $l=1.5e-08 $layer=POLY_cond $X=14.795 $Y=1.515
+ $X2=14.81 $Y2=1.515
r219 78 79 62.997 $w=3.29e-07 $l=4.3e-07 $layer=POLY_cond $X=14.365 $Y=1.515
+ $X2=14.795 $Y2=1.515
r220 77 78 2.19757 $w=3.29e-07 $l=1.5e-08 $layer=POLY_cond $X=14.35 $Y=1.515
+ $X2=14.365 $Y2=1.515
r221 74 75 18.3131 $w=3.29e-07 $l=1.25e-07 $layer=POLY_cond $X=13.81 $Y=1.515
+ $X2=13.935 $Y2=1.515
r222 73 74 44.6839 $w=3.29e-07 $l=3.05e-07 $layer=POLY_cond $X=13.505 $Y=1.515
+ $X2=13.81 $Y2=1.515
r223 66 68 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.21 $Y=2.26
+ $X2=8.21 $Y2=2.355
r224 62 64 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.54 $Y=0.72
+ $X2=6.705 $Y2=0.72
r225 59 77 27.8359 $w=3.29e-07 $l=1.9e-07 $layer=POLY_cond $X=14.16 $Y=1.515
+ $X2=14.35 $Y2=1.515
r226 59 75 32.9635 $w=3.29e-07 $l=2.25e-07 $layer=POLY_cond $X=14.16 $Y=1.515
+ $X2=13.935 $Y2=1.515
r227 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14.16
+ $Y=1.515 $X2=14.16 $Y2=1.515
r228 56 73 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=13.48 $Y=1.515
+ $X2=13.505 $Y2=1.515
r229 56 71 17.5805 $w=3.29e-07 $l=1.2e-07 $layer=POLY_cond $X=13.48 $Y=1.515
+ $X2=13.36 $Y2=1.515
r230 55 58 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.48 $Y=1.515
+ $X2=14.16 $Y2=1.515
r231 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.48
+ $Y=1.515 $X2=13.48 $Y2=1.515
r232 53 55 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=13.385 $Y=1.515
+ $X2=13.48 $Y2=1.515
r233 52 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.3 $Y=1.35
+ $X2=13.385 $Y2=1.515
r234 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=13.3 $Y=0.84
+ $X2=13.3 $Y2=1.35
r235 50 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.125 $Y=0.755
+ $X2=12.04 $Y2=0.755
r236 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.215 $Y=0.755
+ $X2=13.3 $Y2=0.84
r237 49 50 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=13.215 $Y=0.755
+ $X2=12.125 $Y2=0.755
r238 47 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.04 $Y=0.84
+ $X2=12.04 $Y2=0.755
r239 47 48 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=12.04 $Y=0.84
+ $X2=12.04 $Y2=2.27
r240 45 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.955 $Y=0.755
+ $X2=12.04 $Y2=0.755
r241 45 46 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=11.955 $Y=0.755
+ $X2=9.895 $Y2=0.755
r242 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.81 $Y=0.67
+ $X2=9.895 $Y2=0.755
r243 43 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.81 $Y=0.425
+ $X2=9.81 $Y2=0.67
r244 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.725 $Y=0.34
+ $X2=9.81 $Y2=0.425
r245 41 42 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=9.725 $Y=0.34
+ $X2=8.535 $Y2=0.34
r246 40 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.375 $Y=2.355
+ $X2=8.21 $Y2=2.355
r247 39 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.955 $Y=2.355
+ $X2=12.04 $Y2=2.27
r248 39 40 233.561 $w=1.68e-07 $l=3.58e-06 $layer=LI1_cond $X=11.955 $Y=2.355
+ $X2=8.375 $Y2=2.355
r249 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.45 $Y=0.425
+ $X2=8.535 $Y2=0.34
r250 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.45 $Y=0.425
+ $X2=8.45 $Y2=0.595
r251 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.365 $Y=0.68
+ $X2=8.45 $Y2=0.595
r252 35 64 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=8.365 $Y=0.68
+ $X2=6.705 $Y2=0.68
r253 31 80 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.81 $Y=1.68
+ $X2=14.81 $Y2=1.515
r254 31 33 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=14.81 $Y=1.68
+ $X2=14.81 $Y2=2.4
r255 28 79 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.795 $Y=1.35
+ $X2=14.795 $Y2=1.515
r256 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.795 $Y=1.35
+ $X2=14.795 $Y2=0.87
r257 25 78 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.365 $Y=1.35
+ $X2=14.365 $Y2=1.515
r258 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.365 $Y=1.35
+ $X2=14.365 $Y2=0.87
r259 21 77 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.35 $Y=1.68
+ $X2=14.35 $Y2=1.515
r260 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=14.35 $Y=1.68
+ $X2=14.35 $Y2=2.4
r261 18 75 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.935 $Y=1.35
+ $X2=13.935 $Y2=1.515
r262 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.935 $Y=1.35
+ $X2=13.935 $Y2=0.87
r263 14 74 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.81 $Y=1.68
+ $X2=13.81 $Y2=1.515
r264 14 16 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=13.81 $Y=1.68
+ $X2=13.81 $Y2=2.4
r265 11 73 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.505 $Y=1.35
+ $X2=13.505 $Y2=1.515
r266 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.505 $Y=1.35
+ $X2=13.505 $Y2=0.87
r267 7 71 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.36 $Y=1.68
+ $X2=13.36 $Y2=1.515
r268 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=13.36 $Y=1.68
+ $X2=13.36 $Y2=2.4
r269 2 66 300 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_PDIFF $count=2 $X=7.575
+ $Y=2.115 $X2=8.21 $Y2=2.26
r270 1 62 182 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.51 $X2=6.54 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%VPWR 1 2 3 4 5 6 7 8 9 30 36 40 46 48 50 55 58
+ 62 63 64 66 71 76 104 108 114 117 124 129 132 136 139 141 145
r167 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r168 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r169 138 139 13.167 $w=4.63e-07 $l=3.15e-07 $layer=LI1_cond $X=11.81 $Y=3.182
+ $X2=12.125 $Y2=3.182
r170 134 138 1.28611 $w=4.63e-07 $l=5e-08 $layer=LI1_cond $X=11.76 $Y=3.182
+ $X2=11.81 $Y2=3.182
r171 134 136 11.8809 $w=4.63e-07 $l=2.65e-07 $layer=LI1_cond $X=11.76 $Y=3.182
+ $X2=11.495 $Y2=3.182
r172 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r173 131 132 12.3953 $w=4.63e-07 $l=2.85e-07 $layer=LI1_cond $X=9.4 $Y=3.182
+ $X2=9.685 $Y2=3.182
r174 127 131 1.02888 $w=4.63e-07 $l=4e-08 $layer=LI1_cond $X=9.36 $Y=3.182
+ $X2=9.4 $Y2=3.182
r175 127 129 11.3664 $w=4.63e-07 $l=2.45e-07 $layer=LI1_cond $X=9.36 $Y=3.182
+ $X2=9.115 $Y2=3.182
r176 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r177 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r178 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r179 117 120 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=1.745 $Y=3.055
+ $X2=1.745 $Y2=3.33
r180 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r181 112 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r182 112 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r183 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r184 109 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.25 $Y=3.33
+ $X2=14.085 $Y2=3.33
r185 109 111 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=14.25 $Y=3.33
+ $X2=14.64 $Y2=3.33
r186 108 144 3.9577 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=14.95 $Y=3.33
+ $X2=15.155 $Y2=3.33
r187 108 111 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.95 $Y=3.33
+ $X2=14.64 $Y2=3.33
r188 107 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r189 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r190 104 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.92 $Y=3.33
+ $X2=14.085 $Y2=3.33
r191 104 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=13.92 $Y=3.33
+ $X2=13.68 $Y2=3.33
r192 103 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r193 103 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r194 102 139 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=12.125 $Y2=3.33
r195 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r196 99 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r197 98 136 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=11.495 $Y2=3.33
r198 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r199 95 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r200 95 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r201 94 132 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.32 $Y=3.33
+ $X2=9.685 $Y2=3.33
r202 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r203 91 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r204 90 129 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=9.115 $Y2=3.33
r205 90 91 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r206 88 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r207 87 90 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=8.88
+ $Y2=3.33
r208 87 88 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r209 85 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=3.33
+ $X2=5.49 $Y2=3.33
r210 85 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.655 $Y=3.33 $X2=6
+ $Y2=3.33
r211 83 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r212 82 83 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r213 80 83 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=5.04 $Y2=3.33
r214 80 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r215 79 82 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=5.04 $Y2=3.33
r216 79 80 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r217 77 120 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.745 $Y2=3.33
r218 77 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.16 $Y2=3.33
r219 76 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.49 $Y2=3.33
r220 76 82 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.325 $Y=3.33
+ $X2=5.04 $Y2=3.33
r221 75 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r222 75 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r224 72 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.69 $Y2=3.33
r225 72 74 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r226 71 120 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.745 $Y2=3.33
r227 71 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r228 69 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r229 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r230 66 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.69 $Y2=3.33
r231 66 68 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r232 64 91 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=8.88 $Y2=3.33
r233 64 88 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=6 $Y2=3.33
r234 62 102 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=12.92 $Y=3.33
+ $X2=12.72 $Y2=3.33
r235 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.92 $Y=3.33
+ $X2=13.085 $Y2=3.33
r236 61 106 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.25 $Y=3.33
+ $X2=13.68 $Y2=3.33
r237 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.25 $Y=3.33
+ $X2=13.085 $Y2=3.33
r238 59 98 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=10.755 $Y=3.33
+ $X2=11.28 $Y2=3.33
r239 58 94 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=10.425 $Y=3.33
+ $X2=10.32 $Y2=3.33
r240 57 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.755 $Y2=3.33
r241 57 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.425 $Y2=3.33
r242 55 57 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=10.59 $Y=3.04
+ $X2=10.59 $Y2=3.33
r243 50 53 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.075 $Y=1.985
+ $X2=15.075 $Y2=2.815
r244 48 144 3.18546 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.155 $Y2=3.33
r245 48 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.075 $Y2=2.815
r246 44 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.085 $Y=3.245
+ $X2=14.085 $Y2=3.33
r247 44 46 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=14.085 $Y=3.245
+ $X2=14.085 $Y2=2.355
r248 40 43 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=13.085 $Y=2.035
+ $X2=13.085 $Y2=2.815
r249 38 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.085 $Y=3.245
+ $X2=13.085 $Y2=3.33
r250 38 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.085 $Y=3.245
+ $X2=13.085 $Y2=2.815
r251 34 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.49 $Y=3.245
+ $X2=5.49 $Y2=3.33
r252 34 36 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.49 $Y=3.245
+ $X2=5.49 $Y2=2.385
r253 30 33 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.135
+ $X2=0.69 $Y2=2.815
r254 28 114 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r255 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.815
r256 9 53 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.9
+ $Y=1.84 $X2=15.035 $Y2=2.815
r257 9 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.9
+ $Y=1.84 $X2=15.035 $Y2=1.985
r258 8 46 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=13.9
+ $Y=1.84 $X2=14.085 $Y2=2.355
r259 7 43 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=12.865
+ $Y=1.84 $X2=13.085 $Y2=2.815
r260 7 40 300 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_PDIFF $count=2 $X=12.865
+ $Y=1.84 $X2=13.085 $Y2=2.035
r261 6 138 600 $w=1.7e-07 $l=1.36754e-06 $layer=licon1_PDIFF $count=1 $X=11.44
+ $Y=1.84 $X2=11.81 $Y2=3.035
r262 5 55 600 $w=1.7e-07 $l=1.30537e-06 $layer=licon1_PDIFF $count=1 $X=10.37
+ $Y=1.84 $X2=10.59 $Y2=3.04
r263 4 131 600 $w=1.7e-07 $l=1.35437e-06 $layer=licon1_PDIFF $count=1 $X=9.06
+ $Y=1.84 $X2=9.4 $Y2=3.035
r264 3 36 300 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=2 $X=5.345
+ $Y=1.84 $X2=5.49 $Y2=2.385
r265 2 117 600 $w=1.7e-07 $l=1.31787e-06 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.81 $X2=1.745 $Y2=3.055
r266 1 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.815
r267 1 30 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_200_74# 1 2 3 4 15 17 19 21 22 23 26 28 29
+ 31 32 35 39 41 42
c110 19 0 5.85186e-20 $X=1.18 $Y=2.135
c111 17 0 1.1782e-19 $X=1.18 $Y=2.63
c112 15 0 1.40087e-19 $X=1.14 $Y=0.515
r113 42 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.33 $Y=2.715 $X2=3.33
+ $Y2=2.795
r114 39 40 8.26042 $w=1.92e-07 $l=1.3e-07 $layer=LI1_cond $X=1.92 $Y=0.895
+ $X2=2.05 $Y2=0.895
r115 33 35 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=3.285 $Y=0.425
+ $X2=3.285 $Y2=0.835
r116 31 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.155 $Y=0.34
+ $X2=3.285 $Y2=0.425
r117 31 32 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.155 $Y=0.34
+ $X2=2.135 $Y2=0.34
r118 30 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=2.715
+ $X2=1.92 $Y2=2.715
r119 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=2.715
+ $X2=3.33 $Y2=2.715
r120 29 30 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.165 $Y=2.715
+ $X2=2.005 $Y2=2.715
r121 28 40 1.44825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.05 $Y=0.79
+ $X2=2.05 $Y2=0.895
r122 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=0.425
+ $X2=2.135 $Y2=0.34
r123 27 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.05 $Y=0.425
+ $X2=2.05 $Y2=0.79
r124 26 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=2.63
+ $X2=1.92 $Y2=2.715
r125 25 39 1.44825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.92 $Y=1 $X2=1.92
+ $Y2=0.895
r126 25 26 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=1.92 $Y=1 $X2=1.92
+ $Y2=2.63
r127 24 38 4.60552 $w=1.7e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.345 $Y=2.715
+ $X2=1.18 $Y2=2.805
r128 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=2.715
+ $X2=1.92 $Y2=2.715
r129 23 24 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.835 $Y=2.715
+ $X2=1.345 $Y2=2.715
r130 21 39 5.05061 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.895
+ $X2=1.92 $Y2=0.895
r131 21 22 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=1.835 $Y=0.895
+ $X2=1.305 $Y2=0.895
r132 17 38 3.16065 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=1.18 $Y=2.63
+ $X2=1.18 $Y2=2.805
r133 17 19 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.18 $Y=2.63
+ $X2=1.18 $Y2=2.135
r134 13 22 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=1.14 $Y=0.79
+ $X2=1.305 $Y2=0.895
r135 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=0.79
+ $X2=1.14 $Y2=0.515
r136 4 45 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=1.81 $X2=3.33 $Y2=2.795
r137 3 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.96 $X2=1.18 $Y2=2.815
r138 3 19 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.96 $X2=1.18 $Y2=2.135
r139 2 35 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.11
+ $Y=0.57 $X2=3.25 $Y2=0.835
r140 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_430_362# 1 2 3 4 14 16 19 21 22 23 26 33 35
c84 23 0 1.26128e-19 $X=4.367 $Y=2.072
c85 21 0 1.75426e-19 $X=4.23 $Y=2.375
c86 16 0 1.11098e-19 $X=2.34 $Y=1.955
r87 31 33 8.2628 $w=2.63e-07 $l=1.9e-07 $layer=LI1_cond $X=4.23 $Y=1.177
+ $X2=4.42 $Y2=1.177
r88 27 33 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.42 $Y=1.31
+ $X2=4.42 $Y2=1.177
r89 27 35 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.42 $Y=1.31
+ $X2=4.42 $Y2=1.935
r90 24 26 7.96233 $w=2.73e-07 $l=1.9e-07 $layer=LI1_cond $X=4.367 $Y=2.29
+ $X2=4.367 $Y2=2.1
r91 23 35 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=4.367 $Y=2.072
+ $X2=4.367 $Y2=1.935
r92 23 26 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=4.367 $Y=2.072
+ $X2=4.367 $Y2=2.1
r93 21 38 5.44791 $w=2.73e-07 $l=1.3e-07 $layer=LI1_cond $X=4.367 $Y=2.375
+ $X2=4.367 $Y2=2.505
r94 21 24 3.5621 $w=2.73e-07 $l=8.5e-08 $layer=LI1_cond $X=4.367 $Y=2.375
+ $X2=4.367 $Y2=2.29
r95 21 22 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=4.23 $Y=2.375
+ $X2=2.505 $Y2=2.375
r96 19 29 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.39 $Y=0.895
+ $X2=2.39 $Y2=1.79
r97 16 29 7.72582 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=1.955
+ $X2=2.34 $Y2=1.79
r98 14 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.34 $Y=2.29
+ $X2=2.505 $Y2=2.375
r99 14 16 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.34 $Y=2.29
+ $X2=2.34 $Y2=1.955
r100 4 38 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.81 $X2=4.315 $Y2=2.505
r101 4 26 600 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.81 $X2=4.315 $Y2=2.1
r102 3 16 300 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=2 $X=2.15
+ $Y=1.81 $X2=2.34 $Y2=1.955
r103 2 31 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.65 $X2=4.23 $Y2=1.135
r104 1 19 182 $w=1.7e-07 $l=5.09166e-07 $layer=licon1_NDIFF $count=1 $X=2.205
+ $Y=0.47 $X2=2.39 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%A_1183_102# 1 2 3 13 14 20 23 26 27 33 34 38
c107 34 0 5.38428e-20 $X=9.36 $Y=1.665
r108 34 41 14.808 $w=2.76e-07 $l=3.35e-07 $layer=LI1_cond $X=9.215 $Y=1.665
+ $X2=9.215 $Y2=2
r109 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r110 30 38 3.00637 $w=2.28e-07 $l=6e-08 $layer=LI1_cond $X=6 $Y=1.665 $X2=6.06
+ $Y2=1.665
r111 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=1.665 $X2=6
+ $Y2=1.665
r112 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=1.665
+ $X2=6 $Y2=1.665
r113 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=9.36 $Y2=1.665
r114 26 27 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=6.145 $Y2=1.665
r115 23 25 9.50985 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.04 $Y=0.68
+ $X2=6.04 $Y2=0.875
r116 18 34 6.87116 $w=2.76e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.13 $Y=1.55
+ $X2=9.215 $Y2=1.665
r117 18 20 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.13 $Y=1.55
+ $X2=9.13 $Y2=1.1
r118 14 41 2.62467 $w=2e-07 $l=1.7e-07 $layer=LI1_cond $X=9.045 $Y=2 $X2=9.215
+ $Y2=2
r119 14 16 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=9.045 $Y=2 $X2=8.745
+ $Y2=2
r120 13 25 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.06 $Y=1.02
+ $X2=6.06 $Y2=0.875
r121 11 38 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.06 $Y=1.55
+ $X2=6.06 $Y2=1.665
r122 11 13 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.06 $Y=1.55
+ $X2=6.06 $Y2=1.02
r123 3 16 600 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=2.115 $X2=8.745 $Y2=2
r124 2 20 182 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=1 $X=8.985
+ $Y=0.6 $X2=9.13 $Y2=1.1
r125 1 23 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=5.915
+ $Y=0.51 $X2=6.04 $Y2=0.68
r126 1 13 182 $w=1.7e-07 $l=5.77971e-07 $layer=licon1_NDIFF $count=1 $X=5.915
+ $Y=0.51 $X2=6.06 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%COUT 1 2 3 4 13 17 23 26 27 30
r46 27 30 4.90119 $w=4.33e-07 $l=1.85e-07 $layer=LI1_cond $X=11.177 $Y=1.85
+ $X2=11.177 $Y2=1.665
r47 27 29 2.73535 $w=4.35e-07 $l=1.25e-07 $layer=LI1_cond $X=11.177 $Y=1.85
+ $X2=11.177 $Y2=1.975
r48 25 30 10.7296 $w=4.33e-07 $l=4.05e-07 $layer=LI1_cond $X=11.177 $Y=1.26
+ $X2=11.177 $Y2=1.665
r49 25 26 1.09397 $w=4.35e-07 $l=1.25e-07 $layer=LI1_cond $X=11.177 $Y=1.26
+ $X2=11.177 $Y2=1.135
r50 21 26 9.00716 $w=2.1e-07 $l=2.18e-07 $layer=LI1_cond $X=11.395 $Y=1.135
+ $X2=11.177 $Y2=1.135
r51 21 23 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=11.395 $Y=1.135
+ $X2=11.62 $Y2=1.135
r52 17 26 9.00716 $w=2.1e-07 $l=2.36155e-07 $layer=LI1_cond $X=10.96 $Y=1.095
+ $X2=11.177 $Y2=1.135
r53 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.96 $Y=1.095
+ $X2=10.64 $Y2=1.095
r54 13 29 4.74857 $w=2.5e-07 $l=2.17e-07 $layer=LI1_cond $X=10.96 $Y=1.975
+ $X2=11.177 $Y2=1.975
r55 13 15 41.7184 $w=2.48e-07 $l=9.05e-07 $layer=LI1_cond $X=10.96 $Y=1.975
+ $X2=10.055 $Y2=1.975
r56 4 29 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=10.99
+ $Y=1.84 $X2=11.125 $Y2=2.015
r57 3 15 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.92
+ $Y=1.84 $X2=10.055 $Y2=2.015
r58 2 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=11.48
+ $Y=0.5 $X2=11.62 $Y2=1.095
r59 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=10.5
+ $Y=0.5 $X2=10.64 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%SUM 1 2 3 4 13 15 19 21 23 24 27 30 34 35 36
+ 37 44
c63 19 0 1.44963e-19 $X=13.72 $Y=0.645
r64 42 44 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=14.587 $Y=2.02
+ $X2=14.587 $Y2=2.035
r65 36 37 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.587 $Y=2.405
+ $X2=14.587 $Y2=2.775
r66 35 42 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=14.587 $Y=1.935
+ $X2=14.587 $Y2=2.02
r67 35 36 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=14.587 $Y=2.07
+ $X2=14.587 $Y2=2.405
r68 35 44 1.20404 $w=3.33e-07 $l=3.5e-08 $layer=LI1_cond $X=14.587 $Y=2.07
+ $X2=14.587 $Y2=2.035
r69 30 35 3.22182 $w=2.92e-07 $l=1.0015e-07 $layer=LI1_cond $X=14.62 $Y=1.85
+ $X2=14.587 $Y2=1.935
r70 29 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.62 $Y=1.18
+ $X2=14.62 $Y2=1.095
r71 29 30 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=14.62 $Y=1.18
+ $X2=14.62 $Y2=1.85
r72 25 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.62 $Y=1.01
+ $X2=14.62 $Y2=1.095
r73 25 27 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=14.62 $Y=1.01
+ $X2=14.62 $Y2=0.645
r74 23 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.495 $Y=1.095
+ $X2=14.62 $Y2=1.095
r75 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.495 $Y=1.095
+ $X2=13.805 $Y2=1.095
r76 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.75 $Y=1.935
+ $X2=13.585 $Y2=1.935
r77 21 35 3.35233 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=14.42 $Y=1.935
+ $X2=14.587 $Y2=1.935
r78 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.42 $Y=1.935
+ $X2=13.75 $Y2=1.935
r79 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.68 $Y=1.01
+ $X2=13.805 $Y2=1.095
r80 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=13.68 $Y=1.01
+ $X2=13.68 $Y2=0.645
r81 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.585 $Y=2.02
+ $X2=13.585 $Y2=1.935
r82 13 15 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=13.585 $Y=2.02
+ $X2=13.585 $Y2=2.815
r83 4 35 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.44
+ $Y=1.84 $X2=14.585 $Y2=2.015
r84 4 37 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=14.44
+ $Y=1.84 $X2=14.585 $Y2=2.815
r85 3 32 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=13.45
+ $Y=1.84 $X2=13.585 $Y2=2.015
r86 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.45
+ $Y=1.84 $X2=13.585 $Y2=2.815
r87 2 34 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=14.44
+ $Y=0.5 $X2=14.58 $Y2=1.095
r88 2 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=14.44
+ $Y=0.5 $X2=14.58 $Y2=0.645
r89 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.58
+ $Y=0.5 $X2=13.72 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_4%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54 58
+ 60 62 65 66 68 69 71 72 74 75 77 78 79 85 108 112 117 123 126 129 133
r161 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r162 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r163 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r164 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r165 121 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r166 121 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=14.16 $Y2=0
r167 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r168 118 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.315 $Y=0
+ $X2=14.15 $Y2=0
r169 118 120 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=14.315 $Y=0
+ $X2=14.64 $Y2=0
r170 117 132 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=14.915 $Y=0
+ $X2=15.137 $Y2=0
r171 117 120 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=14.915 $Y=0
+ $X2=14.64 $Y2=0
r172 116 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r173 116 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r174 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r175 113 126 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=13.375 $Y=0
+ $X2=13.205 $Y2=0
r176 113 115 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.375 $Y=0
+ $X2=13.68 $Y2=0
r177 112 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.985 $Y=0
+ $X2=14.15 $Y2=0
r178 112 115 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.985 $Y=0
+ $X2=13.68 $Y2=0
r179 111 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r180 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r181 108 126 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=13.035 $Y=0
+ $X2=13.205 $Y2=0
r182 108 110 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.035 $Y=0
+ $X2=12.72 $Y2=0
r183 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r184 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r185 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r186 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r187 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.8 $Y2=0
r188 100 101 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r189 97 100 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=9.84
+ $Y2=0
r190 97 98 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r191 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r192 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r193 92 95 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r194 92 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r195 91 94 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r196 91 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r197 89 123 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=1.665 $Y2=0
r198 89 91 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=2.16 $Y2=0
r199 88 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r200 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 85 123 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=1.665 $Y2=0
r202 85 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r203 83 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r204 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r205 79 101 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=9.84 $Y2=0
r206 79 98 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=7.68 $Y=0 $X2=5.04
+ $Y2=0
r207 77 106 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.965 $Y=0
+ $X2=11.76 $Y2=0
r208 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.965 $Y=0
+ $X2=12.13 $Y2=0
r209 76 110 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.72 $Y2=0
r210 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.13 $Y2=0
r211 74 103 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=0
+ $X2=10.8 $Y2=0
r212 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=0
+ $X2=11.13 $Y2=0
r213 73 106 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=11.295 $Y=0
+ $X2=11.76 $Y2=0
r214 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.295 $Y=0
+ $X2=11.13 $Y2=0
r215 71 100 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=9.84 $Y2=0
r216 71 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=10.19 $Y2=0
r217 70 103 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.8 $Y2=0
r218 70 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.19 $Y2=0
r219 68 94 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.56
+ $Y2=0
r220 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.75
+ $Y2=0
r221 67 97 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=5.04 $Y2=0
r222 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.915 $Y=0 $X2=4.75
+ $Y2=0
r223 65 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r224 65 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r225 64 87 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.2
+ $Y2=0
r226 64 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r227 60 132 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.08 $Y=0.085
+ $X2=15.137 $Y2=0
r228 60 62 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=15.08 $Y=0.085
+ $X2=15.08 $Y2=0.645
r229 56 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.15 $Y=0.085
+ $X2=14.15 $Y2=0
r230 56 58 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=14.15 $Y=0.085
+ $X2=14.15 $Y2=0.7
r231 52 126 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0
r232 52 54 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0.335
r233 48 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0
r234 48 50 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0.335
r235 44 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.13 $Y=0.085
+ $X2=11.13 $Y2=0
r236 44 46 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=11.13 $Y=0.085
+ $X2=11.13 $Y2=0.335
r237 40 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.19 $Y=0.085
+ $X2=10.19 $Y2=0
r238 40 42 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=10.19 $Y=0.085
+ $X2=10.19 $Y2=0.335
r239 36 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0
r240 36 38 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0.37
r241 32 123 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0
r242 32 34 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.665 $Y=0.085
+ $X2=1.665 $Y2=0.455
r243 28 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r244 28 30 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.495
r245 9 62 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=14.87
+ $Y=0.5 $X2=15.08 $Y2=0.645
r246 8 58 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=14.01
+ $Y=0.5 $X2=14.15 $Y2=0.7
r247 7 54 182 $w=1.7e-07 $l=3.60347e-07 $layer=licon1_NDIFF $count=1 $X=12.98
+ $Y=0.6 $X2=13.205 $Y2=0.335
r248 6 50 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=11.91
+ $Y=0.5 $X2=12.13 $Y2=0.335
r249 5 46 182 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=1 $X=10.93
+ $Y=0.5 $X2=11.13 $Y2=0.335
r250 4 42 182 $w=1.7e-07 $l=7.712e-07 $layer=licon1_NDIFF $count=1 $X=9.5 $Y=0.6
+ $X2=10.15 $Y2=0.335
r251 3 38 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.225 $X2=4.75 $Y2=0.37
r252 2 34 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.31 $X2=1.705 $Y2=0.455
r253 1 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends


* File: sky130_fd_sc_ms__o211ai_1.pxi.spice
* Created: Wed Sep  2 12:20:32 2020
* 
x_PM_SKY130_FD_SC_MS__O211AI_1%A1 N_A1_M1004_g N_A1_M1006_g A1 N_A1_c_52_n
+ N_A1_c_53_n PM_SKY130_FD_SC_MS__O211AI_1%A1
x_PM_SKY130_FD_SC_MS__O211AI_1%A2 N_A2_M1005_g N_A2_M1000_g A2 A2 A2 A2
+ N_A2_c_81_n A2 PM_SKY130_FD_SC_MS__O211AI_1%A2
x_PM_SKY130_FD_SC_MS__O211AI_1%B1 N_B1_M1001_g N_B1_M1003_g B1 B1 B1
+ N_B1_c_122_n B1 PM_SKY130_FD_SC_MS__O211AI_1%B1
x_PM_SKY130_FD_SC_MS__O211AI_1%C1 N_C1_M1007_g N_C1_M1002_g C1 N_C1_c_160_n
+ N_C1_c_161_n PM_SKY130_FD_SC_MS__O211AI_1%C1
x_PM_SKY130_FD_SC_MS__O211AI_1%VPWR N_VPWR_M1004_s N_VPWR_M1003_d N_VPWR_c_192_n
+ N_VPWR_c_193_n N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_196_n VPWR
+ N_VPWR_c_197_n N_VPWR_c_191_n PM_SKY130_FD_SC_MS__O211AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O211AI_1%Y N_Y_M1007_d N_Y_M1005_d N_Y_M1002_d N_Y_c_226_n
+ N_Y_c_227_n N_Y_c_228_n N_Y_c_229_n N_Y_c_224_n N_Y_c_231_n Y Y N_Y_c_225_n
+ PM_SKY130_FD_SC_MS__O211AI_1%Y
x_PM_SKY130_FD_SC_MS__O211AI_1%A_31_74# N_A_31_74#_M1006_s N_A_31_74#_M1000_d
+ N_A_31_74#_c_270_n N_A_31_74#_c_271_n N_A_31_74#_c_272_n N_A_31_74#_c_273_n
+ PM_SKY130_FD_SC_MS__O211AI_1%A_31_74#
x_PM_SKY130_FD_SC_MS__O211AI_1%VGND N_VGND_M1006_d N_VGND_c_296_n VGND
+ N_VGND_c_297_n N_VGND_c_298_n N_VGND_c_299_n N_VGND_c_300_n
+ PM_SKY130_FD_SC_MS__O211AI_1%VGND
cc_1 VNB N_A1_M1004_g 0.00188936f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A1_M1006_g 0.0310333f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A1_c_52_n 0.0050357f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_A1_c_53_n 0.0591131f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_5 VNB N_A2_M1005_g 0.00186418f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_6 VNB N_A2_M1000_g 0.0224026f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_7 VNB A2 0.0130937f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A2_c_81_n 0.0286147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A2 4.83307e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1001_g 0.024159f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_11 VNB N_B1_M1003_g 0.00196134f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_12 VNB B1 0.00339768f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB B1 0.00548062f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_14 VNB N_B1_c_122_n 0.0287823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C1_M1002_g 0.00715508f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_16 VNB C1 0.00370468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C1_c_160_n 0.0358943f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_18 VNB N_C1_c_161_n 0.0236718f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_19 VNB N_VPWR_c_191_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_224_n 0.0310722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_225_n 0.0239756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_31_74#_c_270_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_A_31_74#_c_271_n 0.00796953f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_24 VNB N_A_31_74#_c_272_n 0.00898165f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_25 VNB N_A_31_74#_c_273_n 0.00260143f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_26 VNB N_VGND_c_296_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_27 VNB N_VGND_c_297_n 0.0197879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_298_n 0.0547577f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_29 VNB N_VGND_c_299_n 0.194045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_300_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_A1_M1004_g 0.0266416f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_32 VPB N_A1_c_52_n 0.00916391f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_33 VPB N_A2_M1005_g 0.0259251f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_34 VPB A2 0.00329461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_B1_M1003_g 0.0255198f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_36 VPB N_C1_M1002_g 0.0286321f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_37 VPB N_VPWR_c_192_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_38 VPB N_VPWR_c_193_n 0.0495887f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_39 VPB N_VPWR_c_194_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_40 VPB N_VPWR_c_195_n 0.0383522f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_41 VPB N_VPWR_c_196_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_197_n 0.0246348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_191_n 0.0657523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_Y_c_226_n 0.00339147f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_45 VPB N_Y_c_227_n 0.00791398f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_46 VPB N_Y_c_228_n 0.00551202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_229_n 0.0542942f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_48 VPB N_Y_c_224_n 0.00725366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_Y_c_231_n 0.0210267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 N_A1_M1004_g N_A2_M1005_g 0.0422488f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_51 N_A1_M1006_g N_A2_M1000_g 0.0278145f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_52 N_A1_c_52_n A2 0.0230252f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_53 N_A1_c_53_n A2 0.00304525f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_54 N_A1_c_52_n N_A2_c_81_n 2.46571e-19 $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_55 N_A1_c_53_n N_A2_c_81_n 0.0422488f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_56 N_A1_M1004_g A2 0.00709248f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A1_c_52_n A2 0.01146f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_58 N_A1_M1004_g N_VPWR_c_193_n 0.00536186f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_59 N_A1_c_52_n N_VPWR_c_193_n 0.0219687f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_60 N_A1_c_53_n N_VPWR_c_193_n 0.00135527f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_61 N_A1_M1004_g N_VPWR_c_195_n 0.00553757f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A1_M1004_g N_VPWR_c_191_n 0.0109222f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A1_M1006_g N_A_31_74#_c_270_n 0.00968761f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A1_M1006_g N_A_31_74#_c_271_n 0.0152697f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_65 N_A1_c_53_n N_A_31_74#_c_271_n 2.07531e-19 $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_66 N_A1_M1006_g N_A_31_74#_c_272_n 0.00206782f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_67 N_A1_c_52_n N_A_31_74#_c_272_n 0.0260039f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_68 N_A1_c_53_n N_A_31_74#_c_272_n 0.00265502f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_69 N_A1_M1006_g N_VGND_c_296_n 0.00539757f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A1_M1006_g N_VGND_c_297_n 0.00434272f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A1_M1006_g N_VGND_c_299_n 0.00824496f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A2_M1000_g N_B1_M1001_g 0.0143797f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A2_M1005_g N_B1_M1003_g 0.0233545f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_74 A2 B1 0.0197279f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A2_c_81_n B1 4.19259e-19 $X=1 $Y=1.465 $X2=0 $Y2=0
cc_76 A2 N_B1_c_122_n 4.1782e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A2_c_81_n N_B1_c_122_n 0.0181621f $X=1 $Y=1.465 $X2=0 $Y2=0
cc_78 N_A2_M1005_g N_VPWR_c_194_n 6.41112e-19 $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A2_M1005_g N_VPWR_c_195_n 0.00553757f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_80 A2 N_VPWR_c_195_n 0.00571228f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_81 N_A2_M1005_g N_VPWR_c_191_n 0.0109172f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_82 A2 N_VPWR_c_191_n 0.00794958f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_83 A2 A_119_368# 0.00907286f $X=0.72 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_84 N_A2_M1005_g N_Y_c_226_n 0.013124f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A2_M1005_g N_Y_c_228_n 0.002111f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_86 A2 N_Y_c_228_n 0.00338979f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A2_c_81_n N_Y_c_228_n 3.16589e-19 $X=1 $Y=1.465 $X2=0 $Y2=0
cc_88 A2 N_Y_c_228_n 0.0062742f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_89 N_A2_M1000_g N_A_31_74#_c_270_n 9.1183e-19 $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A2_M1000_g N_A_31_74#_c_271_n 0.0128142f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_91 A2 N_A_31_74#_c_271_n 0.041574f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A2_c_81_n N_A_31_74#_c_271_n 0.00127414f $X=1 $Y=1.465 $X2=0 $Y2=0
cc_93 N_A2_M1000_g N_A_31_74#_c_273_n 4.33993e-19 $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A2_M1000_g N_VGND_c_296_n 0.00956268f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A2_M1000_g N_VGND_c_298_n 0.00383152f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A2_M1000_g N_VGND_c_299_n 0.00757954f $X=1.015 $Y=0.74 $X2=0 $Y2=0
cc_97 B1 N_C1_M1002_g 0.00176701f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_B1_c_122_n N_C1_M1002_g 0.0307679f $X=1.57 $Y=1.465 $X2=0 $Y2=0
cc_99 B1 C1 0.00880658f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_100 B1 C1 0.0192202f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B1_c_122_n C1 2.81336e-19 $X=1.57 $Y=1.465 $X2=0 $Y2=0
cc_102 B1 N_C1_c_160_n 0.00153306f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_122_n N_C1_c_160_n 0.0132056f $X=1.57 $Y=1.465 $X2=0 $Y2=0
cc_104 N_B1_M1001_g N_C1_c_161_n 0.0233562f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_105 B1 N_C1_c_161_n 0.00938955f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_106 N_B1_M1003_g N_VPWR_c_194_n 0.0177256f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_107 N_B1_M1003_g N_VPWR_c_195_n 0.00460063f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_108 N_B1_M1003_g N_VPWR_c_191_n 0.009107f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_109 N_B1_M1003_g N_Y_c_226_n 0.0142201f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_110 N_B1_M1003_g N_Y_c_227_n 0.0174033f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_111 B1 N_Y_c_227_n 0.0250894f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B1_c_122_n N_Y_c_227_n 0.00263385f $X=1.57 $Y=1.465 $X2=0 $Y2=0
cc_113 B1 N_Y_c_228_n 0.00421666f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B1_c_122_n N_Y_c_228_n 0.00136199f $X=1.57 $Y=1.465 $X2=0 $Y2=0
cc_115 N_B1_M1003_g N_Y_c_229_n 9.77239e-19 $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_116 B1 N_Y_c_225_n 0.0338432f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_117 B1 N_A_31_74#_c_271_n 0.0016373f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 N_B1_M1001_g N_A_31_74#_c_273_n 8.38786e-19 $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_119 N_B1_M1001_g N_VGND_c_296_n 6.58032e-19 $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_120 N_B1_M1001_g N_VGND_c_298_n 0.00461464f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_121 B1 N_VGND_c_298_n 0.00653424f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_122 N_B1_M1001_g N_VGND_c_299_n 0.00910985f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_123 B1 N_VGND_c_299_n 0.00794958f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_124 B1 A_311_74# 0.0161056f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_125 N_C1_M1002_g N_VPWR_c_194_n 0.00398325f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_126 N_C1_M1002_g N_VPWR_c_197_n 0.005209f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_127 N_C1_M1002_g N_VPWR_c_191_n 0.00986479f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_128 N_C1_M1002_g N_Y_c_227_n 0.013639f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_129 C1 N_Y_c_227_n 0.0124525f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_130 N_C1_c_160_n N_Y_c_227_n 5.07644e-19 $X=2.14 $Y=1.385 $X2=0 $Y2=0
cc_131 N_C1_M1002_g N_Y_c_229_n 0.0148712f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_132 N_C1_M1002_g N_Y_c_224_n 0.00713608f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_133 C1 N_Y_c_224_n 0.0188818f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_134 N_C1_c_160_n N_Y_c_224_n 0.00681233f $X=2.14 $Y=1.385 $X2=0 $Y2=0
cc_135 N_C1_c_161_n N_Y_c_224_n 0.00339074f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_136 N_C1_M1002_g N_Y_c_231_n 0.00189161f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_137 C1 N_Y_c_231_n 0.00619061f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_138 N_C1_c_160_n N_Y_c_231_n 5.21084e-19 $X=2.14 $Y=1.385 $X2=0 $Y2=0
cc_139 C1 N_Y_c_225_n 0.0192616f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_140 N_C1_c_160_n N_Y_c_225_n 0.00108316f $X=2.14 $Y=1.385 $X2=0 $Y2=0
cc_141 N_C1_c_161_n N_Y_c_225_n 0.0112973f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_142 N_C1_c_161_n N_VGND_c_298_n 0.00377174f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_143 N_C1_c_161_n N_VGND_c_299_n 0.00628921f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_144 N_VPWR_c_194_n N_Y_c_226_n 0.0485389f $X=1.87 $Y=2.305 $X2=0 $Y2=0
cc_145 N_VPWR_c_195_n N_Y_c_226_n 0.0146357f $X=1.705 $Y=3.33 $X2=0 $Y2=0
cc_146 N_VPWR_c_191_n N_Y_c_226_n 0.0121141f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_M1003_d N_Y_c_227_n 0.00218982f $X=1.735 $Y=1.84 $X2=0 $Y2=0
cc_148 N_VPWR_c_194_n N_Y_c_227_n 0.0189268f $X=1.87 $Y=2.305 $X2=0 $Y2=0
cc_149 N_VPWR_c_194_n N_Y_c_229_n 0.0350101f $X=1.87 $Y=2.305 $X2=0 $Y2=0
cc_150 N_VPWR_c_197_n N_Y_c_229_n 0.0250349f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_c_191_n N_Y_c_229_n 0.0206536f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_152 N_Y_c_228_n N_A_31_74#_c_271_n 0.00821726f $X=1.455 $Y=1.885 $X2=0 $Y2=0
cc_153 N_Y_c_225_n N_VGND_c_298_n 0.0216534f $X=2.682 $Y=0.725 $X2=0 $Y2=0
cc_154 N_Y_c_225_n N_VGND_c_299_n 0.0246737f $X=2.682 $Y=0.725 $X2=0 $Y2=0
cc_155 N_A_31_74#_c_271_n N_VGND_M1006_d 0.00256964f $X=1.145 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_31_74#_c_270_n N_VGND_c_296_n 0.0169251f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_157 N_A_31_74#_c_271_n N_VGND_c_296_n 0.0201026f $X=1.145 $Y=1.045 $X2=0
+ $Y2=0
cc_158 N_A_31_74#_c_273_n N_VGND_c_296_n 0.0161397f $X=1.23 $Y=0.515 $X2=0 $Y2=0
cc_159 N_A_31_74#_c_270_n N_VGND_c_297_n 0.0145639f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_160 N_A_31_74#_c_273_n N_VGND_c_298_n 0.011066f $X=1.23 $Y=0.515 $X2=0 $Y2=0
cc_161 N_A_31_74#_c_270_n N_VGND_c_299_n 0.0119984f $X=0.3 $Y=0.515 $X2=0 $Y2=0
cc_162 N_A_31_74#_c_273_n N_VGND_c_299_n 0.00915947f $X=1.23 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o2111a_1.pxi.spice
* Created: Wed Sep  2 12:17:36 2020
* 
x_PM_SKY130_FD_SC_MS__O2111A_1%A_82_48# N_A_82_48#_M1011_s N_A_82_48#_M1008_d
+ N_A_82_48#_M1002_d N_A_82_48#_M1007_g N_A_82_48#_M1003_g N_A_82_48#_c_74_n
+ N_A_82_48#_c_75_n N_A_82_48#_c_86_p N_A_82_48#_c_129_p N_A_82_48#_c_76_n
+ N_A_82_48#_c_103_p N_A_82_48#_c_77_n N_A_82_48#_c_78_n N_A_82_48#_c_82_n
+ N_A_82_48#_c_83_n N_A_82_48#_c_79_n PM_SKY130_FD_SC_MS__O2111A_1%A_82_48#
x_PM_SKY130_FD_SC_MS__O2111A_1%D1 N_D1_M1008_g N_D1_c_154_n N_D1_M1011_g
+ N_D1_c_155_n D1 N_D1_c_157_n N_D1_c_158_n PM_SKY130_FD_SC_MS__O2111A_1%D1
x_PM_SKY130_FD_SC_MS__O2111A_1%C1 N_C1_M1005_g N_C1_M1000_g C1 C1 C1 C1
+ N_C1_c_201_n PM_SKY130_FD_SC_MS__O2111A_1%C1
x_PM_SKY130_FD_SC_MS__O2111A_1%B1 N_B1_M1001_g N_B1_M1002_g B1 N_B1_c_241_n
+ N_B1_c_242_n PM_SKY130_FD_SC_MS__O2111A_1%B1
x_PM_SKY130_FD_SC_MS__O2111A_1%A2 N_A2_M1004_g N_A2_M1010_g A2 N_A2_c_276_n
+ PM_SKY130_FD_SC_MS__O2111A_1%A2
x_PM_SKY130_FD_SC_MS__O2111A_1%A1 N_A1_M1009_g N_A1_M1006_g A1 N_A1_c_309_n
+ N_A1_c_310_n PM_SKY130_FD_SC_MS__O2111A_1%A1
x_PM_SKY130_FD_SC_MS__O2111A_1%X N_X_M1007_s N_X_M1003_s N_X_c_333_n N_X_c_334_n
+ X X X X N_X_c_335_n PM_SKY130_FD_SC_MS__O2111A_1%X
x_PM_SKY130_FD_SC_MS__O2111A_1%VPWR N_VPWR_M1003_d N_VPWR_M1005_d N_VPWR_M1006_d
+ N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n VPWR
+ N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n
+ N_VPWR_c_356_n PM_SKY130_FD_SC_MS__O2111A_1%VPWR
x_PM_SKY130_FD_SC_MS__O2111A_1%VGND N_VGND_M1007_d N_VGND_M1004_d N_VGND_c_405_n
+ N_VGND_c_406_n VGND N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n PM_SKY130_FD_SC_MS__O2111A_1%VGND
x_PM_SKY130_FD_SC_MS__O2111A_1%A_471_74# N_A_471_74#_M1001_d N_A_471_74#_M1009_d
+ N_A_471_74#_c_449_n N_A_471_74#_c_450_n N_A_471_74#_c_451_n
+ N_A_471_74#_c_452_n PM_SKY130_FD_SC_MS__O2111A_1%A_471_74#
cc_1 VNB N_A_82_48#_M1003_g 0.00705046f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_82_48#_c_74_n 0.00153124f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.07
cc_3 VNB N_A_82_48#_c_75_n 0.0174507f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.295
cc_4 VNB N_A_82_48#_c_76_n 0.0112873f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.515
cc_5 VNB N_A_82_48#_c_77_n 0.00538141f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_6 VNB N_A_82_48#_c_78_n 0.0371751f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_7 VNB N_A_82_48#_c_79_n 0.0234345f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.22
cc_8 VNB N_D1_c_154_n 0.0165545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D1_c_155_n 0.0324276f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_10 VNB D1 0.00165832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_11 VNB N_D1_c_157_n 0.0135906f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.55
cc_12 VNB N_D1_c_158_n 0.0135632f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.295
cc_13 VNB N_C1_M1000_g 0.0335784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB C1 0.0022543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C1_c_201_n 0.0136808f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.155
cc_16 VNB N_B1_M1001_g 0.0291183f $X=-0.19 $Y=-0.245 $X2=2.48 $Y2=2.065
cc_17 VNB N_B1_c_241_n 0.0199345f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_18 VNB N_B1_c_242_n 0.00796532f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_19 VNB N_A2_M1004_g 0.0311844f $X=-0.19 $Y=-0.245 $X2=2.48 $Y2=2.065
cc_20 VNB A2 0.00520679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_276_n 0.0185676f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_22 VNB N_A1_M1009_g 0.0314484f $X=-0.19 $Y=-0.245 $X2=2.48 $Y2=2.065
cc_23 VNB N_A1_M1006_g 0.00185508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_309_n 0.0585543f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_25 VNB N_A1_c_310_n 0.00488709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_333_n 0.0235276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_334_n 0.00489291f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_28 VNB N_X_c_335_n 0.0284024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_356_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_405_n 0.0135318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_406_n 0.00975957f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_32 VNB N_VGND_c_407_n 0.0169946f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.55
cc_33 VNB N_VGND_c_408_n 0.0574108f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.155
cc_34 VNB N_VGND_c_409_n 0.0196288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_410_n 0.249202f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.295
cc_36 VNB N_VGND_c_411_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_37 VNB N_VGND_c_412_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.157
cc_38 VNB N_A_471_74#_c_449_n 0.00335011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_471_74#_c_450_n 0.0131391f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_40 VNB N_A_471_74#_c_451_n 0.0095993f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_41 VNB N_A_471_74#_c_452_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_42 VPB N_A_82_48#_M1003_g 0.0291513f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_43 VPB N_A_82_48#_c_74_n 0.00314065f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.07
cc_44 VPB N_A_82_48#_c_82_n 0.00301947f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=2.24
cc_45 VPB N_A_82_48#_c_83_n 0.00402851f $X=-0.19 $Y=1.66 $X2=2.7 $Y2=2.21
cc_46 VPB N_D1_M1008_g 0.0248898f $X=-0.19 $Y=1.66 $X2=2.48 $Y2=2.065
cc_47 VPB D1 0.00142441f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_48 VPB N_D1_c_157_n 0.020819f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.55
cc_49 VPB N_C1_M1005_g 0.0247775f $X=-0.19 $Y=1.66 $X2=2.48 $Y2=2.065
cc_50 VPB C1 0.00139918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_C1_c_201_n 0.026223f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.155
cc_52 VPB N_B1_M1002_g 0.0344197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_B1_c_241_n 0.00899022f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_54 VPB N_B1_c_242_n 0.00470511f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.55
cc_55 VPB N_A2_M1010_g 0.0212788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB A2 0.01111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A2_c_276_n 0.00898898f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_58 VPB N_A1_M1006_g 0.0316355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A1_c_310_n 0.0072578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB X 0.0128625f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_61 VPB X 0.0411673f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.21
cc_62 VPB N_X_c_335_n 0.00749244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_357_n 0.0112316f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_64 VPB N_VPWR_c_358_n 0.0174828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_359_n 0.0118719f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=2.07
cc_66 VPB N_VPWR_c_360_n 0.0511896f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.295
cc_67 VPB N_VPWR_c_361_n 0.0189953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_362_n 0.0229347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_363_n 0.0331177f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_70 VPB N_VPWR_c_364_n 0.00632158f $X=-0.19 $Y=1.66 $X2=2.7 $Y2=2.21
cc_71 VPB N_VPWR_c_365_n 0.0105532f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.55
cc_72 VPB N_VPWR_c_356_n 0.08535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 N_A_82_48#_M1003_g N_D1_M1008_g 0.0158764f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_74 N_A_82_48#_c_74_n N_D1_M1008_g 0.00381516f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_75 N_A_82_48#_c_86_p N_D1_M1008_g 0.013707f $X=1.195 $Y=2.155 $X2=0 $Y2=0
cc_76 N_A_82_48#_c_82_n N_D1_M1008_g 0.0135158f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_77 N_A_82_48#_c_76_n N_D1_c_154_n 0.0190115f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_78 N_A_82_48#_c_75_n N_D1_c_155_n 0.005455f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_79 N_A_82_48#_c_76_n N_D1_c_155_n 0.00458903f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_80 N_A_82_48#_c_78_n N_D1_c_155_n 0.00826486f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_81 N_A_82_48#_c_79_n N_D1_c_155_n 4.52431e-19 $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_82 N_A_82_48#_c_74_n D1 0.0203563f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_83 N_A_82_48#_c_75_n D1 0.0260844f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_84 N_A_82_48#_c_86_p D1 0.0111593f $X=1.195 $Y=2.155 $X2=0 $Y2=0
cc_85 N_A_82_48#_c_82_n D1 0.00809383f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_86 N_A_82_48#_M1003_g N_D1_c_157_n 0.00725163f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_82_48#_c_74_n N_D1_c_157_n 0.00250307f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_88 N_A_82_48#_c_75_n N_D1_c_157_n 0.00133731f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_89 N_A_82_48#_c_82_n N_D1_c_157_n 6.57128e-19 $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_90 N_A_82_48#_c_75_n N_D1_c_158_n 0.00357242f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_91 N_A_82_48#_c_77_n N_D1_c_158_n 0.00325742f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_92 N_A_82_48#_c_103_p N_C1_M1005_g 0.0165888f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_93 N_A_82_48#_c_82_n N_C1_M1005_g 8.7706e-19 $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_94 N_A_82_48#_c_75_n C1 0.0111966f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_95 N_A_82_48#_c_76_n C1 0.0488331f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_96 N_A_82_48#_c_103_p C1 0.0233095f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_97 N_A_82_48#_c_103_p N_C1_c_201_n 0.00470945f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_98 N_A_82_48#_c_103_p N_B1_M1002_g 0.0199368f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_99 N_A_82_48#_c_83_n N_B1_M1002_g 0.00432128f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_100 N_A_82_48#_c_103_p N_B1_c_241_n 5.76756e-19 $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_101 N_A_82_48#_c_103_p N_B1_c_242_n 0.0215212f $X=2.535 $Y=2.157 $X2=0 $Y2=0
cc_102 N_A_82_48#_c_83_n N_A2_M1010_g 0.0193168f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_103 N_A_82_48#_c_83_n A2 0.00743045f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_104 N_A_82_48#_c_83_n N_A2_c_276_n 6.25105e-19 $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_105 N_A_82_48#_c_83_n N_A1_M1006_g 0.00249225f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_106 N_A_82_48#_c_79_n N_X_c_333_n 4.44442e-19 $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A_82_48#_M1003_g X 0.0036289f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_82_48#_c_74_n X 0.0101424f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_109 N_A_82_48#_c_77_n X 4.42944e-19 $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_110 N_A_82_48#_c_78_n X 2.17346e-19 $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_82_48#_M1003_g X 0.0147265f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_82_48#_M1003_g N_X_c_335_n 0.00601455f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_82_48#_c_74_n N_X_c_335_n 0.0122487f $X=0.7 $Y=2.07 $X2=0 $Y2=0
cc_114 N_A_82_48#_c_77_n N_X_c_335_n 0.02563f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_115 N_A_82_48#_c_79_n N_X_c_335_n 0.013355f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_116 N_A_82_48#_c_74_n N_VPWR_M1003_d 0.00434847f $X=0.7 $Y=2.07 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_82_48#_c_86_p N_VPWR_M1003_d 0.0118004f $X=1.195 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_82_48#_c_129_p N_VPWR_M1003_d 0.00271221f $X=0.785 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_82_48#_c_103_p N_VPWR_M1005_d 0.0147749f $X=2.535 $Y=2.157 $X2=0
+ $Y2=0
cc_120 N_A_82_48#_M1003_g N_VPWR_c_357_n 0.00431748f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_82_48#_c_86_p N_VPWR_c_357_n 0.0128995f $X=1.195 $Y=2.155 $X2=0 $Y2=0
cc_122 N_A_82_48#_c_129_p N_VPWR_c_357_n 0.0119464f $X=0.785 $Y=2.155 $X2=0
+ $Y2=0
cc_123 N_A_82_48#_c_82_n N_VPWR_c_357_n 0.0297393f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_124 N_A_82_48#_c_103_p N_VPWR_c_358_n 0.0321113f $X=2.535 $Y=2.157 $X2=0
+ $Y2=0
cc_125 N_A_82_48#_c_82_n N_VPWR_c_358_n 0.00139434f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_126 N_A_82_48#_c_83_n N_VPWR_c_358_n 0.00127335f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_127 N_A_82_48#_c_83_n N_VPWR_c_360_n 0.0258836f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_128 N_A_82_48#_M1003_g N_VPWR_c_361_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_82_48#_c_82_n N_VPWR_c_362_n 0.0118983f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_130 N_A_82_48#_c_83_n N_VPWR_c_363_n 0.0118983f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_131 N_A_82_48#_M1003_g N_VPWR_c_356_n 0.00990469f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_82_48#_c_82_n N_VPWR_c_356_n 0.0116774f $X=1.36 $Y=2.24 $X2=0 $Y2=0
cc_133 N_A_82_48#_c_83_n N_VPWR_c_356_n 0.0116774f $X=2.7 $Y=2.21 $X2=0 $Y2=0
cc_134 N_A_82_48#_c_75_n N_VGND_c_405_n 0.00658384f $X=1.08 $Y=1.295 $X2=0 $Y2=0
cc_135 N_A_82_48#_c_76_n N_VGND_c_405_n 0.0477412f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_136 N_A_82_48#_c_77_n N_VGND_c_405_n 0.019655f $X=0.61 $Y=1.295 $X2=0 $Y2=0
cc_137 N_A_82_48#_c_78_n N_VGND_c_405_n 0.00140455f $X=0.6 $Y=1.385 $X2=0 $Y2=0
cc_138 N_A_82_48#_c_79_n N_VGND_c_405_n 0.0156276f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_139 N_A_82_48#_c_79_n N_VGND_c_407_n 0.00383152f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A_82_48#_c_76_n N_VGND_c_408_n 0.011066f $X=1.245 $Y=0.515 $X2=0 $Y2=0
cc_141 N_A_82_48#_c_76_n N_VGND_c_410_n 0.00915947f $X=1.245 $Y=0.515 $X2=0
+ $Y2=0
cc_142 N_A_82_48#_c_79_n N_VGND_c_410_n 0.00761163f $X=0.587 $Y=1.22 $X2=0 $Y2=0
cc_143 N_D1_c_154_n N_C1_M1000_g 0.0705403f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_144 N_D1_c_158_n N_C1_M1000_g 0.0043485f $X=1.17 $Y=1.55 $X2=0 $Y2=0
cc_145 N_D1_c_154_n C1 0.0181159f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_146 N_D1_c_155_n C1 0.00518893f $X=1.53 $Y=1.26 $X2=0 $Y2=0
cc_147 D1 C1 0.0209972f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_148 N_D1_c_157_n C1 0.0010797f $X=1.17 $Y=1.715 $X2=0 $Y2=0
cc_149 N_D1_c_158_n C1 0.00464587f $X=1.17 $Y=1.55 $X2=0 $Y2=0
cc_150 N_D1_M1008_g N_C1_c_201_n 0.0176293f $X=1.135 $Y=2.485 $X2=0 $Y2=0
cc_151 N_D1_c_155_n N_C1_c_201_n 0.00343303f $X=1.53 $Y=1.26 $X2=0 $Y2=0
cc_152 D1 N_C1_c_201_n 0.00112962f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_153 N_D1_c_157_n N_C1_c_201_n 0.0192424f $X=1.17 $Y=1.715 $X2=0 $Y2=0
cc_154 N_D1_M1008_g X 9.5413e-19 $X=1.135 $Y=2.485 $X2=0 $Y2=0
cc_155 N_D1_M1008_g N_VPWR_c_357_n 0.00830324f $X=1.135 $Y=2.485 $X2=0 $Y2=0
cc_156 N_D1_M1008_g N_VPWR_c_362_n 0.00616627f $X=1.135 $Y=2.485 $X2=0 $Y2=0
cc_157 N_D1_M1008_g N_VPWR_c_356_n 0.00634024f $X=1.135 $Y=2.485 $X2=0 $Y2=0
cc_158 N_D1_c_154_n N_VGND_c_405_n 0.00361162f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_159 N_D1_c_154_n N_VGND_c_408_n 0.0039925f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_160 N_D1_c_154_n N_VGND_c_410_n 0.00702246f $X=1.53 $Y=1.185 $X2=0 $Y2=0
cc_161 N_C1_M1000_g N_B1_M1001_g 0.0599213f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_162 C1 N_B1_M1001_g 0.00363173f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_163 N_C1_M1005_g N_B1_M1002_g 0.019596f $X=1.635 $Y=2.485 $X2=0 $Y2=0
cc_164 C1 N_B1_M1002_g 6.51483e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_165 N_C1_c_201_n N_B1_M1002_g 0.00617601f $X=1.89 $Y=1.735 $X2=0 $Y2=0
cc_166 N_C1_M1000_g N_B1_c_241_n 0.0200714f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_167 C1 N_B1_c_241_n 2.77362e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_168 N_C1_M1000_g N_B1_c_242_n 0.0025595f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_169 C1 N_B1_c_242_n 0.0296056f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_170 N_C1_M1005_g N_VPWR_c_358_n 0.00805335f $X=1.635 $Y=2.485 $X2=0 $Y2=0
cc_171 N_C1_M1005_g N_VPWR_c_362_n 0.00645549f $X=1.635 $Y=2.485 $X2=0 $Y2=0
cc_172 N_C1_M1005_g N_VPWR_c_356_n 0.00634024f $X=1.635 $Y=2.485 $X2=0 $Y2=0
cc_173 N_C1_M1000_g N_VGND_c_408_n 0.0039925f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_174 C1 N_VGND_c_408_n 0.00851294f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_175 N_C1_M1000_g N_VGND_c_410_n 0.00696958f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_176 C1 N_VGND_c_410_n 0.0108483f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_177 C1 A_321_74# 0.00133334f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_178 C1 N_A_471_74#_c_451_n 0.0030385f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_179 N_B1_M1001_g N_A2_M1004_g 0.0179083f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_M1002_g N_A2_M1010_g 0.0305507f $X=2.39 $Y=2.485 $X2=0 $Y2=0
cc_181 N_B1_c_241_n A2 4.13845e-19 $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_182 N_B1_c_242_n A2 0.0249368f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_183 N_B1_c_241_n N_A2_c_276_n 0.0214219f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B1_c_242_n N_A2_c_276_n 4.14478e-19 $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_185 N_B1_M1002_g N_VPWR_c_358_n 0.00813216f $X=2.39 $Y=2.485 $X2=0 $Y2=0
cc_186 N_B1_M1002_g N_VPWR_c_363_n 0.00645549f $X=2.39 $Y=2.485 $X2=0 $Y2=0
cc_187 N_B1_M1002_g N_VPWR_c_356_n 0.00634024f $X=2.39 $Y=2.485 $X2=0 $Y2=0
cc_188 N_B1_M1001_g N_VGND_c_408_n 0.00461464f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B1_M1001_g N_VGND_c_410_n 0.00909821f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B1_M1001_g N_A_471_74#_c_449_n 8.94767e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B1_M1001_g N_A_471_74#_c_451_n 3.11521e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_192 N_B1_c_241_n N_A_471_74#_c_451_n 0.00307668f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B1_c_242_n N_A_471_74#_c_451_n 0.00722443f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A2_M1004_g N_A1_M1009_g 0.0277451f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A2_M1010_g N_A1_M1006_g 0.067526f $X=2.925 $Y=2.405 $X2=0 $Y2=0
cc_196 A2 N_A1_c_309_n 0.00293932f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A2_c_276_n N_A1_c_309_n 0.0204011f $X=2.88 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A2_M1004_g N_A1_c_310_n 5.08722e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_199 A2 N_A1_c_310_n 0.0299012f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A2_c_276_n N_A1_c_310_n 2.31792e-19 $X=2.88 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A2_M1010_g N_VPWR_c_360_n 0.00347972f $X=2.925 $Y=2.405 $X2=0 $Y2=0
cc_202 N_A2_M1010_g N_VPWR_c_363_n 0.00616627f $X=2.925 $Y=2.405 $X2=0 $Y2=0
cc_203 N_A2_M1010_g N_VPWR_c_356_n 0.00634024f $X=2.925 $Y=2.405 $X2=0 $Y2=0
cc_204 N_A2_M1004_g N_VGND_c_406_n 0.0036453f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A2_M1004_g N_VGND_c_408_n 0.00461464f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A2_M1004_g N_VGND_c_410_n 0.00909258f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A2_M1004_g N_A_471_74#_c_449_n 5.32432e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A2_M1004_g N_A_471_74#_c_450_n 0.0144173f $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_209 A2 N_A_471_74#_c_450_n 0.0270243f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A2_c_276_n N_A_471_74#_c_450_n 0.00424874f $X=2.88 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A2_M1004_g N_A_471_74#_c_452_n 6.2684e-19 $X=2.79 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A1_M1006_g N_VPWR_c_360_n 0.0237438f $X=3.345 $Y=2.405 $X2=0 $Y2=0
cc_213 N_A1_c_309_n N_VPWR_c_360_n 0.00152096f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_214 N_A1_c_310_n N_VPWR_c_360_n 0.0266029f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_215 N_A1_M1006_g N_VPWR_c_363_n 0.00536686f $X=3.345 $Y=2.405 $X2=0 $Y2=0
cc_216 N_A1_M1006_g N_VPWR_c_356_n 0.00531876f $X=3.345 $Y=2.405 $X2=0 $Y2=0
cc_217 N_A1_M1009_g N_VGND_c_406_n 0.00572341f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1009_g N_VGND_c_409_n 0.00434272f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_M1009_g N_VGND_c_410_n 0.00824797f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_M1009_g N_A_471_74#_c_450_n 0.017525f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_c_309_n N_A_471_74#_c_450_n 0.00240334f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_222 N_A1_c_310_n N_A_471_74#_c_450_n 0.0264387f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_223 N_A1_M1009_g N_A_471_74#_c_452_n 0.00977408f $X=3.33 $Y=0.74 $X2=0 $Y2=0
cc_224 X N_VPWR_c_357_n 0.0223717f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_225 X N_VPWR_c_361_n 0.0154414f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_226 X N_VPWR_c_356_n 0.0127129f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_227 N_X_c_333_n N_VGND_c_405_n 0.0254628f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_228 N_X_c_333_n N_VGND_c_407_n 0.0115164f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_229 N_X_c_333_n N_VGND_c_410_n 0.00953044f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_230 N_VGND_c_406_n N_A_471_74#_c_449_n 0.00158095f $X=3.045 $Y=0.57 $X2=0
+ $Y2=0
cc_231 N_VGND_c_408_n N_A_471_74#_c_449_n 0.0146357f $X=2.88 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_410_n N_A_471_74#_c_449_n 0.0121141f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_M1004_d N_A_471_74#_c_450_n 0.00318135f $X=2.865 $Y=0.37 $X2=0
+ $Y2=0
cc_234 N_VGND_c_406_n N_A_471_74#_c_450_n 0.022455f $X=3.045 $Y=0.57 $X2=0 $Y2=0
cc_235 N_VGND_c_406_n N_A_471_74#_c_452_n 0.0173003f $X=3.045 $Y=0.57 $X2=0
+ $Y2=0
cc_236 N_VGND_c_409_n N_A_471_74#_c_452_n 0.0145639f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_410_n N_A_471_74#_c_452_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o21bai_2.pex.spice
* Created: Fri Aug 28 17:56:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21BAI_2%B1_N 3 7 9 15 16
r33 14 16 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.625 $Y=1.515
+ $X2=0.7 $Y2=1.515
r34 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.515 $X2=0.625 $Y2=1.515
r35 11 14 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.625 $Y2=1.515
r36 9 15 4.60977 $w=3.73e-07 $l=1.5e-07 $layer=LI1_cond $X=0.647 $Y=1.665
+ $X2=0.647 $Y2=1.515
r37 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.7 $Y=1.68 $X2=0.7
+ $Y2=1.515
r38 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.7 $Y=1.68 $X2=0.7
+ $Y2=2.34
r39 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r40 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%A_27_74# 1 2 9 11 13 16 18 20 21 24 28 34
+ 36 40 43 45 46
c86 16 0 1.41978e-19 $X=1.92 $Y=2.4
r87 45 46 7.85017 $w=5.23e-07 $l=8.5e-08 $layer=LI1_cond $X=0.377 $Y=2.035
+ $X2=0.377 $Y2=1.95
r88 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.385 $X2=1.195 $Y2=1.385
r89 38 40 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.195 $Y=1.18
+ $X2=1.195 $Y2=1.385
r90 37 43 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.095
+ $X2=0.24 $Y2=1.095
r91 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.03 $Y=1.095
+ $X2=1.195 $Y2=1.18
r92 36 37 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.03 $Y=1.095
+ $X2=0.365 $Y2=1.095
r93 32 45 4.03249 $w=5.23e-07 $l=1.77e-07 $layer=LI1_cond $X=0.377 $Y=2.212
+ $X2=0.377 $Y2=2.035
r94 32 34 11.4596 $w=5.23e-07 $l=5.03e-07 $layer=LI1_cond $X=0.377 $Y=2.212
+ $X2=0.377 $Y2=2.715
r95 30 43 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=1.18
+ $X2=0.24 $Y2=1.095
r96 30 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.2 $Y=1.18 $X2=0.2
+ $Y2=1.95
r97 26 43 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.01 $X2=0.24
+ $Y2=1.095
r98 26 28 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r99 23 24 67.5114 $w=3.07e-07 $l=4.3e-07 $layer=POLY_cond $X=1.485 $Y=1.385
+ $X2=1.915 $Y2=1.385
r100 22 23 2.35505 $w=3.07e-07 $l=1.5e-08 $layer=POLY_cond $X=1.47 $Y=1.385
+ $X2=1.485 $Y2=1.385
r101 21 41 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.38 $Y=1.385
+ $X2=1.195 $Y2=1.385
r102 21 22 13.4516 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.38 $Y=1.385
+ $X2=1.47 $Y2=1.385
r103 18 24 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.22
+ $X2=1.915 $Y2=1.385
r104 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.915 $Y=1.22
+ $X2=1.915 $Y2=0.74
r105 14 24 0.785016 $w=3.07e-07 $l=5e-09 $layer=POLY_cond $X=1.92 $Y=1.385
+ $X2=1.915 $Y2=1.385
r106 14 16 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=1.92 $Y=1.525
+ $X2=1.92 $Y2=2.4
r107 11 23 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.485 $Y2=1.385
r108 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.485 $Y2=0.74
r109 7 22 15.2536 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=1.55
+ $X2=1.47 $Y2=1.385
r110 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.47 $Y=1.55 $X2=1.47
+ $Y2=2.4
r111 2 45 400 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=1.84 $X2=0.475 $Y2=2.035
r112 2 34 400 $w=1.7e-07 $l=9.49342e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=1.84 $X2=0.475 $Y2=2.715
r113 1 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%A1 3 7 11 15 19 20 22 23 25 31 32 37
c85 7 0 1.89662e-19 $X=2.46 $Y=2.4
c86 3 0 1.9405e-19 $X=2.415 $Y=0.74
r87 35 37 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.6 $Y=1.65 $X2=3.6
+ $Y2=1.665
r88 31 34 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.89 $Y=1.485
+ $X2=3.89 $Y2=1.65
r89 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.89 $Y=1.485
+ $X2=3.89 $Y2=1.32
r90 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.485 $X2=3.89 $Y2=1.485
r91 25 32 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.6 $Y=1.485
+ $X2=3.89 $Y2=1.485
r92 25 35 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.485 $X2=3.6
+ $Y2=1.65
r93 25 37 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=3.6 $Y=1.7 $X2=3.6
+ $Y2=1.665
r94 24 25 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.6 $Y=1.95 $X2=3.6
+ $Y2=1.7
r95 22 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.6 $Y2=1.95
r96 22 23 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=2.58 $Y2=2.035
r97 20 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.515
+ $X2=2.415 $Y2=1.68
r98 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.515 $X2=2.415 $Y2=1.515
r99 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=1.95
+ $X2=2.58 $Y2=2.035
r100 17 19 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.415 $Y=1.95
+ $X2=2.415 $Y2=1.515
r101 15 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.805 $Y=0.74
+ $X2=3.805 $Y2=1.32
r102 11 34 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.815 $Y=2.4
+ $X2=3.815 $Y2=1.65
r103 7 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.46 $Y=2.4 $X2=2.46
+ $Y2=1.68
r104 1 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.515
r105 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%A2 3 7 11 15 17 24 26
c55 24 0 1.21621e-19 $X=3.03 $Y=1.515
r56 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.36 $Y=1.515
+ $X2=3.375 $Y2=1.515
r57 23 25 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.03 $Y=1.515
+ $X2=3.36 $Y2=1.515
r58 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.515 $X2=3.03 $Y2=1.515
r59 21 23 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=2.945 $Y=1.515
+ $X2=3.03 $Y2=1.515
r60 19 21 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.91 $Y=1.515
+ $X2=2.945 $Y2=1.515
r61 17 24 4.16546 $w=4.13e-07 $l=1.5e-07 $layer=LI1_cond $X=3.027 $Y=1.665
+ $X2=3.027 $Y2=1.515
r62 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.35
+ $X2=3.375 $Y2=1.515
r63 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.375 $Y=1.35
+ $X2=3.375 $Y2=0.74
r64 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=1.68
+ $X2=3.36 $Y2=1.515
r65 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.36 $Y=1.68 $X2=3.36
+ $Y2=2.4
r66 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=1.35
+ $X2=2.945 $Y2=1.515
r67 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.945 $Y=1.35
+ $X2=2.945 $Y2=0.74
r68 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.68
+ $X2=2.91 $Y2=1.515
r69 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.91 $Y=1.68 $X2=2.91
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%VPWR 1 2 3 12 18 20 22 26 28 33 38 47 50 54
r56 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 39 50 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.165 $Y2=3.33
r64 39 41 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 38 53 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.137 $Y2=3.33
r66 38 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r70 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 33 50 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.98 $Y=3.33
+ $X2=2.165 $Y2=3.33
r72 33 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r73 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r74 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 28 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r76 28 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 26 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 22 25 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.08 $Y=1.985
+ $X2=4.08 $Y2=2.815
r81 20 53 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.137 $Y2=3.33
r82 20 25 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=2.815
r83 16 50 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=3.33
r84 16 18 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=2.815
r85 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.17 $Y=1.985
+ $X2=1.17 $Y2=2.815
r86 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r87 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.815
r88 3 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=2.815
r89 3 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=1.985
r90 2 18 600 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.84 $X2=2.165 $Y2=2.815
r91 1 15 400 $w=1.7e-07 $l=1.1494e-06 $layer=licon1_PDIFF $count=1 $X=0.79
+ $Y=1.84 $X2=1.17 $Y2=2.815
r92 1 12 400 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=1 $X=0.79
+ $Y=1.84 $X2=1.17 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%Y 1 2 3 12 16 18 20 24 25 26 27 42
c43 16 0 1.9405e-19 $X=1.7 $Y=0.8
r44 32 42 1.78887 $w=3.33e-07 $l=5.2e-08 $layer=LI1_cond $X=1.697 $Y=1.347
+ $X2=1.697 $Y2=1.295
r45 26 27 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=1.697 $Y=1.665
+ $X2=1.697 $Y2=1.985
r46 25 42 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=1.697 $Y=1.278
+ $X2=1.697 $Y2=1.295
r47 25 40 4.13832 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=1.697 $Y=1.278
+ $X2=1.697 $Y2=1.18
r48 25 26 10.3892 $w=3.33e-07 $l=3.02e-07 $layer=LI1_cond $X=1.697 $Y=1.363
+ $X2=1.697 $Y2=1.665
r49 25 32 0.550421 $w=3.33e-07 $l=1.6e-08 $layer=LI1_cond $X=1.697 $Y=1.363
+ $X2=1.697 $Y2=1.347
r50 23 27 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=1.697 $Y=2.29
+ $X2=1.697 $Y2=1.985
r51 23 24 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=1.697 $Y=2.29
+ $X2=1.697 $Y2=2.375
r52 20 22 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=3.135 $Y=2.46 $X2=3.135
+ $Y2=2.51
r53 19 24 3.35233 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.865 $Y=2.375
+ $X2=1.697 $Y2=2.375
r54 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.05 $Y=2.375
+ $X2=3.135 $Y2=2.46
r55 18 19 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=3.05 $Y=2.375
+ $X2=1.865 $Y2=2.375
r56 16 40 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=1.74 $Y=0.8 $X2=1.74
+ $Y2=1.18
r57 10 24 3.22182 $w=2.92e-07 $l=1.03899e-07 $layer=LI1_cond $X=1.655 $Y=2.46
+ $X2=1.697 $Y2=2.375
r58 10 12 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=1.655 $Y=2.46
+ $X2=1.655 $Y2=2.815
r59 3 22 600 $w=1.7e-07 $l=7.34405e-07 $layer=licon1_PDIFF $count=1 $X=3 $Y=1.84
+ $X2=3.135 $Y2=2.51
r60 2 27 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.56
+ $Y=1.84 $X2=1.695 $Y2=1.985
r61 2 12 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.84 $X2=1.695 $Y2=2.815
r62 1 16 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%A_510_368# 1 2 7 11 14
c27 14 0 1.41978e-19 $X=2.685 $Y=2.805
c28 7 0 6.80408e-20 $X=3.42 $Y=2.99
r29 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.685 $Y=2.805
+ $X2=2.685 $Y2=2.99
r30 9 11 18.2327 $w=3.33e-07 $l=5.3e-07 $layer=LI1_cond $X=3.587 $Y=2.905
+ $X2=3.587 $Y2=2.375
r31 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=2.99
+ $X2=2.685 $Y2=2.99
r32 7 9 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=3.42 $Y=2.99
+ $X2=3.587 $Y2=2.905
r33 7 8 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.42 $Y=2.99 $X2=2.85
+ $Y2=2.99
r34 2 11 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.45
+ $Y=1.84 $X2=3.585 $Y2=2.375
r35 1 14 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.84 $X2=2.685 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48 51
+ 54
r54 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r58 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r59 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.59
+ $Y2=0
r60 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=4.08
+ $Y2=0
r61 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r62 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r63 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.7
+ $Y2=0
r65 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.12
+ $Y2=0
r66 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.59
+ $Y2=0
r67 37 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.12
+ $Y2=0
r68 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r69 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r70 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r71 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r72 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r73 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.7
+ $Y2=0
r74 29 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.16
+ $Y2=0
r75 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r76 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r78 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r79 22 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r80 22 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r81 22 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r82 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0
r83 18 20 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0.645
r84 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0
r85 14 16 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0.675
r86 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r87 10 12 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.675
r88 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.37 $X2=3.59 $Y2=0.645
r89 2 16 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.37 $X2=2.7 $Y2=0.675
r90 1 12 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__O21BAI_2%A_225_74# 1 2 3 4 15 17 18 22 23 24 27 29
+ 33 35
r64 31 33 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.06 $Y=0.98
+ $X2=4.06 $Y2=0.515
r65 30 35 5.16603 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.245 $Y=1.065
+ $X2=3.16 $Y2=1.08
r66 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.935 $Y=1.065
+ $X2=4.06 $Y2=0.98
r67 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.935 $Y=1.065
+ $X2=3.245 $Y2=1.065
r68 25 35 1.34256 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.16 $Y=0.98 $X2=3.16
+ $Y2=1.08
r69 25 27 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.16 $Y=0.98
+ $X2=3.16 $Y2=0.515
r70 23 35 5.16603 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.075 $Y=1.095
+ $X2=3.16 $Y2=1.08
r71 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.075 $Y=1.095
+ $X2=2.365 $Y2=1.095
r72 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.2 $Y=1.01
+ $X2=2.365 $Y2=1.095
r73 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.2 $Y=1.01 $X2=2.2
+ $Y2=0.515
r74 19 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.2 $Y=0.425 $X2=2.2
+ $Y2=0.515
r75 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=2.2 $Y2=0.425
r76 17 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=1.435 $Y2=0.34
r77 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.27 $Y=0.425
+ $X2=1.435 $Y2=0.34
r78 13 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.27 $Y=0.425
+ $X2=1.27 $Y2=0.675
r79 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
r80 3 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.02
+ $Y=0.37 $X2=3.16 $Y2=0.515
r81 2 22 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.2 $Y2=0.515
r82 1 15 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.675
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 X a_162_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_586_94# A2_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VGND a_162_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_162_48# B2 a_1009_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_820_392# a_586_94# a_162_48# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VPWR A1_N a_586_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_1009_74# B2 a_162_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 X a_162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR B2 a_820_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VPWR a_162_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 VGND a_586_94# a_162_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_1009_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 VPWR B1 a_820_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 VPWR a_162_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 VGND B1 a_1009_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_162_48# a_586_94# a_820_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 a_820_392# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X17 VGND A1_N a_586_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 X a_162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_820_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X20 X a_162_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_586_368# A2_N a_586_94# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 VGND a_162_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__ebufn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__ebufn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.500000 1.795000 1.830000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.435300 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.500000 0.835000 1.830000 ;
        RECT 0.665000 1.830000 0.835000 2.420000 ;
        RECT 0.665000 2.420000 2.195000 2.590000 ;
        RECT 1.865000 2.340000 2.195000 2.420000 ;
        RECT 1.865000 2.590000 2.195000 3.010000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.350000 3.755000 1.130000 ;
        RECT 3.235000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.085000  0.455000 0.530000 1.150000 ;
      RECT 0.085000  1.150000 2.200000 1.320000 ;
      RECT 0.085000  1.320000 0.255000 2.000000 ;
      RECT 0.085000  2.000000 0.445000 2.880000 ;
      RECT 0.650000  2.760000 0.980000 3.245000 ;
      RECT 0.700000  0.085000 0.985000 0.850000 ;
      RECT 1.155000  0.455000 1.450000 0.810000 ;
      RECT 1.155000  0.810000 2.660000 0.980000 ;
      RECT 1.185000  2.000000 2.135000 2.170000 ;
      RECT 1.185000  2.170000 1.695000 2.250000 ;
      RECT 1.870000  1.320000 2.200000 1.340000 ;
      RECT 1.965000  1.710000 3.065000 1.880000 ;
      RECT 1.965000  1.880000 2.135000 2.000000 ;
      RECT 2.365000  2.050000 2.695000 3.245000 ;
      RECT 2.390000  0.085000 2.720000 0.640000 ;
      RECT 2.460000  0.980000 2.660000 1.320000 ;
      RECT 2.460000  1.320000 3.415000 1.650000 ;
      RECT 2.460000  1.650000 3.065000 1.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_ms__ebufn_1
END LIBRARY

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a21boi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.430000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.430000 3.715000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.490000 7.555000 1.820000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.500800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.700000 0.770000 1.810000 0.940000 ;
        RECT 0.700000 0.940000 0.950000 1.130000 ;
        RECT 1.480000 0.940000 1.810000 1.090000 ;
        RECT 1.480000 1.090000 5.720000 1.150000 ;
        RECT 1.480000 1.150000 4.745000 1.260000 ;
        RECT 3.965000 1.260000 4.745000 1.780000 ;
        RECT 4.165000 1.780000 4.745000 1.820000 ;
        RECT 4.165000 1.820000 5.395000 1.990000 ;
        RECT 4.165000 1.990000 4.495000 2.735000 ;
        RECT 4.575000 0.980000 5.720000 1.090000 ;
        RECT 4.610000 0.350000 4.860000 0.980000 ;
        RECT 5.065000 1.990000 5.395000 2.735000 ;
        RECT 5.470000 0.350000 5.720000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  1.950000 3.995000 2.120000 ;
      RECT 0.115000  2.120000 0.365000 2.980000 ;
      RECT 0.190000  0.350000 2.160000 0.600000 ;
      RECT 0.190000  0.600000 0.520000 1.130000 ;
      RECT 0.565000  2.290000 0.895000 3.245000 ;
      RECT 1.095000  2.120000 1.265000 2.980000 ;
      RECT 1.465000  2.290000 1.795000 3.245000 ;
      RECT 1.990000  0.600000 2.160000 0.750000 ;
      RECT 1.990000  0.750000 3.960000 0.920000 ;
      RECT 1.995000  1.820000 2.165000 1.950000 ;
      RECT 1.995000  2.120000 2.165000 2.980000 ;
      RECT 2.340000  0.085000 2.670000 0.580000 ;
      RECT 2.365000  2.290000 2.615000 3.245000 ;
      RECT 2.815000  2.120000 3.145000 2.980000 ;
      RECT 2.850000  0.510000 3.020000 0.750000 ;
      RECT 3.200000  0.085000 3.530000 0.580000 ;
      RECT 3.345000  2.290000 3.515000 3.245000 ;
      RECT 3.710000  0.510000 3.960000 0.750000 ;
      RECT 3.715000  2.120000 3.995000 2.905000 ;
      RECT 3.715000  2.905000 5.845000 3.075000 ;
      RECT 4.180000  0.085000 4.430000 0.880000 ;
      RECT 4.665000  2.160000 4.895000 2.905000 ;
      RECT 4.915000  1.320000 6.195000 1.650000 ;
      RECT 5.040000  0.085000 5.290000 0.810000 ;
      RECT 5.565000  1.820000 5.845000 2.905000 ;
      RECT 5.900000  0.085000 6.230000 0.980000 ;
      RECT 6.025000  1.150000 6.660000 1.320000 ;
      RECT 6.025000  1.650000 6.195000 1.990000 ;
      RECT 6.025000  1.990000 6.815000 2.160000 ;
      RECT 6.035000  2.330000 6.365000 3.245000 ;
      RECT 6.400000  0.350000 6.660000 1.150000 ;
      RECT 6.535000  2.160000 6.815000 2.980000 ;
      RECT 7.015000  2.100000 7.265000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_ms__a21boi_4
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR C1 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=2.262e+12p pd=1.704e+07u as=1e+12p ps=8e+06u
M1001 X a_83_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=1.5521e+12p ps=1.276e+07u
M1002 VPWR A1 a_1341_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.8e+11p ps=5.36e+06u
M1003 a_83_244# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1341_392# A2 a_1034_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.015e+12p ps=8.03e+06u
M1005 a_1341_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_564_78# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.02922e+12p pd=9.63e+06u as=0p ps=0u
M1007 a_651_78# B1 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=6.88e+11p pd=4.71e+06u as=0p ps=0u
M1008 a_83_244# A3 a_1034_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_83_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=8.12e+11p pd=5.93e+06u as=0p ps=0u
M1010 X a_83_244# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_83_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1034_392# A3 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_83_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_83_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_564_78# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1034_392# A2 a_1341_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_83_244# C1 a_651_78# VNB nlowvt w=640000u l=150000u
+  ad=3.4395e+11p pd=2.59e+06u as=0p ps=0u
M1018 VPWR a_83_244# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_83_244# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B1 a_83_244# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_564_78# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A2 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_651_78# C1 a_83_244# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A3 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_83_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_564_78# B1 a_651_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A1 a_564_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

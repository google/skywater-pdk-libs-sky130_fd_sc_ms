* File: sky130_fd_sc_ms__xnor3_2.spice
* Created: Fri Aug 28 18:18:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xnor3_2.pex.spice"
.subckt sky130_fd_sc_ms__xnor3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_83_247#_M1012_g N_A_27_373#_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1010 N_A_83_247#_M1010_d N_A_M1010_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.12 AS=0.1152 PD=1.015 PS=1 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75000.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_329_81#_M1018_d N_B_M1018_g N_A_83_247#_M1010_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.144664 AS=0.12 PD=1.44906 PS=1.015 NRD=0 NRS=17.808 M=1 R=4.26667
+ SA=75001.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_A_27_373#_M1004_d N_A_397_21#_M1004_g N_A_329_81#_M1018_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0817019 AS=0.0949358 PD=0.792453 PS=0.950943 NRD=0
+ NRS=48.864 M=1 R=2.8 SA=75000.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_335_373#_M1003_d N_B_M1003_g N_A_27_373#_M1004_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.124498 PD=0.99 PS=1.20755 NRD=2.808 NRS=14.988 M=1
+ R=4.26667 SA=75001 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1002 N_A_83_247#_M1002_d N_A_397_21#_M1002_g N_A_335_373#_M1003_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.3525 AS=0.112 PD=2.83 PS=0.99 NRD=92.952 NRS=10.308 M=1
+ R=4.26667 SA=75001.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1016 N_VGND_M1016_d N_B_M1016_g N_A_397_21#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3368 AS=0.2109 PD=2.67 PS=2.05 NRD=64.884 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1023 N_A_1057_74#_M1023_d N_A_1027_48#_M1023_g N_A_329_81#_M1023_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_335_373#_M1019_d N_C_M1019_g N_A_1057_74#_M1023_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1013_d N_C_M1013_g N_A_1027_48#_M1013_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.276711 AS=0.1197 PD=1.33603 PS=1.41 NRD=172.524 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_1057_74#_M1009_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.487539 PD=1.02 PS=2.35397 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75000.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_X_M1009_d N_A_1057_74#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_A_83_247#_M1015_g N_A_27_373#_M1015_s VPB PSHORT L=0.18
+ W=1 AD=0.18 AS=0.28 PD=1.36 PS=2.56 NRD=1.9503 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1022 N_A_83_247#_M1022_d N_A_M1022_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=1
+ AD=0.187826 AS=0.18 PD=1.47826 PS=1.36 NRD=0.9653 NRS=13.7703 M=1 R=5.55556
+ SA=90000.7 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1000 N_A_335_373#_M1000_d N_B_M1000_g N_A_83_247#_M1022_d VPB PSHORT L=0.18
+ W=0.84 AD=0.185141 AS=0.157774 PD=1.44162 PS=1.24174 NRD=36.3465 NRS=18.1634
+ M=1 R=4.66667 SA=90001.3 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1011 N_A_27_373#_M1011_d N_A_397_21#_M1011_g N_A_335_373#_M1000_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.0928 AS=0.141059 PD=0.93 PS=1.09838 NRD=4.6098 NRS=0 M=1
+ R=3.55556 SA=90001.9 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1014 N_A_329_81#_M1014_d N_B_M1014_g N_A_27_373#_M1011_d VPB PSHORT L=0.18
+ W=0.64 AD=0.123849 AS=0.0928 PD=1.03784 PS=0.93 NRD=26.9299 NRS=0 M=1
+ R=3.55556 SA=90002.3 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1001 N_A_83_247#_M1001_d N_A_397_21#_M1001_g N_A_329_81#_M1014_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.364 AS=0.162551 PD=2.86 PS=1.36216 NRD=88.7091 NRS=0 M=1
+ R=4.66667 SA=90002.2 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1021 N_VPWR_M1021_d N_B_M1021_g N_A_397_21#_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.4214 AS=0.308 PD=3.12 PS=2.79 NRD=14.0658 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.3 A=0.2016 P=2.6 MULT=1
MM1005 N_A_1057_74#_M1005_d N_A_1027_48#_M1005_g N_A_335_373#_M1005_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.201225 AS=0.231 PD=1.405 PS=2.23 NRD=18.7544 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1007 N_A_329_81#_M1007_d N_C_M1007_g N_A_1057_74#_M1005_d VPB PSHORT L=0.18
+ W=0.84 AD=0.231 AS=0.201225 PD=2.23 PS=1.405 NRD=0 NRS=19.9167 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1020 N_VPWR_M1020_d N_C_M1020_g N_A_1027_48#_M1020_s VPB PSHORT L=0.18 W=0.64
+ AD=0.165236 AS=0.176 PD=1.17818 PS=1.83 NRD=70.7821 NRS=0 M=1 R=3.55556
+ SA=90000.2 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1006 N_X_M1006_d N_A_1057_74#_M1006_g N_VPWR_M1020_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.289164 PD=1.39 PS=2.06182 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1006_d N_A_1057_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
c_100 VNB 0 7.64129e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__xnor3_2.pxi.spice"
*
.ends
*
*

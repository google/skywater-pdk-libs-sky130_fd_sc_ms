* File: sky130_fd_sc_ms__dfrbp_2.pxi.spice
* Created: Wed Sep  2 12:02:49 2020
* 
x_PM_SKY130_FD_SC_MS__DFRBP_2%D N_D_M1036_g N_D_M1012_g N_D_c_266_n N_D_c_267_n
+ N_D_c_268_n D D N_D_c_270_n PM_SKY130_FD_SC_MS__DFRBP_2%D
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_298_294# N_A_298_294#_M1006_d
+ N_A_298_294#_M1011_s N_A_298_294#_M1024_d N_A_298_294#_M1023_g
+ N_A_298_294#_M1031_g N_A_298_294#_c_297_n N_A_298_294#_c_298_n
+ N_A_298_294#_c_299_n N_A_298_294#_c_300_n N_A_298_294#_c_301_n
+ N_A_298_294#_c_302_n N_A_298_294#_c_342_p N_A_298_294#_c_303_n
+ N_A_298_294#_c_304_n N_A_298_294#_c_305_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_298_294#
x_PM_SKY130_FD_SC_MS__DFRBP_2%RESET_B N_RESET_B_M1004_g N_RESET_B_M1037_g
+ N_RESET_B_c_403_n N_RESET_B_c_404_n N_RESET_B_M1011_g N_RESET_B_M1028_g
+ N_RESET_B_M1002_g N_RESET_B_M1021_g N_RESET_B_c_408_n N_RESET_B_c_409_n
+ N_RESET_B_c_410_n N_RESET_B_c_411_n N_RESET_B_c_412_n RESET_B
+ N_RESET_B_c_413_n N_RESET_B_c_414_n N_RESET_B_c_415_n N_RESET_B_c_416_n
+ N_RESET_B_c_417_n N_RESET_B_c_418_n PM_SKY130_FD_SC_MS__DFRBP_2%RESET_B
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_334_119# N_A_334_119#_M1031_d
+ N_A_334_119#_M1025_d N_A_334_119#_M1023_d N_A_334_119#_M1027_s
+ N_A_334_119#_M1015_g N_A_334_119#_c_607_n N_A_334_119#_M1013_g
+ N_A_334_119#_c_609_n N_A_334_119#_c_610_n N_A_334_119#_c_611_n
+ N_A_334_119#_c_612_n N_A_334_119#_c_647_n N_A_334_119#_c_635_n
+ N_A_334_119#_c_613_n N_A_334_119#_c_614_n N_A_334_119#_c_615_n
+ N_A_334_119#_c_616_n N_A_334_119#_c_617_n N_A_334_119#_c_618_n
+ N_A_334_119#_c_619_n N_A_334_119#_c_702_p N_A_334_119#_c_620_n
+ N_A_334_119#_c_621_n N_A_334_119#_c_622_n N_A_334_119#_c_623_n
+ N_A_334_119#_c_624_n N_A_334_119#_c_625_n N_A_334_119#_c_626_n
+ N_A_334_119#_c_627_n N_A_334_119#_c_628_n N_A_334_119#_c_629_n
+ N_A_334_119#_c_630_n N_A_334_119#_c_631_n N_A_334_119#_c_632_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_334_119#
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_818_418# N_A_818_418#_M1029_s
+ N_A_818_418#_M1034_s N_A_818_418#_M1026_g N_A_818_418#_M1032_g
+ N_A_818_418#_c_830_n N_A_818_418#_M1025_g N_A_818_418#_M1005_g
+ N_A_818_418#_c_832_n N_A_818_418#_c_833_n N_A_818_418#_c_834_n
+ N_A_818_418#_c_835_n N_A_818_418#_c_845_n N_A_818_418#_c_846_n
+ N_A_818_418#_c_847_n N_A_818_418#_c_848_n N_A_818_418#_c_849_n
+ N_A_818_418#_c_850_n N_A_818_418#_c_836_n N_A_818_418#_c_837_n
+ N_A_818_418#_c_838_n N_A_818_418#_c_839_n N_A_818_418#_c_854_n
+ N_A_818_418#_c_840_n N_A_818_418#_c_841_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_818_418#
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_728_331# N_A_728_331#_M1007_d
+ N_A_728_331#_M1009_d N_A_728_331#_M1024_g N_A_728_331#_M1006_g
+ N_A_728_331#_c_988_n N_A_728_331#_c_989_n N_A_728_331#_M1029_g
+ N_A_728_331#_M1034_g N_A_728_331#_c_999_n N_A_728_331#_M1017_g
+ N_A_728_331#_c_1001_n N_A_728_331#_M1027_g N_A_728_331#_c_992_n
+ N_A_728_331#_c_1002_n N_A_728_331#_c_1089_n N_A_728_331#_c_993_n
+ N_A_728_331#_c_1003_n N_A_728_331#_c_1024_n N_A_728_331#_c_994_n
+ N_A_728_331#_c_995_n N_A_728_331#_c_996_n N_A_728_331#_c_1027_n
+ N_A_728_331#_c_1006_n N_A_728_331#_c_1007_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_728_331#
x_PM_SKY130_FD_SC_MS__DFRBP_2%CLK N_CLK_c_1149_n N_CLK_M1007_g N_CLK_M1009_g CLK
+ N_CLK_c_1151_n PM_SKY130_FD_SC_MS__DFRBP_2%CLK
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_1800_291# N_A_1800_291#_M1018_d
+ N_A_1800_291#_M1002_d N_A_1800_291#_M1014_g N_A_1800_291#_c_1191_n
+ N_A_1800_291#_M1008_g N_A_1800_291#_c_1192_n N_A_1800_291#_c_1193_n
+ N_A_1800_291#_c_1194_n N_A_1800_291#_c_1229_n N_A_1800_291#_c_1233_p
+ N_A_1800_291#_c_1195_n N_A_1800_291#_c_1216_n N_A_1800_291#_c_1202_n
+ N_A_1800_291#_c_1196_n N_A_1800_291#_c_1197_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_1800_291#
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_1586_149# N_A_1586_149#_M1017_d
+ N_A_1586_149#_M1027_d N_A_1586_149#_M1018_g N_A_1586_149#_M1019_g
+ N_A_1586_149#_M1030_g N_A_1586_149#_c_1285_n N_A_1586_149#_M1010_g
+ N_A_1586_149#_M1035_g N_A_1586_149#_c_1286_n N_A_1586_149#_M1033_g
+ N_A_1586_149#_M1020_g N_A_1586_149#_M1022_g N_A_1586_149#_c_1303_n
+ N_A_1586_149#_c_1296_n N_A_1586_149#_c_1288_n N_A_1586_149#_c_1289_n
+ N_A_1586_149#_c_1298_n N_A_1586_149#_c_1290_n N_A_1586_149#_c_1291_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_1586_149#
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_2366_352# N_A_2366_352#_M1022_d
+ N_A_2366_352#_M1020_d N_A_2366_352#_M1000_g N_A_2366_352#_M1001_g
+ N_A_2366_352#_M1003_g N_A_2366_352#_M1016_g N_A_2366_352#_c_1423_n
+ N_A_2366_352#_c_1430_n N_A_2366_352#_c_1424_n N_A_2366_352#_c_1425_n
+ N_A_2366_352#_c_1426_n PM_SKY130_FD_SC_MS__DFRBP_2%A_2366_352#
x_PM_SKY130_FD_SC_MS__DFRBP_2%VPWR N_VPWR_M1036_s N_VPWR_M1004_d N_VPWR_M1011_d
+ N_VPWR_M1034_d N_VPWR_M1014_d N_VPWR_M1019_d N_VPWR_M1035_s N_VPWR_M1000_s
+ N_VPWR_M1003_s N_VPWR_c_1481_n N_VPWR_c_1482_n N_VPWR_c_1483_n N_VPWR_c_1484_n
+ N_VPWR_c_1485_n N_VPWR_c_1486_n N_VPWR_c_1487_n N_VPWR_c_1488_n
+ N_VPWR_c_1489_n N_VPWR_c_1490_n N_VPWR_c_1491_n N_VPWR_c_1492_n
+ N_VPWR_c_1493_n N_VPWR_c_1494_n N_VPWR_c_1495_n VPWR N_VPWR_c_1496_n
+ N_VPWR_c_1497_n N_VPWR_c_1498_n N_VPWR_c_1499_n N_VPWR_c_1500_n
+ N_VPWR_c_1501_n N_VPWR_c_1502_n N_VPWR_c_1503_n N_VPWR_c_1504_n
+ N_VPWR_c_1480_n PM_SKY130_FD_SC_MS__DFRBP_2%VPWR
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_70_74# N_A_70_74#_M1012_s N_A_70_74#_M1006_s
+ N_A_70_74#_M1036_d N_A_70_74#_M1026_d N_A_70_74#_c_1629_n N_A_70_74#_c_1634_n
+ N_A_70_74#_c_1635_n N_A_70_74#_c_1636_n N_A_70_74#_c_1637_n
+ N_A_70_74#_c_1638_n N_A_70_74#_c_1639_n N_A_70_74#_c_1640_n
+ N_A_70_74#_c_1641_n N_A_70_74#_c_1642_n N_A_70_74#_c_1643_n
+ N_A_70_74#_c_1644_n N_A_70_74#_c_1630_n N_A_70_74#_c_1631_n
+ N_A_70_74#_c_1646_n N_A_70_74#_c_1647_n N_A_70_74#_c_1632_n
+ N_A_70_74#_c_1649_n N_A_70_74#_c_1633_n PM_SKY130_FD_SC_MS__DFRBP_2%A_70_74#
x_PM_SKY130_FD_SC_MS__DFRBP_2%Q_N N_Q_N_M1010_s N_Q_N_M1030_d N_Q_N_c_1785_n
+ N_Q_N_c_1783_n Q_N PM_SKY130_FD_SC_MS__DFRBP_2%Q_N
x_PM_SKY130_FD_SC_MS__DFRBP_2%Q N_Q_M1001_d N_Q_M1000_d N_Q_c_1815_n
+ N_Q_c_1816_n N_Q_c_1812_n Q N_Q_c_1814_n Q PM_SKY130_FD_SC_MS__DFRBP_2%Q
x_PM_SKY130_FD_SC_MS__DFRBP_2%VGND N_VGND_M1037_d N_VGND_M1028_s N_VGND_M1029_d
+ N_VGND_M1008_d N_VGND_M1010_d N_VGND_M1033_d N_VGND_M1001_s N_VGND_M1016_s
+ N_VGND_c_1843_n N_VGND_c_1844_n N_VGND_c_1845_n N_VGND_c_1846_n
+ N_VGND_c_1847_n N_VGND_c_1848_n N_VGND_c_1849_n N_VGND_c_1850_n
+ N_VGND_c_1851_n N_VGND_c_1852_n N_VGND_c_1853_n N_VGND_c_1854_n
+ N_VGND_c_1855_n N_VGND_c_1856_n N_VGND_c_1857_n N_VGND_c_1858_n
+ N_VGND_c_1859_n VGND N_VGND_c_1860_n N_VGND_c_1861_n N_VGND_c_1862_n
+ N_VGND_c_1863_n N_VGND_c_1864_n N_VGND_c_1865_n N_VGND_c_1866_n
+ N_VGND_c_1867_n PM_SKY130_FD_SC_MS__DFRBP_2%VGND
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_614_81# N_A_614_81#_M1015_d N_A_614_81#_M1032_d
+ N_A_614_81#_c_1989_n N_A_614_81#_c_1990_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_614_81#
x_PM_SKY130_FD_SC_MS__DFRBP_2%A_1499_149# N_A_1499_149#_M1017_s
+ N_A_1499_149#_M1008_s N_A_1499_149#_c_2013_n N_A_1499_149#_c_2014_n
+ N_A_1499_149#_c_2015_n N_A_1499_149#_c_2016_n
+ PM_SKY130_FD_SC_MS__DFRBP_2%A_1499_149#
cc_1 VNB N_D_M1036_g 0.00700378f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=2.17
cc_2 VNB N_D_c_266_n 0.0210189f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_3 VNB N_D_c_267_n 0.0283274f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.05
cc_4 VNB N_D_c_268_n 0.0320517f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.57
cc_5 VNB D 0.0402073f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_D_c_270_n 0.02563f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.065
cc_7 VNB N_A_298_294#_M1031_g 0.021236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_298_294#_c_297_n 0.00685382f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.065
cc_9 VNB N_A_298_294#_c_298_n 0.00484772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_298_294#_c_299_n 0.0297732f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.065
cc_11 VNB N_A_298_294#_c_300_n 0.00387465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_298_294#_c_301_n 0.019696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_298_294#_c_302_n 0.00642483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_298_294#_c_303_n 0.00334726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_298_294#_c_304_n 0.00112476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_298_294#_c_305_n 3.53072e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_RESET_B_M1037_g 0.0431384f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.05
cc_18 VNB N_RESET_B_c_403_n 0.113795f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_19 VNB N_RESET_B_c_404_n 0.0123083f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.05
cc_20 VNB N_RESET_B_M1011_g 0.0323751f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_21 VNB N_RESET_B_M1028_g 0.0495583f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.065
cc_22 VNB N_RESET_B_M1021_g 0.0431388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_RESET_B_c_408_n 0.00884897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_RESET_B_c_409_n 0.00143791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_RESET_B_c_410_n 0.0404656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_RESET_B_c_411_n 0.00181538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_RESET_B_c_412_n 0.0015362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_RESET_B_c_413_n 0.0204572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_RESET_B_c_414_n 0.0015645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_RESET_B_c_415_n 0.0277655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_RESET_B_c_416_n 0.00462831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_c_417_n 0.0165198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_418_n 0.00386078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_334_119#_c_607_n 0.0270185f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.065
cc_35 VNB N_A_334_119#_M1013_g 0.0234715f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.925
cc_36 VNB N_A_334_119#_c_609_n 0.0156643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_334_119#_c_610_n 0.0113755f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.065
cc_38 VNB N_A_334_119#_c_611_n 0.00231808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_334_119#_c_612_n 0.0109602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_334_119#_c_613_n 0.0114601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_334_119#_c_614_n 0.0112194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_334_119#_c_615_n 0.00387155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_334_119#_c_616_n 0.0371118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_334_119#_c_617_n 0.00225927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_334_119#_c_618_n 0.00311976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_334_119#_c_619_n 0.00704603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_334_119#_c_620_n 0.0035579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_334_119#_c_621_n 0.00153929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_334_119#_c_622_n 0.0293297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_334_119#_c_623_n 0.00355388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_334_119#_c_624_n 0.0273514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_334_119#_c_625_n 0.0270442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_334_119#_c_626_n 0.0108619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_334_119#_c_627_n 0.00314018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_334_119#_c_628_n 0.00175721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_334_119#_c_629_n 0.00402758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_334_119#_c_630_n 8.59793e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_334_119#_c_631_n 0.00230646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_334_119#_c_632_n 0.0506314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_818_418#_M1032_g 0.040937f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_61 VNB N_A_818_418#_c_830_n 0.0204366f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.065
cc_62 VNB N_A_818_418#_M1005_g 0.00292692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_818_418#_c_832_n 0.0115671f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_64 VNB N_A_818_418#_c_833_n 0.0168787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_818_418#_c_834_n 0.0222244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_818_418#_c_835_n 0.0117883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_818_418#_c_836_n 6.24838e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_818_418#_c_837_n 0.00117943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_818_418#_c_838_n 0.0420897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_818_418#_c_839_n 0.00139432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_818_418#_c_840_n 0.00520919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_818_418#_c_841_n 0.0492961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_728_331#_M1024_g 0.0220127f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_74 VNB N_A_728_331#_M1006_g 0.0615892f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_75 VNB N_A_728_331#_c_988_n 0.111851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_728_331#_c_989_n 0.0102577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_728_331#_M1029_g 0.0143554f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.925
cc_78 VNB N_A_728_331#_M1017_g 0.0439787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_728_331#_c_992_n 0.0147343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_728_331#_c_993_n 0.00412543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_728_331#_c_994_n 0.0664706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_728_331#_c_995_n 0.00496454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_728_331#_c_996_n 0.00414255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_CLK_c_1149_n 0.0206637f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.57
cc_85 VNB CLK 0.00912873f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.05
cc_86 VNB N_CLK_c_1151_n 0.0389791f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.325
cc_87 VNB N_A_1800_291#_c_1191_n 0.0185916f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_88 VNB N_A_1800_291#_c_1192_n 0.0210915f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.065
cc_89 VNB N_A_1800_291#_c_1193_n 0.00103268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1800_291#_c_1194_n 0.0178538f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.065
cc_91 VNB N_A_1800_291#_c_1195_n 0.00794995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1800_291#_c_1196_n 0.00950159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1800_291#_c_1197_n 0.0271658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1586_149#_M1018_g 0.021266f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_95 VNB N_A_1586_149#_M1019_g 0.001735f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_96 VNB N_A_1586_149#_c_1285_n 0.0164413f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.065
cc_97 VNB N_A_1586_149#_c_1286_n 0.0144188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1586_149#_M1022_g 0.0229039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1586_149#_c_1288_n 0.00303624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1586_149#_c_1289_n 0.02459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1586_149#_c_1290_n 0.00358249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1586_149#_c_1291_n 0.151718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2366_352#_M1000_g 0.00188649f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_104 VNB N_A_2366_352#_M1001_g 0.0234349f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_105 VNB N_A_2366_352#_M1003_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.065
cc_106 VNB N_A_2366_352#_M1016_g 0.0265988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2366_352#_c_1423_n 0.00718732f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.065
cc_108 VNB N_A_2366_352#_c_1424_n 0.0169817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2366_352#_c_1425_n 0.0109542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2366_352#_c_1426_n 0.0767803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VPWR_c_1480_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_70_74#_c_1629_n 0.0104114f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_113 VNB N_A_70_74#_c_1630_n 0.00974934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_70_74#_c_1631_n 0.00594127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_70_74#_c_1632_n 0.00708308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_70_74#_c_1633_n 0.00977141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_Q_N_c_1783_n 0.00215184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB Q_N 5.1574e-19 $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=1.065
cc_119 VNB N_Q_c_1812_n 0.00335076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB Q 0.00448002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_Q_c_1814_n 0.00232136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1843_n 0.00898475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1844_n 0.00823049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1845_n 0.00652305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1846_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1847_n 0.00782424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1848_n 0.00524489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1849_n 0.0168886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1850_n 0.0103919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1851_n 0.0515355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1852_n 0.0185105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1853_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1854_n 0.071262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1855_n 0.00477852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1856_n 0.0835402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1857_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1858_n 0.0311181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1859_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1860_n 0.0337099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1861_n 0.0171743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1862_n 0.0188091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1863_n 0.0189106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1864_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1865_n 0.00632462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1866_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1867_n 0.735357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_614_81#_c_1989_n 0.0302536f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.58
cc_148 VNB N_A_614_81#_c_1990_n 0.0209611f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_149 VNB N_A_1499_149#_c_2013_n 0.00155523f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.9
cc_150 VNB N_A_1499_149#_c_2014_n 0.00899648f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.325
cc_151 VNB N_A_1499_149#_c_2015_n 0.00304708f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=1.57
cc_152 VNB N_A_1499_149#_c_2016_n 0.00653449f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_153 VPB N_D_M1036_g 0.0359018f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=2.17
cc_154 VPB N_A_298_294#_M1023_g 0.0245122f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.57
cc_155 VPB N_A_298_294#_c_297_n 0.0037484f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.065
cc_156 VPB N_A_298_294#_c_298_n 0.0017434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_298_294#_c_299_n 0.0194737f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.065
cc_158 VPB N_A_298_294#_c_300_n 0.00841927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_298_294#_c_302_n 0.00715762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_M1004_g 0.0219322f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=2.17
cc_161 VPB N_RESET_B_M1011_g 0.0268402f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.84
cc_162 VPB N_RESET_B_M1002_g 0.0259413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_408_n 0.00496561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_RESET_B_c_409_n 0.00720642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_RESET_B_c_410_n 0.0255385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_RESET_B_c_412_n 0.00230825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_RESET_B_c_413_n 0.0117937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_RESET_B_c_414_n 8.04582e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_RESET_B_c_417_n 0.0106231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_RESET_B_c_418_n 0.00189077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_334_119#_M1013_g 0.0221265f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.925
cc_172 VPB N_A_334_119#_c_611_n 0.00230449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_334_119#_c_635_n 0.00186364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_334_119#_c_628_n 0.00164564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_818_418#_M1026_g 0.0225511f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_176 VPB N_A_818_418#_M1005_g 0.0314026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_818_418#_c_835_n 0.00234699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_818_418#_c_845_n 0.00704052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_818_418#_c_846_n 0.0129394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_818_418#_c_847_n 0.0127007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_818_418#_c_848_n 0.00903971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_818_418#_c_849_n 0.0163995f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_818_418#_c_850_n 0.00534806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_818_418#_c_836_n 0.00284699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_818_418#_c_838_n 0.0193237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_818_418#_c_839_n 0.00504835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_818_418#_c_854_n 0.00436524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_728_331#_M1024_g 0.0200078f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_189 VPB N_A_728_331#_M1034_g 0.0305135f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.065
cc_190 VPB N_A_728_331#_c_999_n 0.0206163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_728_331#_M1017_g 0.00409839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_728_331#_c_1001_n 0.0349666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_728_331#_c_1002_n 0.003561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_728_331#_c_1003_n 0.00527774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_728_331#_c_994_n 0.0234418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_728_331#_c_995_n 8.76898e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_728_331#_c_1006_n 0.0017718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_728_331#_c_1007_n 0.0502965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_CLK_M1009_g 0.0286372f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=0.58
cc_200 VPB CLK 0.00114738f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.05
cc_201 VPB N_CLK_c_1151_n 0.00742415f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.325
cc_202 VPB N_A_1800_291#_M1014_g 0.0244967f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_203 VPB N_A_1800_291#_c_1193_n 0.00188652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1800_291#_c_1194_n 0.0125985f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.065
cc_205 VPB N_A_1800_291#_c_1195_n 0.00132863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1800_291#_c_1202_n 0.0104085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1586_149#_M1019_g 0.0331259f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.84
cc_208 VPB N_A_1586_149#_M1030_g 0.0215451f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.065
cc_209 VPB N_A_1586_149#_M1035_g 0.0220266f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_210 VPB N_A_1586_149#_M1020_g 0.0245043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1586_149#_c_1296_n 0.00819726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1586_149#_c_1288_n 0.00167495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1586_149#_c_1298_n 0.00176994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1586_149#_c_1291_n 0.0260122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_2366_352#_M1000_g 0.0250255f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_216 VPB N_A_2366_352#_M1003_g 0.0273944f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.065
cc_217 VPB N_A_2366_352#_c_1423_n 0.0138067f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.065
cc_218 VPB N_A_2366_352#_c_1430_n 0.014366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1481_n 0.0213265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1482_n 0.0551816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1483_n 0.0105202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1484_n 0.0722425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1485_n 0.0598931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1486_n 0.0300013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1487_n 0.0169533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1488_n 0.017583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1489_n 0.0281037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1490_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1491_n 0.0684935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1492_n 0.014661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1493_n 0.00780095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1494_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1495_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1496_n 0.0359062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1497_n 0.0763038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1498_n 0.0257899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1499_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1500_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1501_n 0.021173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1502_n 0.00689862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1503_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1504_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1480_n 0.212063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_70_74#_c_1634_n 0.00421024f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.065
cc_245 VPB N_A_70_74#_c_1635_n 0.00261742f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.925
cc_246 VPB N_A_70_74#_c_1636_n 0.00694245f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.065
cc_247 VPB N_A_70_74#_c_1637_n 0.00554076f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_248 VPB N_A_70_74#_c_1638_n 0.0231501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_70_74#_c_1639_n 4.17542e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_70_74#_c_1640_n 0.00645712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_70_74#_c_1641_n 8.66945e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_70_74#_c_1642_n 5.45555e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_70_74#_c_1643_n 0.0116901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_70_74#_c_1644_n 0.00217659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_70_74#_c_1631_n 0.00660484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_70_74#_c_1646_n 0.0116401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_70_74#_c_1647_n 0.00592749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_70_74#_c_1632_n 0.00217358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_70_74#_c_1649_n 0.00107725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_Q_N_c_1785_n 0.00438419f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_261 VPB N_Q_c_1815_n 0.00412671f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.9
cc_262 VPB N_Q_c_1816_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=1.325
cc_263 VPB N_Q_c_1812_n 0.00148895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 N_D_M1036_g N_RESET_B_M1004_g 0.0152952f $X=0.62 $Y=2.17 $X2=0 $Y2=0
cc_265 N_D_c_267_n N_RESET_B_M1037_g 0.0240229f $X=0.5 $Y=1.05 $X2=0 $Y2=0
cc_266 N_D_c_270_n N_RESET_B_M1037_g 0.0161854f $X=0.385 $Y=1.065 $X2=0 $Y2=0
cc_267 N_D_c_266_n N_RESET_B_c_404_n 0.0240229f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_268 N_D_c_268_n N_RESET_B_c_413_n 0.0171542f $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_269 N_D_c_268_n N_RESET_B_c_414_n 2.85099e-19 $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_270 N_D_M1036_g N_VPWR_c_1482_n 0.0042749f $X=0.62 $Y=2.17 $X2=0 $Y2=0
cc_271 N_D_c_268_n N_VPWR_c_1482_n 0.00205106f $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_272 D N_VPWR_c_1482_n 0.0195039f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_273 N_D_M1036_g N_VPWR_c_1492_n 0.00523095f $X=0.62 $Y=2.17 $X2=0 $Y2=0
cc_274 N_D_c_266_n N_A_70_74#_c_1629_n 0.00857082f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_275 N_D_c_267_n N_A_70_74#_c_1629_n 0.00462754f $X=0.5 $Y=1.05 $X2=0 $Y2=0
cc_276 D N_A_70_74#_c_1629_n 0.0156724f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_277 N_D_M1036_g N_A_70_74#_c_1634_n 0.00228068f $X=0.62 $Y=2.17 $X2=0 $Y2=0
cc_278 N_D_M1036_g N_A_70_74#_c_1635_n 0.0068046f $X=0.62 $Y=2.17 $X2=0 $Y2=0
cc_279 N_D_M1036_g N_A_70_74#_c_1632_n 0.0176322f $X=0.62 $Y=2.17 $X2=0 $Y2=0
cc_280 N_D_c_266_n N_A_70_74#_c_1632_n 0.0100763f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_281 N_D_c_267_n N_A_70_74#_c_1632_n 0.00567785f $X=0.5 $Y=1.05 $X2=0 $Y2=0
cc_282 N_D_c_268_n N_A_70_74#_c_1632_n 0.00556586f $X=0.465 $Y=1.57 $X2=0 $Y2=0
cc_283 D N_A_70_74#_c_1632_n 0.0551626f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_284 N_D_c_270_n N_A_70_74#_c_1632_n 0.00633941f $X=0.385 $Y=1.065 $X2=0 $Y2=0
cc_285 N_D_c_266_n N_VGND_c_1860_n 0.00296902f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_286 N_D_c_266_n N_VGND_c_1867_n 0.00367527f $X=0.5 $Y=0.9 $X2=0 $Y2=0
cc_287 D N_VGND_c_1867_n 0.00842173f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_288 N_A_298_294#_c_297_n N_RESET_B_M1004_g 0.0252019f $X=1.58 $Y=1.635 $X2=0
+ $Y2=0
cc_289 N_A_298_294#_M1031_g N_RESET_B_M1037_g 0.021518f $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_290 N_A_298_294#_M1031_g N_RESET_B_c_403_n 0.0101626f $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_291 N_A_298_294#_c_298_n N_RESET_B_M1011_g 0.00477445f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_292 N_A_298_294#_c_299_n N_RESET_B_M1011_g 0.00105273f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_293 N_A_298_294#_c_300_n N_RESET_B_M1011_g 0.010321f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_294 N_A_298_294#_c_301_n N_RESET_B_M1011_g 0.0185237f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_295 N_A_298_294#_c_297_n N_RESET_B_c_408_n 3.65631e-19 $X=1.58 $Y=1.635 $X2=0
+ $Y2=0
cc_296 N_A_298_294#_c_298_n N_RESET_B_c_408_n 0.0162655f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_297 N_A_298_294#_c_299_n N_RESET_B_c_408_n 0.00403772f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_298 N_A_298_294#_c_302_n N_RESET_B_c_408_n 0.0122088f $X=2.435 $Y=2.03 $X2=0
+ $Y2=0
cc_299 N_A_298_294#_c_301_n N_RESET_B_c_410_n 0.0243589f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_300 N_A_298_294#_c_303_n N_RESET_B_c_410_n 0.0190818f $X=4.002 $Y=1.945 $X2=0
+ $Y2=0
cc_301 N_A_298_294#_c_304_n N_RESET_B_c_410_n 0.00433885f $X=3.955 $Y=2.03 $X2=0
+ $Y2=0
cc_302 N_A_298_294#_c_305_n N_RESET_B_c_410_n 0.00550817f $X=4.05 $Y=1.44 $X2=0
+ $Y2=0
cc_303 N_A_298_294#_c_298_n N_RESET_B_c_411_n 6.49536e-19 $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_304 N_A_298_294#_c_301_n N_RESET_B_c_411_n 0.00789264f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_305 N_A_298_294#_M1031_g N_RESET_B_c_413_n 0.00107375f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_306 N_A_298_294#_c_297_n N_RESET_B_c_413_n 0.0201922f $X=1.58 $Y=1.635 $X2=0
+ $Y2=0
cc_307 N_A_298_294#_c_297_n N_RESET_B_c_414_n 8.3331e-19 $X=1.58 $Y=1.635 $X2=0
+ $Y2=0
cc_308 N_A_298_294#_M1031_g N_RESET_B_c_415_n 3.7765e-19 $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_309 N_A_298_294#_c_298_n N_RESET_B_c_415_n 4.89963e-19 $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_310 N_A_298_294#_c_299_n N_RESET_B_c_415_n 0.0184325f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_311 N_A_298_294#_c_301_n N_RESET_B_c_415_n 8.73334e-19 $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_312 N_A_298_294#_c_302_n N_RESET_B_c_415_n 0.00223986f $X=2.435 $Y=2.03 $X2=0
+ $Y2=0
cc_313 N_A_298_294#_c_298_n N_RESET_B_c_416_n 0.01583f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_314 N_A_298_294#_c_299_n N_RESET_B_c_416_n 0.00119402f $X=1.99 $Y=1.635 $X2=0
+ $Y2=0
cc_315 N_A_298_294#_c_302_n N_RESET_B_c_416_n 0.0235047f $X=2.435 $Y=2.03 $X2=0
+ $Y2=0
cc_316 N_A_298_294#_c_302_n N_A_334_119#_M1023_d 0.00352076f $X=2.435 $Y=2.03
+ $X2=0 $Y2=0
cc_317 N_A_298_294#_c_301_n N_A_334_119#_M1013_g 0.0132418f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_318 N_A_298_294#_c_342_p N_A_334_119#_M1013_g 0.00120833f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_319 N_A_298_294#_M1023_g N_A_334_119#_c_611_n 0.0134753f $X=1.58 $Y=2.46
+ $X2=0 $Y2=0
cc_320 N_A_298_294#_M1031_g N_A_334_119#_c_611_n 0.00924782f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_321 N_A_298_294#_c_297_n N_A_334_119#_c_611_n 0.0098523f $X=1.58 $Y=1.635
+ $X2=0 $Y2=0
cc_322 N_A_298_294#_c_298_n N_A_334_119#_c_611_n 0.0333361f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_323 N_A_298_294#_c_300_n N_A_334_119#_c_611_n 0.00534183f $X=2.35 $Y=2.57
+ $X2=0 $Y2=0
cc_324 N_A_298_294#_c_302_n N_A_334_119#_c_611_n 0.0132849f $X=2.435 $Y=2.03
+ $X2=0 $Y2=0
cc_325 N_A_298_294#_M1031_g N_A_334_119#_c_612_n 0.0106156f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_326 N_A_298_294#_M1023_g N_A_334_119#_c_647_n 0.00569928f $X=1.58 $Y=2.46
+ $X2=0 $Y2=0
cc_327 N_A_298_294#_M1023_g N_A_334_119#_c_635_n 6.83967e-19 $X=1.58 $Y=2.46
+ $X2=0 $Y2=0
cc_328 N_A_298_294#_c_299_n N_A_334_119#_c_635_n 0.0034741f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_329 N_A_298_294#_c_300_n N_A_334_119#_c_635_n 0.0120221f $X=2.35 $Y=2.57
+ $X2=0 $Y2=0
cc_330 N_A_298_294#_c_302_n N_A_334_119#_c_635_n 0.0102734f $X=2.435 $Y=2.03
+ $X2=0 $Y2=0
cc_331 N_A_298_294#_M1031_g N_A_334_119#_c_614_n 0.0123248f $X=1.595 $Y=0.965
+ $X2=0 $Y2=0
cc_332 N_A_298_294#_c_298_n N_A_334_119#_c_614_n 0.0253273f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_333 N_A_298_294#_c_299_n N_A_334_119#_c_614_n 0.00801172f $X=1.99 $Y=1.635
+ $X2=0 $Y2=0
cc_334 N_A_298_294#_c_301_n N_A_334_119#_c_630_n 0.021845f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_335 N_A_298_294#_c_305_n N_A_334_119#_c_630_n 0.00328107f $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_336 N_A_298_294#_c_301_n N_A_334_119#_c_632_n 0.00855282f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_337 N_A_298_294#_c_305_n N_A_334_119#_c_632_n 0.00106934f $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_338 N_A_298_294#_c_342_p N_A_818_418#_M1026_g 0.00830557f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_339 N_A_298_294#_c_303_n N_A_818_418#_M1032_g 0.00241812f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_340 N_A_298_294#_c_304_n N_A_818_418#_M1032_g 0.00133552f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_341 N_A_298_294#_c_342_p N_A_818_418#_c_832_n 0.00358646f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_342 N_A_298_294#_c_304_n N_A_818_418#_c_832_n 0.00149325f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_343 N_A_298_294#_c_305_n N_A_818_418#_c_832_n 3.65173e-19 $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_344 N_A_298_294#_c_301_n N_A_728_331#_M1024_g 0.0130291f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_345 N_A_298_294#_c_342_p N_A_728_331#_M1024_g 0.0128349f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_346 N_A_298_294#_c_303_n N_A_728_331#_M1024_g 0.00367203f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_347 N_A_298_294#_c_304_n N_A_728_331#_M1024_g 0.00312435f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_348 N_A_298_294#_c_303_n N_A_728_331#_M1006_g 0.00100194f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_349 N_A_298_294#_c_305_n N_A_728_331#_M1006_g 0.00895915f $X=4.05 $Y=1.44
+ $X2=0 $Y2=0
cc_350 N_A_298_294#_c_303_n N_A_728_331#_c_992_n 0.00470135f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_351 N_A_298_294#_c_304_n N_A_728_331#_c_992_n 0.00324895f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_352 N_A_298_294#_M1023_g N_VPWR_c_1493_n 0.00325836f $X=1.58 $Y=2.46 $X2=0
+ $Y2=0
cc_353 N_A_298_294#_M1023_g N_VPWR_c_1496_n 0.00363213f $X=1.58 $Y=2.46 $X2=0
+ $Y2=0
cc_354 N_A_298_294#_M1023_g N_VPWR_c_1480_n 0.00459536f $X=1.58 $Y=2.46 $X2=0
+ $Y2=0
cc_355 N_A_298_294#_M1023_g N_A_70_74#_c_1634_n 5.18041e-19 $X=1.58 $Y=2.46
+ $X2=0 $Y2=0
cc_356 N_A_298_294#_M1023_g N_A_70_74#_c_1635_n 0.0033814f $X=1.58 $Y=2.46 $X2=0
+ $Y2=0
cc_357 N_A_298_294#_M1023_g N_A_70_74#_c_1636_n 0.0100494f $X=1.58 $Y=2.46 $X2=0
+ $Y2=0
cc_358 N_A_298_294#_M1023_g N_A_70_74#_c_1638_n 0.00109206f $X=1.58 $Y=2.46
+ $X2=0 $Y2=0
cc_359 N_A_298_294#_c_300_n N_A_70_74#_c_1638_n 0.01889f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_360 N_A_298_294#_c_301_n N_A_70_74#_c_1640_n 0.0555839f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_361 N_A_298_294#_c_342_p N_A_70_74#_c_1640_n 0.0105352f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_362 N_A_298_294#_c_300_n N_A_70_74#_c_1641_n 0.0127294f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_363 N_A_298_294#_c_301_n N_A_70_74#_c_1641_n 0.0133351f $X=3.79 $Y=2.03 $X2=0
+ $Y2=0
cc_364 N_A_298_294#_c_342_p N_A_70_74#_c_1642_n 0.0151126f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_365 N_A_298_294#_c_342_p N_A_70_74#_c_1643_n 0.0204496f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_366 N_A_298_294#_c_305_n N_A_70_74#_c_1630_n 0.0169762f $X=4.05 $Y=1.44 $X2=0
+ $Y2=0
cc_367 N_A_298_294#_c_342_p N_A_70_74#_c_1631_n 0.0202223f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_368 N_A_298_294#_c_303_n N_A_70_74#_c_1631_n 0.0221864f $X=4.002 $Y=1.945
+ $X2=0 $Y2=0
cc_369 N_A_298_294#_c_304_n N_A_70_74#_c_1631_n 0.0127253f $X=3.955 $Y=2.03
+ $X2=0 $Y2=0
cc_370 N_A_298_294#_c_305_n N_A_70_74#_c_1631_n 0.0124256f $X=4.05 $Y=1.44 $X2=0
+ $Y2=0
cc_371 N_A_298_294#_c_342_p N_A_70_74#_c_1646_n 0.0127893f $X=3.955 $Y=2.57
+ $X2=0 $Y2=0
cc_372 N_A_298_294#_M1023_g N_A_70_74#_c_1649_n 0.0192136f $X=1.58 $Y=2.46 $X2=0
+ $Y2=0
cc_373 N_A_298_294#_c_300_n N_A_70_74#_c_1649_n 0.0044788f $X=2.35 $Y=2.57 $X2=0
+ $Y2=0
cc_374 N_A_298_294#_c_301_n N_A_70_74#_c_1633_n 0.00484801f $X=3.79 $Y=2.03
+ $X2=0 $Y2=0
cc_375 N_A_298_294#_M1031_g N_VGND_c_1843_n 0.0028854f $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_376 N_A_298_294#_M1031_g N_VGND_c_1844_n 8.31286e-19 $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_377 N_A_298_294#_M1031_g N_VGND_c_1867_n 7.88961e-19 $X=1.595 $Y=0.965 $X2=0
+ $Y2=0
cc_378 N_RESET_B_M1028_g N_A_334_119#_c_607_n 0.0171459f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_379 N_RESET_B_c_415_n N_A_334_119#_c_607_n 0.00381284f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_380 N_RESET_B_c_416_n N_A_334_119#_c_607_n 2.21753e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_381 N_RESET_B_M1011_g N_A_334_119#_M1013_g 0.0190315f $X=2.575 $Y=2.635 $X2=0
+ $Y2=0
cc_382 N_RESET_B_M1028_g N_A_334_119#_c_609_n 0.0348579f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_383 N_RESET_B_M1004_g N_A_334_119#_c_611_n 0.00243148f $X=1.07 $Y=2.17 $X2=0
+ $Y2=0
cc_384 N_RESET_B_M1037_g N_A_334_119#_c_611_n 0.00103829f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_385 N_RESET_B_c_408_n N_A_334_119#_c_611_n 0.0226342f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_386 N_RESET_B_c_409_n N_A_334_119#_c_611_n 0.00266791f $X=1.345 $Y=1.665
+ $X2=0 $Y2=0
cc_387 N_RESET_B_c_413_n N_A_334_119#_c_611_n 8.14073e-19 $X=1.115 $Y=1.615
+ $X2=0 $Y2=0
cc_388 N_RESET_B_c_414_n N_A_334_119#_c_611_n 0.023733f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_389 N_RESET_B_M1037_g N_A_334_119#_c_612_n 6.06377e-19 $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_390 N_RESET_B_c_403_n N_A_334_119#_c_612_n 0.00739262f $X=2.53 $Y=0.18 $X2=0
+ $Y2=0
cc_391 N_RESET_B_M1028_g N_A_334_119#_c_612_n 0.00635203f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_392 N_RESET_B_c_408_n N_A_334_119#_c_635_n 0.00472163f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_393 N_RESET_B_M1028_g N_A_334_119#_c_613_n 0.0172211f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_394 N_RESET_B_c_408_n N_A_334_119#_c_613_n 0.00885452f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_395 N_RESET_B_c_411_n N_A_334_119#_c_613_n 0.00142776f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_396 N_RESET_B_c_415_n N_A_334_119#_c_613_n 0.00395315f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_397 N_RESET_B_c_416_n N_A_334_119#_c_613_n 0.0175537f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_398 N_RESET_B_M1037_g N_A_334_119#_c_614_n 2.77273e-19 $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_399 N_RESET_B_M1028_g N_A_334_119#_c_614_n 0.00376661f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_400 N_RESET_B_c_408_n N_A_334_119#_c_614_n 0.00922151f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_401 N_RESET_B_M1028_g N_A_334_119#_c_615_n 0.00614625f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_402 N_RESET_B_M1028_g N_A_334_119#_c_617_n 0.00157742f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_403 N_RESET_B_M1028_g N_A_334_119#_c_618_n 0.00489643f $X=2.605 $Y=0.615
+ $X2=0 $Y2=0
cc_404 N_RESET_B_c_410_n N_A_334_119#_c_618_n 0.00204418f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_405 N_RESET_B_c_415_n N_A_334_119#_c_618_n 2.34651e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_406 N_RESET_B_c_416_n N_A_334_119#_c_618_n 0.008544f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_407 N_RESET_B_c_410_n N_A_334_119#_c_626_n 0.0139858f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_408 N_RESET_B_c_410_n N_A_334_119#_c_627_n 0.00558182f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_409 N_RESET_B_c_410_n N_A_334_119#_c_628_n 0.0242285f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_410 N_RESET_B_c_410_n N_A_334_119#_c_629_n 0.00503259f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_411 N_RESET_B_c_411_n N_A_334_119#_c_629_n 0.00118193f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_412 N_RESET_B_c_410_n N_A_334_119#_c_630_n 0.0217894f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_413 N_RESET_B_c_411_n N_A_334_119#_c_630_n 0.00230201f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_414 N_RESET_B_c_415_n N_A_334_119#_c_630_n 3.31881e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_415 N_RESET_B_c_416_n N_A_334_119#_c_630_n 0.0149803f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_416 N_RESET_B_M1011_g N_A_334_119#_c_632_n 0.00419637f $X=2.575 $Y=2.635
+ $X2=0 $Y2=0
cc_417 N_RESET_B_c_410_n N_A_334_119#_c_632_n 0.00756058f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_418 N_RESET_B_c_415_n N_A_334_119#_c_632_n 0.0168959f $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_419 N_RESET_B_c_416_n N_A_334_119#_c_632_n 8.2739e-19 $X=2.55 $Y=1.61 $X2=0
+ $Y2=0
cc_420 N_RESET_B_c_410_n N_A_818_418#_M1032_g 0.00702513f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_421 N_RESET_B_c_410_n N_A_818_418#_M1005_g 0.00255598f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_422 N_RESET_B_c_410_n N_A_818_418#_c_832_n 0.00175829f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_423 N_RESET_B_c_410_n N_A_818_418#_c_833_n 0.0108262f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_424 N_RESET_B_c_410_n N_A_818_418#_c_834_n 0.00323944f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_425 N_RESET_B_c_410_n N_A_818_418#_c_835_n 0.0319081f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_426 N_RESET_B_c_410_n N_A_818_418#_c_836_n 0.0156071f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_427 N_RESET_B_c_410_n N_A_818_418#_c_837_n 0.015652f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_428 N_RESET_B_c_410_n N_A_818_418#_c_839_n 0.0164077f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_429 N_RESET_B_c_410_n N_A_818_418#_c_840_n 0.0142935f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_430 N_RESET_B_c_410_n N_A_818_418#_c_841_n 0.0052628f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_431 N_RESET_B_c_410_n N_A_728_331#_M1006_g 0.00214871f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_432 N_RESET_B_c_410_n N_A_728_331#_M1034_g 0.00815231f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_433 N_RESET_B_c_410_n N_A_728_331#_c_999_n 0.00996207f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_434 N_RESET_B_c_410_n N_A_728_331#_M1017_g 0.00279101f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_435 N_RESET_B_c_410_n N_A_728_331#_c_1001_n 0.00829884f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_436 N_RESET_B_c_410_n N_A_728_331#_c_992_n 0.00419627f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_437 N_RESET_B_c_410_n N_A_728_331#_c_1002_n 0.0132491f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_438 N_RESET_B_c_410_n N_A_728_331#_c_993_n 6.34002e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_439 N_RESET_B_c_410_n N_A_728_331#_c_1024_n 0.033043f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_440 N_RESET_B_c_410_n N_A_728_331#_c_994_n 0.0112673f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_441 N_RESET_B_c_410_n N_A_728_331#_c_995_n 0.0200477f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_442 N_RESET_B_c_410_n N_A_728_331#_c_1027_n 0.0404507f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_443 N_RESET_B_c_410_n N_A_728_331#_c_1007_n 0.00622674f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_444 N_RESET_B_c_410_n N_CLK_M1009_g 0.00315336f $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_445 N_RESET_B_c_410_n CLK 0.023017f $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_446 N_RESET_B_c_410_n N_CLK_c_1151_n 0.00911865f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_447 N_RESET_B_M1002_g N_A_1800_291#_M1014_g 0.0150607f $X=9.77 $Y=2.155 $X2=0
+ $Y2=0
cc_448 N_RESET_B_M1021_g N_A_1800_291#_c_1191_n 0.0189671f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_449 N_RESET_B_M1002_g N_A_1800_291#_c_1193_n 0.00327579f $X=9.77 $Y=2.155
+ $X2=0 $Y2=0
cc_450 N_RESET_B_c_410_n N_A_1800_291#_c_1193_n 0.0212822f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_451 N_RESET_B_c_412_n N_A_1800_291#_c_1193_n 4.42853e-19 $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_452 N_RESET_B_c_417_n N_A_1800_291#_c_1193_n 5.04651e-19 $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_453 N_RESET_B_c_418_n N_A_1800_291#_c_1193_n 0.0185283f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_454 N_RESET_B_c_410_n N_A_1800_291#_c_1194_n 0.00455672f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_455 N_RESET_B_c_417_n N_A_1800_291#_c_1194_n 0.0211533f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_456 N_RESET_B_c_418_n N_A_1800_291#_c_1194_n 0.00111757f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_457 N_RESET_B_M1021_g N_A_1800_291#_c_1195_n 6.13047e-19 $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_458 N_RESET_B_c_412_n N_A_1800_291#_c_1195_n 0.0057125f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_459 N_RESET_B_c_418_n N_A_1800_291#_c_1195_n 0.00751959f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_460 N_RESET_B_M1002_g N_A_1800_291#_c_1216_n 0.0132475f $X=9.77 $Y=2.155
+ $X2=0 $Y2=0
cc_461 N_RESET_B_c_410_n N_A_1800_291#_c_1216_n 0.0101524f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_462 N_RESET_B_c_412_n N_A_1800_291#_c_1216_n 0.00804058f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_463 N_RESET_B_c_417_n N_A_1800_291#_c_1216_n 0.00301383f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_464 N_RESET_B_c_418_n N_A_1800_291#_c_1216_n 0.0234256f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_465 N_RESET_B_M1002_g N_A_1800_291#_c_1202_n 0.00757071f $X=9.77 $Y=2.155
+ $X2=0 $Y2=0
cc_466 N_RESET_B_M1021_g N_A_1800_291#_c_1196_n 0.00122306f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_467 N_RESET_B_M1021_g N_A_1800_291#_c_1197_n 0.0129042f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_417_n N_A_1800_291#_c_1197_n 2.59732e-19 $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_469 N_RESET_B_M1021_g N_A_1586_149#_M1018_g 0.0677574f $X=9.795 $Y=0.58 $X2=0
+ $Y2=0
cc_470 N_RESET_B_M1002_g N_A_1586_149#_M1019_g 0.0157555f $X=9.77 $Y=2.155 $X2=0
+ $Y2=0
cc_471 N_RESET_B_c_417_n N_A_1586_149#_M1019_g 0.0112352f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_410_n N_A_1586_149#_c_1303_n 0.0116802f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_473 N_RESET_B_c_410_n N_A_1586_149#_c_1288_n 0.0176982f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_474 N_RESET_B_M1021_g N_A_1586_149#_c_1289_n 0.0209819f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_475 N_RESET_B_c_410_n N_A_1586_149#_c_1289_n 0.017962f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_476 N_RESET_B_c_412_n N_A_1586_149#_c_1289_n 0.00291677f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_477 N_RESET_B_c_417_n N_A_1586_149#_c_1289_n 0.00422011f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_418_n N_A_1586_149#_c_1289_n 0.0280535f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_410_n N_A_1586_149#_c_1298_n 0.011953f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_480 N_RESET_B_M1021_g N_A_1586_149#_c_1291_n 0.0112352f $X=9.795 $Y=0.58
+ $X2=0 $Y2=0
cc_481 N_RESET_B_c_412_n N_A_1586_149#_c_1291_n 0.00422393f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_418_n N_A_1586_149#_c_1291_n 0.00318809f $X=9.705 $Y=1.615
+ $X2=0 $Y2=0
cc_483 N_RESET_B_M1011_g N_VPWR_c_1483_n 0.00111111f $X=2.575 $Y=2.635 $X2=0
+ $Y2=0
cc_484 N_RESET_B_M1002_g N_VPWR_c_1485_n 0.00405738f $X=9.77 $Y=2.155 $X2=0
+ $Y2=0
cc_485 N_RESET_B_c_410_n N_VPWR_c_1485_n 2.52709e-19 $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_486 N_RESET_B_M1004_g N_VPWR_c_1492_n 3.78197e-19 $X=1.07 $Y=2.17 $X2=0 $Y2=0
cc_487 N_RESET_B_M1011_g N_VPWR_c_1496_n 9.00187e-19 $X=2.575 $Y=2.635 $X2=0
+ $Y2=0
cc_488 N_RESET_B_M1002_g N_VPWR_c_1480_n 0.00461881f $X=9.77 $Y=2.155 $X2=0
+ $Y2=0
cc_489 N_RESET_B_M1037_g N_A_70_74#_c_1629_n 0.00192882f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_490 N_RESET_B_M1004_g N_A_70_74#_c_1634_n 0.0047611f $X=1.07 $Y=2.17 $X2=0
+ $Y2=0
cc_491 N_RESET_B_c_413_n N_A_70_74#_c_1634_n 0.00133324f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_492 N_RESET_B_M1004_g N_A_70_74#_c_1635_n 0.00932127f $X=1.07 $Y=2.17 $X2=0
+ $Y2=0
cc_493 N_RESET_B_M1004_g N_A_70_74#_c_1636_n 0.00659052f $X=1.07 $Y=2.17 $X2=0
+ $Y2=0
cc_494 N_RESET_B_M1011_g N_A_70_74#_c_1638_n 0.0118011f $X=2.575 $Y=2.635 $X2=0
+ $Y2=0
cc_495 N_RESET_B_M1011_g N_A_70_74#_c_1639_n 0.016483f $X=2.575 $Y=2.635 $X2=0
+ $Y2=0
cc_496 N_RESET_B_M1011_g N_A_70_74#_c_1641_n 0.00647474f $X=2.575 $Y=2.635 $X2=0
+ $Y2=0
cc_497 N_RESET_B_c_410_n N_A_70_74#_c_1630_n 0.0107306f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_498 N_RESET_B_c_410_n N_A_70_74#_c_1631_n 0.0218579f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_499 N_RESET_B_M1004_g N_A_70_74#_c_1632_n 0.00187008f $X=1.07 $Y=2.17 $X2=0
+ $Y2=0
cc_500 N_RESET_B_M1037_g N_A_70_74#_c_1632_n 0.00934166f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_501 N_RESET_B_c_409_n N_A_70_74#_c_1632_n 0.00155586f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_502 N_RESET_B_c_413_n N_A_70_74#_c_1632_n 0.0021837f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_503 N_RESET_B_c_414_n N_A_70_74#_c_1632_n 0.0230072f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_504 N_RESET_B_c_410_n N_A_70_74#_c_1633_n 0.0110159f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_505 N_RESET_B_M1037_g N_VGND_c_1843_n 0.00804421f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_506 N_RESET_B_c_403_n N_VGND_c_1843_n 0.0231021f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_507 N_RESET_B_c_413_n N_VGND_c_1843_n 0.00246294f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_414_n N_VGND_c_1843_n 0.00589903f $X=1.115 $Y=1.615 $X2=0
+ $Y2=0
cc_509 N_RESET_B_c_403_n N_VGND_c_1844_n 0.0228038f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_510 N_RESET_B_M1028_g N_VGND_c_1844_n 0.00790765f $X=2.605 $Y=0.615 $X2=0
+ $Y2=0
cc_511 N_RESET_B_M1021_g N_VGND_c_1846_n 0.0101946f $X=9.795 $Y=0.58 $X2=0 $Y2=0
cc_512 N_RESET_B_c_403_n N_VGND_c_1852_n 0.0211705f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_513 N_RESET_B_c_403_n N_VGND_c_1854_n 0.00564095f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_514 N_RESET_B_M1021_g N_VGND_c_1858_n 0.00383152f $X=9.795 $Y=0.58 $X2=0
+ $Y2=0
cc_515 N_RESET_B_c_404_n N_VGND_c_1860_n 0.00600995f $X=1.14 $Y=0.18 $X2=0 $Y2=0
cc_516 N_RESET_B_c_403_n N_VGND_c_1867_n 0.0377703f $X=2.53 $Y=0.18 $X2=0 $Y2=0
cc_517 N_RESET_B_c_404_n N_VGND_c_1867_n 0.0112887f $X=1.14 $Y=0.18 $X2=0 $Y2=0
cc_518 N_RESET_B_M1021_g N_VGND_c_1867_n 0.0075694f $X=9.795 $Y=0.58 $X2=0 $Y2=0
cc_519 N_RESET_B_c_410_n N_A_614_81#_c_1990_n 0.0159116f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_520 N_RESET_B_c_410_n N_A_1499_149#_c_2013_n 4.58014e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_334_119#_c_619_n N_A_818_418#_M1029_s 0.00227252f $X=5.15 $Y=0.66
+ $X2=-0.19 $Y2=-0.245
cc_522 N_A_334_119#_c_702_p N_A_818_418#_M1029_s 0.0027085f $X=6.025 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_523 N_A_334_119#_c_620_n N_A_818_418#_M1029_s 0.00199188f $X=5.235 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_524 N_A_334_119#_c_625_n N_A_818_418#_c_830_n 0.0119277f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_525 N_A_334_119#_c_702_p N_A_818_418#_c_835_n 0.0105363f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_526 N_A_334_119#_c_620_n N_A_818_418#_c_835_n 0.0124528f $X=5.235 $Y=0.745
+ $X2=0 $Y2=0
cc_527 N_A_334_119#_c_628_n N_A_818_418#_c_847_n 0.0123434f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_528 N_A_334_119#_c_628_n N_A_818_418#_c_848_n 0.00909361f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_529 N_A_334_119#_M1027_s N_A_818_418#_c_849_n 0.00366073f $X=7.665 $Y=1.945
+ $X2=0 $Y2=0
cc_530 N_A_334_119#_c_628_n N_A_818_418#_c_849_n 0.0123303f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_531 N_A_334_119#_c_628_n N_A_818_418#_c_836_n 0.0499795f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_532 N_A_334_119#_c_624_n N_A_818_418#_c_840_n 0.0024581f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_533 N_A_334_119#_c_626_n N_A_818_418#_c_840_n 0.0147826f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_534 N_A_334_119#_c_628_n N_A_818_418#_c_840_n 0.00609504f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_535 N_A_334_119#_M1013_g N_A_728_331#_M1024_g 0.0412924f $X=3.34 $Y=2.635
+ $X2=0 $Y2=0
cc_536 N_A_334_119#_c_610_n N_A_728_331#_M1006_g 0.007711f $X=3.012 $Y=1.05
+ $X2=0 $Y2=0
cc_537 N_A_334_119#_c_616_n N_A_728_331#_M1006_g 0.00252325f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_538 N_A_334_119#_c_618_n N_A_728_331#_M1006_g 7.95442e-19 $X=3.01 $Y=1.555
+ $X2=0 $Y2=0
cc_539 N_A_334_119#_c_630_n N_A_728_331#_M1006_g 2.86655e-19 $X=3.09 $Y=1.68
+ $X2=0 $Y2=0
cc_540 N_A_334_119#_c_632_n N_A_728_331#_M1006_g 0.00556159f $X=3.34 $Y=1.68
+ $X2=0 $Y2=0
cc_541 N_A_334_119#_c_616_n N_A_728_331#_c_988_n 0.0575563f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_542 N_A_334_119#_c_702_p N_A_728_331#_c_988_n 0.00157743f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_543 N_A_334_119#_c_609_n N_A_728_331#_c_989_n 0.00720262f $X=3.012 $Y=0.9
+ $X2=0 $Y2=0
cc_544 N_A_334_119#_c_616_n N_A_728_331#_c_989_n 0.0074164f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_545 N_A_334_119#_c_616_n N_A_728_331#_M1029_g 2.14932e-19 $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_546 N_A_334_119#_c_619_n N_A_728_331#_M1029_g 0.00722282f $X=5.15 $Y=0.66
+ $X2=0 $Y2=0
cc_547 N_A_334_119#_c_702_p N_A_728_331#_M1029_g 0.0190035f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_548 N_A_334_119#_c_621_n N_A_728_331#_M1029_g 0.00429098f $X=6.11 $Y=0.66
+ $X2=0 $Y2=0
cc_549 N_A_334_119#_c_628_n N_A_728_331#_c_999_n 0.00926793f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_550 N_A_334_119#_c_624_n N_A_728_331#_M1017_g 0.00510454f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_551 N_A_334_119#_c_625_n N_A_728_331#_M1017_g 9.86678e-19 $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_552 N_A_334_119#_c_626_n N_A_728_331#_M1017_g 0.00939999f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_553 N_A_334_119#_c_628_n N_A_728_331#_M1017_g 0.00547121f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_554 N_A_334_119#_c_628_n N_A_728_331#_c_1001_n 0.0073511f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_555 N_A_334_119#_c_630_n N_A_728_331#_c_992_n 3.90209e-19 $X=3.09 $Y=1.68
+ $X2=0 $Y2=0
cc_556 N_A_334_119#_c_632_n N_A_728_331#_c_992_n 0.0412924f $X=3.34 $Y=1.68
+ $X2=0 $Y2=0
cc_557 N_A_334_119#_c_626_n N_A_728_331#_c_1003_n 0.00320602f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_558 N_A_334_119#_c_627_n N_A_728_331#_c_1003_n 0.00513005f $X=7.385 $Y=1.44
+ $X2=0 $Y2=0
cc_559 N_A_334_119#_c_628_n N_A_728_331#_c_1003_n 0.0223244f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_560 N_A_334_119#_c_702_p N_A_728_331#_c_1024_n 0.0191238f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_561 N_A_334_119#_c_702_p N_A_728_331#_c_994_n 0.0116618f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_562 N_A_334_119#_c_702_p N_A_728_331#_c_996_n 0.0151771f $X=6.025 $Y=0.745
+ $X2=0 $Y2=0
cc_563 N_A_334_119#_c_621_n N_A_728_331#_c_996_n 0.001895f $X=6.11 $Y=0.66 $X2=0
+ $Y2=0
cc_564 N_A_334_119#_c_622_n N_A_728_331#_c_996_n 0.0322868f $X=7.215 $Y=0.34
+ $X2=0 $Y2=0
cc_565 N_A_334_119#_c_624_n N_A_728_331#_c_996_n 0.0206296f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_566 N_A_334_119#_c_628_n N_A_728_331#_c_1006_n 0.00241743f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_567 N_A_334_119#_c_626_n N_A_728_331#_c_1007_n 0.00851598f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_568 N_A_334_119#_c_627_n N_A_728_331#_c_1007_n 0.00337292f $X=7.385 $Y=1.44
+ $X2=0 $Y2=0
cc_569 N_A_334_119#_c_628_n N_A_728_331#_c_1007_n 0.0010833f $X=7.795 $Y=2.09
+ $X2=0 $Y2=0
cc_570 N_A_334_119#_c_702_p N_CLK_c_1149_n 9.69516e-19 $X=6.025 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_571 N_A_334_119#_c_621_n N_CLK_c_1149_n 0.0063257f $X=6.11 $Y=0.66 $X2=-0.19
+ $Y2=-0.245
cc_572 N_A_334_119#_c_622_n N_CLK_c_1149_n 0.00861985f $X=7.215 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_573 N_A_334_119#_c_624_n N_CLK_c_1149_n 0.0091992f $X=7.3 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_574 N_A_334_119#_c_624_n CLK 0.0138701f $X=7.3 $Y=1.355 $X2=0 $Y2=0
cc_575 N_A_334_119#_c_627_n CLK 0.0150422f $X=7.385 $Y=1.44 $X2=0 $Y2=0
cc_576 N_A_334_119#_c_628_n CLK 0.00323555f $X=7.795 $Y=2.09 $X2=0 $Y2=0
cc_577 N_A_334_119#_c_627_n N_CLK_c_1151_n 0.00108413f $X=7.385 $Y=1.44 $X2=0
+ $Y2=0
cc_578 N_A_334_119#_c_625_n N_A_1800_291#_c_1191_n 0.00175601f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_579 N_A_334_119#_M1025_d N_A_1586_149#_c_1303_n 0.00571341f $X=8.405 $Y=0.425
+ $X2=0 $Y2=0
cc_580 N_A_334_119#_M1025_d N_A_1586_149#_c_1290_n 0.0013268f $X=8.405 $Y=0.425
+ $X2=0 $Y2=0
cc_581 N_A_334_119#_M1013_g N_VPWR_c_1483_n 0.00321759f $X=3.34 $Y=2.635 $X2=0
+ $Y2=0
cc_582 N_A_334_119#_M1013_g N_VPWR_c_1484_n 0.00413068f $X=3.34 $Y=2.635 $X2=0
+ $Y2=0
cc_583 N_A_334_119#_M1013_g N_VPWR_c_1480_n 0.00390913f $X=3.34 $Y=2.635 $X2=0
+ $Y2=0
cc_584 N_A_334_119#_c_611_n N_A_70_74#_c_1634_n 0.00560265f $X=1.57 $Y=2.285
+ $X2=0 $Y2=0
cc_585 N_A_334_119#_c_647_n N_A_70_74#_c_1636_n 0.00876016f $X=1.655 $Y=2.37
+ $X2=0 $Y2=0
cc_586 N_A_334_119#_M1023_d N_A_70_74#_c_1638_n 0.0034154f $X=1.67 $Y=1.96 $X2=0
+ $Y2=0
cc_587 N_A_334_119#_c_635_n N_A_70_74#_c_1638_n 0.00696584f $X=1.805 $Y=2.37
+ $X2=0 $Y2=0
cc_588 N_A_334_119#_M1013_g N_A_70_74#_c_1639_n 0.001637f $X=3.34 $Y=2.635 $X2=0
+ $Y2=0
cc_589 N_A_334_119#_M1013_g N_A_70_74#_c_1640_n 0.0140935f $X=3.34 $Y=2.635
+ $X2=0 $Y2=0
cc_590 N_A_334_119#_M1013_g N_A_70_74#_c_1642_n 0.0100927f $X=3.34 $Y=2.635
+ $X2=0 $Y2=0
cc_591 N_A_334_119#_M1013_g N_A_70_74#_c_1644_n 0.00267271f $X=3.34 $Y=2.635
+ $X2=0 $Y2=0
cc_592 N_A_334_119#_c_611_n N_A_70_74#_c_1632_n 0.00906065f $X=1.57 $Y=2.285
+ $X2=0 $Y2=0
cc_593 N_A_334_119#_M1023_d N_A_70_74#_c_1649_n 0.00898705f $X=1.67 $Y=1.96
+ $X2=0 $Y2=0
cc_594 N_A_334_119#_c_647_n N_A_70_74#_c_1649_n 0.00397928f $X=1.655 $Y=2.37
+ $X2=0 $Y2=0
cc_595 N_A_334_119#_c_635_n N_A_70_74#_c_1649_n 0.00473461f $X=1.805 $Y=2.37
+ $X2=0 $Y2=0
cc_596 N_A_334_119#_c_610_n N_A_70_74#_c_1633_n 0.00441246f $X=3.012 $Y=1.05
+ $X2=0 $Y2=0
cc_597 N_A_334_119#_c_615_n N_A_70_74#_c_1633_n 0.00314822f $X=2.79 $Y=1.015
+ $X2=0 $Y2=0
cc_598 N_A_334_119#_c_618_n N_A_70_74#_c_1633_n 0.0114522f $X=3.01 $Y=1.555
+ $X2=0 $Y2=0
cc_599 N_A_334_119#_c_629_n N_A_70_74#_c_1633_n 0.0106126f $X=3.01 $Y=1.1 $X2=0
+ $Y2=0
cc_600 N_A_334_119#_c_632_n N_A_70_74#_c_1633_n 0.00282478f $X=3.34 $Y=1.68
+ $X2=0 $Y2=0
cc_601 N_A_334_119#_c_702_p N_VGND_M1029_d 0.0205914f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_602 N_A_334_119#_c_621_n N_VGND_M1029_d 0.00621489f $X=6.11 $Y=0.66 $X2=0
+ $Y2=0
cc_603 N_A_334_119#_c_612_n N_VGND_c_1843_n 0.0314529f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_604 N_A_334_119#_c_609_n N_VGND_c_1844_n 2.1461e-19 $X=3.012 $Y=0.9 $X2=0
+ $Y2=0
cc_605 N_A_334_119#_c_612_n N_VGND_c_1844_n 0.0289901f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_606 N_A_334_119#_c_613_n N_VGND_c_1844_n 0.0194224f $X=2.705 $Y=1.1 $X2=0
+ $Y2=0
cc_607 N_A_334_119#_c_617_n N_VGND_c_1844_n 0.0133176f $X=2.875 $Y=0.34 $X2=0
+ $Y2=0
cc_608 N_A_334_119#_c_616_n N_VGND_c_1845_n 0.00787195f $X=5.065 $Y=0.34 $X2=0
+ $Y2=0
cc_609 N_A_334_119#_c_619_n N_VGND_c_1845_n 0.00291186f $X=5.15 $Y=0.66 $X2=0
+ $Y2=0
cc_610 N_A_334_119#_c_702_p N_VGND_c_1845_n 0.0190193f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_611 N_A_334_119#_c_621_n N_VGND_c_1845_n 0.00491053f $X=6.11 $Y=0.66 $X2=0
+ $Y2=0
cc_612 N_A_334_119#_c_623_n N_VGND_c_1845_n 0.0145006f $X=6.195 $Y=0.34 $X2=0
+ $Y2=0
cc_613 N_A_334_119#_c_625_n N_VGND_c_1846_n 0.00292246f $X=8.615 $Y=0.34 $X2=0
+ $Y2=0
cc_614 N_A_334_119#_c_612_n N_VGND_c_1852_n 0.0146228f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_615 N_A_334_119#_c_609_n N_VGND_c_1854_n 9.15902e-19 $X=3.012 $Y=0.9 $X2=0
+ $Y2=0
cc_616 N_A_334_119#_c_616_n N_VGND_c_1854_n 0.153051f $X=5.065 $Y=0.34 $X2=0
+ $Y2=0
cc_617 N_A_334_119#_c_617_n N_VGND_c_1854_n 0.0121867f $X=2.875 $Y=0.34 $X2=0
+ $Y2=0
cc_618 N_A_334_119#_c_702_p N_VGND_c_1854_n 0.0051071f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_619 N_A_334_119#_c_702_p N_VGND_c_1856_n 0.00279509f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_620 N_A_334_119#_c_622_n N_VGND_c_1856_n 0.0656484f $X=7.215 $Y=0.34 $X2=0
+ $Y2=0
cc_621 N_A_334_119#_c_623_n N_VGND_c_1856_n 0.0120335f $X=6.195 $Y=0.34 $X2=0
+ $Y2=0
cc_622 N_A_334_119#_c_625_n N_VGND_c_1856_n 0.0895608f $X=8.615 $Y=0.34 $X2=0
+ $Y2=0
cc_623 N_A_334_119#_c_631_n N_VGND_c_1856_n 0.0121867f $X=7.3 $Y=0.34 $X2=0
+ $Y2=0
cc_624 N_A_334_119#_M1025_d N_VGND_c_1867_n 0.00257669f $X=8.405 $Y=0.425 $X2=0
+ $Y2=0
cc_625 N_A_334_119#_c_612_n N_VGND_c_1867_n 0.010799f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_626 N_A_334_119#_c_616_n N_VGND_c_1867_n 0.0889116f $X=5.065 $Y=0.34 $X2=0
+ $Y2=0
cc_627 N_A_334_119#_c_617_n N_VGND_c_1867_n 0.00660921f $X=2.875 $Y=0.34 $X2=0
+ $Y2=0
cc_628 N_A_334_119#_c_702_p N_VGND_c_1867_n 0.0161016f $X=6.025 $Y=0.745 $X2=0
+ $Y2=0
cc_629 N_A_334_119#_c_622_n N_VGND_c_1867_n 0.0383417f $X=7.215 $Y=0.34 $X2=0
+ $Y2=0
cc_630 N_A_334_119#_c_623_n N_VGND_c_1867_n 0.00658039f $X=6.195 $Y=0.34 $X2=0
+ $Y2=0
cc_631 N_A_334_119#_c_625_n N_VGND_c_1867_n 0.052445f $X=8.615 $Y=0.34 $X2=0
+ $Y2=0
cc_632 N_A_334_119#_c_631_n N_VGND_c_1867_n 0.00660921f $X=7.3 $Y=0.34 $X2=0
+ $Y2=0
cc_633 N_A_334_119#_c_615_n A_536_81# 0.00157084f $X=2.79 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_634 N_A_334_119#_c_616_n N_A_614_81#_M1015_d 0.00277417f $X=5.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_635 N_A_334_119#_c_609_n N_A_614_81#_c_1989_n 0.00242033f $X=3.012 $Y=0.9
+ $X2=0 $Y2=0
cc_636 N_A_334_119#_c_616_n N_A_614_81#_c_1989_n 0.127151f $X=5.065 $Y=0.34
+ $X2=0 $Y2=0
cc_637 N_A_334_119#_c_619_n N_A_614_81#_c_1989_n 0.00545207f $X=5.15 $Y=0.66
+ $X2=0 $Y2=0
cc_638 N_A_334_119#_c_620_n N_A_614_81#_c_1989_n 0.00983818f $X=5.235 $Y=0.745
+ $X2=0 $Y2=0
cc_639 N_A_334_119#_c_629_n N_A_614_81#_c_1989_n 0.00184287f $X=3.01 $Y=1.1
+ $X2=0 $Y2=0
cc_640 N_A_334_119#_c_620_n N_A_614_81#_c_1990_n 0.00559801f $X=5.235 $Y=0.745
+ $X2=0 $Y2=0
cc_641 N_A_334_119#_c_624_n N_A_1499_149#_c_2013_n 0.0310557f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_642 N_A_334_119#_c_626_n N_A_1499_149#_c_2013_n 0.0133791f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_643 N_A_334_119#_M1025_d N_A_1499_149#_c_2014_n 0.00704081f $X=8.405 $Y=0.425
+ $X2=0 $Y2=0
cc_644 N_A_334_119#_c_625_n N_A_1499_149#_c_2014_n 0.0689604f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_645 N_A_334_119#_c_626_n N_A_1499_149#_c_2014_n 0.00378293f $X=7.71 $Y=1.44
+ $X2=0 $Y2=0
cc_646 N_A_334_119#_c_624_n N_A_1499_149#_c_2015_n 0.0143225f $X=7.3 $Y=1.355
+ $X2=0 $Y2=0
cc_647 N_A_334_119#_c_625_n N_A_1499_149#_c_2015_n 0.0132852f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_648 N_A_334_119#_c_625_n N_A_1499_149#_c_2016_n 0.00562463f $X=8.615 $Y=0.34
+ $X2=0 $Y2=0
cc_649 N_A_818_418#_c_847_n N_A_728_331#_M1009_d 0.00762356f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_650 N_A_818_418#_M1032_g N_A_728_331#_M1024_g 0.00720264f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_651 N_A_818_418#_c_832_n N_A_728_331#_M1024_g 0.0255473f $X=4.215 $Y=2.165
+ $X2=0 $Y2=0
cc_652 N_A_818_418#_M1032_g N_A_728_331#_M1006_g 0.0191869f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_653 N_A_818_418#_M1032_g N_A_728_331#_c_988_n 0.00194711f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_654 N_A_818_418#_c_835_n N_A_728_331#_c_988_n 4.78794e-19 $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_655 N_A_818_418#_c_835_n N_A_728_331#_M1029_g 0.0172164f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_656 N_A_818_418#_c_835_n N_A_728_331#_M1034_g 0.00313167f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_657 N_A_818_418#_c_845_n N_A_728_331#_M1034_g 0.00828611f $X=5.605 $Y=2.425
+ $X2=0 $Y2=0
cc_658 N_A_818_418#_c_846_n N_A_728_331#_M1034_g 0.0112382f $X=5.62 $Y=2.815
+ $X2=0 $Y2=0
cc_659 N_A_818_418#_c_847_n N_A_728_331#_M1034_g 0.0159172f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_660 N_A_818_418#_c_838_n N_A_728_331#_M1034_g 0.00418573f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_661 N_A_818_418#_c_839_n N_A_728_331#_M1034_g 0.00909396f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_662 N_A_818_418#_c_854_n N_A_728_331#_M1034_g 4.64231e-19 $X=5.605 $Y=2.51
+ $X2=0 $Y2=0
cc_663 N_A_818_418#_c_830_n N_A_728_331#_M1017_g 0.017713f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_664 N_A_818_418#_M1005_g N_A_728_331#_M1017_g 0.00179297f $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_665 N_A_818_418#_c_836_n N_A_728_331#_M1017_g 9.47689e-19 $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_666 N_A_818_418#_c_840_n N_A_728_331#_M1017_g 0.0029963f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_667 N_A_818_418#_c_841_n N_A_728_331#_M1017_g 0.00522227f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_668 N_A_818_418#_M1005_g N_A_728_331#_c_1001_n 0.0110263f $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_669 N_A_818_418#_c_848_n N_A_728_331#_c_1001_n 0.00278374f $X=7.41 $Y=2.905
+ $X2=0 $Y2=0
cc_670 N_A_818_418#_c_849_n N_A_728_331#_c_1001_n 0.0153683f $X=8.05 $Y=2.99
+ $X2=0 $Y2=0
cc_671 N_A_818_418#_c_836_n N_A_728_331#_c_1001_n 0.03443f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_672 N_A_818_418#_c_840_n N_A_728_331#_c_1001_n 3.50893e-19 $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_673 N_A_818_418#_c_835_n N_A_728_331#_c_1002_n 0.00408409f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_674 N_A_818_418#_c_847_n N_A_728_331#_c_1089_n 0.00999472f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_675 N_A_818_418#_c_839_n N_A_728_331#_c_1089_n 0.0180713f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_676 N_A_818_418#_c_847_n N_A_728_331#_c_1003_n 0.027879f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_677 N_A_818_418#_c_835_n N_A_728_331#_c_1024_n 0.0251507f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_678 N_A_818_418#_c_839_n N_A_728_331#_c_1024_n 0.0104391f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_679 N_A_818_418#_c_835_n N_A_728_331#_c_994_n 0.0119567f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_680 N_A_818_418#_c_839_n N_A_728_331#_c_994_n 0.00909499f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_681 N_A_818_418#_c_847_n N_A_728_331#_c_1027_n 0.0208991f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_682 N_A_818_418#_c_847_n N_A_728_331#_c_1006_n 0.0211506f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_683 N_A_818_418#_c_847_n N_A_728_331#_c_1007_n 0.00761439f $X=7.315 $Y=2.51
+ $X2=0 $Y2=0
cc_684 N_A_818_418#_c_847_n N_CLK_M1009_g 0.0176081f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_685 N_A_818_418#_c_848_n N_CLK_M1009_g 0.00714171f $X=7.41 $Y=2.905 $X2=0
+ $Y2=0
cc_686 N_A_818_418#_c_850_n N_CLK_M1009_g 0.00464142f $X=7.505 $Y=2.99 $X2=0
+ $Y2=0
cc_687 N_A_818_418#_M1005_g N_A_1800_291#_M1014_g 0.0371377f $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_688 N_A_818_418#_c_841_n N_A_1800_291#_c_1193_n 5.09728e-19 $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_689 N_A_818_418#_c_841_n N_A_1800_291#_c_1194_n 0.0212366f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_690 N_A_818_418#_M1005_g N_A_1800_291#_c_1229_n 2.32678e-19 $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_691 N_A_818_418#_c_841_n N_A_1800_291#_c_1197_n 0.00528894f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_692 N_A_818_418#_c_849_n N_A_1586_149#_M1027_d 0.00180442f $X=8.05 $Y=2.99
+ $X2=0 $Y2=0
cc_693 N_A_818_418#_c_836_n N_A_1586_149#_M1027_d 0.0211382f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_694 N_A_818_418#_c_830_n N_A_1586_149#_c_1303_n 0.010471f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_695 N_A_818_418#_c_840_n N_A_1586_149#_c_1303_n 0.0325809f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_696 N_A_818_418#_c_841_n N_A_1586_149#_c_1303_n 0.0100601f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_697 N_A_818_418#_M1005_g N_A_1586_149#_c_1296_n 0.00709662f $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_698 N_A_818_418#_c_836_n N_A_1586_149#_c_1296_n 0.0217185f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_699 N_A_818_418#_c_830_n N_A_1586_149#_c_1288_n 2.62577e-19 $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_700 N_A_818_418#_M1005_g N_A_1586_149#_c_1288_n 0.00810399f $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_701 N_A_818_418#_c_836_n N_A_1586_149#_c_1288_n 0.00843187f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_702 N_A_818_418#_c_840_n N_A_1586_149#_c_1288_n 0.0242956f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_703 N_A_818_418#_c_841_n N_A_1586_149#_c_1288_n 0.00983263f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_704 N_A_818_418#_M1005_g N_A_1586_149#_c_1298_n 0.0124997f $X=8.7 $Y=2.155
+ $X2=0 $Y2=0
cc_705 N_A_818_418#_c_836_n N_A_1586_149#_c_1298_n 0.0133994f $X=8.135 $Y=2.905
+ $X2=0 $Y2=0
cc_706 N_A_818_418#_c_840_n N_A_1586_149#_c_1298_n 0.00496924f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_707 N_A_818_418#_c_841_n N_A_1586_149#_c_1298_n 0.00381709f $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_708 N_A_818_418#_c_830_n N_A_1586_149#_c_1290_n 0.00560477f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_709 N_A_818_418#_c_847_n N_VPWR_M1034_d 0.0167442f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_710 N_A_818_418#_M1026_g N_VPWR_c_1484_n 8.82486e-19 $X=4.18 $Y=2.635 $X2=0
+ $Y2=0
cc_711 N_A_818_418#_c_846_n N_VPWR_c_1484_n 0.0158876f $X=5.62 $Y=2.815 $X2=0
+ $Y2=0
cc_712 N_A_818_418#_c_847_n N_VPWR_c_1484_n 0.00237224f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_713 N_A_818_418#_c_847_n N_VPWR_c_1497_n 0.0108267f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_714 N_A_818_418#_c_849_n N_VPWR_c_1497_n 0.046643f $X=8.05 $Y=2.99 $X2=0
+ $Y2=0
cc_715 N_A_818_418#_c_850_n N_VPWR_c_1497_n 0.013574f $X=7.505 $Y=2.99 $X2=0
+ $Y2=0
cc_716 N_A_818_418#_c_846_n N_VPWR_c_1501_n 0.0077782f $X=5.62 $Y=2.815 $X2=0
+ $Y2=0
cc_717 N_A_818_418#_c_847_n N_VPWR_c_1501_n 0.0396821f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_718 N_A_818_418#_M1005_g N_VPWR_c_1480_n 0.00461881f $X=8.7 $Y=2.155 $X2=0
+ $Y2=0
cc_719 N_A_818_418#_c_846_n N_VPWR_c_1480_n 0.0130823f $X=5.62 $Y=2.815 $X2=0
+ $Y2=0
cc_720 N_A_818_418#_c_847_n N_VPWR_c_1480_n 0.0273027f $X=7.315 $Y=2.51 $X2=0
+ $Y2=0
cc_721 N_A_818_418#_c_849_n N_VPWR_c_1480_n 0.0269839f $X=8.05 $Y=2.99 $X2=0
+ $Y2=0
cc_722 N_A_818_418#_c_850_n N_VPWR_c_1480_n 0.00737799f $X=7.505 $Y=2.99 $X2=0
+ $Y2=0
cc_723 N_A_818_418#_M1026_g N_A_70_74#_c_1643_n 0.013201f $X=4.18 $Y=2.635 $X2=0
+ $Y2=0
cc_724 N_A_818_418#_c_832_n N_A_70_74#_c_1643_n 4.87905e-19 $X=4.215 $Y=2.165
+ $X2=0 $Y2=0
cc_725 N_A_818_418#_M1032_g N_A_70_74#_c_1630_n 0.00741469f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_726 N_A_818_418#_M1026_g N_A_70_74#_c_1631_n 0.00397916f $X=4.18 $Y=2.635
+ $X2=0 $Y2=0
cc_727 N_A_818_418#_M1032_g N_A_70_74#_c_1631_n 0.0268581f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_728 N_A_818_418#_c_832_n N_A_70_74#_c_1631_n 0.00336914f $X=4.215 $Y=2.165
+ $X2=0 $Y2=0
cc_729 N_A_818_418#_c_833_n N_A_70_74#_c_1631_n 5.73127e-19 $X=4.81 $Y=2.075
+ $X2=0 $Y2=0
cc_730 N_A_818_418#_c_834_n N_A_70_74#_c_1631_n 0.0103062f $X=4.645 $Y=2.075
+ $X2=0 $Y2=0
cc_731 N_A_818_418#_c_835_n N_A_70_74#_c_1631_n 0.00560911f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_732 N_A_818_418#_c_837_n N_A_70_74#_c_1631_n 0.0256551f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_733 N_A_818_418#_c_839_n N_A_70_74#_c_1631_n 0.00236354f $X=5.62 $Y=2.005
+ $X2=0 $Y2=0
cc_734 N_A_818_418#_M1026_g N_A_70_74#_c_1646_n 0.0034344f $X=4.18 $Y=2.635
+ $X2=0 $Y2=0
cc_735 N_A_818_418#_c_832_n N_A_70_74#_c_1646_n 7.19263e-19 $X=4.215 $Y=2.165
+ $X2=0 $Y2=0
cc_736 N_A_818_418#_c_834_n N_A_70_74#_c_1647_n 0.0126159f $X=4.645 $Y=2.075
+ $X2=0 $Y2=0
cc_737 N_A_818_418#_c_846_n N_A_70_74#_c_1647_n 0.00966629f $X=5.62 $Y=2.815
+ $X2=0 $Y2=0
cc_738 N_A_818_418#_c_837_n N_A_70_74#_c_1647_n 0.0185116f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_739 N_A_818_418#_c_854_n N_A_70_74#_c_1647_n 0.00506182f $X=5.605 $Y=2.51
+ $X2=0 $Y2=0
cc_740 N_A_818_418#_c_830_n N_VGND_c_1856_n 8.63546e-19 $X=8.33 $Y=1.275 $X2=0
+ $Y2=0
cc_741 N_A_818_418#_M1032_g N_A_614_81#_c_1989_n 4.73936e-19 $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_742 N_A_818_418#_M1032_g N_A_614_81#_c_1990_n 0.00301077f $X=4.265 $Y=1.37
+ $X2=0 $Y2=0
cc_743 N_A_818_418#_c_833_n N_A_614_81#_c_1990_n 0.00492069f $X=4.81 $Y=2.075
+ $X2=0 $Y2=0
cc_744 N_A_818_418#_c_835_n N_A_614_81#_c_1990_n 0.0435989f $X=5.26 $Y=1.085
+ $X2=0 $Y2=0
cc_745 N_A_818_418#_c_837_n N_A_614_81#_c_1990_n 0.00853807f $X=5.15 $Y=2.075
+ $X2=0 $Y2=0
cc_746 N_A_818_418#_c_830_n N_A_1499_149#_c_2014_n 0.0127492f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_747 N_A_818_418#_c_841_n N_A_1499_149#_c_2014_n 5.41658e-19 $X=8.455 $Y=1.44
+ $X2=0 $Y2=0
cc_748 N_A_818_418#_c_830_n N_A_1499_149#_c_2016_n 0.00461776f $X=8.33 $Y=1.275
+ $X2=0 $Y2=0
cc_749 N_A_728_331#_c_993_n N_CLK_c_1149_n 0.0170252f $X=6.45 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_750 N_A_728_331#_c_996_n N_CLK_c_1149_n 0.0182609f $X=6.795 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_751 N_A_728_331#_M1034_g N_CLK_M1009_g 0.0224592f $X=5.845 $Y=2.4 $X2=0 $Y2=0
cc_752 N_A_728_331#_c_1002_n N_CLK_M1009_g 0.00313147f $X=6.18 $Y=1.84 $X2=0
+ $Y2=0
cc_753 N_A_728_331#_c_1027_n N_CLK_M1009_g 0.0154827f $X=6.705 $Y=2.047 $X2=0
+ $Y2=0
cc_754 N_A_728_331#_c_1006_n N_CLK_M1009_g 0.00586452f $X=7.035 $Y=2.047 $X2=0
+ $Y2=0
cc_755 N_A_728_331#_c_1007_n N_CLK_M1009_g 0.00863215f $X=7.34 $Y=1.795 $X2=0
+ $Y2=0
cc_756 N_A_728_331#_M1007_d CLK 0.00277495f $X=6.655 $Y=0.49 $X2=0 $Y2=0
cc_757 N_A_728_331#_c_993_n CLK 0.00994406f $X=6.45 $Y=1.34 $X2=0 $Y2=0
cc_758 N_A_728_331#_c_994_n CLK 2.34167e-19 $X=6.1 $Y=1.505 $X2=0 $Y2=0
cc_759 N_A_728_331#_c_995_n CLK 0.0259649f $X=6.45 $Y=1.505 $X2=0 $Y2=0
cc_760 N_A_728_331#_c_996_n CLK 0.0173596f $X=6.795 $Y=0.8 $X2=0 $Y2=0
cc_761 N_A_728_331#_c_1006_n CLK 0.0206329f $X=7.035 $Y=2.047 $X2=0 $Y2=0
cc_762 N_A_728_331#_c_994_n N_CLK_c_1151_n 0.0161568f $X=6.1 $Y=1.505 $X2=0
+ $Y2=0
cc_763 N_A_728_331#_c_995_n N_CLK_c_1151_n 0.00638468f $X=6.45 $Y=1.505 $X2=0
+ $Y2=0
cc_764 N_A_728_331#_c_996_n N_CLK_c_1151_n 0.00126242f $X=6.795 $Y=0.8 $X2=0
+ $Y2=0
cc_765 N_A_728_331#_c_1006_n N_CLK_c_1151_n 0.00158298f $X=7.035 $Y=2.047 $X2=0
+ $Y2=0
cc_766 N_A_728_331#_M1017_g N_A_1586_149#_c_1303_n 0.00269433f $X=7.855 $Y=0.955
+ $X2=0 $Y2=0
cc_767 N_A_728_331#_c_1001_n N_A_1586_149#_c_1303_n 0.00159115f $X=8.02 $Y=1.87
+ $X2=0 $Y2=0
cc_768 N_A_728_331#_c_1001_n N_A_1586_149#_c_1296_n 8.74828e-19 $X=8.02 $Y=1.87
+ $X2=0 $Y2=0
cc_769 N_A_728_331#_c_1001_n N_A_1586_149#_c_1298_n 5.63311e-19 $X=8.02 $Y=1.87
+ $X2=0 $Y2=0
cc_770 N_A_728_331#_c_1089_n N_VPWR_M1034_d 0.00889138f $X=6.265 $Y=2.005 $X2=0
+ $Y2=0
cc_771 N_A_728_331#_c_1027_n N_VPWR_M1034_d 0.00668832f $X=6.705 $Y=2.047 $X2=0
+ $Y2=0
cc_772 N_A_728_331#_M1024_g N_VPWR_c_1484_n 8.82486e-19 $X=3.73 $Y=2.635 $X2=0
+ $Y2=0
cc_773 N_A_728_331#_M1034_g N_VPWR_c_1484_n 0.00396012f $X=5.845 $Y=2.4 $X2=0
+ $Y2=0
cc_774 N_A_728_331#_c_1001_n N_VPWR_c_1497_n 0.00349658f $X=8.02 $Y=1.87 $X2=0
+ $Y2=0
cc_775 N_A_728_331#_M1034_g N_VPWR_c_1501_n 0.00556935f $X=5.845 $Y=2.4 $X2=0
+ $Y2=0
cc_776 N_A_728_331#_M1034_g N_VPWR_c_1480_n 0.00514497f $X=5.845 $Y=2.4 $X2=0
+ $Y2=0
cc_777 N_A_728_331#_c_1001_n N_VPWR_c_1480_n 0.00432848f $X=8.02 $Y=1.87 $X2=0
+ $Y2=0
cc_778 N_A_728_331#_M1024_g N_A_70_74#_c_1640_n 0.00137531f $X=3.73 $Y=2.635
+ $X2=0 $Y2=0
cc_779 N_A_728_331#_M1024_g N_A_70_74#_c_1642_n 0.00552805f $X=3.73 $Y=2.635
+ $X2=0 $Y2=0
cc_780 N_A_728_331#_M1024_g N_A_70_74#_c_1643_n 0.0125659f $X=3.73 $Y=2.635
+ $X2=0 $Y2=0
cc_781 N_A_728_331#_M1006_g N_A_70_74#_c_1630_n 0.0123257f $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_782 N_A_728_331#_c_992_n N_A_70_74#_c_1630_n 9.00795e-19 $X=3.775 $Y=1.805
+ $X2=0 $Y2=0
cc_783 N_A_728_331#_M1006_g N_A_70_74#_c_1631_n 7.75671e-19 $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_784 N_A_728_331#_M1006_g N_A_70_74#_c_1633_n 0.00370416f $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_785 N_A_728_331#_c_992_n N_A_70_74#_c_1633_n 0.00142161f $X=3.775 $Y=1.805
+ $X2=0 $Y2=0
cc_786 N_A_728_331#_c_993_n N_VGND_M1029_d 0.0103537f $X=6.45 $Y=1.34 $X2=0
+ $Y2=0
cc_787 N_A_728_331#_c_996_n N_VGND_M1029_d 0.00927667f $X=6.795 $Y=0.8 $X2=0
+ $Y2=0
cc_788 N_A_728_331#_c_988_n N_VGND_c_1845_n 0.00688197f $X=5.4 $Y=0.34 $X2=0
+ $Y2=0
cc_789 N_A_728_331#_c_988_n N_VGND_c_1854_n 0.00849616f $X=5.4 $Y=0.34 $X2=0
+ $Y2=0
cc_790 N_A_728_331#_c_989_n N_VGND_c_1854_n 0.0095216f $X=3.91 $Y=0.34 $X2=0
+ $Y2=0
cc_791 N_A_728_331#_c_988_n N_VGND_c_1867_n 0.0107407f $X=5.4 $Y=0.34 $X2=0
+ $Y2=0
cc_792 N_A_728_331#_M1006_g N_A_614_81#_c_1989_n 0.0139459f $X=3.835 $Y=1.37
+ $X2=0 $Y2=0
cc_793 N_A_728_331#_c_988_n N_A_614_81#_c_1989_n 0.00598631f $X=5.4 $Y=0.34
+ $X2=0 $Y2=0
cc_794 N_A_728_331#_M1029_g N_A_614_81#_c_1989_n 5.30126e-19 $X=5.475 $Y=0.86
+ $X2=0 $Y2=0
cc_795 N_A_728_331#_M1029_g N_A_614_81#_c_1990_n 0.00494998f $X=5.475 $Y=0.86
+ $X2=0 $Y2=0
cc_796 N_A_728_331#_c_999_n N_A_1499_149#_c_2013_n 2.85935e-19 $X=7.78 $Y=1.795
+ $X2=0 $Y2=0
cc_797 N_A_728_331#_M1017_g N_A_1499_149#_c_2013_n 0.0010439f $X=7.855 $Y=0.955
+ $X2=0 $Y2=0
cc_798 N_A_728_331#_M1017_g N_A_1499_149#_c_2014_n 0.0130579f $X=7.855 $Y=0.955
+ $X2=0 $Y2=0
cc_799 N_CLK_M1009_g N_VPWR_c_1497_n 0.00403892f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_800 N_CLK_M1009_g N_VPWR_c_1501_n 0.00596951f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_801 N_CLK_M1009_g N_VPWR_c_1480_n 0.00531308f $X=6.645 $Y=2.4 $X2=0 $Y2=0
cc_802 N_CLK_c_1149_n N_VGND_c_1845_n 2.58254e-19 $X=6.58 $Y=1.34 $X2=0 $Y2=0
cc_803 N_CLK_c_1149_n N_VGND_c_1856_n 7.26245e-19 $X=6.58 $Y=1.34 $X2=0 $Y2=0
cc_804 N_A_1800_291#_c_1195_n N_A_1586_149#_M1018_g 0.00518619f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_805 N_A_1800_291#_c_1196_n N_A_1586_149#_M1018_g 0.00799557f $X=10.59
+ $Y=0.557 $X2=0 $Y2=0
cc_806 N_A_1800_291#_c_1233_p N_A_1586_149#_M1019_g 0.0174444f $X=10.505
+ $Y=2.035 $X2=0 $Y2=0
cc_807 N_A_1800_291#_c_1195_n N_A_1586_149#_M1019_g 0.00533899f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_808 N_A_1800_291#_c_1202_n N_A_1586_149#_M1019_g 0.00832431f $X=10.16
+ $Y=2.167 $X2=0 $Y2=0
cc_809 N_A_1800_291#_c_1233_p N_A_1586_149#_M1030_g 0.00446702f $X=10.505
+ $Y=2.035 $X2=0 $Y2=0
cc_810 N_A_1800_291#_c_1195_n N_A_1586_149#_M1030_g 0.00706145f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_811 N_A_1800_291#_c_1202_n N_A_1586_149#_M1030_g 5.26076e-19 $X=10.16
+ $Y=2.167 $X2=0 $Y2=0
cc_812 N_A_1800_291#_c_1195_n N_A_1586_149#_c_1285_n 0.00115321f $X=10.59
+ $Y=1.95 $X2=0 $Y2=0
cc_813 N_A_1800_291#_M1014_g N_A_1586_149#_c_1296_n 0.0011673f $X=9.12 $Y=2.155
+ $X2=0 $Y2=0
cc_814 N_A_1800_291#_c_1229_n N_A_1586_149#_c_1296_n 9.30394e-19 $X=9.33
+ $Y=2.035 $X2=0 $Y2=0
cc_815 N_A_1800_291#_M1014_g N_A_1586_149#_c_1288_n 7.81006e-19 $X=9.12 $Y=2.155
+ $X2=0 $Y2=0
cc_816 N_A_1800_291#_c_1193_n N_A_1586_149#_c_1288_n 0.0338518f $X=9.165 $Y=1.62
+ $X2=0 $Y2=0
cc_817 N_A_1800_291#_c_1194_n N_A_1586_149#_c_1288_n 0.00180678f $X=9.165
+ $Y=1.62 $X2=0 $Y2=0
cc_818 N_A_1800_291#_c_1197_n N_A_1586_149#_c_1288_n 0.00374138f $X=9.165
+ $Y=1.455 $X2=0 $Y2=0
cc_819 N_A_1800_291#_c_1192_n N_A_1586_149#_c_1289_n 0.0167639f $X=9.365 $Y=0.94
+ $X2=0 $Y2=0
cc_820 N_A_1800_291#_c_1193_n N_A_1586_149#_c_1289_n 0.0181585f $X=9.165 $Y=1.62
+ $X2=0 $Y2=0
cc_821 N_A_1800_291#_c_1194_n N_A_1586_149#_c_1289_n 0.00346941f $X=9.165
+ $Y=1.62 $X2=0 $Y2=0
cc_822 N_A_1800_291#_c_1195_n N_A_1586_149#_c_1289_n 0.0259151f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_823 N_A_1800_291#_c_1196_n N_A_1586_149#_c_1289_n 0.00784134f $X=10.59
+ $Y=0.557 $X2=0 $Y2=0
cc_824 N_A_1800_291#_c_1197_n N_A_1586_149#_c_1289_n 0.01522f $X=9.165 $Y=1.455
+ $X2=0 $Y2=0
cc_825 N_A_1800_291#_M1014_g N_A_1586_149#_c_1298_n 0.00105096f $X=9.12 $Y=2.155
+ $X2=0 $Y2=0
cc_826 N_A_1800_291#_c_1193_n N_A_1586_149#_c_1298_n 0.00190034f $X=9.165
+ $Y=1.62 $X2=0 $Y2=0
cc_827 N_A_1800_291#_c_1229_n N_A_1586_149#_c_1298_n 0.0123059f $X=9.33 $Y=2.035
+ $X2=0 $Y2=0
cc_828 N_A_1800_291#_c_1233_p N_A_1586_149#_c_1291_n 0.00356911f $X=10.505
+ $Y=2.035 $X2=0 $Y2=0
cc_829 N_A_1800_291#_c_1195_n N_A_1586_149#_c_1291_n 0.0303375f $X=10.59 $Y=1.95
+ $X2=0 $Y2=0
cc_830 N_A_1800_291#_c_1196_n N_A_1586_149#_c_1291_n 0.00670663f $X=10.59
+ $Y=0.557 $X2=0 $Y2=0
cc_831 N_A_1800_291#_c_1229_n N_VPWR_M1014_d 6.8564e-19 $X=9.33 $Y=2.035 $X2=0
+ $Y2=0
cc_832 N_A_1800_291#_c_1216_n N_VPWR_M1014_d 0.00751611f $X=9.83 $Y=2.167 $X2=0
+ $Y2=0
cc_833 N_A_1800_291#_c_1233_p N_VPWR_M1019_d 0.00524314f $X=10.505 $Y=2.035
+ $X2=0 $Y2=0
cc_834 N_A_1800_291#_c_1195_n N_VPWR_M1019_d 0.00219613f $X=10.59 $Y=1.95 $X2=0
+ $Y2=0
cc_835 N_A_1800_291#_M1014_g N_VPWR_c_1485_n 0.00415305f $X=9.12 $Y=2.155 $X2=0
+ $Y2=0
cc_836 N_A_1800_291#_c_1194_n N_VPWR_c_1485_n 2.42318e-19 $X=9.165 $Y=1.62 $X2=0
+ $Y2=0
cc_837 N_A_1800_291#_c_1229_n N_VPWR_c_1485_n 0.00546648f $X=9.33 $Y=2.035 $X2=0
+ $Y2=0
cc_838 N_A_1800_291#_c_1216_n N_VPWR_c_1485_n 0.023051f $X=9.83 $Y=2.167 $X2=0
+ $Y2=0
cc_839 N_A_1800_291#_c_1202_n N_VPWR_c_1485_n 0.0037186f $X=10.16 $Y=2.167 $X2=0
+ $Y2=0
cc_840 N_A_1800_291#_c_1233_p N_VPWR_c_1486_n 0.0211944f $X=10.505 $Y=2.035
+ $X2=0 $Y2=0
cc_841 N_A_1800_291#_c_1202_n N_VPWR_c_1486_n 0.00370987f $X=10.16 $Y=2.167
+ $X2=0 $Y2=0
cc_842 N_A_1800_291#_M1014_g N_VPWR_c_1480_n 0.00461881f $X=9.12 $Y=2.155 $X2=0
+ $Y2=0
cc_843 N_A_1800_291#_c_1195_n N_Q_N_c_1785_n 0.0178706f $X=10.59 $Y=1.95 $X2=0
+ $Y2=0
cc_844 N_A_1800_291#_c_1195_n Q_N 0.0206203f $X=10.59 $Y=1.95 $X2=0 $Y2=0
cc_845 N_A_1800_291#_c_1191_n N_VGND_c_1846_n 0.00904236f $X=9.365 $Y=0.865
+ $X2=0 $Y2=0
cc_846 N_A_1800_291#_c_1196_n N_VGND_c_1846_n 0.0127168f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_847 N_A_1800_291#_c_1195_n N_VGND_c_1847_n 0.0247783f $X=10.59 $Y=1.95 $X2=0
+ $Y2=0
cc_848 N_A_1800_291#_c_1196_n N_VGND_c_1847_n 0.0333158f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_849 N_A_1800_291#_c_1191_n N_VGND_c_1856_n 0.00383152f $X=9.365 $Y=0.865
+ $X2=0 $Y2=0
cc_850 N_A_1800_291#_c_1196_n N_VGND_c_1858_n 0.0200848f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_851 N_A_1800_291#_c_1191_n N_VGND_c_1867_n 0.00762539f $X=9.365 $Y=0.865
+ $X2=0 $Y2=0
cc_852 N_A_1800_291#_c_1192_n N_VGND_c_1867_n 0.00141224f $X=9.365 $Y=0.94 $X2=0
+ $Y2=0
cc_853 N_A_1800_291#_c_1196_n N_VGND_c_1867_n 0.0169453f $X=10.59 $Y=0.557 $X2=0
+ $Y2=0
cc_854 N_A_1800_291#_c_1191_n N_A_1499_149#_c_2016_n 7.31217e-19 $X=9.365
+ $Y=0.865 $X2=0 $Y2=0
cc_855 N_A_1800_291#_c_1192_n N_A_1499_149#_c_2016_n 0.00244996f $X=9.365
+ $Y=0.94 $X2=0 $Y2=0
cc_856 N_A_1586_149#_M1020_g N_A_2366_352#_c_1423_n 0.00959603f $X=11.74 $Y=2.26
+ $X2=0 $Y2=0
cc_857 N_A_1586_149#_c_1291_n N_A_2366_352#_c_1423_n 0.0183752f $X=11.74
+ $Y=1.267 $X2=0 $Y2=0
cc_858 N_A_1586_149#_M1020_g N_A_2366_352#_c_1430_n 0.0211078f $X=11.74 $Y=2.26
+ $X2=0 $Y2=0
cc_859 N_A_1586_149#_M1022_g N_A_2366_352#_c_1424_n 0.00874126f $X=12.05 $Y=0.69
+ $X2=0 $Y2=0
cc_860 N_A_1586_149#_c_1291_n N_A_2366_352#_c_1426_n 0.0054628f $X=11.74
+ $Y=1.267 $X2=0 $Y2=0
cc_861 N_A_1586_149#_c_1296_n N_VPWR_c_1485_n 0.00147567f $X=8.475 $Y=2.155
+ $X2=0 $Y2=0
cc_862 N_A_1586_149#_M1019_g N_VPWR_c_1486_n 0.0037152f $X=10.22 $Y=2.155 $X2=0
+ $Y2=0
cc_863 N_A_1586_149#_M1030_g N_VPWR_c_1486_n 0.0136841f $X=10.755 $Y=2.32 $X2=0
+ $Y2=0
cc_864 N_A_1586_149#_M1035_g N_VPWR_c_1486_n 5.14339e-19 $X=11.205 $Y=2.32 $X2=0
+ $Y2=0
cc_865 N_A_1586_149#_c_1291_n N_VPWR_c_1486_n 3.38899e-19 $X=11.74 $Y=1.267
+ $X2=0 $Y2=0
cc_866 N_A_1586_149#_M1030_g N_VPWR_c_1487_n 0.00519349f $X=10.755 $Y=2.32 $X2=0
+ $Y2=0
cc_867 N_A_1586_149#_M1035_g N_VPWR_c_1487_n 0.00519349f $X=11.205 $Y=2.32 $X2=0
+ $Y2=0
cc_868 N_A_1586_149#_M1030_g N_VPWR_c_1488_n 6.8825e-19 $X=10.755 $Y=2.32 $X2=0
+ $Y2=0
cc_869 N_A_1586_149#_M1035_g N_VPWR_c_1488_n 0.0205757f $X=11.205 $Y=2.32 $X2=0
+ $Y2=0
cc_870 N_A_1586_149#_M1020_g N_VPWR_c_1488_n 0.00892026f $X=11.74 $Y=2.26 $X2=0
+ $Y2=0
cc_871 N_A_1586_149#_c_1291_n N_VPWR_c_1488_n 0.00495468f $X=11.74 $Y=1.267
+ $X2=0 $Y2=0
cc_872 N_A_1586_149#_M1020_g N_VPWR_c_1489_n 0.00359304f $X=11.74 $Y=2.26 $X2=0
+ $Y2=0
cc_873 N_A_1586_149#_M1020_g N_VPWR_c_1498_n 0.00534617f $X=11.74 $Y=2.26 $X2=0
+ $Y2=0
cc_874 N_A_1586_149#_M1019_g N_VPWR_c_1480_n 0.00461881f $X=10.22 $Y=2.155 $X2=0
+ $Y2=0
cc_875 N_A_1586_149#_M1030_g N_VPWR_c_1480_n 0.00524044f $X=10.755 $Y=2.32 $X2=0
+ $Y2=0
cc_876 N_A_1586_149#_M1035_g N_VPWR_c_1480_n 0.00524044f $X=11.205 $Y=2.32 $X2=0
+ $Y2=0
cc_877 N_A_1586_149#_M1020_g N_VPWR_c_1480_n 0.00581878f $X=11.74 $Y=2.26 $X2=0
+ $Y2=0
cc_878 N_A_1586_149#_c_1298_n A_1758_389# 0.00310111f $X=8.81 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_879 N_A_1586_149#_M1030_g N_Q_N_c_1785_n 0.00148016f $X=10.755 $Y=2.32 $X2=0
+ $Y2=0
cc_880 N_A_1586_149#_M1035_g N_Q_N_c_1785_n 0.00374516f $X=11.205 $Y=2.32 $X2=0
+ $Y2=0
cc_881 N_A_1586_149#_c_1291_n N_Q_N_c_1785_n 0.0067137f $X=11.74 $Y=1.267 $X2=0
+ $Y2=0
cc_882 N_A_1586_149#_c_1285_n N_Q_N_c_1783_n 0.00521369f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_883 N_A_1586_149#_c_1286_n N_Q_N_c_1783_n 2.74318e-19 $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_884 N_A_1586_149#_c_1285_n Q_N 0.00609559f $X=11.145 $Y=1.185 $X2=0 $Y2=0
cc_885 N_A_1586_149#_c_1286_n Q_N 0.0143409f $X=11.575 $Y=1.185 $X2=0 $Y2=0
cc_886 N_A_1586_149#_M1022_g Q_N 0.00393154f $X=12.05 $Y=0.69 $X2=0 $Y2=0
cc_887 N_A_1586_149#_c_1291_n Q_N 0.0829724f $X=11.74 $Y=1.267 $X2=0 $Y2=0
cc_888 N_A_1586_149#_M1018_g N_VGND_c_1846_n 0.00157764f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_889 N_A_1586_149#_c_1289_n N_VGND_c_1846_n 0.0192815f $X=10.245 $Y=1.1 $X2=0
+ $Y2=0
cc_890 N_A_1586_149#_M1018_g N_VGND_c_1847_n 0.00300622f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_891 N_A_1586_149#_c_1285_n N_VGND_c_1847_n 0.00400592f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_892 N_A_1586_149#_c_1291_n N_VGND_c_1847_n 0.00510356f $X=11.74 $Y=1.267
+ $X2=0 $Y2=0
cc_893 N_A_1586_149#_c_1285_n N_VGND_c_1848_n 4.16356e-19 $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_894 N_A_1586_149#_c_1286_n N_VGND_c_1848_n 0.00689813f $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_895 N_A_1586_149#_M1022_g N_VGND_c_1848_n 0.00197289f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_896 N_A_1586_149#_c_1291_n N_VGND_c_1848_n 7.47495e-19 $X=11.74 $Y=1.267
+ $X2=0 $Y2=0
cc_897 N_A_1586_149#_M1022_g N_VGND_c_1849_n 0.00293008f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_898 N_A_1586_149#_M1018_g N_VGND_c_1858_n 0.00433162f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_899 N_A_1586_149#_c_1285_n N_VGND_c_1861_n 0.00434272f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_900 N_A_1586_149#_c_1286_n N_VGND_c_1861_n 0.00383152f $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_901 N_A_1586_149#_M1022_g N_VGND_c_1862_n 0.00461464f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_902 N_A_1586_149#_M1018_g N_VGND_c_1867_n 0.00822018f $X=10.155 $Y=0.58 $X2=0
+ $Y2=0
cc_903 N_A_1586_149#_c_1285_n N_VGND_c_1867_n 0.00825283f $X=11.145 $Y=1.185
+ $X2=0 $Y2=0
cc_904 N_A_1586_149#_c_1286_n N_VGND_c_1867_n 0.0036906f $X=11.575 $Y=1.185
+ $X2=0 $Y2=0
cc_905 N_A_1586_149#_M1022_g N_VGND_c_1867_n 0.00912757f $X=12.05 $Y=0.69 $X2=0
+ $Y2=0
cc_906 N_A_1586_149#_M1017_d N_A_1499_149#_c_2014_n 0.0042087f $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_907 N_A_1586_149#_c_1303_n N_A_1499_149#_c_2014_n 0.0461856f $X=8.725 $Y=1.02
+ $X2=0 $Y2=0
cc_908 N_A_1586_149#_c_1289_n N_A_1499_149#_c_2014_n 0.00709406f $X=10.245
+ $Y=1.1 $X2=0 $Y2=0
cc_909 N_A_1586_149#_c_1290_n N_A_1499_149#_c_2014_n 0.0142962f $X=8.81 $Y=1.1
+ $X2=0 $Y2=0
cc_910 N_A_1586_149#_c_1289_n N_A_1499_149#_c_2016_n 0.0203727f $X=10.245 $Y=1.1
+ $X2=0 $Y2=0
cc_911 N_A_2366_352#_c_1423_n N_VPWR_c_1488_n 0.00617394f $X=12.1 $Y=1.945 $X2=0
+ $Y2=0
cc_912 N_A_2366_352#_c_1430_n N_VPWR_c_1488_n 0.0233044f $X=12.06 $Y=2.615 $X2=0
+ $Y2=0
cc_913 N_A_2366_352#_M1000_g N_VPWR_c_1489_n 0.00546761f $X=12.915 $Y=2.4 $X2=0
+ $Y2=0
cc_914 N_A_2366_352#_c_1423_n N_VPWR_c_1489_n 0.0106305f $X=12.1 $Y=1.945 $X2=0
+ $Y2=0
cc_915 N_A_2366_352#_c_1430_n N_VPWR_c_1489_n 0.0706466f $X=12.06 $Y=2.615 $X2=0
+ $Y2=0
cc_916 N_A_2366_352#_c_1425_n N_VPWR_c_1489_n 0.0261101f $X=12.8 $Y=1.465 $X2=0
+ $Y2=0
cc_917 N_A_2366_352#_c_1426_n N_VPWR_c_1489_n 0.00389761f $X=13.365 $Y=1.465
+ $X2=0 $Y2=0
cc_918 N_A_2366_352#_M1003_g N_VPWR_c_1491_n 0.00546761f $X=13.365 $Y=2.4 $X2=0
+ $Y2=0
cc_919 N_A_2366_352#_c_1426_n N_VPWR_c_1491_n 0.00152598f $X=13.365 $Y=1.465
+ $X2=0 $Y2=0
cc_920 N_A_2366_352#_c_1430_n N_VPWR_c_1498_n 0.00996859f $X=12.06 $Y=2.615
+ $X2=0 $Y2=0
cc_921 N_A_2366_352#_M1000_g N_VPWR_c_1499_n 0.005209f $X=12.915 $Y=2.4 $X2=0
+ $Y2=0
cc_922 N_A_2366_352#_M1003_g N_VPWR_c_1499_n 0.005209f $X=13.365 $Y=2.4 $X2=0
+ $Y2=0
cc_923 N_A_2366_352#_M1000_g N_VPWR_c_1480_n 0.00986727f $X=12.915 $Y=2.4 $X2=0
+ $Y2=0
cc_924 N_A_2366_352#_M1003_g N_VPWR_c_1480_n 0.00985497f $X=13.365 $Y=2.4 $X2=0
+ $Y2=0
cc_925 N_A_2366_352#_c_1430_n N_VPWR_c_1480_n 0.0131729f $X=12.06 $Y=2.615 $X2=0
+ $Y2=0
cc_926 N_A_2366_352#_c_1423_n Q_N 0.0130882f $X=12.1 $Y=1.945 $X2=0 $Y2=0
cc_927 N_A_2366_352#_c_1424_n Q_N 0.0259548f $X=12.265 $Y=0.515 $X2=0 $Y2=0
cc_928 N_A_2366_352#_M1000_g N_Q_c_1815_n 0.0036649f $X=12.915 $Y=2.4 $X2=0
+ $Y2=0
cc_929 N_A_2366_352#_M1003_g N_Q_c_1815_n 0.00215936f $X=13.365 $Y=2.4 $X2=0
+ $Y2=0
cc_930 N_A_2366_352#_c_1426_n N_Q_c_1815_n 0.0018941f $X=13.365 $Y=1.465 $X2=0
+ $Y2=0
cc_931 N_A_2366_352#_M1000_g N_Q_c_1816_n 0.0127634f $X=12.915 $Y=2.4 $X2=0
+ $Y2=0
cc_932 N_A_2366_352#_M1003_g N_Q_c_1816_n 0.0127634f $X=13.365 $Y=2.4 $X2=0
+ $Y2=0
cc_933 N_A_2366_352#_M1000_g N_Q_c_1812_n 0.00411176f $X=12.915 $Y=2.4 $X2=0
+ $Y2=0
cc_934 N_A_2366_352#_M1001_g N_Q_c_1812_n 0.00405899f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_935 N_A_2366_352#_M1003_g N_Q_c_1812_n 0.00903338f $X=13.365 $Y=2.4 $X2=0
+ $Y2=0
cc_936 N_A_2366_352#_M1016_g N_Q_c_1812_n 0.0040077f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_937 N_A_2366_352#_c_1425_n N_Q_c_1812_n 0.0249855f $X=12.8 $Y=1.465 $X2=0
+ $Y2=0
cc_938 N_A_2366_352#_c_1426_n N_Q_c_1812_n 0.0262103f $X=13.365 $Y=1.465 $X2=0
+ $Y2=0
cc_939 N_A_2366_352#_M1001_g Q 0.00327512f $X=13.01 $Y=0.74 $X2=0 $Y2=0
cc_940 N_A_2366_352#_M1016_g Q 0.00323247f $X=13.44 $Y=0.74 $X2=0 $Y2=0
cc_941 N_A_2366_352#_M1001_g N_Q_c_1814_n 0.00838251f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_942 N_A_2366_352#_M1016_g N_Q_c_1814_n 0.00821863f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_943 N_A_2366_352#_c_1424_n N_VGND_c_1848_n 0.00157123f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_944 N_A_2366_352#_M1001_g N_VGND_c_1849_n 0.00610844f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_945 N_A_2366_352#_c_1424_n N_VGND_c_1849_n 0.0562664f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_946 N_A_2366_352#_c_1425_n N_VGND_c_1849_n 0.0209312f $X=12.8 $Y=1.465 $X2=0
+ $Y2=0
cc_947 N_A_2366_352#_c_1426_n N_VGND_c_1849_n 0.00589713f $X=13.365 $Y=1.465
+ $X2=0 $Y2=0
cc_948 N_A_2366_352#_M1016_g N_VGND_c_1851_n 0.00618831f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_949 N_A_2366_352#_c_1424_n N_VGND_c_1862_n 0.0130739f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_950 N_A_2366_352#_M1001_g N_VGND_c_1863_n 0.00433834f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_951 N_A_2366_352#_M1016_g N_VGND_c_1863_n 0.00433834f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_952 N_A_2366_352#_M1001_g N_VGND_c_1867_n 0.00824977f $X=13.01 $Y=0.74 $X2=0
+ $Y2=0
cc_953 N_A_2366_352#_M1016_g N_VGND_c_1867_n 0.00823359f $X=13.44 $Y=0.74 $X2=0
+ $Y2=0
cc_954 N_A_2366_352#_c_1424_n N_VGND_c_1867_n 0.0108215f $X=12.265 $Y=0.515
+ $X2=0 $Y2=0
cc_955 N_VPWR_c_1482_n N_A_70_74#_c_1634_n 0.036541f $X=0.345 $Y=2.17 $X2=0
+ $Y2=0
cc_956 N_VPWR_M1004_d N_A_70_74#_c_1636_n 0.00994687f $X=0.135 $Y=2.81 $X2=0
+ $Y2=0
cc_957 N_VPWR_c_1492_n N_A_70_74#_c_1636_n 0.0312655f $X=1.21 $Y=3.19 $X2=0
+ $Y2=0
cc_958 N_VPWR_c_1496_n N_A_70_74#_c_1636_n 0.0030955f $X=2.945 $Y=3.33 $X2=0
+ $Y2=0
cc_959 N_VPWR_c_1480_n N_A_70_74#_c_1636_n 0.00699554f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_960 N_VPWR_c_1482_n N_A_70_74#_c_1637_n 0.0152343f $X=0.345 $Y=2.17 $X2=0
+ $Y2=0
cc_961 N_VPWR_c_1492_n N_A_70_74#_c_1637_n 0.0271618f $X=1.21 $Y=3.19 $X2=0
+ $Y2=0
cc_962 N_VPWR_c_1480_n N_A_70_74#_c_1637_n 0.00204634f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_963 N_VPWR_c_1483_n N_A_70_74#_c_1638_n 0.0147094f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_964 N_VPWR_c_1496_n N_A_70_74#_c_1638_n 0.0656248f $X=2.945 $Y=3.33 $X2=0
+ $Y2=0
cc_965 N_VPWR_c_1480_n N_A_70_74#_c_1638_n 0.0378114f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_966 N_VPWR_M1011_d N_A_70_74#_c_1639_n 0.00463987f $X=2.665 $Y=2.425 $X2=0
+ $Y2=0
cc_967 N_VPWR_c_1483_n N_A_70_74#_c_1639_n 0.0209842f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_968 N_VPWR_M1011_d N_A_70_74#_c_1640_n 0.00947326f $X=2.665 $Y=2.425 $X2=0
+ $Y2=0
cc_969 N_VPWR_c_1483_n N_A_70_74#_c_1640_n 0.0200956f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_970 N_VPWR_c_1483_n N_A_70_74#_c_1642_n 0.0118091f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_971 N_VPWR_c_1484_n N_A_70_74#_c_1643_n 0.0485775f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_972 N_VPWR_c_1480_n N_A_70_74#_c_1643_n 0.0283783f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_973 N_VPWR_c_1483_n N_A_70_74#_c_1644_n 0.0144269f $X=3.03 $Y=2.79 $X2=0
+ $Y2=0
cc_974 N_VPWR_c_1484_n N_A_70_74#_c_1644_n 0.0121867f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_975 N_VPWR_c_1480_n N_A_70_74#_c_1644_n 0.00660921f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_976 N_VPWR_c_1484_n N_A_70_74#_c_1646_n 0.0125688f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_977 N_VPWR_c_1480_n N_A_70_74#_c_1646_n 0.00710542f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_978 N_VPWR_c_1484_n N_A_70_74#_c_1647_n 0.0118092f $X=5.99 $Y=3.33 $X2=0
+ $Y2=0
cc_979 N_VPWR_c_1480_n N_A_70_74#_c_1647_n 0.0155687f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_980 N_VPWR_c_1482_n N_A_70_74#_c_1632_n 7.16831e-19 $X=0.345 $Y=2.17 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1493_n N_A_70_74#_c_1649_n 0.00879319f $X=1.435 $Y=3.19 $X2=0
+ $Y2=0
cc_982 N_VPWR_c_1496_n N_A_70_74#_c_1649_n 0.0114644f $X=2.945 $Y=3.33 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1480_n N_A_70_74#_c_1649_n 0.00617045f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_984 N_VPWR_c_1486_n N_Q_N_c_1785_n 0.0207342f $X=10.53 $Y=2.375 $X2=0 $Y2=0
cc_985 N_VPWR_c_1487_n N_Q_N_c_1785_n 0.0056634f $X=11.265 $Y=3.33 $X2=0 $Y2=0
cc_986 N_VPWR_c_1488_n N_Q_N_c_1785_n 0.0394917f $X=11.43 $Y=1.905 $X2=0 $Y2=0
cc_987 N_VPWR_c_1480_n N_Q_N_c_1785_n 0.00589694f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_988 N_VPWR_c_1488_n Q_N 0.0257228f $X=11.43 $Y=1.905 $X2=0 $Y2=0
cc_989 N_VPWR_c_1489_n N_Q_c_1815_n 0.0450694f $X=12.64 $Y=1.985 $X2=0 $Y2=0
cc_990 N_VPWR_c_1491_n N_Q_c_1815_n 0.0450694f $X=13.64 $Y=1.985 $X2=0 $Y2=0
cc_991 N_VPWR_c_1499_n N_Q_c_1816_n 0.0144623f $X=13.475 $Y=3.33 $X2=0 $Y2=0
cc_992 N_VPWR_c_1480_n N_Q_c_1816_n 0.0118344f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_993 N_A_70_74#_c_1640_n A_686_485# 3.01779e-19 $X=3.365 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_994 N_A_70_74#_c_1642_n A_686_485# 0.00392104f $X=3.45 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_995 N_A_70_74#_c_1629_n A_156_74# 0.00286631f $X=0.685 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_996 N_A_70_74#_c_1632_n A_156_74# 0.00153008f $X=0.845 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_997 N_A_70_74#_c_1632_n N_VGND_c_1843_n 0.00990285f $X=0.845 $Y=1.95 $X2=0
+ $Y2=0
cc_998 N_A_70_74#_c_1629_n N_VGND_c_1860_n 0.0167633f $X=0.685 $Y=0.515 $X2=0
+ $Y2=0
cc_999 N_A_70_74#_c_1629_n N_VGND_c_1867_n 0.0179018f $X=0.685 $Y=0.515 $X2=0
+ $Y2=0
cc_1000 N_A_70_74#_c_1631_n N_A_614_81#_M1032_d 0.00447556f $X=4.39 $Y=2.41
+ $X2=0 $Y2=0
cc_1001 N_A_70_74#_c_1630_n N_A_614_81#_c_1989_n 0.0576187f $X=4.305 $Y=1.02
+ $X2=0 $Y2=0
cc_1002 N_A_70_74#_c_1633_n N_A_614_81#_c_1989_n 0.0300095f $X=3.53 $Y=1.02
+ $X2=0 $Y2=0
cc_1003 N_A_70_74#_c_1630_n N_A_614_81#_c_1990_n 0.0147455f $X=4.305 $Y=1.02
+ $X2=0 $Y2=0
cc_1004 N_A_70_74#_c_1631_n N_A_614_81#_c_1990_n 0.0371597f $X=4.39 $Y=2.41
+ $X2=0 $Y2=0
cc_1005 Q_N N_VGND_M1033_d 0.00584895f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1006 N_Q_N_c_1783_n N_VGND_c_1847_n 0.0151654f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1007 Q_N N_VGND_c_1847_n 0.00847611f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1008 N_Q_N_c_1783_n N_VGND_c_1848_n 0.010186f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1009 Q_N N_VGND_c_1848_n 0.0165497f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1010 N_Q_N_c_1783_n N_VGND_c_1861_n 0.0114405f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1011 N_Q_N_c_1783_n N_VGND_c_1867_n 0.00941304f $X=11.36 $Y=0.515 $X2=0 $Y2=0
cc_1012 Q_N N_VGND_c_1867_n 0.00714657f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1013 N_Q_c_1814_n N_VGND_c_1849_n 0.0308594f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1014 N_Q_c_1814_n N_VGND_c_1851_n 0.0323079f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1015 N_Q_c_1814_n N_VGND_c_1863_n 0.0157615f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1016 N_Q_c_1814_n N_VGND_c_1867_n 0.0120285f $X=13.225 $Y=0.495 $X2=0 $Y2=0
cc_1017 N_VGND_c_1856_n N_A_1499_149#_c_2014_n 0.0040788f $X=9.415 $Y=0 $X2=0
+ $Y2=0
cc_1018 N_VGND_c_1867_n N_A_1499_149#_c_2014_n 0.00820175f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1019 N_VGND_c_1846_n N_A_1499_149#_c_2016_n 0.0139893f $X=9.58 $Y=0.555 $X2=0
+ $Y2=0
cc_1020 N_VGND_c_1856_n N_A_1499_149#_c_2016_n 0.0106808f $X=9.415 $Y=0 $X2=0
+ $Y2=0
cc_1021 N_VGND_c_1867_n N_A_1499_149#_c_2016_n 0.00901185f $X=13.68 $Y=0 $X2=0
+ $Y2=0

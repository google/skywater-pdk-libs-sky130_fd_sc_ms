* File: sky130_fd_sc_ms__o311a_2.spice
* Created: Wed Sep  2 12:24:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o311a_2.pex.spice"
.subckt sky130_fd_sc_ms__o311a_2  VNB VPB C1 B1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1001 A_135_74# N_C1_M1001_g N_A_32_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0999 AS=0.2701 PD=1.01 PS=2.21 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1013 N_A_219_74#_M1013_d N_B1_M1013_g A_135_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0999 PD=1.13 PS=1.01 NRD=17.832 NRS=12.972 M=1 R=4.93333
+ SA=75000.7 SB=75003 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A3_M1002_g N_A_219_74#_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2487 AS=0.1443 PD=1.49 PS=1.13 NRD=45.576 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1000 N_A_219_74#_M1000_d N_A2_M1000_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2487 PD=1.02 PS=1.49 NRD=0 NRS=45.576 M=1 R=4.93333 SA=75002
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_219_74#_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.16465 AS=0.1036 PD=1.185 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_A_32_74#_M1005_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.16465 PD=1.02 PS=1.185 NRD=0 NRS=15.396 M=1 R=4.93333 SA=75003
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1005_d N_A_32_74#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2775 PD=1.02 PS=2.23 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75003.4
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_C1_M1007_g N_A_32_74#_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.28 PD=1.39 PS=2.56 NRD=18.715 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1006 N_A_32_74#_M1006_d N_B1_M1006_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1
+ AD=0.18566 AS=0.195 PD=1.39623 PS=1.39 NRD=17.0602 NRS=2.9353 M=1 R=5.55556
+ SA=90000.8 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1010 A_363_368# N_A3_M1010_g N_A_32_74#_M1006_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1344 AS=0.20794 PD=1.36 PS=1.56377 NRD=11.426 NRS=0 M=1 R=6.22222
+ SA=90001.2 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1003 A_447_368# N_A2_M1003_g A_363_368# VPB PSHORT L=0.18 W=1.12 AD=0.2016
+ AS=0.1344 PD=1.48 PS=1.36 NRD=21.9852 NRS=11.426 M=1 R=6.22222 SA=90001.6
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_447_368# VPB PSHORT L=0.18 W=1.12 AD=0.2268
+ AS=0.2016 PD=1.525 PS=1.48 NRD=0 NRS=21.9852 M=1 R=6.22222 SA=90002.1
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1011_d N_A_32_74#_M1011_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2268 PD=1.39 PS=1.525 NRD=0 NRS=22.852 M=1 R=6.22222 SA=90002.7
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1011_d N_A_32_74#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__o311a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o221a_2.pex.spice
* Created: Wed Sep  2 12:22:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O221A_2%C1 3 5 7 8 15
r29 14 15 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=0.505 $Y=1.385
+ $X2=0.75 $Y2=1.385
r30 11 14 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.385
+ $X2=0.505 $Y2=1.385
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r32 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r33 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.75 $Y=1.22
+ $X2=0.75 $Y2=1.385
r34 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.75 $Y=1.22 $X2=0.75
+ $Y2=0.74
r35 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.385
r36 1 3 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%B1 3 5 7 8 12 13
c40 3 0 5.3557e-20 $X=1.245 $Y=0.74
r41 11 13 2.6679 $w=2.71e-07 $l=1.5e-08 $layer=POLY_cond $X=1.23 $Y=1.537
+ $X2=1.245 $Y2=1.537
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.515 $X2=1.23 $Y2=1.515
r43 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=1.515
r44 5 13 60.4723 $w=2.71e-07 $l=4.23698e-07 $layer=POLY_cond $X=1.585 $Y=1.725
+ $X2=1.245 $Y2=1.537
r45 5 7 164.683 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=1.585 $Y=1.725
+ $X2=1.585 $Y2=2.34
r46 1 13 16.5906 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.245 $Y=1.35
+ $X2=1.245 $Y2=1.537
r47 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.245 $Y=1.35
+ $X2=1.245 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%B2 1 3 4 8 14 15 19 21
c41 8 0 9.70842e-20 $X=2.005 $Y=2.34
c42 1 0 1.67816e-19 $X=1.75 $Y=1.185
r43 19 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.515
+ $X2=2.08 $Y2=1.68
r44 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.515 $X2=2.08 $Y2=1.515
r45 15 20 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.08
+ $Y2=1.565
r46 14 20 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=2.08
+ $Y2=1.565
r47 8 21 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.005 $Y=2.34
+ $X2=2.005 $Y2=1.68
r48 4 10 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.08 $Y=1.26 $X2=1.75
+ $Y2=1.26
r49 4 19 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.08 $Y=1.335 $X2=2.08
+ $Y2=1.515
r50 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.185
+ $X2=1.75 $Y2=1.26
r51 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.75 $Y=1.185
+ $X2=1.75 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%A2 3 7 9 12 13
c34 13 0 9.70842e-20 $X=2.65 $Y=1.515
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.515
+ $X2=2.65 $Y2=1.68
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.515
+ $X2=2.65 $Y2=1.35
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.515 $X2=2.65 $Y2=1.515
r38 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=1.515
r39 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.74 $Y=0.74 $X2=2.74
+ $Y2=1.35
r40 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.575 $Y=2.34
+ $X2=2.575 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%A1 3 7 9 12 13
c43 3 0 1.17819e-19 $X=3.145 $Y=2.34
r44 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.515
+ $X2=3.22 $Y2=1.68
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.515
+ $X2=3.22 $Y2=1.35
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.515 $X2=3.22 $Y2=1.515
r47 9 13 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=3.195 $Y=1.665
+ $X2=3.195 $Y2=1.515
r48 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.17 $Y=0.74 $X2=3.17
+ $Y2=1.35
r49 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.145 $Y=2.34
+ $X2=3.145 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%A_27_368# 1 2 3 12 16 18 22 26 28 31 35 38
+ 39 43 45 48 53 54 56 60 63
r118 63 64 31.0318 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.395
+ $X2=3.765 $Y2=1.32
r119 61 66 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.485
+ $X2=3.765 $Y2=1.65
r120 61 63 15.2746 $w=3.4e-07 $l=9e-08 $layer=POLY_cond $X=3.765 $Y=1.485
+ $X2=3.765 $Y2=1.395
r121 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.485 $X2=3.76 $Y2=1.485
r122 57 60 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.65 $Y=1.485
+ $X2=3.76 $Y2=1.485
r123 52 53 5.41145 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.97
+ $X2=0.775 $Y2=1.97
r124 50 52 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.97
+ $X2=0.69 $Y2=1.97
r125 47 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.65 $Y=1.65
+ $X2=3.65 $Y2=1.485
r126 47 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.65 $Y=1.65 $X2=3.65
+ $Y2=1.95
r127 46 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.035
+ $X2=2.23 $Y2=2.035
r128 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.565 $Y=2.035
+ $X2=3.65 $Y2=1.95
r129 45 46 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.565 $Y=2.035
+ $X2=2.395 $Y2=2.035
r130 41 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.035
r131 41 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.375
r132 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=2.035
+ $X2=2.23 $Y2=2.035
r133 39 53 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.065 $Y=2.035
+ $X2=0.775 $Y2=2.035
r134 38 52 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=1.82 $X2=0.69
+ $Y2=1.97
r135 38 54 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.69 $Y=1.82
+ $X2=0.69 $Y2=1.01
r136 33 54 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=0.572 $Y=0.808
+ $X2=0.572 $Y2=1.01
r137 33 35 8.33743 $w=4.03e-07 $l=2.93e-07 $layer=LI1_cond $X=0.572 $Y=0.808
+ $X2=0.572 $Y2=0.515
r138 29 50 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=1.97
r139 29 31 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.695
r140 24 28 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=4.295 $Y=1.47
+ $X2=4.24 $Y2=1.395
r141 24 26 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=4.295 $Y=1.47
+ $X2=4.295 $Y2=2.4
r142 20 28 18.8402 $w=1.65e-07 $l=1.04283e-07 $layer=POLY_cond $X=4.17 $Y=1.32
+ $X2=4.24 $Y2=1.395
r143 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.17 $Y=1.32
+ $X2=4.17 $Y2=0.74
r144 19 63 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.935 $Y=1.395
+ $X2=3.765 $Y2=1.395
r145 18 28 6.66866 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.095 $Y=1.395
+ $X2=4.24 $Y2=1.395
r146 18 19 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.095 $Y=1.395
+ $X2=3.935 $Y2=1.395
r147 16 66 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.845 $Y=2.4
+ $X2=3.845 $Y2=1.65
r148 12 64 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.74 $Y=0.74
+ $X2=3.74 $Y2=1.32
r149 3 56 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.84 $X2=2.23 $Y2=2.035
r150 3 43 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.84 $X2=2.23 $Y2=2.375
r151 2 50 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r152 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.695
r153 1 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.39
+ $Y=0.37 $X2=0.535 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%VPWR 1 2 3 12 16 20 22 26 28 33 41 47 50 54
r48 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r52 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 42 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=3.33
+ $X2=3.57 $Y2=3.33
r55 42 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 41 53 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.617 $Y2=3.33
r57 41 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 36 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 34 47 15.5867 $w=1.7e-07 $l=4.55e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.07 $Y2=3.33
r64 34 36 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.57 $Y2=3.33
r66 33 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 31 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 28 47 15.5867 $w=1.7e-07 $l=4.55e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.07 $Y2=3.33
r70 28 30 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 26 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 26 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 22 25 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.56 $Y=1.985
+ $X2=4.56 $Y2=2.815
r74 20 53 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.617 $Y2=3.33
r75 20 25 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.56 $Y2=2.815
r76 16 19 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.57 $Y=2.455
+ $X2=3.57 $Y2=2.815
r77 14 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=3.33
r78 14 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.815
r79 10 47 3.36946 $w=9.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r80 10 12 11.6637 $w=9.08e-07 $l=8.7e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.375
r81 3 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.815
r82 3 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=1.985
r83 2 19 600 $w=1.7e-07 $l=1.13015e-06 $layer=licon1_PDIFF $count=1 $X=3.235
+ $Y=1.84 $X2=3.57 $Y2=2.815
r84 2 16 600 $w=1.7e-07 $l=7.64362e-07 $layer=licon1_PDIFF $count=1 $X=3.235
+ $Y=1.84 $X2=3.57 $Y2=2.455
r85 1 12 150 $w=1.7e-07 $l=9.97246e-07 $layer=licon1_PDIFF $count=4 $X=0.595
+ $Y=1.84 $X2=1.36 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%X 1 2 9 14 15 16 17 23 29
c35 14 0 1.17819e-19 $X=4.07 $Y=1.985
r36 21 29 0.805779 $w=4.73e-07 $l=3.2e-08 $layer=LI1_cond $X=4.027 $Y=0.893
+ $X2=4.027 $Y2=0.925
r37 17 31 9.71933 $w=4.73e-07 $l=1.79e-07 $layer=LI1_cond $X=4.027 $Y=0.951
+ $X2=4.027 $Y2=1.13
r38 17 29 0.654696 $w=4.73e-07 $l=2.6e-08 $layer=LI1_cond $X=4.027 $Y=0.951
+ $X2=4.027 $Y2=0.925
r39 17 21 0.679876 $w=4.73e-07 $l=2.7e-08 $layer=LI1_cond $X=4.027 $Y=0.866
+ $X2=4.027 $Y2=0.893
r40 16 17 7.83117 $w=4.73e-07 $l=3.11e-07 $layer=LI1_cond $X=4.027 $Y=0.555
+ $X2=4.027 $Y2=0.866
r41 16 23 1.00722 $w=4.73e-07 $l=4e-08 $layer=LI1_cond $X=4.027 $Y=0.555
+ $X2=4.027 $Y2=0.515
r42 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.18 $Y=1.82 $X2=4.18
+ $Y2=1.13
r43 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=1.985
+ $X2=4.085 $Y2=1.82
r44 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=4.085 $Y=2 $X2=4.085
+ $Y2=1.985
r45 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=4.085 $Y=2 $X2=4.085
+ $Y2=2.815
r46 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.84 $X2=4.07 $Y2=1.985
r47 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.84 $X2=4.07 $Y2=2.815
r48 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.815
+ $Y=0.37 $X2=3.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%A_165_74# 1 2 9 12 13
r26 13 16 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.965 $Y=0.435
+ $X2=1.965 $Y2=0.665
r27 10 12 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.435
+ $X2=1.03 $Y2=0.435
r28 9 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=0.435
+ $X2=1.965 $Y2=0.435
r29 9 10 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.8 $Y=0.435
+ $X2=1.115 $Y2=0.435
r30 2 16 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.37 $X2=1.965 $Y2=0.665
r31 1 12 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=0.825
+ $Y=0.37 $X2=1.03 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%A_264_74# 1 2 7 11 14
c35 14 0 1.67816e-19 $X=1.495 $Y=0.965
c36 7 0 5.3557e-20 $X=2.87 $Y=1.095
r37 14 16 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=1.457 $Y=0.965
+ $X2=1.457 $Y2=1.095
r38 9 11 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.995 $Y=1.01
+ $X2=2.995 $Y2=0.515
r39 8 16 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=1.62 $Y=1.095
+ $X2=1.457 $Y2=1.095
r40 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.87 $Y=1.095
+ $X2=2.995 $Y2=1.01
r41 7 8 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.87 $Y=1.095
+ $X2=1.62 $Y2=1.095
r42 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.515
r43 1 14 182 $w=1.7e-07 $l=6.76868e-07 $layer=licon1_NDIFF $count=1 $X=1.32
+ $Y=0.37 $X2=1.495 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__O221A_2%VGND 1 2 3 12 16 18 20 23 24 26 27 28 40 46
r54 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r55 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r56 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 40 45 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.617
+ $Y2=0
r58 40 42 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.08
+ $Y2=0
r59 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r60 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 32 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r63 31 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r64 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 28 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r66 28 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r67 26 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.12
+ $Y2=0
r68 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.455
+ $Y2=0
r69 25 42 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=4.08
+ $Y2=0
r70 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.455
+ $Y2=0
r71 23 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r72 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.525
+ $Y2=0
r73 22 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=3.12
+ $Y2=0
r74 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.525
+ $Y2=0
r75 18 45 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.617 $Y2=0
r76 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.515
r77 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0
r78 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0.515
r79 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0
r80 10 12 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0.665
r81 3 20 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=4.245
+ $Y=0.37 $X2=4.52 $Y2=0.515
r82 2 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.245
+ $Y=0.37 $X2=3.455 $Y2=0.515
r83 1 12 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.37 $X2=2.525 $Y2=0.665
.ends


* File: sky130_fd_sc_ms__maj3_1.pxi.spice
* Created: Fri Aug 28 17:38:46 2020
* 
x_PM_SKY130_FD_SC_MS__MAJ3_1%A_84_74# N_A_84_74#_M1004_d N_A_84_74#_M1008_d
+ N_A_84_74#_M1010_d N_A_84_74#_M1003_d N_A_84_74#_M1002_g N_A_84_74#_M1001_g
+ N_A_84_74#_c_70_n N_A_84_74#_c_71_n N_A_84_74#_c_72_n N_A_84_74#_c_80_n
+ N_A_84_74#_c_73_n N_A_84_74#_c_117_p N_A_84_74#_c_74_n N_A_84_74#_c_108_p
+ N_A_84_74#_c_82_n N_A_84_74#_c_83_n N_A_84_74#_c_75_n N_A_84_74#_c_96_p
+ N_A_84_74#_c_76_n N_A_84_74#_c_77_n PM_SKY130_FD_SC_MS__MAJ3_1%A_84_74#
x_PM_SKY130_FD_SC_MS__MAJ3_1%B N_B_M1004_g N_B_M1010_g N_B_c_186_n N_B_M1013_g
+ N_B_M1009_g B N_B_c_187_n N_B_c_188_n PM_SKY130_FD_SC_MS__MAJ3_1%B
x_PM_SKY130_FD_SC_MS__MAJ3_1%C N_C_M1007_g N_C_M1012_g N_C_M1008_g N_C_M1003_g
+ N_C_c_236_n N_C_c_237_n C N_C_c_238_n N_C_c_239_n N_C_c_240_n N_C_c_241_n
+ PM_SKY130_FD_SC_MS__MAJ3_1%C
x_PM_SKY130_FD_SC_MS__MAJ3_1%A N_A_M1011_g N_A_c_297_n N_A_M1006_g N_A_c_299_n
+ N_A_c_300_n N_A_M1005_g N_A_c_302_n N_A_M1000_g A N_A_c_305_n N_A_c_306_n
+ PM_SKY130_FD_SC_MS__MAJ3_1%A
x_PM_SKY130_FD_SC_MS__MAJ3_1%X N_X_M1002_s N_X_M1001_s N_X_c_369_n N_X_c_370_n X
+ X X N_X_c_371_n PM_SKY130_FD_SC_MS__MAJ3_1%X
x_PM_SKY130_FD_SC_MS__MAJ3_1%VPWR N_VPWR_M1001_d N_VPWR_M1012_d N_VPWR_c_391_n
+ N_VPWR_c_392_n VPWR N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_390_n
+ N_VPWR_c_396_n N_VPWR_c_397_n PM_SKY130_FD_SC_MS__MAJ3_1%VPWR
x_PM_SKY130_FD_SC_MS__MAJ3_1%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_c_436_n
+ N_VGND_c_437_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_438_n N_VGND_c_439_n
+ VGND N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n
+ PM_SKY130_FD_SC_MS__MAJ3_1%VGND
cc_1 VNB N_A_84_74#_c_70_n 0.00825211f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.175
cc_2 VNB N_A_84_74#_c_71_n 0.00591492f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.175
cc_3 VNB N_A_84_74#_c_72_n 0.00347054f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=0.745
cc_4 VNB N_A_84_74#_c_73_n 0.00257431f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.95
cc_5 VNB N_A_84_74#_c_74_n 9.46947e-19 $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.175
cc_6 VNB N_A_84_74#_c_75_n 0.0269145f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_7 VNB N_A_84_74#_c_76_n 0.0172793f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.05
cc_8 VNB N_A_84_74#_c_77_n 0.0215805f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.35
cc_9 VNB N_B_M1004_g 0.021382f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.92
cc_10 VNB N_B_c_186_n 0.0152338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_187_n 0.00195337f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=0.745
cc_12 VNB N_B_c_188_n 0.026819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_236_n 0.0121979f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.4
cc_14 VNB N_C_c_237_n 0.0216658f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.4
cc_15 VNB N_C_c_238_n 0.0222716f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=0.745
cc_16 VNB N_C_c_239_n 0.0134552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_c_240_n 0.0207444f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.775
cc_18 VNB N_C_c_241_n 0.00130225f $X=-0.19 $Y=-0.245 $X2=3.395 $Y2=2.035
cc_19 VNB N_A_M1011_g 0.0285172f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=1.92
cc_20 VNB N_A_c_297_n 0.00564537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_M1006_g 0.0117219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_299_n 0.115517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_300_n 0.011606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_M1005_g 0.0107186f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.87
cc_25 VNB N_A_c_302_n 0.00493571f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.87
cc_26 VNB N_A_M1000_g 0.00711931f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.4
cc_27 VNB A 0.0240534f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.12
cc_28 VNB N_A_c_305_n 0.0540726f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.775
cc_29 VNB N_A_c_306_n 0.0129204f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.175
cc_30 VNB N_X_c_369_n 0.0241167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_370_n 0.00713231f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_32 VNB N_X_c_371_n 0.0221111f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.26
cc_33 VNB N_VPWR_c_390_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.37 $Y2=1.175
cc_34 VNB N_VGND_c_436_n 0.0108282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_437_n 0.0136584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_438_n 0.0381259f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.4
cc_37 VNB N_VGND_c_439_n 0.00229531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_440_n 0.0195478f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.09
cc_39 VNB N_VGND_c_441_n 0.0337601f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=2.775
cc_40 VNB N_VGND_c_442_n 0.221862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_443_n 0.00603779f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_42 VPB N_A_84_74#_M1001_g 0.0281595f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_43 VPB N_A_84_74#_c_71_n 0.00269398f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.175
cc_44 VPB N_A_84_74#_c_80_n 0.00300211f $X=-0.19 $Y=1.66 $X2=1.73 $Y2=2.775
cc_45 VPB N_A_84_74#_c_73_n 0.00217743f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.95
cc_46 VPB N_A_84_74#_c_82_n 0.00861803f $X=-0.19 $Y=1.66 $X2=3.56 $Y2=2.12
cc_47 VPB N_A_84_74#_c_83_n 0.0339166f $X=-0.19 $Y=1.66 $X2=3.56 $Y2=2.775
cc_48 VPB N_A_84_74#_c_75_n 0.00581463f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_49 VPB N_B_M1010_g 0.0204622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_B_M1009_g 0.0195924f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.87
cc_51 VPB N_B_c_187_n 0.0102481f $X=-0.19 $Y=1.66 $X2=1.645 $Y2=0.745
cc_52 VPB N_B_c_188_n 0.0132668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_C_M1012_g 0.0208372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_C_M1003_g 0.028852f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_55 VPB N_C_c_236_n 0.00701532f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_56 VPB N_C_c_237_n 0.0111038f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_57 VPB N_C_c_238_n 0.0115828f $X=-0.19 $Y=1.66 $X2=1.645 $Y2=0.745
cc_58 VPB N_C_c_241_n 0.00301732f $X=-0.19 $Y=1.66 $X2=3.395 $Y2=2.035
cc_59 VPB N_A_M1006_g 0.0255797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_M1000_g 0.0251826f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_61 VPB X 0.0503518f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.87
cc_62 VPB N_X_c_371_n 0.00919581f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.26
cc_63 VPB N_VPWR_c_391_n 0.00788465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_392_n 0.0069838f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.4
cc_65 VPB N_VPWR_c_393_n 0.0435374f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=1.175
cc_66 VPB N_VPWR_c_394_n 0.0315964f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.95
cc_67 VPB N_VPWR_c_390_n 0.0999658f $X=-0.19 $Y=1.66 $X2=3.37 $Y2=1.175
cc_68 VPB N_VPWR_c_396_n 0.0263192f $X=-0.19 $Y=1.66 $X2=2.065 $Y2=2.035
cc_69 VPB N_VPWR_c_397_n 0.00776418f $X=-0.19 $Y=1.66 $X2=3.56 $Y2=2.775
cc_70 N_A_84_74#_c_70_n N_B_M1004_g 0.0106503f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_71 N_A_84_74#_c_72_n N_B_M1004_g 0.00928072f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_72 N_A_84_74#_c_73_n N_B_M1004_g 9.50889e-19 $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_73 N_A_84_74#_c_74_n N_B_M1004_g 0.00112012f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_74 N_A_84_74#_c_80_n N_B_M1010_g 2.93395e-19 $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_75 N_A_84_74#_c_73_n N_B_M1010_g 9.53185e-19 $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_76 N_A_84_74#_c_72_n N_B_c_186_n 0.00347549f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_77 N_A_84_74#_c_73_n N_B_c_186_n 0.00527567f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_78 N_A_84_74#_c_74_n N_B_c_186_n 0.0145888f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_79 N_A_84_74#_c_80_n N_B_M1009_g 0.0157105f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_80 N_A_84_74#_c_73_n N_B_M1009_g 0.00551729f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_81 N_A_84_74#_c_96_p N_B_M1009_g 0.0138418f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_82 N_A_84_74#_M1001_g N_B_c_187_n 4.8198e-19 $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_84_74#_c_70_n N_B_c_187_n 0.0453726f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_84 N_A_84_74#_c_71_n N_B_c_187_n 0.0136497f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_85 N_A_84_74#_c_73_n N_B_c_187_n 0.0221901f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_86 N_A_84_74#_c_75_n N_B_c_187_n 2.4932e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A_84_74#_c_96_p N_B_c_187_n 0.00788943f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_88 N_A_84_74#_c_73_n N_B_c_188_n 0.0107607f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_89 N_A_84_74#_c_74_n N_B_c_188_n 0.00563521f $X=2.065 $Y=1.175 $X2=0 $Y2=0
cc_90 N_A_84_74#_c_96_p N_B_c_188_n 0.00413935f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_91 N_A_84_74#_c_80_n N_C_M1012_g 0.00265691f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_92 N_A_84_74#_c_73_n N_C_M1012_g 0.00283072f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_93 N_A_84_74#_c_108_p N_C_M1012_g 0.0164957f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_84_74#_c_108_p N_C_M1003_g 0.012823f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_95 N_A_84_74#_c_82_n N_C_M1003_g 0.0012593f $X=3.56 $Y=2.12 $X2=0 $Y2=0
cc_96 N_A_84_74#_c_83_n N_C_M1003_g 0.0160401f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_97 N_A_84_74#_c_108_p N_C_c_236_n 0.0380714f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_84_74#_c_82_n N_C_c_236_n 0.0121815f $X=3.56 $Y=2.12 $X2=0 $Y2=0
cc_99 N_A_84_74#_c_76_n N_C_c_236_n 0.0137699f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_100 N_A_84_74#_c_82_n N_C_c_237_n 0.00332066f $X=3.56 $Y=2.12 $X2=0 $Y2=0
cc_101 N_A_84_74#_c_76_n N_C_c_237_n 0.0040945f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_102 N_A_84_74#_c_117_p N_C_c_238_n 0.00505145f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_103 N_A_84_74#_c_108_p N_C_c_238_n 8.78225e-19 $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_104 N_A_84_74#_c_73_n N_C_c_239_n 0.0042291f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_105 N_A_84_74#_c_117_p N_C_c_239_n 0.0131284f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_106 N_A_84_74#_c_117_p N_C_c_240_n 0.00928007f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_107 N_A_84_74#_c_76_n N_C_c_240_n 0.00674358f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_108 N_A_84_74#_c_73_n N_C_c_241_n 0.0228143f $X=1.98 $Y=1.95 $X2=0 $Y2=0
cc_109 N_A_84_74#_c_117_p N_C_c_241_n 0.0728496f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_110 N_A_84_74#_c_108_p N_C_c_241_n 0.0335591f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A_84_74#_c_70_n N_A_M1011_g 0.0179891f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_112 N_A_84_74#_c_71_n N_A_M1011_g 0.0055338f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_113 N_A_84_74#_c_72_n N_A_M1011_g 0.00182632f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_114 N_A_84_74#_c_77_n N_A_M1011_g 0.0199957f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_115 N_A_84_74#_c_70_n N_A_c_297_n 9.05238e-19 $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_116 N_A_84_74#_c_75_n N_A_c_297_n 0.0197603f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A_84_74#_M1001_g N_A_M1006_g 0.0132905f $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_84_74#_c_72_n N_A_c_299_n 0.00612247f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_119 N_A_84_74#_c_117_p N_A_M1005_g 0.0124955f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_120 N_A_84_74#_c_76_n N_A_M1005_g 0.00116861f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_121 N_A_84_74#_c_108_p N_A_M1000_g 0.0171007f $X=3.395 $Y=2.035 $X2=0 $Y2=0
cc_122 N_A_84_74#_c_83_n N_A_M1000_g 0.00266928f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_123 N_A_84_74#_c_76_n A 0.0178486f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_124 N_A_84_74#_c_117_p N_A_c_306_n 0.0147496f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_125 N_A_84_74#_c_76_n N_A_c_306_n 0.00467871f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_126 N_A_84_74#_c_77_n N_X_c_369_n 0.00692086f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_84_74#_c_71_n N_X_c_370_n 0.00152814f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_128 N_A_84_74#_c_77_n N_X_c_370_n 0.00300451f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_129 N_A_84_74#_M1001_g X 0.0151561f $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A_84_74#_c_71_n X 0.00361172f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_131 N_A_84_74#_M1001_g N_X_c_371_n 0.00402233f $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_84_74#_c_71_n N_X_c_371_n 0.0303017f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_133 N_A_84_74#_c_77_n N_X_c_371_n 0.0100022f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_134 N_A_84_74#_c_108_p N_VPWR_M1012_d 0.00503584f $X=3.395 $Y=2.035 $X2=0
+ $Y2=0
cc_135 N_A_84_74#_M1001_g N_VPWR_c_391_n 0.00396119f $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_84_74#_c_71_n N_VPWR_c_391_n 0.00648751f $X=0.785 $Y=1.175 $X2=0
+ $Y2=0
cc_137 N_A_84_74#_c_80_n N_VPWR_c_391_n 0.0256573f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_138 N_A_84_74#_c_75_n N_VPWR_c_391_n 5.65558e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A_84_74#_c_96_p N_VPWR_c_391_n 0.00572303f $X=1.73 $Y=2.095 $X2=0 $Y2=0
cc_140 N_A_84_74#_c_80_n N_VPWR_c_392_n 0.0192019f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_141 N_A_84_74#_c_108_p N_VPWR_c_392_n 0.0232055f $X=3.395 $Y=2.035 $X2=0
+ $Y2=0
cc_142 N_A_84_74#_c_83_n N_VPWR_c_392_n 0.0187356f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_143 N_A_84_74#_c_80_n N_VPWR_c_393_n 0.0125236f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_144 N_A_84_74#_c_83_n N_VPWR_c_394_n 0.0125236f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_145 N_A_84_74#_M1001_g N_VPWR_c_390_n 0.00990615f $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_84_74#_c_80_n N_VPWR_c_390_n 0.0117917f $X=1.73 $Y=2.775 $X2=0 $Y2=0
cc_147 N_A_84_74#_c_83_n N_VPWR_c_390_n 0.0117917f $X=3.56 $Y=2.775 $X2=0 $Y2=0
cc_148 N_A_84_74#_M1001_g N_VPWR_c_396_n 0.005209f $X=0.55 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_84_74#_c_108_p A_409_384# 0.0096152f $X=3.395 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_84_74#_c_108_p A_601_384# 0.00621497f $X=3.395 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_84_74#_c_70_n N_VGND_M1002_d 0.00132837f $X=1.48 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_84_74#_c_71_n N_VGND_M1002_d 0.00248319f $X=0.785 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_84_74#_c_117_p N_VGND_M1007_d 0.00661484f $X=3.37 $Y=1.175 $X2=0
+ $Y2=0
cc_154 N_A_84_74#_c_70_n N_VGND_c_436_n 0.0112589f $X=1.48 $Y=1.175 $X2=0 $Y2=0
cc_155 N_A_84_74#_c_71_n N_VGND_c_436_n 0.0135036f $X=0.785 $Y=1.175 $X2=0 $Y2=0
cc_156 N_A_84_74#_c_72_n N_VGND_c_436_n 0.0105579f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_157 N_A_84_74#_c_75_n N_VGND_c_436_n 5.99498e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A_84_74#_c_77_n N_VGND_c_436_n 0.00580418f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_159 N_A_84_74#_c_72_n N_VGND_c_437_n 0.00420212f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_160 N_A_84_74#_c_117_p N_VGND_c_453_n 0.00820442f $X=3.37 $Y=1.175 $X2=0
+ $Y2=0
cc_161 N_A_84_74#_c_117_p N_VGND_c_454_n 0.02198f $X=3.37 $Y=1.175 $X2=0 $Y2=0
cc_162 N_A_84_74#_c_76_n N_VGND_c_454_n 0.00216203f $X=3.535 $Y=1.05 $X2=0 $Y2=0
cc_163 N_A_84_74#_c_72_n N_VGND_c_438_n 0.00725358f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_164 N_A_84_74#_c_77_n N_VGND_c_440_n 0.00467453f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_165 N_A_84_74#_c_72_n N_VGND_c_442_n 0.00890448f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_166 N_A_84_74#_c_77_n N_VGND_c_442_n 0.00505379f $X=0.587 $Y=1.35 $X2=0 $Y2=0
cc_167 N_A_84_74#_c_70_n A_223_120# 0.0048076f $X=1.48 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A_84_74#_c_117_p A_403_136# 0.0096152f $X=3.37 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_84_74#_c_117_p A_595_136# 0.00453974f $X=3.37 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_170 N_B_M1009_g N_C_M1012_g 0.0671297f $X=1.955 $Y=2.42 $X2=0 $Y2=0
cc_171 N_B_c_188_n N_C_c_238_n 0.0209073f $X=1.955 $Y=1.595 $X2=0 $Y2=0
cc_172 N_B_c_186_n N_C_c_239_n 0.0451321f $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_173 N_B_c_188_n N_C_c_241_n 3.74525e-19 $X=1.955 $Y=1.595 $X2=0 $Y2=0
cc_174 N_B_M1004_g N_A_M1011_g 0.0437821f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_175 N_B_M1004_g N_A_c_297_n 0.0143837f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_176 N_B_M1010_g N_A_M1006_g 0.0675302f $X=1.475 $Y=2.42 $X2=0 $Y2=0
cc_177 N_B_c_187_n N_A_M1006_g 0.0130461f $X=1.52 $Y=1.595 $X2=0 $Y2=0
cc_178 N_B_c_188_n N_A_M1006_g 0.0143837f $X=1.955 $Y=1.595 $X2=0 $Y2=0
cc_179 N_B_M1004_g N_A_c_299_n 0.0103098f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_180 N_B_c_186_n N_A_c_299_n 0.00746712f $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_181 N_B_M1010_g N_VPWR_c_391_n 0.00334491f $X=1.475 $Y=2.42 $X2=0 $Y2=0
cc_182 N_B_M1009_g N_VPWR_c_392_n 0.00236707f $X=1.955 $Y=2.42 $X2=0 $Y2=0
cc_183 N_B_M1010_g N_VPWR_c_393_n 0.00658449f $X=1.475 $Y=2.42 $X2=0 $Y2=0
cc_184 N_B_M1009_g N_VPWR_c_393_n 0.00628513f $X=1.955 $Y=2.42 $X2=0 $Y2=0
cc_185 N_B_M1010_g N_VPWR_c_390_n 0.00639697f $X=1.475 $Y=2.42 $X2=0 $Y2=0
cc_186 N_B_M1009_g N_VPWR_c_390_n 0.00639697f $X=1.955 $Y=2.42 $X2=0 $Y2=0
cc_187 N_B_M1004_g N_VGND_c_436_n 0.00147743f $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_188 N_B_c_186_n N_VGND_c_437_n 7.10756e-19 $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_189 N_B_c_186_n N_VGND_c_453_n 5.65853e-19 $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_190 N_B_M1004_g N_VGND_c_442_n 9.33152e-19 $X=1.43 $Y=0.92 $X2=0 $Y2=0
cc_191 N_B_c_186_n N_VGND_c_442_n 9.5708e-19 $X=1.94 $Y=1.43 $X2=0 $Y2=0
cc_192 N_C_c_239_n N_A_c_299_n 0.00683881f $X=2.435 $Y=1.4 $X2=0 $Y2=0
cc_193 N_C_c_239_n N_A_M1005_g 0.0240392f $X=2.435 $Y=1.4 $X2=0 $Y2=0
cc_194 N_C_c_236_n N_A_c_302_n 0.00424265f $X=3.41 $Y=1.595 $X2=0 $Y2=0
cc_195 N_C_c_238_n N_A_c_302_n 0.0234781f $X=2.45 $Y=1.595 $X2=0 $Y2=0
cc_196 N_C_c_240_n N_A_c_302_n 0.0444619f $X=3.41 $Y=1.43 $X2=0 $Y2=0
cc_197 N_C_M1012_g N_A_M1000_g 0.0201707f $X=2.375 $Y=2.42 $X2=0 $Y2=0
cc_198 N_C_c_236_n N_A_M1000_g 0.0125533f $X=3.41 $Y=1.595 $X2=0 $Y2=0
cc_199 N_C_c_237_n N_A_M1000_g 0.0444619f $X=3.41 $Y=1.595 $X2=0 $Y2=0
cc_200 N_C_c_241_n N_A_M1000_g 5.65769e-19 $X=2.755 $Y=1.605 $X2=0 $Y2=0
cc_201 N_C_c_240_n A 0.00384087f $X=3.41 $Y=1.43 $X2=0 $Y2=0
cc_202 N_C_c_239_n N_A_c_305_n 0.00110103f $X=2.435 $Y=1.4 $X2=0 $Y2=0
cc_203 N_C_c_240_n N_A_c_305_n 0.040752f $X=3.41 $Y=1.43 $X2=0 $Y2=0
cc_204 N_C_c_240_n N_A_c_306_n 0.00756106f $X=3.41 $Y=1.43 $X2=0 $Y2=0
cc_205 N_C_M1012_g N_VPWR_c_392_n 0.0171423f $X=2.375 $Y=2.42 $X2=0 $Y2=0
cc_206 N_C_M1003_g N_VPWR_c_392_n 0.0023091f $X=3.335 $Y=2.42 $X2=0 $Y2=0
cc_207 N_C_M1012_g N_VPWR_c_393_n 0.00547402f $X=2.375 $Y=2.42 $X2=0 $Y2=0
cc_208 N_C_M1003_g N_VPWR_c_394_n 0.00628513f $X=3.335 $Y=2.42 $X2=0 $Y2=0
cc_209 N_C_M1012_g N_VPWR_c_390_n 0.00536634f $X=2.375 $Y=2.42 $X2=0 $Y2=0
cc_210 N_C_M1003_g N_VPWR_c_390_n 0.00639697f $X=3.335 $Y=2.42 $X2=0 $Y2=0
cc_211 N_C_c_239_n N_VGND_c_437_n 0.00678491f $X=2.435 $Y=1.4 $X2=0 $Y2=0
cc_212 N_C_c_239_n N_VGND_c_453_n 0.00784325f $X=2.435 $Y=1.4 $X2=0 $Y2=0
cc_213 N_C_c_240_n N_VGND_c_454_n 6.83236e-19 $X=3.41 $Y=1.43 $X2=0 $Y2=0
cc_214 N_C_c_240_n N_VGND_c_441_n 4.78105e-19 $X=3.41 $Y=1.43 $X2=0 $Y2=0
cc_215 N_C_c_239_n N_VGND_c_442_n 3.25407e-19 $X=2.435 $Y=1.4 $X2=0 $Y2=0
cc_216 N_A_M1011_g N_X_c_369_n 8.44714e-19 $X=1.04 $Y=0.92 $X2=0 $Y2=0
cc_217 N_A_M1006_g X 6.64279e-19 $X=1.055 $Y=2.42 $X2=0 $Y2=0
cc_218 N_A_M1006_g N_VPWR_c_391_n 0.0237312f $X=1.055 $Y=2.42 $X2=0 $Y2=0
cc_219 N_A_M1000_g N_VPWR_c_392_n 0.0159666f $X=2.915 $Y=2.42 $X2=0 $Y2=0
cc_220 N_A_M1006_g N_VPWR_c_393_n 0.00565692f $X=1.055 $Y=2.42 $X2=0 $Y2=0
cc_221 N_A_M1000_g N_VPWR_c_394_n 0.00602273f $X=2.915 $Y=2.42 $X2=0 $Y2=0
cc_222 N_A_M1006_g N_VPWR_c_390_n 0.00554404f $X=1.055 $Y=2.42 $X2=0 $Y2=0
cc_223 N_A_M1000_g N_VPWR_c_390_n 0.00589942f $X=2.915 $Y=2.42 $X2=0 $Y2=0
cc_224 N_A_M1011_g N_VGND_c_436_n 0.0223799f $X=1.04 $Y=0.92 $X2=0 $Y2=0
cc_225 N_A_c_300_n N_VGND_c_436_n 0.00786053f $X=1.115 $Y=0.185 $X2=0 $Y2=0
cc_226 N_A_c_299_n N_VGND_c_437_n 0.0157239f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_227 N_A_M1005_g N_VGND_c_437_n 0.0029973f $X=2.9 $Y=1 $X2=0 $Y2=0
cc_228 N_A_c_305_n N_VGND_c_437_n 0.00210171f $X=2.81 $Y=0.185 $X2=0 $Y2=0
cc_229 N_A_c_306_n N_VGND_c_437_n 0.0249987f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_230 N_A_c_299_n N_VGND_c_454_n 0.00129982f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_231 N_A_M1005_g N_VGND_c_454_n 0.00645394f $X=2.9 $Y=1 $X2=0 $Y2=0
cc_232 N_A_c_305_n N_VGND_c_454_n 0.00419722f $X=2.81 $Y=0.185 $X2=0 $Y2=0
cc_233 N_A_c_306_n N_VGND_c_454_n 0.0125685f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_234 N_A_c_300_n N_VGND_c_438_n 0.0430809f $X=1.115 $Y=0.185 $X2=0 $Y2=0
cc_235 N_A_c_299_n N_VGND_c_441_n 0.0122079f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_236 N_A_c_306_n N_VGND_c_441_n 0.0712235f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_237 N_A_c_299_n N_VGND_c_442_n 0.0536057f $X=2.645 $Y=0.185 $X2=0 $Y2=0
cc_238 N_A_c_300_n N_VGND_c_442_n 0.00750358f $X=1.115 $Y=0.185 $X2=0 $Y2=0
cc_239 N_A_c_305_n N_VGND_c_442_n 0.0102245f $X=2.81 $Y=0.185 $X2=0 $Y2=0
cc_240 N_A_c_306_n N_VGND_c_442_n 0.0393319f $X=3.485 $Y=0.462 $X2=0 $Y2=0
cc_241 X N_VPWR_c_391_n 0.0406301f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_242 X N_VPWR_c_390_n 0.0147443f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_243 X N_VPWR_c_396_n 0.0178955f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_244 N_X_c_369_n N_VGND_c_436_n 0.0171569f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_245 N_X_c_369_n N_VGND_c_440_n 0.0103924f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_246 N_X_c_369_n N_VGND_c_442_n 0.0121284f $X=0.28 $Y=0.645 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o21a_4.pxi.spice
* Created: Wed Sep  2 12:21:43 2020
* 
x_PM_SKY130_FD_SC_MS__O21A_4%A2 N_A2_M1011_g N_A2_M1003_g N_A2_M1004_g
+ N_A2_M1013_g A2 N_A2_c_104_n N_A2_c_105_n PM_SKY130_FD_SC_MS__O21A_4%A2
x_PM_SKY130_FD_SC_MS__O21A_4%A1 N_A1_c_153_n N_A1_M1014_g N_A1_M1015_g
+ N_A1_c_156_n N_A1_c_157_n N_A1_M1016_g N_A1_M1018_g A1 N_A1_c_160_n
+ PM_SKY130_FD_SC_MS__O21A_4%A1
x_PM_SKY130_FD_SC_MS__O21A_4%B1 N_B1_M1010_g N_B1_M1000_g N_B1_M1019_g
+ N_B1_M1008_g B1 B1 N_B1_c_221_n PM_SKY130_FD_SC_MS__O21A_4%B1
x_PM_SKY130_FD_SC_MS__O21A_4%A_219_387# N_A_219_387#_M1010_s
+ N_A_219_387#_M1011_d N_A_219_387#_M1000_d N_A_219_387#_M1007_g
+ N_A_219_387#_c_271_n N_A_219_387#_M1001_g N_A_219_387#_M1009_g
+ N_A_219_387#_c_273_n N_A_219_387#_M1002_g N_A_219_387#_c_285_n
+ N_A_219_387#_M1012_g N_A_219_387#_c_274_n N_A_219_387#_M1005_g
+ N_A_219_387#_c_286_n N_A_219_387#_M1017_g N_A_219_387#_c_275_n
+ N_A_219_387#_M1006_g N_A_219_387#_c_290_n N_A_219_387#_c_276_n
+ N_A_219_387#_c_277_n N_A_219_387#_c_278_n N_A_219_387#_c_312_n
+ N_A_219_387#_c_279_n N_A_219_387#_c_280_n N_A_219_387#_c_292_n
+ N_A_219_387#_c_288_n N_A_219_387#_c_281_n N_A_219_387#_c_282_n
+ PM_SKY130_FD_SC_MS__O21A_4%A_219_387#
x_PM_SKY130_FD_SC_MS__O21A_4%VPWR N_VPWR_M1014_d N_VPWR_M1016_d N_VPWR_M1008_s
+ N_VPWR_M1009_s N_VPWR_M1017_s N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n
+ N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n
+ N_VPWR_c_423_n VPWR N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n
+ N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_414_n PM_SKY130_FD_SC_MS__O21A_4%VPWR
x_PM_SKY130_FD_SC_MS__O21A_4%A_119_387# N_A_119_387#_M1014_s
+ N_A_119_387#_M1013_s N_A_119_387#_c_486_n N_A_119_387#_c_484_n
+ N_A_119_387#_c_485_n N_A_119_387#_c_492_n
+ PM_SKY130_FD_SC_MS__O21A_4%A_119_387#
x_PM_SKY130_FD_SC_MS__O21A_4%X N_X_M1001_s N_X_M1005_s N_X_M1007_d N_X_M1012_d
+ N_X_c_508_n N_X_c_518_n N_X_c_504_n N_X_c_509_n N_X_c_510_n N_X_c_532_n
+ N_X_c_511_n N_X_c_505_n N_X_c_506_n N_X_c_545_n X PM_SKY130_FD_SC_MS__O21A_4%X
x_PM_SKY130_FD_SC_MS__O21A_4%A_27_125# N_A_27_125#_M1015_s N_A_27_125#_M1003_d
+ N_A_27_125#_M1018_s N_A_27_125#_M1019_d N_A_27_125#_c_575_n
+ N_A_27_125#_c_576_n N_A_27_125#_c_577_n N_A_27_125#_c_578_n
+ N_A_27_125#_c_579_n N_A_27_125#_c_580_n N_A_27_125#_c_581_n
+ N_A_27_125#_c_582_n N_A_27_125#_c_583_n N_A_27_125#_c_584_n
+ PM_SKY130_FD_SC_MS__O21A_4%A_27_125#
x_PM_SKY130_FD_SC_MS__O21A_4%VGND N_VGND_M1015_d N_VGND_M1004_s N_VGND_M1001_d
+ N_VGND_M1002_d N_VGND_M1006_d N_VGND_c_642_n N_VGND_c_643_n N_VGND_c_644_n
+ N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n VGND N_VGND_c_648_n
+ N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n N_VGND_c_653_n
+ N_VGND_c_654_n N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n
+ PM_SKY130_FD_SC_MS__O21A_4%VGND
cc_1 VNB N_A2_M1003_g 0.0186294f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.945
cc_2 VNB N_A2_M1004_g 0.0202457f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.945
cc_3 VNB N_A2_c_104_n 0.00175162f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_4 VNB N_A2_c_105_n 0.0305957f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.61
cc_5 VNB N_A1_c_153_n 0.00868929f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.775
cc_6 VNB N_A1_M1014_g 0.0194277f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.435
cc_7 VNB N_A1_M1015_g 0.0364999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_156_n 0.108819f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.445
cc_9 VNB N_A1_c_157_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.945
cc_10 VNB N_A1_M1018_g 0.0331968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A1 0.0046028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_160_n 0.0170803f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_13 VNB N_B1_M1010_g 0.0191682f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.435
cc_14 VNB N_B1_M1019_g 0.0205347f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.945
cc_15 VNB B1 0.0021003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_221_n 0.0321688f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.61
cc_17 VNB N_A_219_387#_M1007_g 0.00685469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_219_387#_c_271_n 0.0198604f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.435
cc_19 VNB N_A_219_387#_M1009_g 0.00622166f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.61
cc_20 VNB N_A_219_387#_c_273_n 0.0164674f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.61
cc_21 VNB N_A_219_387#_c_274_n 0.0166181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_219_387#_c_275_n 0.021272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_219_387#_c_276_n 0.00200913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_219_387#_c_277_n 0.00762265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_219_387#_c_278_n 0.00269748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_219_387#_c_279_n 0.00169712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_219_387#_c_280_n 0.00982261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_219_387#_c_281_n 0.00906033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_219_387#_c_282_n 0.140899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_414_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_504_n 0.00215307f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.61
cc_32 VNB N_X_c_505_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_506_n 0.00177379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.00943489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_125#_c_575_n 0.022896f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.435
cc_36 VNB N_A_27_125#_c_576_n 0.00568431f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_37 VNB N_A_27_125#_c_577_n 0.0125745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_125#_c_578_n 0.00206719f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.61
cc_39 VNB N_A_27_125#_c_579_n 0.00867474f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_40 VNB N_A_27_125#_c_580_n 8.44865e-19 $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.61
cc_41 VNB N_A_27_125#_c_581_n 0.0214365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_125#_c_582_n 0.00249092f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.665
cc_43 VNB N_A_27_125#_c_583_n 0.00923286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_125#_c_584_n 0.00177457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_642_n 0.00825723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_643_n 0.00930184f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_47 VNB N_VGND_c_644_n 0.0149193f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.61
cc_48 VNB N_VGND_c_645_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.665
cc_49 VNB N_VGND_c_646_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_647_n 0.0425996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_648_n 0.0191172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_649_n 0.0160823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_650_n 0.0403231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_651_n 0.017175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_652_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_653_n 0.00446116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_654_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_655_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_656_n 0.00668318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_657_n 0.320652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VPB N_A2_M1011_g 0.0200827f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.435
cc_62 VPB N_A2_M1013_g 0.0201673f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.435
cc_63 VPB N_A2_c_104_n 0.0047247f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_64 VPB N_A2_c_105_n 0.0177568f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.61
cc_65 VPB N_A1_M1014_g 0.0369551f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.435
cc_66 VPB N_A1_M1016_g 0.0217514f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.775
cc_67 VPB A1 0.00434418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A1_c_160_n 0.0110334f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_69 VPB N_B1_M1000_g 0.022836f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.945
cc_70 VPB N_B1_M1008_g 0.0243126f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.435
cc_71 VPB B1 0.00518591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_B1_c_221_n 0.0195848f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.61
cc_73 VPB N_A_219_387#_M1007_g 0.0243751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_219_387#_M1009_g 0.0225257f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.61
cc_75 VPB N_A_219_387#_c_285_n 0.0171241f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_76 VPB N_A_219_387#_c_286_n 0.0195136f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.665
cc_77 VPB N_A_219_387#_c_279_n 0.00445481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_219_387#_c_288_n 0.00378636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_219_387#_c_282_n 0.0140383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_415_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_416_n 0.055333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_417_n 0.0173751f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_83 VPB N_VPWR_c_418_n 0.0205087f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.61
cc_84 VPB N_VPWR_c_419_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_420_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_421_n 0.0513896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_422_n 0.0217043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_423_n 0.00920679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_424_n 0.039459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_425_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_426_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_427_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_428_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_414_n 0.0835591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_119_387#_c_484_n 0.00746603f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.775
cc_96 VPB N_A_119_387#_c_485_n 0.00324772f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.435
cc_97 VPB N_X_c_508_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.435
cc_98 VPB N_X_c_509_n 0.00283613f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_99 VPB N_X_c_510_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_100 VPB N_X_c_511_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB X 0.00923524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 N_A2_M1003_g N_A1_c_153_n 0.00461814f $X=1 $Y=0.945 $X2=-0.19 $Y2=-0.245
cc_103 N_A2_M1011_g N_A1_M1014_g 0.0116075f $X=1.005 $Y=2.435 $X2=0 $Y2=0
cc_104 N_A2_c_104_n N_A1_M1014_g 0.00227822f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_105 N_A2_c_105_n N_A1_M1014_g 0.0199852f $X=1.455 $Y=1.61 $X2=0 $Y2=0
cc_106 N_A2_M1003_g N_A1_M1015_g 0.0205891f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_107 N_A2_M1003_g N_A1_c_156_n 0.00894529f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_108 N_A2_M1004_g N_A1_c_156_n 0.00895007f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_109 N_A2_M1013_g N_A1_M1016_g 0.0234251f $X=1.455 $Y=2.435 $X2=0 $Y2=0
cc_110 N_A2_M1004_g N_A1_M1018_g 0.0222303f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_111 N_A2_c_104_n A1 0.0177636f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_112 N_A2_c_105_n A1 0.00145483f $X=1.455 $Y=1.61 $X2=0 $Y2=0
cc_113 N_A2_c_104_n N_A1_c_160_n 3.92399e-19 $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_114 N_A2_c_105_n N_A1_c_160_n 0.0177602f $X=1.455 $Y=1.61 $X2=0 $Y2=0
cc_115 N_A2_M1013_g N_A_219_387#_c_290_n 0.0136543f $X=1.455 $Y=2.435 $X2=0
+ $Y2=0
cc_116 N_A2_c_104_n N_A_219_387#_c_290_n 0.00780011f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_117 N_A2_M1011_g N_A_219_387#_c_292_n 0.0109711f $X=1.005 $Y=2.435 $X2=0
+ $Y2=0
cc_118 N_A2_M1013_g N_A_219_387#_c_292_n 0.0104072f $X=1.455 $Y=2.435 $X2=0
+ $Y2=0
cc_119 N_A2_c_104_n N_A_219_387#_c_292_n 0.0231394f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_120 N_A2_c_105_n N_A_219_387#_c_292_n 7.01268e-19 $X=1.455 $Y=1.61 $X2=0
+ $Y2=0
cc_121 N_A2_M1011_g N_VPWR_c_416_n 4.51712e-19 $X=1.005 $Y=2.435 $X2=0 $Y2=0
cc_122 N_A2_M1011_g N_VPWR_c_424_n 0.00113339f $X=1.005 $Y=2.435 $X2=0 $Y2=0
cc_123 N_A2_M1013_g N_VPWR_c_424_n 0.00113339f $X=1.455 $Y=2.435 $X2=0 $Y2=0
cc_124 N_A2_c_104_n N_A_119_387#_c_486_n 0.00217105f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_125 N_A2_c_105_n N_A_119_387#_c_486_n 2.00459e-19 $X=1.455 $Y=1.61 $X2=0
+ $Y2=0
cc_126 N_A2_M1011_g N_A_119_387#_c_484_n 0.0155346f $X=1.005 $Y=2.435 $X2=0
+ $Y2=0
cc_127 N_A2_M1013_g N_A_119_387#_c_484_n 0.0157584f $X=1.455 $Y=2.435 $X2=0
+ $Y2=0
cc_128 N_A2_M1003_g N_A_27_125#_c_575_n 8.14629e-19 $X=1 $Y=0.945 $X2=0 $Y2=0
cc_129 N_A2_M1003_g N_A_27_125#_c_576_n 0.0125078f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_130 N_A2_c_104_n N_A_27_125#_c_576_n 0.0216324f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_131 N_A2_c_105_n N_A_27_125#_c_576_n 6.26462e-19 $X=1.455 $Y=1.61 $X2=0 $Y2=0
cc_132 N_A2_M1004_g N_A_27_125#_c_578_n 0.00735846f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_133 N_A2_M1004_g N_A_27_125#_c_579_n 0.0116092f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_134 N_A2_c_104_n N_A_27_125#_c_579_n 0.0088782f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_135 N_A2_c_105_n N_A_27_125#_c_579_n 0.001253f $X=1.455 $Y=1.61 $X2=0 $Y2=0
cc_136 N_A2_M1004_g N_A_27_125#_c_580_n 8.55081e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_137 N_A2_M1004_g N_A_27_125#_c_584_n 8.39256e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_138 N_A2_c_104_n N_A_27_125#_c_584_n 0.0210722f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_139 N_A2_c_105_n N_A_27_125#_c_584_n 7.84649e-19 $X=1.455 $Y=1.61 $X2=0 $Y2=0
cc_140 N_A2_M1003_g N_VGND_c_642_n 0.00763474f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_141 N_A2_M1004_g N_VGND_c_642_n 4.4191e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_142 N_A2_M1004_g N_VGND_c_643_n 0.00378934f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_143 N_A2_M1003_g N_VGND_c_657_n 7.97988e-19 $X=1 $Y=0.945 $X2=0 $Y2=0
cc_144 N_A2_M1004_g N_VGND_c_657_n 9.49986e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_145 N_A1_M1018_g N_B1_M1010_g 0.0145764f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_146 N_A1_M1016_g N_B1_M1000_g 0.0241429f $X=1.955 $Y=2.435 $X2=0 $Y2=0
cc_147 A1 B1 0.0227747f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A1_c_160_n B1 2.18718e-19 $X=1.96 $Y=1.61 $X2=0 $Y2=0
cc_149 A1 N_B1_c_221_n 0.00413574f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A1_c_160_n N_B1_c_221_n 0.0182242f $X=1.96 $Y=1.61 $X2=0 $Y2=0
cc_151 N_A1_M1016_g N_A_219_387#_c_290_n 0.0169721f $X=1.955 $Y=2.435 $X2=0
+ $Y2=0
cc_152 A1 N_A_219_387#_c_290_n 0.0321436f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A1_c_160_n N_A_219_387#_c_290_n 7.92341e-19 $X=1.96 $Y=1.61 $X2=0 $Y2=0
cc_154 N_A1_M1016_g N_A_219_387#_c_292_n 6.68293e-19 $X=1.955 $Y=2.435 $X2=0
+ $Y2=0
cc_155 N_A1_M1016_g N_A_219_387#_c_288_n 8.03883e-19 $X=1.955 $Y=2.435 $X2=0
+ $Y2=0
cc_156 N_A1_M1014_g N_VPWR_c_416_n 0.017686f $X=0.505 $Y=2.435 $X2=0 $Y2=0
cc_157 N_A1_M1016_g N_VPWR_c_417_n 0.00526268f $X=1.955 $Y=2.435 $X2=0 $Y2=0
cc_158 N_A1_M1014_g N_VPWR_c_424_n 0.00558361f $X=0.505 $Y=2.435 $X2=0 $Y2=0
cc_159 N_A1_M1016_g N_VPWR_c_424_n 0.00578564f $X=1.955 $Y=2.435 $X2=0 $Y2=0
cc_160 N_A1_M1014_g N_VPWR_c_414_n 0.00541439f $X=0.505 $Y=2.435 $X2=0 $Y2=0
cc_161 N_A1_M1016_g N_VPWR_c_414_n 0.00537853f $X=1.955 $Y=2.435 $X2=0 $Y2=0
cc_162 N_A1_M1016_g N_A_119_387#_c_484_n 0.00400061f $X=1.955 $Y=2.435 $X2=0
+ $Y2=0
cc_163 N_A1_M1014_g N_A_119_387#_c_485_n 0.00122724f $X=0.505 $Y=2.435 $X2=0
+ $Y2=0
cc_164 N_A1_M1016_g N_A_119_387#_c_492_n 0.00787532f $X=1.955 $Y=2.435 $X2=0
+ $Y2=0
cc_165 N_A1_M1015_g N_A_27_125#_c_575_n 0.00756074f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_166 N_A1_c_153_n N_A_27_125#_c_576_n 0.00116345f $X=0.505 $Y=1.43 $X2=0 $Y2=0
cc_167 N_A1_M1015_g N_A_27_125#_c_576_n 0.0152942f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_168 N_A1_M1015_g N_A_27_125#_c_577_n 0.00167997f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_169 N_A1_c_156_n N_A_27_125#_c_578_n 0.00449567f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_170 N_A1_M1018_g N_A_27_125#_c_578_n 8.40186e-19 $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_171 N_A1_M1018_g N_A_27_125#_c_579_n 0.0126915f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_172 A1 N_A_27_125#_c_579_n 0.0380956f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A1_c_160_n N_A_27_125#_c_579_n 0.0043465f $X=1.96 $Y=1.61 $X2=0 $Y2=0
cc_174 N_A1_M1018_g N_A_27_125#_c_580_n 0.0113517f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_175 N_A1_M1018_g N_A_27_125#_c_582_n 0.00615508f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_176 N_A1_M1015_g N_VGND_c_642_n 0.0151444f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_177 N_A1_c_156_n N_VGND_c_642_n 0.0235422f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_178 N_A1_c_156_n N_VGND_c_643_n 0.0235859f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_179 N_A1_M1018_g N_VGND_c_643_n 0.00876868f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_180 N_A1_c_157_n N_VGND_c_648_n 0.00730708f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_181 N_A1_c_156_n N_VGND_c_649_n 0.0187698f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_182 N_A1_c_156_n N_VGND_c_650_n 0.00719493f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_183 N_A1_c_156_n N_VGND_c_657_n 0.0361523f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_184 N_A1_c_157_n N_VGND_c_657_n 0.0101958f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_185 N_B1_c_221_n N_A_219_387#_M1007_g 0.0207569f $X=3.025 $Y=1.61 $X2=0 $Y2=0
cc_186 N_B1_M1000_g N_A_219_387#_c_290_n 0.0153407f $X=2.495 $Y=2.355 $X2=0
+ $Y2=0
cc_187 B1 N_A_219_387#_c_290_n 0.0083868f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_188 N_B1_M1019_g N_A_219_387#_c_276_n 0.011831f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_189 N_B1_M1019_g N_A_219_387#_c_277_n 0.012382f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_190 B1 N_A_219_387#_c_277_n 0.0306534f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_191 N_B1_c_221_n N_A_219_387#_c_277_n 0.00486294f $X=3.025 $Y=1.61 $X2=0
+ $Y2=0
cc_192 N_B1_M1010_g N_A_219_387#_c_278_n 0.00229365f $X=2.44 $Y=0.945 $X2=0
+ $Y2=0
cc_193 N_B1_M1019_g N_A_219_387#_c_278_n 0.00147096f $X=2.87 $Y=0.945 $X2=0
+ $Y2=0
cc_194 B1 N_A_219_387#_c_278_n 0.0206608f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_195 N_B1_c_221_n N_A_219_387#_c_278_n 0.00283411f $X=3.025 $Y=1.61 $X2=0
+ $Y2=0
cc_196 N_B1_M1008_g N_A_219_387#_c_312_n 0.0185742f $X=3.025 $Y=2.355 $X2=0
+ $Y2=0
cc_197 B1 N_A_219_387#_c_312_n 0.021363f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_198 N_B1_M1008_g N_A_219_387#_c_279_n 0.00344322f $X=3.025 $Y=2.355 $X2=0
+ $Y2=0
cc_199 B1 N_A_219_387#_c_279_n 0.0193018f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_200 N_B1_c_221_n N_A_219_387#_c_279_n 6.43806e-19 $X=3.025 $Y=1.61 $X2=0
+ $Y2=0
cc_201 N_B1_M1000_g N_A_219_387#_c_288_n 0.0113021f $X=2.495 $Y=2.355 $X2=0
+ $Y2=0
cc_202 N_B1_M1008_g N_A_219_387#_c_288_n 0.00379271f $X=3.025 $Y=2.355 $X2=0
+ $Y2=0
cc_203 B1 N_A_219_387#_c_288_n 0.0246587f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_204 N_B1_c_221_n N_A_219_387#_c_288_n 0.00131617f $X=3.025 $Y=1.61 $X2=0
+ $Y2=0
cc_205 N_B1_M1019_g N_A_219_387#_c_281_n 0.0021086f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_206 B1 N_A_219_387#_c_281_n 0.00318495f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_207 N_B1_c_221_n N_A_219_387#_c_281_n 0.00192995f $X=3.025 $Y=1.61 $X2=0
+ $Y2=0
cc_208 N_B1_M1019_g N_A_219_387#_c_282_n 0.0043112f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_209 N_B1_c_221_n N_A_219_387#_c_282_n 0.00393369f $X=3.025 $Y=1.61 $X2=0
+ $Y2=0
cc_210 N_B1_M1000_g N_VPWR_c_417_n 0.00424048f $X=2.495 $Y=2.355 $X2=0 $Y2=0
cc_211 N_B1_M1008_g N_VPWR_c_418_n 0.00794402f $X=3.025 $Y=2.355 $X2=0 $Y2=0
cc_212 N_B1_M1000_g N_VPWR_c_422_n 0.00530844f $X=2.495 $Y=2.355 $X2=0 $Y2=0
cc_213 N_B1_M1008_g N_VPWR_c_422_n 0.00545019f $X=3.025 $Y=2.355 $X2=0 $Y2=0
cc_214 N_B1_M1000_g N_VPWR_c_414_n 0.00587053f $X=2.495 $Y=2.355 $X2=0 $Y2=0
cc_215 N_B1_M1008_g N_VPWR_c_414_n 0.00587053f $X=3.025 $Y=2.355 $X2=0 $Y2=0
cc_216 N_B1_M1010_g N_A_27_125#_c_579_n 0.00248344f $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_217 N_B1_M1010_g N_A_27_125#_c_580_n 0.00918561f $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_218 N_B1_M1019_g N_A_27_125#_c_580_n 4.92416e-19 $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_219 N_B1_M1010_g N_A_27_125#_c_581_n 0.00582977f $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_220 N_B1_M1019_g N_A_27_125#_c_581_n 0.00661564f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_221 N_B1_M1019_g N_A_27_125#_c_583_n 0.0108881f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_222 N_B1_M1010_g N_VGND_c_650_n 2.28708e-19 $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_223 N_A_219_387#_c_290_n N_VPWR_M1016_d 0.00595171f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_224 N_A_219_387#_c_312_n N_VPWR_M1008_s 0.012555f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_225 N_A_219_387#_c_279_n N_VPWR_M1008_s 0.00216561f $X=3.49 $Y=1.95 $X2=0
+ $Y2=0
cc_226 N_A_219_387#_c_290_n N_VPWR_c_417_n 0.0200142f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_227 N_A_219_387#_c_288_n N_VPWR_c_417_n 0.0197393f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_228 N_A_219_387#_M1007_g N_VPWR_c_418_n 0.0112138f $X=3.755 $Y=2.4 $X2=0
+ $Y2=0
cc_229 N_A_219_387#_c_312_n N_VPWR_c_418_n 0.032724f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_230 N_A_219_387#_c_288_n N_VPWR_c_418_n 0.00127803f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_231 N_A_219_387#_M1009_g N_VPWR_c_419_n 0.00343717f $X=4.205 $Y=2.4 $X2=0
+ $Y2=0
cc_232 N_A_219_387#_c_285_n N_VPWR_c_419_n 0.00203999f $X=4.755 $Y=1.76 $X2=0
+ $Y2=0
cc_233 N_A_219_387#_c_286_n N_VPWR_c_421_n 0.00394849f $X=5.205 $Y=1.76 $X2=0
+ $Y2=0
cc_234 N_A_219_387#_c_288_n N_VPWR_c_422_n 0.00826067f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_235 N_A_219_387#_M1007_g N_VPWR_c_425_n 0.005209f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A_219_387#_M1009_g N_VPWR_c_425_n 0.005209f $X=4.205 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_219_387#_c_285_n N_VPWR_c_426_n 0.005209f $X=4.755 $Y=1.76 $X2=0
+ $Y2=0
cc_238 N_A_219_387#_c_286_n N_VPWR_c_426_n 0.005209f $X=5.205 $Y=1.76 $X2=0
+ $Y2=0
cc_239 N_A_219_387#_M1007_g N_VPWR_c_414_n 0.00987399f $X=3.755 $Y=2.4 $X2=0
+ $Y2=0
cc_240 N_A_219_387#_M1009_g N_VPWR_c_414_n 0.00982526f $X=4.205 $Y=2.4 $X2=0
+ $Y2=0
cc_241 N_A_219_387#_c_285_n N_VPWR_c_414_n 0.00982526f $X=4.755 $Y=1.76 $X2=0
+ $Y2=0
cc_242 N_A_219_387#_c_286_n N_VPWR_c_414_n 0.00985497f $X=5.205 $Y=1.76 $X2=0
+ $Y2=0
cc_243 N_A_219_387#_c_288_n N_VPWR_c_414_n 0.0106835f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_244 N_A_219_387#_c_290_n N_A_119_387#_M1013_s 0.00638791f $X=2.565 $Y=2.035
+ $X2=0 $Y2=0
cc_245 N_A_219_387#_M1011_d N_A_119_387#_c_484_n 0.00165831f $X=1.095 $Y=1.935
+ $X2=0 $Y2=0
cc_246 N_A_219_387#_c_292_n N_A_119_387#_c_484_n 0.0159318f $X=1.23 $Y=2.115
+ $X2=0 $Y2=0
cc_247 N_A_219_387#_c_290_n N_A_119_387#_c_492_n 0.0189268f $X=2.565 $Y=2.035
+ $X2=0 $Y2=0
cc_248 N_A_219_387#_M1007_g N_X_c_508_n 0.0206522f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_219_387#_M1009_g N_X_c_508_n 0.0151125f $X=4.205 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_219_387#_c_285_n N_X_c_508_n 4.58171e-19 $X=4.755 $Y=1.76 $X2=0 $Y2=0
cc_251 N_A_219_387#_c_312_n N_X_c_508_n 0.0107656f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_252 N_A_219_387#_c_279_n N_X_c_508_n 0.00334168f $X=3.49 $Y=1.95 $X2=0 $Y2=0
cc_253 N_A_219_387#_c_271_n N_X_c_518_n 0.00219545f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_254 N_A_219_387#_c_280_n N_X_c_518_n 0.0190038f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_255 N_A_219_387#_c_282_n N_X_c_518_n 6.9034e-19 $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_256 N_A_219_387#_c_271_n N_X_c_504_n 0.00638907f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_257 N_A_219_387#_c_273_n N_X_c_504_n 4.40427e-19 $X=4.37 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A_219_387#_M1009_g N_X_c_509_n 0.0134861f $X=4.205 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A_219_387#_c_285_n N_X_c_509_n 0.0102903f $X=4.755 $Y=1.76 $X2=0 $Y2=0
cc_260 N_A_219_387#_c_280_n N_X_c_509_n 0.0482544f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_261 N_A_219_387#_c_282_n N_X_c_509_n 0.00859809f $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_262 N_A_219_387#_M1007_g N_X_c_510_n 0.00408731f $X=3.755 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A_219_387#_M1009_g N_X_c_510_n 0.00228751f $X=4.205 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_219_387#_c_279_n N_X_c_510_n 0.0103981f $X=3.49 $Y=1.95 $X2=0 $Y2=0
cc_265 N_A_219_387#_c_280_n N_X_c_510_n 0.0278089f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_266 N_A_219_387#_c_282_n N_X_c_510_n 0.00245159f $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_267 N_A_219_387#_c_273_n N_X_c_532_n 0.0097547f $X=4.37 $Y=1.22 $X2=0 $Y2=0
cc_268 N_A_219_387#_c_274_n N_X_c_532_n 0.0132906f $X=4.835 $Y=1.22 $X2=0 $Y2=0
cc_269 N_A_219_387#_c_280_n N_X_c_532_n 0.0363197f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_270 N_A_219_387#_c_282_n N_X_c_532_n 8.33715e-19 $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_271 N_A_219_387#_M1009_g N_X_c_511_n 4.58171e-19 $X=4.205 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A_219_387#_c_285_n N_X_c_511_n 0.0151125f $X=4.755 $Y=1.76 $X2=0 $Y2=0
cc_273 N_A_219_387#_c_286_n N_X_c_511_n 0.0157899f $X=5.205 $Y=1.76 $X2=0 $Y2=0
cc_274 N_A_219_387#_c_274_n N_X_c_505_n 3.92313e-19 $X=4.835 $Y=1.22 $X2=0 $Y2=0
cc_275 N_A_219_387#_c_275_n N_X_c_505_n 3.92313e-19 $X=5.265 $Y=1.22 $X2=0 $Y2=0
cc_276 N_A_219_387#_c_274_n N_X_c_506_n 0.00185803f $X=4.835 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A_219_387#_c_275_n N_X_c_506_n 0.00228347f $X=5.265 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A_219_387#_c_280_n N_X_c_506_n 0.0285354f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_279 N_A_219_387#_c_282_n N_X_c_506_n 0.0249566f $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_280 N_A_219_387#_M1009_g N_X_c_545_n 6.05255e-19 $X=4.205 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A_219_387#_c_285_n N_X_c_545_n 0.00126234f $X=4.755 $Y=1.76 $X2=0 $Y2=0
cc_282 N_A_219_387#_c_286_n N_X_c_545_n 0.0062293f $X=5.205 $Y=1.76 $X2=0 $Y2=0
cc_283 N_A_219_387#_c_282_n N_X_c_545_n 0.0185479f $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_284 N_A_219_387#_c_286_n X 0.00745034f $X=5.205 $Y=1.76 $X2=0 $Y2=0
cc_285 N_A_219_387#_c_282_n X 0.0156723f $X=5.205 $Y=1.49 $X2=0 $Y2=0
cc_286 N_A_219_387#_c_277_n N_A_27_125#_M1019_d 0.00396376f $X=3.405 $Y=1.26
+ $X2=0 $Y2=0
cc_287 N_A_219_387#_c_290_n N_A_27_125#_c_579_n 0.00993827f $X=2.565 $Y=2.035
+ $X2=0 $Y2=0
cc_288 N_A_219_387#_c_278_n N_A_27_125#_c_579_n 0.00444516f $X=2.82 $Y=1.26
+ $X2=0 $Y2=0
cc_289 N_A_219_387#_c_276_n N_A_27_125#_c_580_n 0.0186128f $X=2.655 $Y=0.77
+ $X2=0 $Y2=0
cc_290 N_A_219_387#_c_276_n N_A_27_125#_c_581_n 0.0195392f $X=2.655 $Y=0.77
+ $X2=0 $Y2=0
cc_291 N_A_219_387#_c_276_n N_A_27_125#_c_583_n 0.0144986f $X=2.655 $Y=0.77
+ $X2=0 $Y2=0
cc_292 N_A_219_387#_c_277_n N_A_27_125#_c_583_n 0.0266632f $X=3.405 $Y=1.26
+ $X2=0 $Y2=0
cc_293 N_A_219_387#_c_271_n N_VGND_c_644_n 0.00340257f $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_294 N_A_219_387#_c_280_n N_VGND_c_644_n 0.0203976f $X=4.63 $Y=1.385 $X2=0
+ $Y2=0
cc_295 N_A_219_387#_c_281_n N_VGND_c_644_n 0.00131156f $X=3.49 $Y=1.362 $X2=0
+ $Y2=0
cc_296 N_A_219_387#_c_282_n N_VGND_c_644_n 0.00174273f $X=5.205 $Y=1.49 $X2=0
+ $Y2=0
cc_297 N_A_219_387#_c_271_n N_VGND_c_645_n 3.93623e-19 $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_298 N_A_219_387#_c_273_n N_VGND_c_645_n 0.00765879f $X=4.37 $Y=1.22 $X2=0
+ $Y2=0
cc_299 N_A_219_387#_c_274_n N_VGND_c_645_n 0.00768892f $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_300 N_A_219_387#_c_275_n N_VGND_c_645_n 4.1905e-19 $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_301 N_A_219_387#_c_274_n N_VGND_c_647_n 4.70441e-19 $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_302 N_A_219_387#_c_275_n N_VGND_c_647_n 0.0150633f $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_303 N_A_219_387#_c_271_n N_VGND_c_651_n 0.00433834f $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_304 N_A_219_387#_c_273_n N_VGND_c_651_n 0.00383152f $X=4.37 $Y=1.22 $X2=0
+ $Y2=0
cc_305 N_A_219_387#_c_274_n N_VGND_c_652_n 0.00383152f $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_306 N_A_219_387#_c_275_n N_VGND_c_652_n 0.00383152f $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_307 N_A_219_387#_c_271_n N_VGND_c_657_n 0.00824977f $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_308 N_A_219_387#_c_273_n N_VGND_c_657_n 0.00382921f $X=4.37 $Y=1.22 $X2=0
+ $Y2=0
cc_309 N_A_219_387#_c_274_n N_VGND_c_657_n 0.00382921f $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_310 N_A_219_387#_c_275_n N_VGND_c_657_n 0.0075754f $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_417_n N_A_119_387#_c_484_n 0.0130139f $X=2.23 $Y=2.455 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_424_n N_A_119_387#_c_484_n 0.0686911f $X=2.065 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_414_n N_A_119_387#_c_484_n 0.0391401f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_416_n N_A_119_387#_c_485_n 0.0129305f $X=0.28 $Y=2.08 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_424_n N_A_119_387#_c_485_n 0.0179217f $X=2.065 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_414_n N_A_119_387#_c_485_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_418_n N_X_c_508_n 0.023149f $X=3.36 $Y=2.465 $X2=0 $Y2=0
cc_318 N_VPWR_c_419_n N_X_c_508_n 0.0353111f $X=4.48 $Y=2.145 $X2=0 $Y2=0
cc_319 N_VPWR_c_425_n N_X_c_508_n 0.0144623f $X=4.315 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_c_414_n N_X_c_508_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_321 N_VPWR_M1009_s N_X_c_509_n 0.00274845f $X=4.295 $Y=1.84 $X2=0 $Y2=0
cc_322 N_VPWR_c_419_n N_X_c_509_n 0.0208278f $X=4.48 $Y=2.145 $X2=0 $Y2=0
cc_323 N_VPWR_c_419_n N_X_c_511_n 0.0353111f $X=4.48 $Y=2.145 $X2=0 $Y2=0
cc_324 N_VPWR_c_421_n N_X_c_511_n 0.0394385f $X=5.48 $Y=2.115 $X2=0 $Y2=0
cc_325 N_VPWR_c_426_n N_X_c_511_n 0.0144623f $X=5.315 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_c_414_n N_X_c_511_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_421_n X 0.0253467f $X=5.48 $Y=2.115 $X2=0 $Y2=0
cc_328 N_VPWR_c_416_n N_A_27_125#_c_577_n 0.0120242f $X=0.28 $Y=2.08 $X2=0 $Y2=0
cc_329 N_A_119_387#_c_486_n N_A_27_125#_c_576_n 0.00607566f $X=0.78 $Y=2.115
+ $X2=0 $Y2=0
cc_330 N_X_c_532_n N_VGND_M1002_d 0.00395842f $X=4.965 $Y=0.92 $X2=0 $Y2=0
cc_331 N_X_c_504_n N_VGND_c_644_n 0.0188059f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_332 N_X_c_504_n N_VGND_c_645_n 0.0136878f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_333 N_X_c_532_n N_VGND_c_645_n 0.0194786f $X=4.965 $Y=0.92 $X2=0 $Y2=0
cc_334 N_X_c_505_n N_VGND_c_645_n 0.0121521f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_335 N_X_c_505_n N_VGND_c_647_n 0.0180696f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_336 N_X_c_506_n N_VGND_c_647_n 0.00516673f $X=5.05 $Y=1.55 $X2=0 $Y2=0
cc_337 X N_VGND_c_647_n 0.0145768f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_338 N_X_c_504_n N_VGND_c_651_n 0.0119488f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_339 N_X_c_505_n N_VGND_c_652_n 0.00749631f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_340 N_X_c_504_n N_VGND_c_657_n 0.00915121f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_341 N_X_c_532_n N_VGND_c_657_n 0.0118272f $X=4.965 $Y=0.92 $X2=0 $Y2=0
cc_342 N_X_c_505_n N_VGND_c_657_n 0.0062048f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_343 N_A_27_125#_c_576_n N_VGND_M1015_d 0.00256188f $X=1.13 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_344 N_A_27_125#_c_579_n N_VGND_M1004_s 0.00397519f $X=2.06 $Y=1.19 $X2=0
+ $Y2=0
cc_345 N_A_27_125#_c_575_n N_VGND_c_642_n 0.0131747f $X=0.28 $Y=0.77 $X2=0 $Y2=0
cc_346 N_A_27_125#_c_576_n N_VGND_c_642_n 0.0213935f $X=1.13 $Y=1.19 $X2=0 $Y2=0
cc_347 N_A_27_125#_c_578_n N_VGND_c_642_n 0.0125829f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_348 N_A_27_125#_c_578_n N_VGND_c_643_n 0.0120942f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_349 N_A_27_125#_c_579_n N_VGND_c_643_n 0.0257093f $X=2.06 $Y=1.19 $X2=0 $Y2=0
cc_350 N_A_27_125#_c_580_n N_VGND_c_643_n 0.0265871f $X=2.225 $Y=0.77 $X2=0
+ $Y2=0
cc_351 N_A_27_125#_c_582_n N_VGND_c_643_n 0.0142636f $X=2.39 $Y=0.35 $X2=0 $Y2=0
cc_352 N_A_27_125#_c_581_n N_VGND_c_644_n 0.0119252f $X=3 $Y=0.35 $X2=0 $Y2=0
cc_353 N_A_27_125#_c_583_n N_VGND_c_644_n 0.0376042f $X=3.165 $Y=0.805 $X2=0
+ $Y2=0
cc_354 N_A_27_125#_c_575_n N_VGND_c_648_n 0.00702137f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_355 N_A_27_125#_c_578_n N_VGND_c_649_n 0.00528099f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_356 N_A_27_125#_c_581_n N_VGND_c_650_n 0.0591825f $X=3 $Y=0.35 $X2=0 $Y2=0
cc_357 N_A_27_125#_c_582_n N_VGND_c_650_n 0.0221635f $X=2.39 $Y=0.35 $X2=0 $Y2=0
cc_358 N_A_27_125#_c_575_n N_VGND_c_657_n 0.0100521f $X=0.28 $Y=0.77 $X2=0 $Y2=0
cc_359 N_A_27_125#_c_578_n N_VGND_c_657_n 0.00668051f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_360 N_A_27_125#_c_581_n N_VGND_c_657_n 0.035558f $X=3 $Y=0.35 $X2=0 $Y2=0
cc_361 N_A_27_125#_c_582_n N_VGND_c_657_n 0.0126536f $X=2.39 $Y=0.35 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dfbbn_1.pxi.spice
* Created: Wed Sep  2 12:02:22 2020
* 
x_PM_SKY130_FD_SC_MS__DFBBN_1%CLK_N N_CLK_N_M1030_g N_CLK_N_M1035_g CLK_N
+ N_CLK_N_c_281_n N_CLK_N_c_282_n PM_SKY130_FD_SC_MS__DFBBN_1%CLK_N
x_PM_SKY130_FD_SC_MS__DFBBN_1%D N_D_M1014_g N_D_M1017_g D D N_D_c_316_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%D
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_474_405# N_A_474_405#_M1020_d
+ N_A_474_405#_M1021_s N_A_474_405#_M1013_d N_A_474_405#_M1010_g
+ N_A_474_405#_M1006_g N_A_474_405#_M1024_g N_A_474_405#_M1007_g
+ N_A_474_405#_c_362_n N_A_474_405#_c_363_n N_A_474_405#_c_364_n
+ N_A_474_405#_c_365_n N_A_474_405#_c_356_n N_A_474_405#_c_357_n
+ N_A_474_405#_c_430_p N_A_474_405#_c_367_n N_A_474_405#_c_368_n
+ N_A_474_405#_c_369_n N_A_474_405#_c_370_n N_A_474_405#_c_371_n
+ N_A_474_405#_c_372_n N_A_474_405#_c_373_n N_A_474_405#_c_358_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_474_405#
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_200_74# N_A_200_74#_M1036_d N_A_200_74#_M1031_d
+ N_A_200_74#_M1015_g N_A_200_74#_M1005_g N_A_200_74#_M1038_g
+ N_A_200_74#_c_533_n N_A_200_74#_M1022_g N_A_200_74#_c_550_n
+ N_A_200_74#_c_534_n N_A_200_74#_c_551_n N_A_200_74#_c_552_n
+ N_A_200_74#_c_553_n N_A_200_74#_c_554_n N_A_200_74#_c_568_n
+ N_A_200_74#_c_535_n N_A_200_74#_c_555_n N_A_200_74#_c_556_n
+ N_A_200_74#_c_536_n N_A_200_74#_c_537_n N_A_200_74#_c_538_n
+ N_A_200_74#_c_539_n N_A_200_74#_c_559_n N_A_200_74#_c_540_n
+ N_A_200_74#_c_541_n N_A_200_74#_c_561_n N_A_200_74#_c_542_n
+ N_A_200_74#_c_573_n N_A_200_74#_c_543_n N_A_200_74#_c_544_n
+ N_A_200_74#_c_545_n N_A_200_74#_c_546_n N_A_200_74#_c_547_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_200_74#
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_595_119# N_A_595_119#_M1001_d
+ N_A_595_119#_M1015_d N_A_595_119#_c_761_n N_A_595_119#_M1021_g
+ N_A_595_119#_M1020_g N_A_595_119#_c_764_n N_A_595_119#_c_781_n
+ N_A_595_119#_c_789_n N_A_595_119#_c_770_n N_A_595_119#_c_765_n
+ N_A_595_119#_c_766_n N_A_595_119#_c_767_n N_A_595_119#_c_768_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_595_119#
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_978_357# N_A_978_357#_M1008_s
+ N_A_978_357#_M1011_s N_A_978_357#_c_867_n N_A_978_357#_M1003_g
+ N_A_978_357#_M1032_g N_A_978_357#_M1034_g N_A_978_357#_M1019_g
+ N_A_978_357#_c_870_n N_A_978_357#_c_871_n N_A_978_357#_c_872_n
+ N_A_978_357#_c_873_n N_A_978_357#_c_874_n N_A_978_357#_c_928_p
+ N_A_978_357#_c_960_p N_A_978_357#_c_875_n N_A_978_357#_c_876_n
+ N_A_978_357#_c_877_n N_A_978_357#_c_878_n N_A_978_357#_c_879_n
+ N_A_978_357#_c_887_n N_A_978_357#_c_888_n N_A_978_357#_c_880_n
+ N_A_978_357#_c_957_p N_A_978_357#_c_881_n N_A_978_357#_c_882_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_978_357#
x_PM_SKY130_FD_SC_MS__DFBBN_1%SET_B N_SET_B_c_1053_n N_SET_B_M1013_g
+ N_SET_B_M1027_g N_SET_B_c_1048_n N_SET_B_M1025_g N_SET_B_M1016_g
+ N_SET_B_c_1055_n N_SET_B_c_1068_n SET_B N_SET_B_c_1051_n N_SET_B_c_1057_n
+ N_SET_B_c_1052_n PM_SKY130_FD_SC_MS__DFBBN_1%SET_B
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_27_74# N_A_27_74#_M1035_s N_A_27_74#_M1030_s
+ N_A_27_74#_M1036_g N_A_27_74#_M1031_g N_A_27_74#_c_1181_n N_A_27_74#_c_1182_n
+ N_A_27_74#_M1001_g N_A_27_74#_c_1184_n N_A_27_74#_c_1198_n N_A_27_74#_c_1199_n
+ N_A_27_74#_c_1200_n N_A_27_74#_M1012_g N_A_27_74#_M1028_g N_A_27_74#_c_1186_n
+ N_A_27_74#_c_1187_n N_A_27_74#_c_1202_n N_A_27_74#_M1018_g N_A_27_74#_c_1188_n
+ N_A_27_74#_c_1204_n N_A_27_74#_c_1189_n N_A_27_74#_c_1206_n
+ N_A_27_74#_c_1207_n N_A_27_74#_c_1190_n N_A_27_74#_c_1191_n
+ N_A_27_74#_c_1192_n N_A_27_74#_c_1221_n N_A_27_74#_c_1193_n
+ N_A_27_74#_c_1194_n N_A_27_74#_c_1195_n N_A_27_74#_c_1196_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_27_74#
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_1534_446# N_A_1534_446#_M1034_d
+ N_A_1534_446#_M1025_s N_A_1534_446#_M1026_d N_A_1534_446#_M1023_g
+ N_A_1534_446#_M1000_g N_A_1534_446#_M1004_g N_A_1534_446#_M1029_g
+ N_A_1534_446#_c_1366_n N_A_1534_446#_c_1367_n N_A_1534_446#_c_1368_n
+ N_A_1534_446#_c_1380_n N_A_1534_446#_M1039_g N_A_1534_446#_c_1369_n
+ N_A_1534_446#_M1002_g N_A_1534_446#_c_1370_n N_A_1534_446#_c_1371_n
+ N_A_1534_446#_c_1381_n N_A_1534_446#_c_1382_n N_A_1534_446#_c_1499_p
+ N_A_1534_446#_c_1383_n N_A_1534_446#_c_1372_n N_A_1534_446#_c_1384_n
+ N_A_1534_446#_c_1385_n N_A_1534_446#_c_1386_n N_A_1534_446#_c_1387_n
+ N_A_1534_446#_c_1388_n N_A_1534_446#_c_1389_n N_A_1534_446#_c_1373_n
+ N_A_1534_446#_c_1374_n N_A_1534_446#_c_1375_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_1534_446#
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_1349_114# N_A_1349_114#_M1028_d
+ N_A_1349_114#_M1038_d N_A_1349_114#_M1033_g N_A_1349_114#_M1026_g
+ N_A_1349_114#_c_1567_n N_A_1349_114#_c_1572_n N_A_1349_114#_c_1573_n
+ N_A_1349_114#_c_1574_n N_A_1349_114#_c_1568_n N_A_1349_114#_c_1576_n
+ N_A_1349_114#_c_1577_n N_A_1349_114#_c_1647_n N_A_1349_114#_c_1578_n
+ N_A_1349_114#_c_1651_n N_A_1349_114#_c_1579_n N_A_1349_114#_c_1580_n
+ N_A_1349_114#_c_1569_n N_A_1349_114#_c_1570_n N_A_1349_114#_c_1583_n
+ N_A_1349_114#_c_1584_n N_A_1349_114#_c_1585_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_1349_114#
x_PM_SKY130_FD_SC_MS__DFBBN_1%RESET_B N_RESET_B_M1011_g N_RESET_B_M1008_g
+ RESET_B N_RESET_B_c_1720_n N_RESET_B_c_1721_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%RESET_B
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_2412_410# N_A_2412_410#_M1002_s
+ N_A_2412_410#_M1039_s N_A_2412_410#_M1037_g N_A_2412_410#_M1009_g
+ N_A_2412_410#_c_1758_n N_A_2412_410#_c_1759_n N_A_2412_410#_c_1760_n
+ N_A_2412_410#_c_1761_n N_A_2412_410#_c_1762_n N_A_2412_410#_c_1763_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_2412_410#
x_PM_SKY130_FD_SC_MS__DFBBN_1%VPWR N_VPWR_M1030_d N_VPWR_M1017_d N_VPWR_M1003_d
+ N_VPWR_M1007_s N_VPWR_M1023_d N_VPWR_M1025_d N_VPWR_M1011_d N_VPWR_M1039_d
+ N_VPWR_c_1813_n N_VPWR_c_1814_n N_VPWR_c_1815_n N_VPWR_c_1816_n
+ N_VPWR_c_1817_n N_VPWR_c_1818_n N_VPWR_c_1819_n N_VPWR_c_1820_n
+ N_VPWR_c_1821_n N_VPWR_c_1822_n VPWR N_VPWR_c_1823_n N_VPWR_c_1824_n
+ N_VPWR_c_1825_n N_VPWR_c_1826_n N_VPWR_c_1827_n N_VPWR_c_1828_n
+ N_VPWR_c_1829_n N_VPWR_c_1812_n N_VPWR_c_1831_n N_VPWR_c_1832_n
+ N_VPWR_c_1833_n N_VPWR_c_1834_n N_VPWR_c_1835_n N_VPWR_c_1836_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%VPWR
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_311_119# N_A_311_119#_M1014_s
+ N_A_311_119#_M1005_d N_A_311_119#_M1017_s N_A_311_119#_M1012_d
+ N_A_311_119#_c_1985_n N_A_311_119#_c_1969_n N_A_311_119#_c_1970_n
+ N_A_311_119#_c_1971_n N_A_311_119#_c_1972_n N_A_311_119#_c_1979_n
+ N_A_311_119#_c_1973_n N_A_311_119#_c_1980_n N_A_311_119#_c_1981_n
+ N_A_311_119#_c_1974_n N_A_311_119#_c_1975_n N_A_311_119#_c_1983_n
+ N_A_311_119#_c_1976_n N_A_311_119#_c_1977_n N_A_311_119#_c_1978_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_311_119#
x_PM_SKY130_FD_SC_MS__DFBBN_1%Q_N N_Q_N_M1029_d N_Q_N_M1004_d N_Q_N_c_2097_n
+ N_Q_N_c_2098_n Q_N Q_N Q_N Q_N N_Q_N_c_2099_n PM_SKY130_FD_SC_MS__DFBBN_1%Q_N
x_PM_SKY130_FD_SC_MS__DFBBN_1%Q N_Q_M1009_d N_Q_M1037_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__DFBBN_1%Q
x_PM_SKY130_FD_SC_MS__DFBBN_1%VGND N_VGND_M1035_d N_VGND_M1014_d N_VGND_M1027_d
+ N_VGND_M1000_d N_VGND_M1008_d N_VGND_M1002_d N_VGND_c_2147_n N_VGND_c_2148_n
+ N_VGND_c_2149_n N_VGND_c_2150_n N_VGND_c_2151_n N_VGND_c_2152_n VGND
+ N_VGND_c_2153_n N_VGND_c_2154_n N_VGND_c_2155_n N_VGND_c_2156_n
+ N_VGND_c_2157_n N_VGND_c_2158_n N_VGND_c_2159_n N_VGND_c_2160_n
+ N_VGND_c_2161_n N_VGND_c_2162_n N_VGND_c_2163_n N_VGND_c_2164_n
+ N_VGND_c_2165_n N_VGND_c_2166_n PM_SKY130_FD_SC_MS__DFBBN_1%VGND
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_867_119# N_A_867_119#_M1020_s
+ N_A_867_119#_M1032_d N_A_867_119#_c_2279_n N_A_867_119#_c_2280_n
+ N_A_867_119#_c_2281_n N_A_867_119#_c_2282_n
+ PM_SKY130_FD_SC_MS__DFBBN_1%A_867_119#
x_PM_SKY130_FD_SC_MS__DFBBN_1%A_1818_76# N_A_1818_76#_M1016_d
+ N_A_1818_76#_M1033_d N_A_1818_76#_c_2315_n N_A_1818_76#_c_2311_n
+ N_A_1818_76#_c_2312_n PM_SKY130_FD_SC_MS__DFBBN_1%A_1818_76#
cc_1 VNB N_CLK_N_M1030_g 0.00192268f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_CLK_N_M1035_g 0.0292041f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_CLK_N_c_281_n 0.016346f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_4 VNB N_CLK_N_c_282_n 0.0441412f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_5 VNB N_D_M1014_g 0.0216814f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_D_M1017_g 0.00955404f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_7 VNB D 0.00815265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D_c_316_n 0.0419609f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.465
cc_9 VNB N_A_474_405#_M1010_g 0.0386017f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_10 VNB N_A_474_405#_M1024_g 0.0371582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_474_405#_c_356_n 0.001941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_474_405#_c_357_n 0.00390787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_474_405#_c_358_n 0.00828115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_200_74#_c_533_n 0.0207162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_200_74#_c_534_n 0.0109425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_200_74#_c_535_n 0.00448218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_200_74#_c_536_n 0.00350452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_200_74#_c_537_n 0.00156732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_200_74#_c_538_n 0.00800419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_200_74#_c_539_n 0.0113538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_200_74#_c_540_n 0.00999574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_200_74#_c_541_n 0.00789892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_200_74#_c_542_n 0.0410328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_200_74#_c_543_n 0.0020871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_200_74#_c_544_n 0.0334343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_200_74#_c_545_n 0.00271411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_200_74#_c_546_n 0.0161806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_200_74#_c_547_n 0.0432725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_595_119#_c_761_n 0.0253592f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_30 VNB N_A_595_119#_M1021_g 0.00607878f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_31 VNB N_A_595_119#_M1020_g 0.0255867f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_32 VNB N_A_595_119#_c_764_n 0.0125574f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.465
cc_33 VNB N_A_595_119#_c_765_n 0.00722226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_595_119#_c_766_n 0.00105081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_595_119#_c_767_n 0.00780945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_595_119#_c_768_n 0.0276674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_978_357#_c_867_n 0.0279397f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_38 VNB N_A_978_357#_M1032_g 0.0200752f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_39 VNB N_A_978_357#_M1019_g 0.00600683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_978_357#_c_870_n 0.0147484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_978_357#_c_871_n 0.00469357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_978_357#_c_872_n 0.044764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_978_357#_c_873_n 0.00290409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_978_357#_c_874_n 0.00330882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_978_357#_c_875_n 0.00430743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_978_357#_c_876_n 0.0320601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_978_357#_c_877_n 9.45324e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_978_357#_c_878_n 0.0128172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_978_357#_c_879_n 0.00393056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_978_357#_c_880_n 4.53958e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_978_357#_c_881_n 0.0026653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_978_357#_c_882_n 0.0144593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_SET_B_M1027_g 0.0344333f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_54 VNB N_SET_B_c_1048_n 0.0354235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SET_B_M1025_g 0.00426394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_SET_B_M1016_g 0.0183433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SET_B_c_1051_n 0.00645524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_1052_n 0.00175833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_74#_M1036_g 0.0194417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_74#_M1031_g 0.00176691f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_61 VNB N_A_27_74#_c_1181_n 0.131917f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_62 VNB N_A_27_74#_c_1182_n 0.0113774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_74#_M1001_g 0.047777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_74#_c_1184_n 0.274447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_27_74#_M1028_g 0.0303562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_27_74#_c_1186_n 0.0403591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_27_74#_c_1187_n 0.0092319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_74#_c_1188_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_27_74#_c_1189_n 0.0182231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_27_74#_c_1190_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_74#_c_1191_n 0.00333636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_27_74#_c_1192_n 0.00916851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_27_74#_c_1193_n 0.00330574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_27_74#_c_1194_n 7.77832e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_27_74#_c_1195_n 0.00267069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_27_74#_c_1196_n 0.0348189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1534_446#_M1000_g 0.0407631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1534_446#_M1004_g 5.51881e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1534_446#_M1029_g 0.0235282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1534_446#_c_1366_n 0.0485932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1534_446#_c_1367_n 0.0152755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1534_446#_c_1368_n 0.0014249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1534_446#_c_1369_n 0.0197433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1534_446#_c_1370_n 0.028512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1534_446#_c_1371_n 0.00915926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1534_446#_c_1372_n 0.0136932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1534_446#_c_1373_n 0.00592654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1534_446#_c_1374_n 0.0250117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1534_446#_c_1375_n 0.00271654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1349_114#_M1033_g 0.0297354f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_91 VNB N_A_1349_114#_c_1567_n 0.00203818f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.465
cc_92 VNB N_A_1349_114#_c_1568_n 0.00622688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1349_114#_c_1569_n 0.00214252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1349_114#_c_1570_n 0.02403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_RESET_B_M1008_g 0.0240606f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_96 VNB N_RESET_B_c_1720_n 0.0300376f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_97 VNB N_RESET_B_c_1721_n 0.00190844f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_98 VNB N_A_2412_410#_M1037_g 0.00565884f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_99 VNB N_A_2412_410#_M1009_g 0.0261447f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_100 VNB N_A_2412_410#_c_1758_n 0.0385407f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.465
cc_101 VNB N_A_2412_410#_c_1759_n 0.0173865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2412_410#_c_1760_n 0.0132214f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_103 VNB N_A_2412_410#_c_1761_n 0.00107535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2412_410#_c_1762_n 0.00316228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2412_410#_c_1763_n 4.95953e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VPWR_c_1812_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_311_119#_c_1969_n 0.00190227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_311_119#_c_1970_n 0.00165852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_311_119#_c_1971_n 0.00763927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_311_119#_c_1972_n 0.00381808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_311_119#_c_1973_n 0.00475828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_311_119#_c_1974_n 0.00554809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_311_119#_c_1975_n 0.00226481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_311_119#_c_1976_n 0.0127551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_311_119#_c_1977_n 0.0115642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_311_119#_c_1978_n 0.0114046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_Q_N_c_2097_n 0.00882806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_118 VNB N_Q_N_c_2098_n 0.00164555f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_119 VNB N_Q_N_c_2099_n 0.00232427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB Q 0.0550644f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_121 VNB N_VGND_c_2147_n 0.00222691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2148_n 0.00951027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2149_n 0.00588277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2150_n 0.010469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2151_n 0.0159801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2152_n 0.00938486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2153_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2154_n 0.0308837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2155_n 0.0788352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2156_n 0.0629314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2157_n 0.0530939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2158_n 0.0334456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2159_n 0.0189533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2160_n 0.679646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2161_n 0.00501873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2162_n 0.00486067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2163_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2164_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2165_n 0.00631189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2166_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_867_119#_c_2279_n 0.00536288f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_142 VNB N_A_867_119#_c_2280_n 0.016861f $X=-0.19 $Y=-0.245 $X2=0.33 $Y2=1.465
cc_143 VNB N_A_867_119#_c_2281_n 0.00260666f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_144 VNB N_A_867_119#_c_2282_n 0.00281812f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.465
cc_145 VNB N_A_1818_76#_c_2311_n 0.00162264f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_146 VNB N_A_1818_76#_c_2312_n 0.0108274f $X=-0.19 $Y=-0.245 $X2=0.33
+ $Y2=1.465
cc_147 VPB N_CLK_N_M1030_g 0.0298346f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_148 VPB N_CLK_N_c_281_n 0.00713456f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_149 VPB N_D_M1017_g 0.0625342f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_150 VPB N_A_474_405#_M1010_g 0.0200101f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_151 VPB N_A_474_405#_M1006_g 0.0205775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_474_405#_M1007_g 0.0229377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_474_405#_c_362_n 0.00179667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_474_405#_c_363_n 0.0221043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_474_405#_c_364_n 0.00131809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_474_405#_c_365_n 0.00505233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_474_405#_c_357_n 0.00409641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_474_405#_c_367_n 0.00771963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_474_405#_c_368_n 0.00775337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_474_405#_c_369_n 0.00127727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_474_405#_c_370_n 0.0289616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_474_405#_c_371_n 0.00559253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_474_405#_c_372_n 0.00211154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_474_405#_c_373_n 4.51177e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_474_405#_c_358_n 0.0285243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_200_74#_M1015_g 0.0202101f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_167 VPB N_A_200_74#_M1038_g 0.0226796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_200_74#_c_550_n 0.0105209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_200_74#_c_551_n 0.0131775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_200_74#_c_552_n 0.00384363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_200_74#_c_553_n 0.00578472f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_200_74#_c_554_n 0.0197982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_200_74#_c_555_n 0.00425894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_200_74#_c_556_n 0.0305688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_200_74#_c_537_n 0.00329882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_200_74#_c_538_n 0.020983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_200_74#_c_559_n 0.00814275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_200_74#_c_540_n 0.00300733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_200_74#_c_561_n 2.50324e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_595_119#_M1021_g 0.0384009f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_181 VPB N_A_595_119#_c_770_n 0.00552057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_595_119#_c_767_n 0.00925066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_595_119#_c_768_n 0.0137598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_978_357#_c_867_n 0.027131f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_185 VPB N_A_978_357#_M1003_g 0.022145f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_186 VPB N_A_978_357#_M1019_g 0.0321529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_978_357#_c_878_n 0.00613775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_978_357#_c_887_n 0.00376829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_978_357#_c_888_n 0.0019404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_978_357#_c_880_n 0.00225867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_SET_B_c_1053_n 0.0199227f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.63
cc_192 VPB N_SET_B_M1025_g 0.0316408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_SET_B_c_1055_n 0.0391381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_SET_B_c_1051_n 0.0433343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_SET_B_c_1057_n 0.00567459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_SET_B_c_1052_n 0.00577004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_27_74#_M1031_g 0.026269f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_198 VPB N_A_27_74#_c_1198_n 0.0382587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_27_74#_c_1199_n 0.00713209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_27_74#_c_1200_n 0.00650961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_27_74#_M1012_g 0.0376292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_27_74#_c_1202_n 0.00604079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_27_74#_M1018_g 0.0522439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_27_74#_c_1204_n 0.0135635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_27_74#_c_1189_n 0.00818693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_27_74#_c_1206_n 0.00805193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_27_74#_c_1207_n 0.0355666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_27_74#_c_1194_n 0.00273859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1534_446#_M1023_g 0.0231195f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_210 VPB N_A_1534_446#_M1000_g 0.0251063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1534_446#_M1004_g 0.0288772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1534_446#_c_1368_n 0.00788536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1534_446#_c_1380_n 0.0452438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1534_446#_c_1381_n 0.00312755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1534_446#_c_1382_n 0.0710835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1534_446#_c_1383_n 0.0167271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1534_446#_c_1384_n 0.00164807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1534_446#_c_1385_n 0.0029931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1534_446#_c_1386_n 0.012225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1534_446#_c_1387_n 0.00136877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1534_446#_c_1388_n 0.0057012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1534_446#_c_1389_n 0.00581392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1349_114#_M1026_g 0.0301341f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_224 VPB N_A_1349_114#_c_1572_n 0.00308817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1349_114#_c_1573_n 0.0111543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1349_114#_c_1574_n 0.00123654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1349_114#_c_1568_n 0.00159665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1349_114#_c_1576_n 0.00633455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1349_114#_c_1577_n 3.20591e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1349_114#_c_1578_n 0.00181786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1349_114#_c_1579_n 0.00772122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1349_114#_c_1580_n 0.00376295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1349_114#_c_1569_n 0.0015543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1349_114#_c_1570_n 0.0116337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1349_114#_c_1583_n 0.00204067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1349_114#_c_1584_n 0.00228549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1349_114#_c_1585_n 0.00124141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_RESET_B_M1011_g 0.025377f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_239 VPB N_RESET_B_c_1720_n 0.00588606f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_240 VPB N_RESET_B_c_1721_n 0.0028981f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=1.465
cc_241 VPB N_A_2412_410#_M1037_g 0.0307754f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_242 VPB N_A_2412_410#_c_1761_n 0.00725299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1813_n 0.00768638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1814_n 0.00829357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1815_n 0.00339119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1816_n 0.00893764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1817_n 0.0228529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1818_n 0.0150484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1819_n 0.0366913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1820_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1821_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1822_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1823_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1824_n 0.0637883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1825_n 0.0448912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1826_n 0.0196646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1827_n 0.0477054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1828_n 0.0329211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1829_n 0.0197489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1812_n 0.178577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1831_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1832_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1833_n 0.0151302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1834_n 0.0139326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1835_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1836_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_311_119#_c_1979_n 0.0102264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_311_119#_c_1980_n 0.0126281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_311_119#_c_1981_n 0.00421304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_311_119#_c_1974_n 0.00994381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_311_119#_c_1983_n 0.00148805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_311_119#_c_1976_n 0.0148406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB Q_N 0.00377032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB Q_N 0.0154093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_Q_N_c_2099_n 0.00191214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB Q 0.0542187f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_277 N_CLK_N_M1030_g N_A_200_74#_c_550_n 6.27877e-19 $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_278 N_CLK_N_M1030_g N_A_27_74#_M1031_g 0.0304239f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_279 N_CLK_N_M1035_g N_A_27_74#_c_1182_n 0.0271107f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_CLK_N_M1030_g N_A_27_74#_c_1206_n 8.8334e-19 $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_CLK_N_c_281_n N_A_27_74#_c_1206_n 0.0248594f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_282 N_CLK_N_c_282_n N_A_27_74#_c_1206_n 0.0011953f $X=0.495 $Y=1.465 $X2=0
+ $Y2=0
cc_283 N_CLK_N_M1030_g N_A_27_74#_c_1207_n 0.0121004f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_284 N_CLK_N_M1035_g N_A_27_74#_c_1190_n 0.00159319f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_CLK_N_M1035_g N_A_27_74#_c_1191_n 0.0145993f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_CLK_N_c_281_n N_A_27_74#_c_1191_n 0.00971403f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_287 N_CLK_N_c_282_n N_A_27_74#_c_1191_n 0.00100672f $X=0.495 $Y=1.465 $X2=0
+ $Y2=0
cc_288 N_CLK_N_c_281_n N_A_27_74#_c_1192_n 0.0209549f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_289 N_CLK_N_c_282_n N_A_27_74#_c_1192_n 0.00158295f $X=0.495 $Y=1.465 $X2=0
+ $Y2=0
cc_290 N_CLK_N_M1030_g N_A_27_74#_c_1221_n 0.0153058f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_291 N_CLK_N_c_281_n N_A_27_74#_c_1221_n 0.00433199f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_292 N_CLK_N_M1035_g N_A_27_74#_c_1193_n 0.00383463f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_CLK_N_M1030_g N_A_27_74#_c_1194_n 0.00491468f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_294 N_CLK_N_c_281_n N_A_27_74#_c_1194_n 0.0113335f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_295 N_CLK_N_c_281_n N_A_27_74#_c_1195_n 0.0267562f $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_296 N_CLK_N_c_282_n N_A_27_74#_c_1195_n 0.00233952f $X=0.495 $Y=1.465 $X2=0
+ $Y2=0
cc_297 N_CLK_N_c_281_n N_A_27_74#_c_1196_n 2.76539e-19 $X=0.33 $Y=1.465 $X2=0
+ $Y2=0
cc_298 N_CLK_N_c_282_n N_A_27_74#_c_1196_n 0.0207882f $X=0.495 $Y=1.465 $X2=0
+ $Y2=0
cc_299 N_CLK_N_M1030_g N_VPWR_c_1813_n 0.0027763f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_300 N_CLK_N_M1030_g N_VPWR_c_1823_n 0.005209f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_301 N_CLK_N_M1030_g N_VPWR_c_1812_n 0.00986083f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_302 N_CLK_N_M1035_g N_VGND_c_2147_n 0.0125189f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_303 N_CLK_N_M1035_g N_VGND_c_2153_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_304 N_CLK_N_M1035_g N_VGND_c_2160_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_305 N_D_M1014_g N_A_474_405#_M1010_g 0.0157832f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_306 N_D_M1017_g N_A_474_405#_M1010_g 0.0174461f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_307 D N_A_474_405#_M1010_g 0.013583f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_308 N_D_c_316_n N_A_474_405#_M1010_g 0.0213648f $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_309 N_D_M1017_g N_A_474_405#_M1006_g 0.0125745f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_310 N_D_M1017_g N_A_474_405#_c_362_n 2.53239e-19 $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_311 N_D_M1017_g N_A_474_405#_c_370_n 0.0156421f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_312 N_D_M1017_g N_A_474_405#_c_371_n 4.06902e-19 $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_313 N_D_M1014_g N_A_200_74#_c_534_n 0.00280927f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_314 N_D_M1017_g N_A_200_74#_c_551_n 0.0116022f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_315 N_D_M1017_g N_A_200_74#_c_553_n 0.0280504f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_316 D N_A_200_74#_c_554_n 0.0471758f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_317 N_D_c_316_n N_A_200_74#_c_554_n 0.00290311f $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_318 N_D_M1017_g N_A_200_74#_c_568_n 0.00803175f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_319 D N_A_200_74#_c_568_n 0.0133696f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_320 N_D_c_316_n N_A_200_74#_c_568_n 5.80967e-19 $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_321 D N_A_200_74#_c_535_n 0.00391807f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_322 N_D_M1017_g N_A_200_74#_c_540_n 0.00451325f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_323 D N_A_200_74#_c_573_n 0.00187865f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_324 D N_A_200_74#_c_545_n 0.0155335f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_325 N_D_M1014_g N_A_27_74#_c_1181_n 0.00999521f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_326 D N_A_27_74#_M1001_g 0.00260483f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_327 N_D_c_316_n N_A_27_74#_c_1196_n 0.00190331f $X=2.09 $Y=1.345 $X2=0 $Y2=0
cc_328 N_D_M1017_g N_VPWR_c_1814_n 0.00180709f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_329 N_D_M1017_g N_VPWR_c_1819_n 0.00115136f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_330 N_D_M1014_g N_A_311_119#_c_1985_n 0.0100459f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_331 D N_A_311_119#_c_1985_n 0.056469f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_332 N_D_c_316_n N_A_311_119#_c_1985_n 0.00624979f $X=2.09 $Y=1.345 $X2=0
+ $Y2=0
cc_333 N_D_M1014_g N_A_311_119#_c_1969_n 8.06126e-19 $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_334 N_D_M1014_g N_A_311_119#_c_1975_n 0.00774165f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_335 N_D_M1017_g N_A_311_119#_c_1983_n 0.00684398f $X=2.01 $Y=2.725 $X2=0
+ $Y2=0
cc_336 N_D_M1014_g N_A_311_119#_c_1976_n 0.0122916f $X=1.915 $Y=0.805 $X2=0
+ $Y2=0
cc_337 N_D_M1017_g N_A_311_119#_c_1976_n 0.0207313f $X=2.01 $Y=2.725 $X2=0 $Y2=0
cc_338 D N_A_311_119#_c_1976_n 0.0262098f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_339 N_D_M1014_g N_VGND_c_2148_n 0.00252054f $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_340 N_D_M1014_g N_VGND_c_2160_n 9.39239e-19 $X=1.915 $Y=0.805 $X2=0 $Y2=0
cc_341 N_A_474_405#_M1006_g N_A_200_74#_M1015_g 0.0362233f $X=2.61 $Y=2.725
+ $X2=0 $Y2=0
cc_342 N_A_474_405#_c_362_n N_A_200_74#_M1015_g 0.00696646f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_343 N_A_474_405#_c_363_n N_A_200_74#_M1015_g 0.0139274f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_344 N_A_474_405#_M1007_g N_A_200_74#_M1038_g 0.044819f $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_345 N_A_474_405#_c_368_n N_A_200_74#_M1038_g 5.44486e-19 $X=6.12 $Y=2.405
+ $X2=0 $Y2=0
cc_346 N_A_474_405#_M1010_g N_A_200_74#_c_553_n 0.00296524f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_347 N_A_474_405#_M1006_g N_A_200_74#_c_553_n 0.00116718f $X=2.61 $Y=2.725
+ $X2=0 $Y2=0
cc_348 N_A_474_405#_c_362_n N_A_200_74#_c_553_n 0.00512783f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_349 N_A_474_405#_c_370_n N_A_200_74#_c_553_n 0.0010945f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_350 N_A_474_405#_c_371_n N_A_200_74#_c_553_n 0.0192184f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_351 N_A_474_405#_M1010_g N_A_200_74#_c_554_n 0.0109769f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_352 N_A_474_405#_c_370_n N_A_200_74#_c_554_n 0.00437059f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_353 N_A_474_405#_c_371_n N_A_200_74#_c_554_n 0.0325651f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_354 N_A_474_405#_M1010_g N_A_200_74#_c_535_n 0.00178535f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_355 N_A_474_405#_M1010_g N_A_200_74#_c_555_n 0.00498597f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_356 N_A_474_405#_c_363_n N_A_200_74#_c_555_n 0.00330156f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_357 N_A_474_405#_c_370_n N_A_200_74#_c_555_n 3.0079e-19 $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_358 N_A_474_405#_c_371_n N_A_200_74#_c_555_n 0.0262565f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_359 N_A_474_405#_c_370_n N_A_200_74#_c_556_n 0.0204794f $X=2.535 $Y=2.19
+ $X2=0 $Y2=0
cc_360 N_A_474_405#_c_371_n N_A_200_74#_c_556_n 0.00217001f $X=2.72 $Y=2.19
+ $X2=0 $Y2=0
cc_361 N_A_474_405#_M1024_g N_A_200_74#_c_536_n 0.00260546f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_362 N_A_474_405#_M1024_g N_A_200_74#_c_537_n 0.00127909f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_363 N_A_474_405#_c_369_n N_A_200_74#_c_537_n 0.0137339f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_364 N_A_474_405#_c_358_n N_A_200_74#_c_537_n 0.00127078f $X=6.41 $Y=1.795
+ $X2=0 $Y2=0
cc_365 N_A_474_405#_M1024_g N_A_200_74#_c_538_n 8.87914e-19 $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_366 N_A_474_405#_c_369_n N_A_200_74#_c_538_n 0.0030664f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_367 N_A_474_405#_c_358_n N_A_200_74#_c_538_n 0.044819f $X=6.41 $Y=1.795 $X2=0
+ $Y2=0
cc_368 N_A_474_405#_M1024_g N_A_200_74#_c_542_n 0.00706397f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_369 N_A_474_405#_c_356_n N_A_200_74#_c_542_n 0.0141949f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_370 N_A_474_405#_c_357_n N_A_200_74#_c_542_n 0.0246337f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_371 N_A_474_405#_c_369_n N_A_200_74#_c_542_n 0.00188756f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_372 N_A_474_405#_c_358_n N_A_200_74#_c_542_n 3.95095e-19 $X=6.41 $Y=1.795
+ $X2=0 $Y2=0
cc_373 N_A_474_405#_M1010_g N_A_200_74#_c_545_n 6.10356e-19 $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_374 N_A_474_405#_c_363_n N_A_595_119#_M1015_d 0.00223709f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_375 N_A_474_405#_c_363_n N_A_595_119#_M1021_g 0.00596153f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_376 N_A_474_405#_c_365_n N_A_595_119#_M1021_g 0.00825489f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_377 N_A_474_405#_c_357_n N_A_595_119#_M1021_g 0.0156987f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_378 N_A_474_405#_c_372_n N_A_595_119#_M1021_g 0.0149444f $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_379 N_A_474_405#_c_356_n N_A_595_119#_M1020_g 0.00833041f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_380 N_A_474_405#_c_357_n N_A_595_119#_M1020_g 0.00448696f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_381 N_A_474_405#_c_357_n N_A_595_119#_c_764_n 0.00646074f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_382 N_A_474_405#_c_362_n N_A_595_119#_c_781_n 0.00862739f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_383 N_A_474_405#_c_363_n N_A_595_119#_c_781_n 0.0258353f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_384 N_A_474_405#_c_362_n N_A_595_119#_c_770_n 0.00561125f $X=2.72 $Y=2.905
+ $X2=0 $Y2=0
cc_385 N_A_474_405#_M1010_g N_A_595_119#_c_766_n 2.98275e-19 $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_386 N_A_474_405#_c_356_n N_A_978_357#_c_867_n 0.00382926f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_387 N_A_474_405#_c_357_n N_A_978_357#_c_867_n 0.0108324f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_388 N_A_474_405#_c_430_p N_A_978_357#_c_867_n 0.002556f $X=5.57 $Y=2.405
+ $X2=0 $Y2=0
cc_389 N_A_474_405#_c_363_n N_A_978_357#_M1003_g 4.61665e-19 $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_390 N_A_474_405#_c_365_n N_A_978_357#_M1003_g 0.00149124f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_391 N_A_474_405#_c_430_p N_A_978_357#_M1003_g 0.0165889f $X=5.57 $Y=2.405
+ $X2=0 $Y2=0
cc_392 N_A_474_405#_c_372_n N_A_978_357#_M1003_g 4.07968e-19 $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_393 N_A_474_405#_c_356_n N_A_978_357#_M1032_g 0.00781472f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_394 N_A_474_405#_c_357_n N_A_978_357#_M1032_g 0.00250793f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_395 N_A_474_405#_M1024_g N_A_978_357#_c_870_n 0.0131218f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_396 N_A_474_405#_c_369_n N_A_978_357#_c_870_n 0.0239932f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_397 N_A_474_405#_c_358_n N_A_978_357#_c_870_n 0.00671783f $X=6.41 $Y=1.795
+ $X2=0 $Y2=0
cc_398 N_A_474_405#_M1024_g N_A_978_357#_c_871_n 0.00762346f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_399 N_A_474_405#_M1024_g N_A_978_357#_c_873_n 3.98045e-19 $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_400 N_A_474_405#_c_356_n N_A_978_357#_c_880_n 0.0106525f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_401 N_A_474_405#_c_357_n N_A_978_357#_c_880_n 0.0243026f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_402 N_A_474_405#_c_430_p N_A_978_357#_c_880_n 0.00612652f $X=5.57 $Y=2.405
+ $X2=0 $Y2=0
cc_403 N_A_474_405#_c_430_p N_SET_B_c_1053_n 0.0120221f $X=5.57 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_404 N_A_474_405#_c_367_n N_SET_B_c_1053_n 8.70751e-19 $X=5.655 $Y=2.815
+ $X2=-0.19 $Y2=-0.245
cc_405 N_A_474_405#_c_369_n N_SET_B_c_1053_n 0.00337195f $X=6.285 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_406 N_A_474_405#_M1024_g N_SET_B_M1027_g 0.0322389f $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_407 N_A_474_405#_c_356_n N_SET_B_M1027_g 5.41739e-19 $X=4.73 $Y=1.165 $X2=0
+ $Y2=0
cc_408 N_A_474_405#_M1007_g N_SET_B_c_1055_n 0.00374287f $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_409 N_A_474_405#_c_368_n N_SET_B_c_1055_n 0.0124917f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_410 N_A_474_405#_c_369_n N_SET_B_c_1055_n 0.0263837f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_411 N_A_474_405#_c_373_n N_SET_B_c_1055_n 0.00435015f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_412 N_A_474_405#_M1013_d N_SET_B_c_1068_n 0.00108665f $X=5.52 $Y=2.12 $X2=0
+ $Y2=0
cc_413 N_A_474_405#_c_357_n N_SET_B_c_1068_n 0.00473289f $X=4.73 $Y=2.305 $X2=0
+ $Y2=0
cc_414 N_A_474_405#_c_430_p N_SET_B_c_1068_n 0.00339232f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_415 N_A_474_405#_c_369_n N_SET_B_c_1068_n 0.00140895f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_416 N_A_474_405#_c_373_n N_SET_B_c_1068_n 0.00151694f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_417 N_A_474_405#_M1007_g N_SET_B_c_1051_n 0.00158978f $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_418 N_A_474_405#_c_368_n N_SET_B_c_1051_n 4.6316e-19 $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_419 N_A_474_405#_c_369_n N_SET_B_c_1051_n 8.65118e-19 $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_420 N_A_474_405#_c_373_n N_SET_B_c_1051_n 0.00360162f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_421 N_A_474_405#_c_358_n N_SET_B_c_1051_n 0.0159875f $X=6.41 $Y=1.795 $X2=0
+ $Y2=0
cc_422 N_A_474_405#_M1013_d N_SET_B_c_1057_n 6.04948e-19 $X=5.52 $Y=2.12 $X2=0
+ $Y2=0
cc_423 N_A_474_405#_M1007_g N_SET_B_c_1057_n 4.50529e-19 $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_424 N_A_474_405#_c_357_n N_SET_B_c_1057_n 0.0108045f $X=4.73 $Y=2.305 $X2=0
+ $Y2=0
cc_425 N_A_474_405#_c_430_p N_SET_B_c_1057_n 0.00604049f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_426 N_A_474_405#_c_368_n N_SET_B_c_1057_n 6.76383e-19 $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_427 N_A_474_405#_c_369_n N_SET_B_c_1057_n 0.0190661f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_428 N_A_474_405#_c_373_n N_SET_B_c_1057_n 0.00902988f $X=5.655 $Y=2.405 $X2=0
+ $Y2=0
cc_429 N_A_474_405#_c_358_n N_SET_B_c_1057_n 0.00112543f $X=6.41 $Y=1.795 $X2=0
+ $Y2=0
cc_430 N_A_474_405#_M1010_g N_A_27_74#_c_1181_n 0.00997995f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_431 N_A_474_405#_M1010_g N_A_27_74#_M1001_g 0.0820849f $X=2.54 $Y=0.805 $X2=0
+ $Y2=0
cc_432 N_A_474_405#_M1024_g N_A_27_74#_c_1184_n 0.0103107f $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_433 N_A_474_405#_c_363_n N_A_27_74#_M1012_g 0.0151536f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_434 N_A_474_405#_c_365_n N_A_27_74#_M1012_g 0.0045774f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_435 N_A_474_405#_M1024_g N_A_27_74#_M1028_g 0.0270157f $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_436 N_A_474_405#_M1007_g N_A_1349_114#_c_1583_n 0.00269135f $X=6.41 $Y=2.54
+ $X2=0 $Y2=0
cc_437 N_A_474_405#_c_368_n N_A_1349_114#_c_1583_n 0.00689183f $X=6.12 $Y=2.405
+ $X2=0 $Y2=0
cc_438 N_A_474_405#_c_369_n N_A_1349_114#_c_1583_n 0.00834933f $X=6.285 $Y=1.795
+ $X2=0 $Y2=0
cc_439 N_A_474_405#_c_430_p N_VPWR_M1003_d 0.00440306f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_440 N_A_474_405#_c_368_n N_VPWR_M1007_s 0.0038728f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_441 N_A_474_405#_c_369_n N_VPWR_M1007_s 0.00370752f $X=6.285 $Y=1.795 $X2=0
+ $Y2=0
cc_442 N_A_474_405#_M1006_g N_VPWR_c_1814_n 0.00128727f $X=2.61 $Y=2.725 $X2=0
+ $Y2=0
cc_443 N_A_474_405#_c_364_n N_VPWR_c_1814_n 0.0124583f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_444 N_A_474_405#_c_370_n N_VPWR_c_1814_n 0.00218674f $X=2.535 $Y=2.19 $X2=0
+ $Y2=0
cc_445 N_A_474_405#_c_371_n N_VPWR_c_1814_n 0.0077177f $X=2.72 $Y=2.19 $X2=0
+ $Y2=0
cc_446 N_A_474_405#_c_363_n N_VPWR_c_1815_n 0.00551465f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_447 N_A_474_405#_c_365_n N_VPWR_c_1815_n 0.00747891f $X=4.365 $Y=2.905 $X2=0
+ $Y2=0
cc_448 N_A_474_405#_c_430_p N_VPWR_c_1815_n 0.0166513f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_449 N_A_474_405#_c_367_n N_VPWR_c_1815_n 0.0112185f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_450 N_A_474_405#_M1007_g N_VPWR_c_1816_n 0.0113495f $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_451 N_A_474_405#_c_367_n N_VPWR_c_1816_n 0.0232836f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_452 N_A_474_405#_c_368_n N_VPWR_c_1816_n 0.0221541f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_453 N_A_474_405#_c_358_n N_VPWR_c_1816_n 4.92424e-19 $X=6.41 $Y=1.795 $X2=0
+ $Y2=0
cc_454 N_A_474_405#_c_367_n N_VPWR_c_1821_n 0.0110419f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_455 N_A_474_405#_M1006_g N_VPWR_c_1824_n 0.00469973f $X=2.61 $Y=2.725 $X2=0
+ $Y2=0
cc_456 N_A_474_405#_c_363_n N_VPWR_c_1824_n 0.113093f $X=4.2 $Y=2.99 $X2=0 $Y2=0
cc_457 N_A_474_405#_c_364_n N_VPWR_c_1824_n 0.0122392f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_458 N_A_474_405#_M1007_g N_VPWR_c_1825_n 0.00460063f $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_459 N_A_474_405#_M1006_g N_VPWR_c_1812_n 0.00412354f $X=2.61 $Y=2.725 $X2=0
+ $Y2=0
cc_460 N_A_474_405#_M1007_g N_VPWR_c_1812_n 0.00608442f $X=6.41 $Y=2.54 $X2=0
+ $Y2=0
cc_461 N_A_474_405#_c_363_n N_VPWR_c_1812_n 0.0650834f $X=4.2 $Y=2.99 $X2=0
+ $Y2=0
cc_462 N_A_474_405#_c_364_n N_VPWR_c_1812_n 0.00661913f $X=2.805 $Y=2.99 $X2=0
+ $Y2=0
cc_463 N_A_474_405#_c_430_p N_VPWR_c_1812_n 0.00685445f $X=5.57 $Y=2.405 $X2=0
+ $Y2=0
cc_464 N_A_474_405#_c_367_n N_VPWR_c_1812_n 0.00915013f $X=5.655 $Y=2.815 $X2=0
+ $Y2=0
cc_465 N_A_474_405#_c_368_n N_VPWR_c_1812_n 0.0112556f $X=6.12 $Y=2.405 $X2=0
+ $Y2=0
cc_466 N_A_474_405#_c_372_n N_VPWR_c_1812_n 0.0155702f $X=4.815 $Y=2.397 $X2=0
+ $Y2=0
cc_467 N_A_474_405#_c_363_n N_A_311_119#_M1012_d 0.00496562f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_468 N_A_474_405#_M1010_g N_A_311_119#_c_1985_n 0.00932917f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_469 N_A_474_405#_M1010_g N_A_311_119#_c_1969_n 0.00804248f $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_470 N_A_474_405#_c_363_n N_A_311_119#_c_1979_n 0.0189745f $X=4.2 $Y=2.99
+ $X2=0 $Y2=0
cc_471 N_A_474_405#_c_365_n N_A_311_119#_c_1979_n 0.0178266f $X=4.365 $Y=2.905
+ $X2=0 $Y2=0
cc_472 N_A_474_405#_c_357_n N_A_311_119#_c_1979_n 0.00455379f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_473 N_A_474_405#_c_372_n N_A_311_119#_c_1979_n 0.0141436f $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_474 N_A_474_405#_M1021_s N_A_311_119#_c_1980_n 0.00237344f $X=4.235 $Y=2.12
+ $X2=0 $Y2=0
cc_475 N_A_474_405#_c_357_n N_A_311_119#_c_1980_n 0.012968f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_476 N_A_474_405#_c_372_n N_A_311_119#_c_1980_n 0.0190248f $X=4.815 $Y=2.397
+ $X2=0 $Y2=0
cc_477 N_A_474_405#_c_357_n N_A_311_119#_c_1974_n 0.0559808f $X=4.73 $Y=2.305
+ $X2=0 $Y2=0
cc_478 N_A_474_405#_M1010_g N_A_311_119#_c_1975_n 8.52988e-19 $X=2.54 $Y=0.805
+ $X2=0 $Y2=0
cc_479 N_A_474_405#_c_356_n N_A_311_119#_c_1978_n 0.0140524f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_480 N_A_474_405#_c_362_n A_540_503# 0.00432929f $X=2.72 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_481 N_A_474_405#_c_363_n A_540_503# 0.00293798f $X=4.2 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_482 N_A_474_405#_c_357_n A_936_424# 0.002337f $X=4.73 $Y=2.305 $X2=-0.19
+ $Y2=-0.245
cc_483 N_A_474_405#_c_430_p A_936_424# 9.90428e-19 $X=5.57 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_484 N_A_474_405#_c_372_n A_936_424# 0.00197235f $X=4.815 $Y=2.397 $X2=-0.19
+ $Y2=-0.245
cc_485 N_A_474_405#_M1010_g N_VGND_c_2148_n 0.00177627f $X=2.54 $Y=0.805 $X2=0
+ $Y2=0
cc_486 N_A_474_405#_M1024_g N_VGND_c_2149_n 0.00898422f $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_487 N_A_474_405#_M1010_g N_VGND_c_2160_n 7.22543e-19 $X=2.54 $Y=0.805 $X2=0
+ $Y2=0
cc_488 N_A_474_405#_M1024_g N_VGND_c_2160_n 7.88961e-19 $X=6.195 $Y=0.87 $X2=0
+ $Y2=0
cc_489 N_A_474_405#_c_356_n N_A_867_119#_c_2280_n 0.0189518f $X=4.73 $Y=1.165
+ $X2=0 $Y2=0
cc_490 N_A_474_405#_M1024_g N_A_867_119#_c_2282_n 2.31893e-19 $X=6.195 $Y=0.87
+ $X2=0 $Y2=0
cc_491 N_A_200_74#_c_542_n N_A_595_119#_M1020_g 0.00360788f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_492 N_A_200_74#_M1015_g N_A_595_119#_c_781_n 0.00314469f $X=3.03 $Y=2.725
+ $X2=0 $Y2=0
cc_493 N_A_200_74#_c_555_n N_A_595_119#_c_781_n 0.00806096f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_494 N_A_200_74#_c_556_n N_A_595_119#_c_781_n 6.62228e-19 $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_495 N_A_200_74#_c_542_n N_A_595_119#_c_789_n 0.00566444f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_496 N_A_200_74#_c_544_n N_A_595_119#_c_789_n 0.00258703f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_497 N_A_200_74#_c_545_n N_A_595_119#_c_789_n 0.010638f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_498 N_A_200_74#_c_546_n N_A_595_119#_c_789_n 0.00975616f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_499 N_A_200_74#_M1015_g N_A_595_119#_c_770_n 0.00135386f $X=3.03 $Y=2.725
+ $X2=0 $Y2=0
cc_500 N_A_200_74#_c_555_n N_A_595_119#_c_770_n 0.0375973f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_501 N_A_200_74#_c_556_n N_A_595_119#_c_770_n 0.00174016f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_502 N_A_200_74#_c_561_n N_A_595_119#_c_770_n 0.00486726f $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_503 N_A_200_74#_c_542_n N_A_595_119#_c_765_n 0.0170584f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_504 N_A_200_74#_c_573_n N_A_595_119#_c_765_n 3.53962e-19 $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_505 N_A_200_74#_c_544_n N_A_595_119#_c_765_n 0.00564507f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_506 N_A_200_74#_c_545_n N_A_595_119#_c_765_n 0.0192812f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_507 N_A_200_74#_c_546_n N_A_595_119#_c_765_n 0.00542458f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_508 N_A_200_74#_c_573_n N_A_595_119#_c_766_n 0.00201621f $X=3.265 $Y=1.295
+ $X2=0 $Y2=0
cc_509 N_A_200_74#_c_544_n N_A_595_119#_c_766_n 0.00145122f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_510 N_A_200_74#_c_545_n N_A_595_119#_c_766_n 0.0187186f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_511 N_A_200_74#_c_546_n N_A_595_119#_c_766_n 0.00905142f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_512 N_A_200_74#_c_535_n N_A_595_119#_c_767_n 0.0130684f $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_513 N_A_200_74#_c_561_n N_A_595_119#_c_767_n 0.0093116f $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_514 N_A_200_74#_c_542_n N_A_595_119#_c_767_n 0.0194182f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_515 N_A_200_74#_c_544_n N_A_595_119#_c_767_n 0.00147136f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_516 N_A_200_74#_c_545_n N_A_595_119#_c_767_n 0.00918903f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_517 N_A_200_74#_c_535_n N_A_595_119#_c_768_n 9.08222e-19 $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_518 N_A_200_74#_c_542_n N_A_595_119#_c_768_n 0.00815904f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_519 N_A_200_74#_c_544_n N_A_595_119#_c_768_n 0.00239727f $X=3.35 $Y=1.29
+ $X2=0 $Y2=0
cc_520 N_A_200_74#_c_542_n N_A_978_357#_c_867_n 0.00434659f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_521 N_A_200_74#_c_542_n N_A_978_357#_M1032_g 0.00705248f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_522 N_A_200_74#_c_536_n N_A_978_357#_c_870_n 0.0120591f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_523 N_A_200_74#_c_542_n N_A_978_357#_c_870_n 0.045746f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_524 N_A_200_74#_c_543_n N_A_978_357#_c_870_n 2.99413e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_525 N_A_200_74#_c_536_n N_A_978_357#_c_871_n 0.00817666f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_526 N_A_200_74#_c_542_n N_A_978_357#_c_871_n 0.0161182f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_527 N_A_200_74#_c_543_n N_A_978_357#_c_871_n 2.5995e-19 $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_528 N_A_200_74#_c_533_n N_A_978_357#_c_872_n 0.00449896f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_529 N_A_200_74#_c_536_n N_A_978_357#_c_872_n 2.41257e-19 $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_530 N_A_200_74#_c_533_n N_A_978_357#_c_874_n 8.23715e-19 $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_531 N_A_200_74#_c_542_n N_A_978_357#_c_880_n 0.0168823f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_532 N_A_200_74#_c_542_n N_SET_B_M1027_g 0.00712937f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_533 N_A_200_74#_M1038_g N_SET_B_c_1055_n 0.00971235f $X=6.8 $Y=2.54 $X2=0
+ $Y2=0
cc_534 N_A_200_74#_c_537_n N_SET_B_c_1055_n 0.0103776f $X=6.875 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_200_74#_c_539_n N_SET_B_c_1055_n 0.00541798f $X=7.775 $Y=1.395 $X2=0
+ $Y2=0
cc_536 N_A_200_74#_c_543_n N_SET_B_c_1055_n 0.0122618f $X=6.96 $Y=1.295 $X2=0
+ $Y2=0
cc_537 N_A_200_74#_c_542_n N_SET_B_c_1068_n 0.0113058f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_538 N_A_200_74#_c_542_n N_SET_B_c_1057_n 0.00178987f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_539 N_A_200_74#_c_534_n N_A_27_74#_M1036_g 0.00206053f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_540 N_A_200_74#_c_540_n N_A_27_74#_M1036_g 0.00235546f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_541 N_A_200_74#_c_550_n N_A_27_74#_M1031_g 0.0126543f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_542 N_A_200_74#_c_552_n N_A_27_74#_M1031_g 0.00494528f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_543 N_A_200_74#_c_559_n N_A_27_74#_M1031_g 0.0031331f $X=1.17 $Y=1.985 $X2=0
+ $Y2=0
cc_544 N_A_200_74#_c_540_n N_A_27_74#_M1031_g 0.00296813f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_545 N_A_200_74#_c_534_n N_A_27_74#_c_1181_n 0.00766647f $X=1.14 $Y=0.515
+ $X2=0 $Y2=0
cc_546 N_A_200_74#_c_535_n N_A_27_74#_M1001_g 0.00420477f $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_547 N_A_200_74#_c_544_n N_A_27_74#_M1001_g 0.0213331f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_548 N_A_200_74#_c_545_n N_A_27_74#_M1001_g 0.00378881f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_549 N_A_200_74#_c_546_n N_A_27_74#_M1001_g 0.0126333f $X=3.35 $Y=1.125 $X2=0
+ $Y2=0
cc_550 N_A_200_74#_c_546_n N_A_27_74#_c_1184_n 0.00882199f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_551 N_A_200_74#_c_535_n N_A_27_74#_c_1198_n 0.00537991f $X=3.107 $Y=1.685
+ $X2=0 $Y2=0
cc_552 N_A_200_74#_c_561_n N_A_27_74#_c_1198_n 0.00745509f $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_553 N_A_200_74#_c_544_n N_A_27_74#_c_1198_n 0.0217028f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_554 N_A_200_74#_c_545_n N_A_27_74#_c_1198_n 0.00215493f $X=3.35 $Y=1.29 $X2=0
+ $Y2=0
cc_555 N_A_200_74#_c_554_n N_A_27_74#_c_1199_n 0.0109949f $X=2.975 $Y=1.77 $X2=0
+ $Y2=0
cc_556 N_A_200_74#_c_556_n N_A_27_74#_c_1199_n 0.0213645f $X=3.075 $Y=2.19 $X2=0
+ $Y2=0
cc_557 N_A_200_74#_c_555_n N_A_27_74#_c_1200_n 3.84179e-19 $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_558 N_A_200_74#_c_556_n N_A_27_74#_c_1200_n 0.0205307f $X=3.075 $Y=2.19 $X2=0
+ $Y2=0
cc_559 N_A_200_74#_M1015_g N_A_27_74#_M1012_g 0.0137018f $X=3.03 $Y=2.725 $X2=0
+ $Y2=0
cc_560 N_A_200_74#_c_536_n N_A_27_74#_M1028_g 0.00117954f $X=6.892 $Y=1.56 $X2=0
+ $Y2=0
cc_561 N_A_200_74#_c_533_n N_A_27_74#_c_1186_n 5.75074e-19 $X=7.98 $Y=1.23 $X2=0
+ $Y2=0
cc_562 N_A_200_74#_c_536_n N_A_27_74#_c_1186_n 0.0132432f $X=6.892 $Y=1.56 $X2=0
+ $Y2=0
cc_563 N_A_200_74#_c_539_n N_A_27_74#_c_1186_n 0.0139078f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_564 N_A_200_74#_c_547_n N_A_27_74#_c_1186_n 0.0213941f $X=7.98 $Y=1.395 $X2=0
+ $Y2=0
cc_565 N_A_200_74#_c_536_n N_A_27_74#_c_1187_n 0.00177344f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_566 N_A_200_74#_c_538_n N_A_27_74#_c_1187_n 0.0168035f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_567 N_A_200_74#_c_542_n N_A_27_74#_c_1187_n 0.00661136f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_568 N_A_200_74#_c_539_n N_A_27_74#_c_1202_n 2.03345e-19 $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_569 N_A_200_74#_M1038_g N_A_27_74#_M1018_g 0.0278203f $X=6.8 $Y=2.54 $X2=0
+ $Y2=0
cc_570 N_A_200_74#_c_555_n N_A_27_74#_c_1204_n 0.00111738f $X=3.075 $Y=2.19
+ $X2=0 $Y2=0
cc_571 N_A_200_74#_c_561_n N_A_27_74#_c_1204_n 2.83685e-19 $X=3.107 $Y=1.77
+ $X2=0 $Y2=0
cc_572 N_A_200_74#_c_537_n N_A_27_74#_c_1189_n 0.00514147f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_573 N_A_200_74#_c_538_n N_A_27_74#_c_1189_n 0.0205564f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_574 N_A_200_74#_c_539_n N_A_27_74#_c_1189_n 0.0118811f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_575 N_A_200_74#_c_550_n N_A_27_74#_c_1207_n 0.00477437f $X=1.17 $Y=2.815
+ $X2=0 $Y2=0
cc_576 N_A_200_74#_c_541_n N_A_27_74#_c_1191_n 0.0014153f $X=1.235 $Y=1.13 $X2=0
+ $Y2=0
cc_577 N_A_200_74#_c_540_n N_A_27_74#_c_1193_n 0.0048959f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_578 N_A_200_74#_c_559_n N_A_27_74#_c_1194_n 0.00575747f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_579 N_A_200_74#_c_540_n N_A_27_74#_c_1194_n 0.0057101f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_580 N_A_200_74#_c_559_n N_A_27_74#_c_1195_n 0.00521925f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_581 N_A_200_74#_c_540_n N_A_27_74#_c_1195_n 0.0251869f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_582 N_A_200_74#_c_541_n N_A_27_74#_c_1195_n 0.00160233f $X=1.235 $Y=1.13
+ $X2=0 $Y2=0
cc_583 N_A_200_74#_c_559_n N_A_27_74#_c_1196_n 0.00309714f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_584 N_A_200_74#_c_540_n N_A_27_74#_c_1196_n 0.00539244f $X=1.21 $Y=1.82 $X2=0
+ $Y2=0
cc_585 N_A_200_74#_c_541_n N_A_27_74#_c_1196_n 0.00266468f $X=1.235 $Y=1.13
+ $X2=0 $Y2=0
cc_586 N_A_200_74#_c_533_n N_A_1534_446#_M1000_g 0.0491204f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_587 N_A_200_74#_c_547_n N_A_1534_446#_c_1382_n 0.00632126f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_588 N_A_200_74#_c_533_n N_A_1349_114#_c_1567_n 0.0216797f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_589 N_A_200_74#_c_536_n N_A_1349_114#_c_1567_n 0.0236508f $X=6.892 $Y=1.56
+ $X2=0 $Y2=0
cc_590 N_A_200_74#_c_539_n N_A_1349_114#_c_1567_n 0.0641468f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_591 N_A_200_74#_c_542_n N_A_1349_114#_c_1567_n 6.67233e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_592 N_A_200_74#_c_543_n N_A_1349_114#_c_1567_n 0.00293315f $X=6.96 $Y=1.295
+ $X2=0 $Y2=0
cc_593 N_A_200_74#_c_547_n N_A_1349_114#_c_1567_n 0.00161335f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_594 N_A_200_74#_M1038_g N_A_1349_114#_c_1572_n 0.0136426f $X=6.8 $Y=2.54
+ $X2=0 $Y2=0
cc_595 N_A_200_74#_c_539_n N_A_1349_114#_c_1573_n 0.033189f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_596 N_A_200_74#_c_547_n N_A_1349_114#_c_1573_n 0.0076278f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_597 N_A_200_74#_c_537_n N_A_1349_114#_c_1574_n 0.015142f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_598 N_A_200_74#_c_538_n N_A_1349_114#_c_1574_n 5.92995e-19 $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_599 N_A_200_74#_c_539_n N_A_1349_114#_c_1574_n 0.0132387f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_600 N_A_200_74#_c_533_n N_A_1349_114#_c_1568_n 0.00868176f $X=7.98 $Y=1.23
+ $X2=0 $Y2=0
cc_601 N_A_200_74#_c_539_n N_A_1349_114#_c_1568_n 0.0289805f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_602 N_A_200_74#_c_547_n N_A_1349_114#_c_1568_n 0.00735633f $X=7.98 $Y=1.395
+ $X2=0 $Y2=0
cc_603 N_A_200_74#_M1038_g N_A_1349_114#_c_1583_n 0.00493484f $X=6.8 $Y=2.54
+ $X2=0 $Y2=0
cc_604 N_A_200_74#_c_537_n N_A_1349_114#_c_1583_n 0.0149737f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_605 N_A_200_74#_c_538_n N_A_1349_114#_c_1583_n 0.00103977f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_606 N_A_200_74#_c_539_n N_A_1349_114#_c_1583_n 0.00347259f $X=7.775 $Y=1.395
+ $X2=0 $Y2=0
cc_607 N_A_200_74#_M1038_g N_A_1349_114#_c_1584_n 0.0022091f $X=6.8 $Y=2.54
+ $X2=0 $Y2=0
cc_608 N_A_200_74#_c_537_n N_A_1349_114#_c_1584_n 0.0023592f $X=6.875 $Y=1.765
+ $X2=0 $Y2=0
cc_609 N_A_200_74#_c_552_n N_VPWR_c_1813_n 0.0101219f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_610 N_A_200_74#_c_551_n N_VPWR_c_1814_n 0.01287f $X=1.955 $Y=2.99 $X2=0 $Y2=0
cc_611 N_A_200_74#_c_554_n N_VPWR_c_1814_n 0.00224848f $X=2.975 $Y=1.77 $X2=0
+ $Y2=0
cc_612 N_A_200_74#_M1038_g N_VPWR_c_1816_n 0.00142207f $X=6.8 $Y=2.54 $X2=0
+ $Y2=0
cc_613 N_A_200_74#_c_551_n N_VPWR_c_1819_n 0.0469143f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_614 N_A_200_74#_c_552_n N_VPWR_c_1819_n 0.0292499f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_615 N_A_200_74#_M1015_g N_VPWR_c_1824_n 0.00113339f $X=3.03 $Y=2.725 $X2=0
+ $Y2=0
cc_616 N_A_200_74#_M1038_g N_VPWR_c_1825_n 0.005209f $X=6.8 $Y=2.54 $X2=0 $Y2=0
cc_617 N_A_200_74#_M1038_g N_VPWR_c_1812_n 0.00983772f $X=6.8 $Y=2.54 $X2=0
+ $Y2=0
cc_618 N_A_200_74#_c_551_n N_VPWR_c_1812_n 0.026904f $X=1.955 $Y=2.99 $X2=0
+ $Y2=0
cc_619 N_A_200_74#_c_552_n N_VPWR_c_1812_n 0.0157973f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_620 N_A_200_74#_c_551_n N_A_311_119#_M1017_s 0.00600243f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_621 N_A_200_74#_c_542_n N_A_311_119#_c_1971_n 0.00551684f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_622 N_A_200_74#_c_542_n N_A_311_119#_c_1972_n 8.77327e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_623 N_A_200_74#_c_546_n N_A_311_119#_c_1972_n 0.00635523f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_624 N_A_200_74#_c_546_n N_A_311_119#_c_1973_n 0.0044168f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_625 N_A_200_74#_c_542_n N_A_311_119#_c_1980_n 0.00532224f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_626 N_A_200_74#_c_542_n N_A_311_119#_c_1981_n 5.75848e-19 $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_627 N_A_200_74#_c_542_n N_A_311_119#_c_1974_n 0.0131302f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_628 N_A_200_74#_c_534_n N_A_311_119#_c_1975_n 0.057087f $X=1.14 $Y=0.515
+ $X2=0 $Y2=0
cc_629 N_A_200_74#_c_551_n N_A_311_119#_c_1983_n 0.0149535f $X=1.955 $Y=2.99
+ $X2=0 $Y2=0
cc_630 N_A_200_74#_c_553_n N_A_311_119#_c_1983_n 0.0234904f $X=2.04 $Y=2.905
+ $X2=0 $Y2=0
cc_631 N_A_200_74#_c_559_n N_A_311_119#_c_1983_n 0.057087f $X=1.17 $Y=1.985
+ $X2=0 $Y2=0
cc_632 N_A_200_74#_c_553_n N_A_311_119#_c_1976_n 0.0347656f $X=2.04 $Y=2.905
+ $X2=0 $Y2=0
cc_633 N_A_200_74#_c_568_n N_A_311_119#_c_1976_n 0.0120098f $X=2.125 $Y=1.77
+ $X2=0 $Y2=0
cc_634 N_A_200_74#_c_541_n N_A_311_119#_c_1976_n 0.057087f $X=1.235 $Y=1.13
+ $X2=0 $Y2=0
cc_635 N_A_200_74#_c_546_n N_A_311_119#_c_1977_n 0.00150382f $X=3.35 $Y=1.125
+ $X2=0 $Y2=0
cc_636 N_A_200_74#_c_542_n N_A_311_119#_c_1978_n 0.0150322f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_637 N_A_200_74#_c_534_n N_VGND_c_2147_n 0.0165395f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_638 N_A_200_74#_c_534_n N_VGND_c_2148_n 0.00758914f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_639 N_A_200_74#_c_542_n N_VGND_c_2149_n 0.00908153f $X=6.815 $Y=1.295 $X2=0
+ $Y2=0
cc_640 N_A_200_74#_c_534_n N_VGND_c_2154_n 0.0159616f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_200_74#_c_534_n N_VGND_c_2160_n 0.0117867f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_642 N_A_200_74#_c_542_n N_A_867_119#_c_2279_n 0.00677876f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_643 N_A_200_74#_c_542_n N_A_867_119#_c_2282_n 0.00908153f $X=6.815 $Y=1.295
+ $X2=0 $Y2=0
cc_644 N_A_595_119#_M1021_g N_A_978_357#_c_867_n 0.0879274f $X=4.59 $Y=2.54
+ $X2=0 $Y2=0
cc_645 N_A_595_119#_M1020_g N_A_978_357#_c_867_n 0.0132724f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_646 N_A_595_119#_M1020_g N_A_978_357#_M1032_g 0.0211547f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_647 N_A_595_119#_M1020_g N_A_978_357#_c_880_n 2.53172e-19 $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_648 N_A_595_119#_c_766_n N_A_27_74#_M1001_g 0.00526053f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_649 N_A_595_119#_c_767_n N_A_27_74#_M1001_g 3.07252e-19 $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_650 N_A_595_119#_M1020_g N_A_27_74#_c_1184_n 0.00897756f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_651 N_A_595_119#_c_770_n N_A_27_74#_c_1198_n 0.00217111f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_652 N_A_595_119#_c_767_n N_A_27_74#_c_1198_n 0.00872687f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_653 N_A_595_119#_c_768_n N_A_27_74#_c_1198_n 0.00390887f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_654 N_A_595_119#_c_770_n N_A_27_74#_c_1200_n 0.00262194f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_655 N_A_595_119#_c_767_n N_A_27_74#_c_1200_n 0.00124794f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_656 N_A_595_119#_c_781_n N_A_27_74#_M1012_g 0.00495591f $X=3.41 $Y=2.65 $X2=0
+ $Y2=0
cc_657 N_A_595_119#_c_770_n N_A_27_74#_M1012_g 0.0109798f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_658 N_A_595_119#_c_770_n N_A_27_74#_c_1204_n 0.0094144f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_659 N_A_595_119#_M1021_g N_VPWR_c_1815_n 0.00122068f $X=4.59 $Y=2.54 $X2=0
+ $Y2=0
cc_660 N_A_595_119#_M1021_g N_VPWR_c_1824_n 0.00517089f $X=4.59 $Y=2.54 $X2=0
+ $Y2=0
cc_661 N_A_595_119#_M1021_g N_VPWR_c_1812_n 0.00538485f $X=4.59 $Y=2.54 $X2=0
+ $Y2=0
cc_662 N_A_595_119#_c_789_n N_A_311_119#_M1005_d 0.00979049f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_663 N_A_595_119#_c_765_n N_A_311_119#_M1005_d 0.00185193f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_664 N_A_595_119#_c_766_n N_A_311_119#_c_1985_n 0.00837589f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_665 N_A_595_119#_c_766_n N_A_311_119#_c_1969_n 0.0159264f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_666 N_A_595_119#_M1020_g N_A_311_119#_c_1971_n 5.72873e-19 $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_667 N_A_595_119#_c_789_n N_A_311_119#_c_1972_n 0.026311f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_668 N_A_595_119#_M1021_g N_A_311_119#_c_1979_n 0.00193765f $X=4.59 $Y=2.54
+ $X2=0 $Y2=0
cc_669 N_A_595_119#_c_781_n N_A_311_119#_c_1979_n 0.0133863f $X=3.41 $Y=2.65
+ $X2=0 $Y2=0
cc_670 N_A_595_119#_c_770_n N_A_311_119#_c_1979_n 0.0314559f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_671 N_A_595_119#_M1020_g N_A_311_119#_c_1973_n 0.00145038f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_672 N_A_595_119#_c_789_n N_A_311_119#_c_1973_n 0.0135471f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_673 N_A_595_119#_c_765_n N_A_311_119#_c_1973_n 0.00286902f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_674 N_A_595_119#_c_761_n N_A_311_119#_c_1980_n 0.00431129f $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_675 N_A_595_119#_M1021_g N_A_311_119#_c_1980_n 0.00414658f $X=4.59 $Y=2.54
+ $X2=0 $Y2=0
cc_676 N_A_595_119#_c_767_n N_A_311_119#_c_1980_n 0.0106373f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_677 N_A_595_119#_c_768_n N_A_311_119#_c_1980_n 9.61154e-19 $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_678 N_A_595_119#_c_770_n N_A_311_119#_c_1981_n 0.0136812f $X=3.495 $Y=2.565
+ $X2=0 $Y2=0
cc_679 N_A_595_119#_c_767_n N_A_311_119#_c_1981_n 0.022168f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_680 N_A_595_119#_c_768_n N_A_311_119#_c_1981_n 0.00125273f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_681 N_A_595_119#_c_761_n N_A_311_119#_c_1974_n 0.0134603f $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_682 N_A_595_119#_M1021_g N_A_311_119#_c_1974_n 0.00723318f $X=4.59 $Y=2.54
+ $X2=0 $Y2=0
cc_683 N_A_595_119#_M1020_g N_A_311_119#_c_1974_n 0.00397984f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_684 N_A_595_119#_c_765_n N_A_311_119#_c_1974_n 0.00632424f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_685 N_A_595_119#_c_767_n N_A_311_119#_c_1974_n 0.0312801f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_686 N_A_595_119#_c_768_n N_A_311_119#_c_1974_n 0.00130314f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_687 N_A_595_119#_c_789_n N_A_311_119#_c_1977_n 0.0057043f $X=3.635 $Y=0.87
+ $X2=0 $Y2=0
cc_688 N_A_595_119#_c_766_n N_A_311_119#_c_1977_n 0.0198509f $X=3.115 $Y=0.775
+ $X2=0 $Y2=0
cc_689 N_A_595_119#_c_761_n N_A_311_119#_c_1978_n 6.95961e-19 $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_690 N_A_595_119#_M1020_g N_A_311_119#_c_1978_n 0.00341236f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_691 N_A_595_119#_c_765_n N_A_311_119#_c_1978_n 0.0137783f $X=3.72 $Y=1.395
+ $X2=0 $Y2=0
cc_692 N_A_595_119#_c_767_n N_A_311_119#_c_1978_n 0.00657374f $X=3.72 $Y=1.595
+ $X2=0 $Y2=0
cc_693 N_A_595_119#_c_768_n N_A_311_119#_c_1978_n 0.00654668f $X=3.975 $Y=1.47
+ $X2=0 $Y2=0
cc_694 N_A_595_119#_c_761_n N_A_867_119#_c_2279_n 0.00352503f $X=4.5 $Y=1.47
+ $X2=0 $Y2=0
cc_695 N_A_595_119#_M1020_g N_A_867_119#_c_2279_n 0.00948034f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_696 N_A_595_119#_M1020_g N_A_867_119#_c_2280_n 0.00159671f $X=4.695 $Y=0.87
+ $X2=0 $Y2=0
cc_697 N_A_978_357#_c_867_n N_SET_B_M1027_g 0.0121481f $X=4.98 $Y=1.935 $X2=0
+ $Y2=0
cc_698 N_A_978_357#_M1032_g N_SET_B_M1027_g 0.0217173f $X=5.195 $Y=0.87 $X2=0
+ $Y2=0
cc_699 N_A_978_357#_c_870_n N_SET_B_M1027_g 0.0122073f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_700 N_A_978_357#_c_880_n N_SET_B_M1027_g 8.00353e-19 $X=5.125 $Y=1.42 $X2=0
+ $Y2=0
cc_701 N_A_978_357#_M1019_g N_SET_B_c_1048_n 7.28982e-19 $X=9.51 $Y=2.46 $X2=0
+ $Y2=0
cc_702 N_A_978_357#_c_928_p N_SET_B_c_1048_n 0.00529741f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_703 N_A_978_357#_c_875_n N_SET_B_c_1048_n 5.89036e-19 $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_704 N_A_978_357#_c_876_n N_SET_B_c_1048_n 0.00828265f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_705 N_A_978_357#_M1019_g N_SET_B_M1025_g 0.0366301f $X=9.51 $Y=2.46 $X2=0
+ $Y2=0
cc_706 N_A_978_357#_c_874_n N_SET_B_M1016_g 0.00329169f $X=8.46 $Y=0.935 $X2=0
+ $Y2=0
cc_707 N_A_978_357#_c_928_p N_SET_B_M1016_g 0.0159922f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_708 N_A_978_357#_c_875_n N_SET_B_M1016_g 0.00354892f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_709 N_A_978_357#_c_876_n N_SET_B_M1016_g 0.0106664f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_710 N_A_978_357#_c_882_n N_SET_B_M1016_g 0.0276447f $X=9.465 $Y=1.23 $X2=0
+ $Y2=0
cc_711 N_A_978_357#_c_870_n N_SET_B_c_1055_n 0.0122852f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_712 N_A_978_357#_M1003_g N_SET_B_c_1068_n 0.00112442f $X=4.98 $Y=2.54 $X2=0
+ $Y2=0
cc_713 N_A_978_357#_c_870_n N_SET_B_c_1068_n 0.00196094f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_714 N_A_978_357#_c_867_n N_SET_B_c_1051_n 0.0121367f $X=4.98 $Y=1.935 $X2=0
+ $Y2=0
cc_715 N_A_978_357#_M1003_g N_SET_B_c_1051_n 0.0372169f $X=4.98 $Y=2.54 $X2=0
+ $Y2=0
cc_716 N_A_978_357#_c_870_n N_SET_B_c_1051_n 0.00797137f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_717 N_A_978_357#_c_880_n N_SET_B_c_1051_n 2.24557e-19 $X=5.125 $Y=1.42 $X2=0
+ $Y2=0
cc_718 N_A_978_357#_c_867_n N_SET_B_c_1057_n 0.00225274f $X=4.98 $Y=1.935 $X2=0
+ $Y2=0
cc_719 N_A_978_357#_M1003_g N_SET_B_c_1057_n 9.72934e-19 $X=4.98 $Y=2.54 $X2=0
+ $Y2=0
cc_720 N_A_978_357#_c_870_n N_SET_B_c_1057_n 0.0279177f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_721 N_A_978_357#_M1019_g N_SET_B_c_1052_n 0.00800402f $X=9.51 $Y=2.46 $X2=0
+ $Y2=0
cc_722 N_A_978_357#_c_928_p N_SET_B_c_1052_n 0.023413f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_723 N_A_978_357#_c_875_n N_SET_B_c_1052_n 0.0162366f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_724 N_A_978_357#_c_876_n N_SET_B_c_1052_n 0.00100533f $X=9.465 $Y=1.395 $X2=0
+ $Y2=0
cc_725 N_A_978_357#_M1032_g N_A_27_74#_c_1184_n 0.00882199f $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_726 N_A_978_357#_c_872_n N_A_27_74#_c_1184_n 4.42178e-19 $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_727 N_A_978_357#_c_873_n N_A_27_74#_c_1184_n 0.00404452f $X=6.485 $Y=0.425
+ $X2=0 $Y2=0
cc_728 N_A_978_357#_c_871_n N_A_27_74#_M1028_g 0.0114165f $X=6.4 $Y=1.335 $X2=0
+ $Y2=0
cc_729 N_A_978_357#_c_872_n N_A_27_74#_M1028_g 0.0169314f $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_730 N_A_978_357#_c_877_n N_A_1534_446#_M1034_d 0.00741937f $X=10.345 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_731 N_A_978_357#_c_957_p N_A_1534_446#_M1034_d 5.75378e-19 $X=9.465 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_732 N_A_978_357#_c_872_n N_A_1534_446#_M1000_g 0.00372402f $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_733 N_A_978_357#_c_874_n N_A_1534_446#_M1000_g 0.0105501f $X=8.46 $Y=0.935
+ $X2=0 $Y2=0
cc_734 N_A_978_357#_c_960_p N_A_1534_446#_M1000_g 0.00726228f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_735 N_A_978_357#_M1019_g N_A_1534_446#_c_1383_n 0.0158548f $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_736 N_A_978_357#_M1008_s N_A_1534_446#_c_1372_n 0.0022485f $X=10.595 $Y=0.745
+ $X2=0 $Y2=0
cc_737 N_A_978_357#_c_876_n N_A_1534_446#_c_1372_n 3.26158e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_738 N_A_978_357#_c_877_n N_A_1534_446#_c_1372_n 0.0428702f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_739 N_A_978_357#_c_879_n N_A_1534_446#_c_1372_n 0.0231179f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_740 N_A_978_357#_c_957_p N_A_1534_446#_c_1372_n 0.00613989f $X=9.465 $Y=1.02
+ $X2=0 $Y2=0
cc_741 N_A_978_357#_c_881_n N_A_1534_446#_c_1372_n 0.0143583f $X=10.43 $Y=1.02
+ $X2=0 $Y2=0
cc_742 N_A_978_357#_c_882_n N_A_1534_446#_c_1372_n 0.00239488f $X=9.465 $Y=1.23
+ $X2=0 $Y2=0
cc_743 N_A_978_357#_M1019_g N_A_1534_446#_c_1384_n 4.90292e-19 $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_744 N_A_978_357#_M1019_g N_A_1534_446#_c_1385_n 8.11218e-19 $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_745 N_A_978_357#_M1011_s N_A_1534_446#_c_1386_n 0.0108749f $X=10.555 $Y=1.84
+ $X2=0 $Y2=0
cc_746 N_A_978_357#_c_887_n N_A_1534_446#_c_1386_n 0.014265f $X=10.515 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_A_978_357#_c_888_n N_A_1534_446#_c_1386_n 0.0200816f $X=10.685 $Y=2.035
+ $X2=0 $Y2=0
cc_748 N_A_978_357#_c_888_n N_A_1534_446#_c_1387_n 0.00713603f $X=10.685
+ $Y=2.035 $X2=0 $Y2=0
cc_749 N_A_978_357#_M1019_g N_A_1534_446#_c_1389_n 7.57297e-19 $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_750 N_A_978_357#_c_879_n N_A_1534_446#_c_1375_n 0.00799877f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_751 N_A_978_357#_c_875_n N_A_1349_114#_M1033_g 0.00458614f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_752 N_A_978_357#_c_876_n N_A_1349_114#_M1033_g 0.0207024f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_753 N_A_978_357#_c_877_n N_A_1349_114#_M1033_g 0.0135044f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_754 N_A_978_357#_c_878_n N_A_1349_114#_M1033_g 0.00822808f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_755 N_A_978_357#_c_882_n N_A_1349_114#_M1033_g 0.0225065f $X=9.465 $Y=1.23
+ $X2=0 $Y2=0
cc_756 N_A_978_357#_c_878_n N_A_1349_114#_M1026_g 9.92444e-19 $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_757 N_A_978_357#_c_887_n N_A_1349_114#_M1026_g 9.17416e-19 $X=10.515 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_A_978_357#_c_871_n N_A_1349_114#_c_1567_n 0.02006f $X=6.4 $Y=1.335
+ $X2=0 $Y2=0
cc_759 N_A_978_357#_c_872_n N_A_1349_114#_c_1567_n 0.108619f $X=8.375 $Y=0.425
+ $X2=0 $Y2=0
cc_760 N_A_978_357#_c_874_n N_A_1349_114#_c_1567_n 0.020128f $X=8.46 $Y=0.935
+ $X2=0 $Y2=0
cc_761 N_A_978_357#_c_960_p N_A_1349_114#_c_1567_n 0.00655524f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_762 N_A_978_357#_c_960_p N_A_1349_114#_c_1568_n 0.00743036f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_763 N_A_978_357#_c_928_p N_A_1349_114#_c_1576_n 4.73677e-19 $X=9.3 $Y=1.02
+ $X2=0 $Y2=0
cc_764 N_A_978_357#_c_960_p N_A_1349_114#_c_1576_n 0.00452026f $X=8.545 $Y=1.02
+ $X2=0 $Y2=0
cc_765 N_A_978_357#_M1019_g N_A_1349_114#_c_1579_n 0.0148839f $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_766 N_A_978_357#_c_875_n N_A_1349_114#_c_1579_n 0.00902113f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_767 N_A_978_357#_c_876_n N_A_1349_114#_c_1579_n 2.83373e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_768 N_A_978_357#_c_887_n N_A_1349_114#_c_1579_n 0.0149788f $X=10.515 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_A_978_357#_c_875_n N_A_1349_114#_c_1580_n 0.0045977f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_770 N_A_978_357#_c_876_n N_A_1349_114#_c_1580_n 6.67297e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_771 N_A_978_357#_M1019_g N_A_1349_114#_c_1569_n 0.00255856f $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_772 N_A_978_357#_c_875_n N_A_1349_114#_c_1569_n 0.00887229f $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_773 N_A_978_357#_c_876_n N_A_1349_114#_c_1569_n 4.87607e-19 $X=9.465 $Y=1.395
+ $X2=0 $Y2=0
cc_774 N_A_978_357#_c_877_n N_A_1349_114#_c_1569_n 0.0143654f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_775 N_A_978_357#_c_878_n N_A_1349_114#_c_1569_n 0.0397228f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_776 N_A_978_357#_M1019_g N_A_1349_114#_c_1570_n 0.0835739f $X=9.51 $Y=2.46
+ $X2=0 $Y2=0
cc_777 N_A_978_357#_c_877_n N_A_1349_114#_c_1570_n 9.39401e-19 $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_778 N_A_978_357#_c_878_n N_A_1349_114#_c_1570_n 0.00303292f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_779 N_A_978_357#_c_878_n N_RESET_B_M1011_g 0.00380857f $X=10.43 $Y=1.95 $X2=0
+ $Y2=0
cc_780 N_A_978_357#_c_888_n N_RESET_B_M1011_g 0.00344428f $X=10.685 $Y=2.035
+ $X2=0 $Y2=0
cc_781 N_A_978_357#_c_878_n N_RESET_B_M1008_g 0.00606104f $X=10.43 $Y=1.95 $X2=0
+ $Y2=0
cc_782 N_A_978_357#_c_879_n N_RESET_B_M1008_g 0.00307743f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_783 N_A_978_357#_c_878_n N_RESET_B_c_1720_n 0.00307165f $X=10.43 $Y=1.95
+ $X2=0 $Y2=0
cc_784 N_A_978_357#_c_879_n N_RESET_B_c_1720_n 0.00101461f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_785 N_A_978_357#_c_888_n N_RESET_B_c_1720_n 6.26988e-19 $X=10.685 $Y=2.035
+ $X2=0 $Y2=0
cc_786 N_A_978_357#_c_878_n N_RESET_B_c_1721_n 0.0327297f $X=10.43 $Y=1.95 $X2=0
+ $Y2=0
cc_787 N_A_978_357#_c_879_n N_RESET_B_c_1721_n 0.00997949f $X=10.725 $Y=1.02
+ $X2=0 $Y2=0
cc_788 N_A_978_357#_c_888_n N_RESET_B_c_1721_n 0.0108099f $X=10.685 $Y=2.035
+ $X2=0 $Y2=0
cc_789 N_A_978_357#_M1003_g N_VPWR_c_1815_n 0.0101853f $X=4.98 $Y=2.54 $X2=0
+ $Y2=0
cc_790 N_A_978_357#_M1003_g N_VPWR_c_1824_n 0.00460063f $X=4.98 $Y=2.54 $X2=0
+ $Y2=0
cc_791 N_A_978_357#_M1019_g N_VPWR_c_1827_n 0.0037725f $X=9.51 $Y=2.46 $X2=0
+ $Y2=0
cc_792 N_A_978_357#_M1003_g N_VPWR_c_1812_n 0.00460366f $X=4.98 $Y=2.54 $X2=0
+ $Y2=0
cc_793 N_A_978_357#_M1019_g N_VPWR_c_1812_n 0.00466339f $X=9.51 $Y=2.46 $X2=0
+ $Y2=0
cc_794 N_A_978_357#_M1019_g N_VPWR_c_1834_n 0.00336105f $X=9.51 $Y=2.46 $X2=0
+ $Y2=0
cc_795 N_A_978_357#_c_874_n N_VGND_M1000_d 0.00296211f $X=8.46 $Y=0.935 $X2=0
+ $Y2=0
cc_796 N_A_978_357#_c_928_p N_VGND_M1000_d 0.01748f $X=9.3 $Y=1.02 $X2=0 $Y2=0
cc_797 N_A_978_357#_c_960_p N_VGND_M1000_d 8.96084e-19 $X=8.545 $Y=1.02 $X2=0
+ $Y2=0
cc_798 N_A_978_357#_c_870_n N_VGND_c_2149_n 0.0112717f $X=6.315 $Y=1.42 $X2=0
+ $Y2=0
cc_799 N_A_978_357#_c_871_n N_VGND_c_2149_n 0.022822f $X=6.4 $Y=1.335 $X2=0
+ $Y2=0
cc_800 N_A_978_357#_c_873_n N_VGND_c_2149_n 0.014852f $X=6.485 $Y=0.425 $X2=0
+ $Y2=0
cc_801 N_A_978_357#_c_872_n N_VGND_c_2150_n 0.0141848f $X=8.375 $Y=0.425 $X2=0
+ $Y2=0
cc_802 N_A_978_357#_c_874_n N_VGND_c_2150_n 0.0187368f $X=8.46 $Y=0.935 $X2=0
+ $Y2=0
cc_803 N_A_978_357#_c_928_p N_VGND_c_2150_n 0.0135869f $X=9.3 $Y=1.02 $X2=0
+ $Y2=0
cc_804 N_A_978_357#_c_872_n N_VGND_c_2156_n 0.08689f $X=8.375 $Y=0.425 $X2=0
+ $Y2=0
cc_805 N_A_978_357#_c_873_n N_VGND_c_2156_n 0.00789578f $X=6.485 $Y=0.425 $X2=0
+ $Y2=0
cc_806 N_A_978_357#_c_882_n N_VGND_c_2157_n 0.00390708f $X=9.465 $Y=1.23 $X2=0
+ $Y2=0
cc_807 N_A_978_357#_c_872_n N_VGND_c_2160_n 0.0724187f $X=8.375 $Y=0.425 $X2=0
+ $Y2=0
cc_808 N_A_978_357#_c_873_n N_VGND_c_2160_n 0.00563471f $X=6.485 $Y=0.425 $X2=0
+ $Y2=0
cc_809 N_A_978_357#_c_882_n N_VGND_c_2160_n 0.00542671f $X=9.465 $Y=1.23 $X2=0
+ $Y2=0
cc_810 N_A_978_357#_M1032_g N_A_867_119#_c_2279_n 7.14713e-19 $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_811 N_A_978_357#_M1032_g N_A_867_119#_c_2280_n 0.00333342f $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_812 N_A_978_357#_M1032_g N_A_867_119#_c_2282_n 0.00432227f $X=5.195 $Y=0.87
+ $X2=0 $Y2=0
cc_813 N_A_978_357#_c_870_n N_A_867_119#_c_2282_n 0.0112717f $X=6.315 $Y=1.42
+ $X2=0 $Y2=0
cc_814 N_A_978_357#_c_871_n A_1254_119# 0.0103426f $X=6.4 $Y=1.335 $X2=-0.19
+ $Y2=-0.245
cc_815 N_A_978_357#_c_928_p N_A_1818_76#_M1016_d 0.00741543f $X=9.3 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_816 N_A_978_357#_c_877_n N_A_1818_76#_M1033_d 0.0117491f $X=10.345 $Y=1.02
+ $X2=0 $Y2=0
cc_817 N_A_978_357#_c_928_p N_A_1818_76#_c_2315_n 0.0139095f $X=9.3 $Y=1.02
+ $X2=0 $Y2=0
cc_818 N_A_978_357#_c_957_p N_A_1818_76#_c_2315_n 0.0011409f $X=9.465 $Y=1.02
+ $X2=0 $Y2=0
cc_819 N_A_978_357#_c_957_p N_A_1818_76#_c_2312_n 0.00383022f $X=9.465 $Y=1.02
+ $X2=0 $Y2=0
cc_820 N_A_978_357#_c_882_n N_A_1818_76#_c_2312_n 0.0101322f $X=9.465 $Y=1.23
+ $X2=0 $Y2=0
cc_821 N_SET_B_M1027_g N_A_27_74#_c_1184_n 0.0103062f $X=5.695 $Y=0.87 $X2=0
+ $Y2=0
cc_822 N_SET_B_c_1055_n N_A_27_74#_c_1187_n 0.00122312f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_823 N_SET_B_c_1055_n N_A_27_74#_M1018_g 0.00264708f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_824 N_SET_B_c_1055_n N_A_1534_446#_M1025_s 0.00787608f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_825 SET_B N_A_1534_446#_M1025_s 7.77338e-19 $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_826 N_SET_B_c_1052_n N_A_1534_446#_M1025_s 8.81142e-19 $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_827 N_SET_B_c_1048_n N_A_1534_446#_M1000_g 0.0140919f $X=8.89 $Y=1.58 $X2=0
+ $Y2=0
cc_828 N_SET_B_M1025_g N_A_1534_446#_M1000_g 0.0256558f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_829 N_SET_B_M1016_g N_A_1534_446#_M1000_g 0.0128657f $X=9.015 $Y=0.75 $X2=0
+ $Y2=0
cc_830 N_SET_B_c_1055_n N_A_1534_446#_M1000_g 0.00213512f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_831 N_SET_B_c_1052_n N_A_1534_446#_M1000_g 0.00350965f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_832 N_SET_B_M1025_g N_A_1534_446#_c_1381_n 0.00430324f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_833 N_SET_B_c_1055_n N_A_1534_446#_c_1381_n 0.0215507f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_834 N_SET_B_c_1055_n N_A_1534_446#_c_1382_n 0.00932486f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_835 N_SET_B_M1025_g N_A_1534_446#_c_1383_n 0.00894343f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_836 N_SET_B_c_1055_n N_A_1534_446#_c_1388_n 0.00557042f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_837 N_SET_B_M1025_g N_A_1534_446#_c_1389_n 0.00533679f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_838 N_SET_B_c_1055_n N_A_1534_446#_c_1389_n 3.27896e-19 $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_839 N_SET_B_c_1055_n N_A_1349_114#_c_1573_n 0.0280202f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_840 N_SET_B_c_1052_n N_A_1349_114#_c_1568_n 0.015133f $X=8.895 $Y=1.415 $X2=0
+ $Y2=0
cc_841 N_SET_B_M1025_g N_A_1349_114#_c_1576_n 6.08562e-19 $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_842 N_SET_B_c_1055_n N_A_1349_114#_c_1576_n 0.00830114f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_843 N_SET_B_c_1052_n N_A_1349_114#_c_1576_n 0.0150352f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_844 N_SET_B_M1025_g N_A_1349_114#_c_1577_n 0.00222502f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_845 N_SET_B_c_1055_n N_A_1349_114#_c_1577_n 0.0177878f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_846 SET_B N_A_1349_114#_c_1577_n 0.00149807f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_847 N_SET_B_c_1052_n N_A_1349_114#_c_1577_n 0.0155322f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_848 N_SET_B_M1025_g N_A_1349_114#_c_1647_n 0.0131845f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_849 N_SET_B_c_1055_n N_A_1349_114#_c_1647_n 0.00762662f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_850 SET_B N_A_1349_114#_c_1647_n 0.00745861f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_851 N_SET_B_c_1052_n N_A_1349_114#_c_1647_n 0.0153864f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_852 N_SET_B_M1025_g N_A_1349_114#_c_1651_n 0.0017557f $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_853 SET_B N_A_1349_114#_c_1651_n 9.78448e-19 $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_854 N_SET_B_M1025_g N_A_1349_114#_c_1580_n 6.25469e-19 $X=8.89 $Y=2.46 $X2=0
+ $Y2=0
cc_855 SET_B N_A_1349_114#_c_1580_n 0.00127852f $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_856 N_SET_B_c_1052_n N_A_1349_114#_c_1580_n 0.0131771f $X=8.895 $Y=1.415
+ $X2=0 $Y2=0
cc_857 N_SET_B_c_1055_n N_A_1349_114#_c_1583_n 0.033757f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_858 N_SET_B_c_1055_n N_A_1349_114#_c_1584_n 0.0129511f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_859 N_SET_B_c_1055_n N_A_1349_114#_c_1585_n 0.00501285f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_860 SET_B N_VPWR_M1025_d 6.16517e-19 $X=8.795 $Y=1.95 $X2=0 $Y2=0
cc_861 N_SET_B_c_1052_n N_VPWR_M1025_d 0.00170278f $X=8.895 $Y=1.415 $X2=0 $Y2=0
cc_862 N_SET_B_c_1053_n N_VPWR_c_1815_n 0.00897656f $X=5.43 $Y=2.025 $X2=0 $Y2=0
cc_863 N_SET_B_c_1053_n N_VPWR_c_1816_n 0.00236023f $X=5.43 $Y=2.025 $X2=0 $Y2=0
cc_864 N_SET_B_c_1055_n N_VPWR_c_1816_n 0.0011193f $X=8.735 $Y=2.035 $X2=0 $Y2=0
cc_865 N_SET_B_c_1053_n N_VPWR_c_1821_n 0.00460063f $X=5.43 $Y=2.025 $X2=0 $Y2=0
cc_866 N_SET_B_M1025_g N_VPWR_c_1826_n 0.00421734f $X=8.89 $Y=2.46 $X2=0 $Y2=0
cc_867 N_SET_B_c_1053_n N_VPWR_c_1812_n 0.00465993f $X=5.43 $Y=2.025 $X2=0 $Y2=0
cc_868 N_SET_B_M1025_g N_VPWR_c_1812_n 0.00638839f $X=8.89 $Y=2.46 $X2=0 $Y2=0
cc_869 N_SET_B_M1025_g N_VPWR_c_1833_n 0.00289754f $X=8.89 $Y=2.46 $X2=0 $Y2=0
cc_870 N_SET_B_M1025_g N_VPWR_c_1834_n 0.00332085f $X=8.89 $Y=2.46 $X2=0 $Y2=0
cc_871 N_SET_B_M1027_g N_VGND_c_2149_n 0.00339793f $X=5.695 $Y=0.87 $X2=0 $Y2=0
cc_872 N_SET_B_M1016_g N_VGND_c_2150_n 0.00301762f $X=9.015 $Y=0.75 $X2=0 $Y2=0
cc_873 N_SET_B_M1016_g N_VGND_c_2157_n 0.00540881f $X=9.015 $Y=0.75 $X2=0 $Y2=0
cc_874 N_SET_B_M1027_g N_VGND_c_2160_n 7.85159e-19 $X=5.695 $Y=0.87 $X2=0 $Y2=0
cc_875 N_SET_B_M1016_g N_VGND_c_2160_n 0.00542671f $X=9.015 $Y=0.75 $X2=0 $Y2=0
cc_876 N_SET_B_M1027_g N_A_867_119#_c_2282_n 0.00901521f $X=5.695 $Y=0.87 $X2=0
+ $Y2=0
cc_877 N_SET_B_M1016_g N_A_1818_76#_c_2315_n 0.00407202f $X=9.015 $Y=0.75 $X2=0
+ $Y2=0
cc_878 N_SET_B_M1016_g N_A_1818_76#_c_2311_n 0.00343135f $X=9.015 $Y=0.75 $X2=0
+ $Y2=0
cc_879 N_A_27_74#_M1018_g N_A_1534_446#_c_1381_n 9.56776e-19 $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_880 N_A_27_74#_M1018_g N_A_1534_446#_c_1382_n 0.0494357f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_881 N_A_27_74#_M1028_g N_A_1349_114#_c_1567_n 0.00450135f $X=6.67 $Y=0.845
+ $X2=0 $Y2=0
cc_882 N_A_27_74#_c_1186_n N_A_1349_114#_c_1567_n 0.00454853f $X=7.25 $Y=1.27
+ $X2=0 $Y2=0
cc_883 N_A_27_74#_M1018_g N_A_1349_114#_c_1572_n 0.0267114f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_884 N_A_27_74#_c_1202_n N_A_1349_114#_c_1573_n 0.00251451f $X=7.34 $Y=1.89
+ $X2=0 $Y2=0
cc_885 N_A_27_74#_M1018_g N_A_1349_114#_c_1573_n 3.96297e-19 $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_886 N_A_27_74#_c_1202_n N_A_1349_114#_c_1574_n 0.00174329f $X=7.34 $Y=1.89
+ $X2=0 $Y2=0
cc_887 N_A_27_74#_c_1189_n N_A_1349_114#_c_1574_n 0.00489714f $X=7.34 $Y=1.8
+ $X2=0 $Y2=0
cc_888 N_A_27_74#_c_1189_n N_A_1349_114#_c_1568_n 0.00358739f $X=7.34 $Y=1.8
+ $X2=0 $Y2=0
cc_889 N_A_27_74#_M1018_g N_A_1349_114#_c_1583_n 0.0113612f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_890 N_A_27_74#_M1018_g N_A_1349_114#_c_1584_n 0.0082087f $X=7.34 $Y=2.75
+ $X2=0 $Y2=0
cc_891 N_A_27_74#_c_1221_n N_VPWR_M1030_d 0.00283002f $X=0.665 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_892 N_A_27_74#_c_1194_n N_VPWR_M1030_d 0.00140562f $X=0.75 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_893 N_A_27_74#_M1031_g N_VPWR_c_1813_n 0.00120619f $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_894 N_A_27_74#_c_1207_n N_VPWR_c_1813_n 0.0233699f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_895 N_A_27_74#_c_1221_n N_VPWR_c_1813_n 0.0134989f $X=0.665 $Y=2.035 $X2=0
+ $Y2=0
cc_896 N_A_27_74#_M1031_g N_VPWR_c_1819_n 0.00517089f $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_897 N_A_27_74#_c_1207_n N_VPWR_c_1823_n 0.014549f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_898 N_A_27_74#_M1012_g N_VPWR_c_1824_n 0.00113339f $X=3.54 $Y=2.725 $X2=0
+ $Y2=0
cc_899 N_A_27_74#_M1018_g N_VPWR_c_1825_n 0.00367944f $X=7.34 $Y=2.75 $X2=0
+ $Y2=0
cc_900 N_A_27_74#_M1031_g N_VPWR_c_1812_n 0.00982721f $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_901 N_A_27_74#_M1018_g N_VPWR_c_1812_n 0.0048881f $X=7.34 $Y=2.75 $X2=0 $Y2=0
cc_902 N_A_27_74#_c_1207_n N_VPWR_c_1812_n 0.0119743f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_903 N_A_27_74#_c_1181_n N_A_311_119#_c_1985_n 0.00187443f $X=2.825 $Y=0.18
+ $X2=0 $Y2=0
cc_904 N_A_27_74#_M1001_g N_A_311_119#_c_1985_n 0.0025009f $X=2.9 $Y=0.805 $X2=0
+ $Y2=0
cc_905 N_A_27_74#_M1001_g N_A_311_119#_c_1969_n 0.00592273f $X=2.9 $Y=0.805
+ $X2=0 $Y2=0
cc_906 N_A_27_74#_c_1181_n N_A_311_119#_c_1970_n 0.00466053f $X=2.825 $Y=0.18
+ $X2=0 $Y2=0
cc_907 N_A_27_74#_c_1184_n N_A_311_119#_c_1971_n 0.00420304f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_908 N_A_27_74#_M1001_g N_A_311_119#_c_1972_n 0.00141636f $X=2.9 $Y=0.805
+ $X2=0 $Y2=0
cc_909 N_A_27_74#_M1012_g N_A_311_119#_c_1979_n 0.0127443f $X=3.54 $Y=2.725
+ $X2=0 $Y2=0
cc_910 N_A_27_74#_c_1200_n N_A_311_119#_c_1981_n 0.00371933f $X=3.54 $Y=2.055
+ $X2=0 $Y2=0
cc_911 N_A_27_74#_M1036_g N_A_311_119#_c_1975_n 0.00135176f $X=0.925 $Y=0.74
+ $X2=0 $Y2=0
cc_912 N_A_27_74#_c_1181_n N_A_311_119#_c_1975_n 0.00517374f $X=2.825 $Y=0.18
+ $X2=0 $Y2=0
cc_913 N_A_27_74#_M1031_g N_A_311_119#_c_1976_n 0.00196459f $X=0.945 $Y=2.4
+ $X2=0 $Y2=0
cc_914 N_A_27_74#_M1001_g N_A_311_119#_c_1977_n 0.0146966f $X=2.9 $Y=0.805 $X2=0
+ $Y2=0
cc_915 N_A_27_74#_c_1184_n N_A_311_119#_c_1977_n 0.0191582f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_916 N_A_27_74#_c_1191_n N_VGND_M1035_d 0.00210254f $X=0.665 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_917 N_A_27_74#_M1036_g N_VGND_c_2147_n 0.0115341f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_918 N_A_27_74#_c_1182_n N_VGND_c_2147_n 0.0075099f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_919 N_A_27_74#_c_1190_n N_VGND_c_2147_n 0.0164982f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_920 N_A_27_74#_c_1191_n N_VGND_c_2147_n 0.0158226f $X=0.665 $Y=1.045 $X2=0
+ $Y2=0
cc_921 N_A_27_74#_c_1195_n N_VGND_c_2147_n 0.00102653f $X=0.96 $Y=1.465 $X2=0
+ $Y2=0
cc_922 N_A_27_74#_c_1181_n N_VGND_c_2148_n 0.0272601f $X=2.825 $Y=0.18 $X2=0
+ $Y2=0
cc_923 N_A_27_74#_M1001_g N_VGND_c_2148_n 8.03294e-19 $X=2.9 $Y=0.805 $X2=0
+ $Y2=0
cc_924 N_A_27_74#_c_1184_n N_VGND_c_2149_n 0.0256899f $X=6.595 $Y=0.18 $X2=0
+ $Y2=0
cc_925 N_A_27_74#_M1028_g N_VGND_c_2149_n 0.003017f $X=6.67 $Y=0.845 $X2=0 $Y2=0
cc_926 N_A_27_74#_c_1190_n N_VGND_c_2153_n 0.011066f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_927 N_A_27_74#_c_1182_n N_VGND_c_2154_n 0.0339223f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_928 N_A_27_74#_c_1181_n N_VGND_c_2155_n 0.0774212f $X=2.825 $Y=0.18 $X2=0
+ $Y2=0
cc_929 N_A_27_74#_c_1184_n N_VGND_c_2156_n 0.016002f $X=6.595 $Y=0.18 $X2=0
+ $Y2=0
cc_930 N_A_27_74#_c_1181_n N_VGND_c_2160_n 0.0441429f $X=2.825 $Y=0.18 $X2=0
+ $Y2=0
cc_931 N_A_27_74#_c_1182_n N_VGND_c_2160_n 0.00749832f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_932 N_A_27_74#_c_1184_n N_VGND_c_2160_n 0.0930344f $X=6.595 $Y=0.18 $X2=0
+ $Y2=0
cc_933 N_A_27_74#_c_1188_n N_VGND_c_2160_n 0.00370846f $X=2.9 $Y=0.18 $X2=0
+ $Y2=0
cc_934 N_A_27_74#_c_1190_n N_VGND_c_2160_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_935 N_A_27_74#_c_1184_n N_A_867_119#_c_2280_n 0.0188768f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_936 N_A_27_74#_c_1184_n N_A_867_119#_c_2281_n 0.00766706f $X=6.595 $Y=0.18
+ $X2=0 $Y2=0
cc_937 N_A_1534_446#_c_1372_n N_A_1349_114#_M1033_g 0.0104522f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_938 N_A_1534_446#_c_1383_n N_A_1349_114#_M1026_g 0.0141382f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_939 N_A_1534_446#_c_1384_n N_A_1349_114#_M1026_g 0.00370477f $X=10.155
+ $Y=2.46 $X2=0 $Y2=0
cc_940 N_A_1534_446#_c_1385_n N_A_1349_114#_M1026_g 0.00313288f $X=10.155
+ $Y=2.63 $X2=0 $Y2=0
cc_941 N_A_1534_446#_M1000_g N_A_1349_114#_c_1567_n 0.00231064f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_942 N_A_1534_446#_M1023_g N_A_1349_114#_c_1572_n 0.00166962f $X=7.76 $Y=2.75
+ $X2=0 $Y2=0
cc_943 N_A_1534_446#_c_1381_n N_A_1349_114#_c_1573_n 0.00898403f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_944 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1573_n 0.00583408f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_945 N_A_1534_446#_M1000_g N_A_1349_114#_c_1568_n 0.0115778f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_946 N_A_1534_446#_M1000_g N_A_1349_114#_c_1576_n 0.0146118f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_947 N_A_1534_446#_c_1381_n N_A_1349_114#_c_1576_n 8.46766e-19 $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_948 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1576_n 0.0027583f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_949 N_A_1534_446#_M1025_s N_A_1349_114#_c_1577_n 0.00318778f $X=8.52 $Y=1.96
+ $X2=0 $Y2=0
cc_950 N_A_1534_446#_M1000_g N_A_1349_114#_c_1577_n 0.00593993f $X=8.37 $Y=0.91
+ $X2=0 $Y2=0
cc_951 N_A_1534_446#_c_1381_n N_A_1349_114#_c_1577_n 0.0153418f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_952 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1577_n 0.00639578f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_953 N_A_1534_446#_M1025_s N_A_1349_114#_c_1647_n 0.00425226f $X=8.52 $Y=1.96
+ $X2=0 $Y2=0
cc_954 N_A_1534_446#_c_1383_n N_A_1349_114#_c_1647_n 0.0105713f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_955 N_A_1534_446#_c_1389_n N_A_1349_114#_c_1647_n 0.0396679f $X=8.83 $Y=2.805
+ $X2=0 $Y2=0
cc_956 N_A_1534_446#_M1025_s N_A_1349_114#_c_1578_n 4.32645e-19 $X=8.52 $Y=1.96
+ $X2=0 $Y2=0
cc_957 N_A_1534_446#_c_1381_n N_A_1349_114#_c_1578_n 0.0142611f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_958 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1578_n 0.00393624f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_959 N_A_1534_446#_c_1388_n N_A_1349_114#_c_1578_n 0.0139859f $X=8.5 $Y=2.805
+ $X2=0 $Y2=0
cc_960 N_A_1534_446#_M1026_d N_A_1349_114#_c_1579_n 0.00266622f $X=10.02 $Y=1.96
+ $X2=0 $Y2=0
cc_961 N_A_1534_446#_c_1383_n N_A_1349_114#_c_1579_n 0.0138021f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_962 N_A_1534_446#_c_1384_n N_A_1349_114#_c_1579_n 0.0109175f $X=10.155
+ $Y=2.46 $X2=0 $Y2=0
cc_963 N_A_1534_446#_c_1384_n N_A_1349_114#_c_1570_n 4.57727e-19 $X=10.155
+ $Y=2.46 $X2=0 $Y2=0
cc_964 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1583_n 0.00166962f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_965 N_A_1534_446#_c_1381_n N_A_1349_114#_c_1584_n 0.0175173f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_966 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1584_n 8.48859e-19 $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_967 N_A_1534_446#_c_1381_n N_A_1349_114#_c_1585_n 0.0118206f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_968 N_A_1534_446#_c_1382_n N_A_1349_114#_c_1585_n 0.00293763f $X=8.055
+ $Y=2.215 $X2=0 $Y2=0
cc_969 N_A_1534_446#_M1004_g N_RESET_B_M1011_g 0.0309566f $X=11.435 $Y=2.4 $X2=0
+ $Y2=0
cc_970 N_A_1534_446#_c_1385_n N_RESET_B_M1011_g 0.00399864f $X=10.155 $Y=2.63
+ $X2=0 $Y2=0
cc_971 N_A_1534_446#_c_1386_n N_RESET_B_M1011_g 0.0203106f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_972 N_A_1534_446#_c_1387_n N_RESET_B_M1011_g 0.0085913f $X=11.3 $Y=2.29 $X2=0
+ $Y2=0
cc_973 N_A_1534_446#_M1029_g N_RESET_B_M1008_g 0.0144563f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_974 N_A_1534_446#_c_1372_n N_RESET_B_M1008_g 0.013621f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_975 N_A_1534_446#_c_1374_n N_RESET_B_M1008_g 0.0174418f $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_976 N_A_1534_446#_c_1375_n N_RESET_B_M1008_g 0.00614026f $X=11.4 $Y=1.32
+ $X2=0 $Y2=0
cc_977 N_A_1534_446#_M1004_g N_RESET_B_c_1720_n 0.00101722f $X=11.435 $Y=2.4
+ $X2=0 $Y2=0
cc_978 N_A_1534_446#_c_1373_n N_RESET_B_c_1720_n 0.00614026f $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_979 N_A_1534_446#_M1004_g N_RESET_B_c_1721_n 3.16946e-19 $X=11.435 $Y=2.4
+ $X2=0 $Y2=0
cc_980 N_A_1534_446#_c_1372_n N_RESET_B_c_1721_n 0.00326943f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_981 N_A_1534_446#_c_1386_n N_RESET_B_c_1721_n 0.0047568f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_982 N_A_1534_446#_c_1373_n N_RESET_B_c_1721_n 0.0302494f $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_983 N_A_1534_446#_c_1374_n N_RESET_B_c_1721_n 3.51317e-19 $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_984 N_A_1534_446#_c_1380_n N_A_2412_410#_M1037_g 0.0176603f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_985 N_A_1534_446#_c_1371_n N_A_2412_410#_M1037_g 0.0021724f $X=12.19 $Y=1.477
+ $X2=0 $Y2=0
cc_986 N_A_1534_446#_c_1367_n N_A_2412_410#_M1009_g 0.00197661f $X=12.19 $Y=1.32
+ $X2=0 $Y2=0
cc_987 N_A_1534_446#_c_1369_n N_A_2412_410#_M1009_g 0.016648f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_988 N_A_1534_446#_c_1367_n N_A_2412_410#_c_1758_n 0.018228f $X=12.19 $Y=1.32
+ $X2=0 $Y2=0
cc_989 N_A_1534_446#_c_1380_n N_A_2412_410#_c_1758_n 3.10137e-19 $X=12.42
+ $Y=1.975 $X2=0 $Y2=0
cc_990 N_A_1534_446#_c_1370_n N_A_2412_410#_c_1758_n 0.00217096f $X=12.465
+ $Y=0.94 $X2=0 $Y2=0
cc_991 N_A_1534_446#_M1029_g N_A_2412_410#_c_1760_n 0.00269951f $X=11.505
+ $Y=0.795 $X2=0 $Y2=0
cc_992 N_A_1534_446#_c_1367_n N_A_2412_410#_c_1760_n 0.00692844f $X=12.19
+ $Y=1.32 $X2=0 $Y2=0
cc_993 N_A_1534_446#_c_1369_n N_A_2412_410#_c_1760_n 0.00313626f $X=12.465
+ $Y=0.865 $X2=0 $Y2=0
cc_994 N_A_1534_446#_c_1370_n N_A_2412_410#_c_1760_n 0.0152083f $X=12.465
+ $Y=0.94 $X2=0 $Y2=0
cc_995 N_A_1534_446#_M1004_g N_A_2412_410#_c_1761_n 0.00170177f $X=11.435 $Y=2.4
+ $X2=0 $Y2=0
cc_996 N_A_1534_446#_c_1366_n N_A_2412_410#_c_1761_n 7.12587e-19 $X=12.115
+ $Y=1.477 $X2=0 $Y2=0
cc_997 N_A_1534_446#_c_1368_n N_A_2412_410#_c_1761_n 0.0053475f $X=12.19
+ $Y=1.825 $X2=0 $Y2=0
cc_998 N_A_1534_446#_c_1380_n N_A_2412_410#_c_1761_n 0.0299248f $X=12.42
+ $Y=1.975 $X2=0 $Y2=0
cc_999 N_A_1534_446#_c_1371_n N_A_2412_410#_c_1761_n 0.00124729f $X=12.19
+ $Y=1.477 $X2=0 $Y2=0
cc_1000 N_A_1534_446#_c_1380_n N_A_2412_410#_c_1762_n 0.00598615f $X=12.42
+ $Y=1.975 $X2=0 $Y2=0
cc_1001 N_A_1534_446#_c_1370_n N_A_2412_410#_c_1762_n 0.00601101f $X=12.465
+ $Y=0.94 $X2=0 $Y2=0
cc_1002 N_A_1534_446#_c_1366_n N_A_2412_410#_c_1763_n 0.00411413f $X=12.115
+ $Y=1.477 $X2=0 $Y2=0
cc_1003 N_A_1534_446#_c_1367_n N_A_2412_410#_c_1763_n 0.00204812f $X=12.19
+ $Y=1.32 $X2=0 $Y2=0
cc_1004 N_A_1534_446#_c_1371_n N_A_2412_410#_c_1763_n 0.00650752f $X=12.19
+ $Y=1.477 $X2=0 $Y2=0
cc_1005 N_A_1534_446#_c_1381_n N_VPWR_M1023_d 0.00278191f $X=8.055 $Y=2.215
+ $X2=0 $Y2=0
cc_1006 N_A_1534_446#_c_1499_p N_VPWR_M1023_d 0.00618434f $X=8.22 $Y=2.715 $X2=0
+ $Y2=0
cc_1007 N_A_1534_446#_c_1388_n N_VPWR_M1023_d 7.35761e-19 $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1008 N_A_1534_446#_c_1383_n N_VPWR_M1025_d 0.00742597f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1009 N_A_1534_446#_c_1386_n N_VPWR_M1011_d 0.00845613f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_1010 N_A_1534_446#_c_1387_n N_VPWR_M1011_d 0.00532651f $X=11.3 $Y=2.29 $X2=0
+ $Y2=0
cc_1011 N_A_1534_446#_M1004_g N_VPWR_c_1817_n 0.0127341f $X=11.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1012 N_A_1534_446#_c_1386_n N_VPWR_c_1817_n 0.0223125f $X=11.215 $Y=2.375
+ $X2=0 $Y2=0
cc_1013 N_A_1534_446#_c_1380_n N_VPWR_c_1818_n 0.00894788f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_1014 N_A_1534_446#_M1023_g N_VPWR_c_1825_n 0.00553757f $X=7.76 $Y=2.75 $X2=0
+ $Y2=0
cc_1015 N_A_1534_446#_c_1383_n N_VPWR_c_1826_n 0.00283252f $X=9.99 $Y=2.715
+ $X2=0 $Y2=0
cc_1016 N_A_1534_446#_c_1388_n N_VPWR_c_1826_n 0.00532338f $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1017 N_A_1534_446#_c_1389_n N_VPWR_c_1826_n 0.0139012f $X=8.83 $Y=2.805 $X2=0
+ $Y2=0
cc_1018 N_A_1534_446#_c_1383_n N_VPWR_c_1827_n 0.0255903f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1019 N_A_1534_446#_M1004_g N_VPWR_c_1828_n 0.00460063f $X=11.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1020 N_A_1534_446#_c_1380_n N_VPWR_c_1828_n 0.00604985f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_1021 N_A_1534_446#_M1023_g N_VPWR_c_1812_n 0.0109372f $X=7.76 $Y=2.75 $X2=0
+ $Y2=0
cc_1022 N_A_1534_446#_M1004_g N_VPWR_c_1812_n 0.00913687f $X=11.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1023 N_A_1534_446#_c_1380_n N_VPWR_c_1812_n 0.00628405f $X=12.42 $Y=1.975
+ $X2=0 $Y2=0
cc_1024 N_A_1534_446#_c_1499_p N_VPWR_c_1812_n 0.00249612f $X=8.22 $Y=2.715
+ $X2=0 $Y2=0
cc_1025 N_A_1534_446#_c_1383_n N_VPWR_c_1812_n 0.0346754f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1026 N_A_1534_446#_c_1388_n N_VPWR_c_1812_n 0.00743467f $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1027 N_A_1534_446#_c_1389_n N_VPWR_c_1812_n 0.0117742f $X=8.83 $Y=2.805 $X2=0
+ $Y2=0
cc_1028 N_A_1534_446#_M1023_g N_VPWR_c_1833_n 0.00501581f $X=7.76 $Y=2.75 $X2=0
+ $Y2=0
cc_1029 N_A_1534_446#_c_1382_n N_VPWR_c_1833_n 0.00108791f $X=8.055 $Y=2.215
+ $X2=0 $Y2=0
cc_1030 N_A_1534_446#_c_1499_p N_VPWR_c_1833_n 0.0254138f $X=8.22 $Y=2.715 $X2=0
+ $Y2=0
cc_1031 N_A_1534_446#_c_1388_n N_VPWR_c_1833_n 0.00362066f $X=8.5 $Y=2.805 $X2=0
+ $Y2=0
cc_1032 N_A_1534_446#_c_1389_n N_VPWR_c_1833_n 6.13556e-19 $X=8.83 $Y=2.805
+ $X2=0 $Y2=0
cc_1033 N_A_1534_446#_c_1383_n N_VPWR_c_1834_n 0.0243858f $X=9.99 $Y=2.715 $X2=0
+ $Y2=0
cc_1034 N_A_1534_446#_c_1389_n N_VPWR_c_1834_n 6.21509e-19 $X=8.83 $Y=2.805
+ $X2=0 $Y2=0
cc_1035 N_A_1534_446#_c_1383_n A_1920_392# 0.00421874f $X=9.99 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1036 N_A_1534_446#_M1029_g N_Q_N_c_2097_n 0.0126598f $X=11.505 $Y=0.795 $X2=0
+ $Y2=0
cc_1037 N_A_1534_446#_c_1370_n N_Q_N_c_2097_n 9.53622e-19 $X=12.465 $Y=0.94
+ $X2=0 $Y2=0
cc_1038 N_A_1534_446#_M1029_g N_Q_N_c_2098_n 0.00219593f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1039 N_A_1534_446#_c_1366_n N_Q_N_c_2098_n 0.00254586f $X=12.115 $Y=1.477
+ $X2=0 $Y2=0
cc_1040 N_A_1534_446#_c_1367_n N_Q_N_c_2098_n 9.53622e-19 $X=12.19 $Y=1.32 $X2=0
+ $Y2=0
cc_1041 N_A_1534_446#_c_1373_n N_Q_N_c_2098_n 0.00203513f $X=11.42 $Y=1.485
+ $X2=0 $Y2=0
cc_1042 N_A_1534_446#_M1004_g Q_N 0.00171244f $X=11.435 $Y=2.4 $X2=0 $Y2=0
cc_1043 N_A_1534_446#_c_1366_n Q_N 0.00531561f $X=12.115 $Y=1.477 $X2=0 $Y2=0
cc_1044 N_A_1534_446#_c_1380_n Q_N 0.00310181f $X=12.42 $Y=1.975 $X2=0 $Y2=0
cc_1045 N_A_1534_446#_c_1387_n Q_N 0.0152769f $X=11.3 $Y=2.29 $X2=0 $Y2=0
cc_1046 N_A_1534_446#_c_1373_n Q_N 6.77959e-19 $X=11.42 $Y=1.485 $X2=0 $Y2=0
cc_1047 N_A_1534_446#_c_1380_n Q_N 0.00133317f $X=12.42 $Y=1.975 $X2=0 $Y2=0
cc_1048 N_A_1534_446#_M1004_g N_Q_N_c_2099_n 0.00116846f $X=11.435 $Y=2.4 $X2=0
+ $Y2=0
cc_1049 N_A_1534_446#_M1029_g N_Q_N_c_2099_n 0.00120695f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1050 N_A_1534_446#_c_1366_n N_Q_N_c_2099_n 0.0218962f $X=12.115 $Y=1.477
+ $X2=0 $Y2=0
cc_1051 N_A_1534_446#_c_1368_n N_Q_N_c_2099_n 7.20579e-19 $X=12.19 $Y=1.825
+ $X2=0 $Y2=0
cc_1052 N_A_1534_446#_c_1387_n N_Q_N_c_2099_n 0.00479229f $X=11.3 $Y=2.29 $X2=0
+ $Y2=0
cc_1053 N_A_1534_446#_c_1373_n N_Q_N_c_2099_n 0.023841f $X=11.42 $Y=1.485 $X2=0
+ $Y2=0
cc_1054 N_A_1534_446#_c_1375_n N_Q_N_c_2099_n 0.00523611f $X=11.4 $Y=1.32 $X2=0
+ $Y2=0
cc_1055 N_A_1534_446#_c_1369_n Q 8.51067e-19 $X=12.465 $Y=0.865 $X2=0 $Y2=0
cc_1056 N_A_1534_446#_c_1372_n N_VGND_M1008_d 0.0100046f $X=11.215 $Y=0.68 $X2=0
+ $Y2=0
cc_1057 N_A_1534_446#_c_1375_n N_VGND_M1008_d 0.00783804f $X=11.4 $Y=1.32 $X2=0
+ $Y2=0
cc_1058 N_A_1534_446#_M1000_g N_VGND_c_2150_n 5.6876e-19 $X=8.37 $Y=0.91 $X2=0
+ $Y2=0
cc_1059 N_A_1534_446#_M1029_g N_VGND_c_2151_n 0.00513051f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1060 N_A_1534_446#_c_1372_n N_VGND_c_2151_n 0.025628f $X=11.215 $Y=0.68 $X2=0
+ $Y2=0
cc_1061 N_A_1534_446#_c_1369_n N_VGND_c_2152_n 0.00549585f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_1062 N_A_1534_446#_M1000_g N_VGND_c_2156_n 3.43662e-19 $X=8.37 $Y=0.91 $X2=0
+ $Y2=0
cc_1063 N_A_1534_446#_c_1372_n N_VGND_c_2157_n 0.0138172f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_1064 N_A_1534_446#_M1029_g N_VGND_c_2158_n 0.00514022f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1065 N_A_1534_446#_c_1369_n N_VGND_c_2158_n 0.00461464f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_1066 N_A_1534_446#_M1029_g N_VGND_c_2160_n 0.00528353f $X=11.505 $Y=0.795
+ $X2=0 $Y2=0
cc_1067 N_A_1534_446#_c_1369_n N_VGND_c_2160_n 0.00913666f $X=12.465 $Y=0.865
+ $X2=0 $Y2=0
cc_1068 N_A_1534_446#_c_1370_n N_VGND_c_2160_n 6.2279e-19 $X=12.465 $Y=0.94
+ $X2=0 $Y2=0
cc_1069 N_A_1534_446#_c_1372_n N_VGND_c_2160_n 0.0239625f $X=11.215 $Y=0.68
+ $X2=0 $Y2=0
cc_1070 N_A_1534_446#_c_1372_n N_A_1818_76#_M1033_d 0.00713159f $X=11.215
+ $Y=0.68 $X2=0 $Y2=0
cc_1071 N_A_1534_446#_M1034_d N_A_1818_76#_c_2312_n 0.00219516f $X=9.52 $Y=0.38
+ $X2=0 $Y2=0
cc_1072 N_A_1534_446#_c_1372_n N_A_1818_76#_c_2312_n 0.0466631f $X=11.215
+ $Y=0.68 $X2=0 $Y2=0
cc_1073 N_A_1349_114#_c_1570_n N_RESET_B_M1011_g 7.7731e-19 $X=10.005 $Y=1.585
+ $X2=0 $Y2=0
cc_1074 N_A_1349_114#_M1033_g N_RESET_B_c_1720_n 6.81196e-19 $X=9.915 $Y=0.75
+ $X2=0 $Y2=0
cc_1075 N_A_1349_114#_c_1570_n N_RESET_B_c_1720_n 0.00419861f $X=10.005 $Y=1.585
+ $X2=0 $Y2=0
cc_1076 N_A_1349_114#_c_1647_n N_VPWR_M1025_d 0.0119567f $X=9.23 $Y=2.375 $X2=0
+ $Y2=0
cc_1077 N_A_1349_114#_c_1651_n N_VPWR_M1025_d 0.00245622f $X=9.315 $Y=2.29 $X2=0
+ $Y2=0
cc_1078 N_A_1349_114#_c_1580_n N_VPWR_M1025_d 0.00140515f $X=9.4 $Y=2.035 $X2=0
+ $Y2=0
cc_1079 N_A_1349_114#_c_1572_n N_VPWR_c_1816_n 0.0101933f $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1080 N_A_1349_114#_c_1572_n N_VPWR_c_1825_n 0.0240985f $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1081 N_A_1349_114#_M1026_g N_VPWR_c_1827_n 0.00421707f $X=9.93 $Y=2.46 $X2=0
+ $Y2=0
cc_1082 N_A_1349_114#_M1026_g N_VPWR_c_1812_n 0.00638115f $X=9.93 $Y=2.46 $X2=0
+ $Y2=0
cc_1083 N_A_1349_114#_c_1572_n N_VPWR_c_1812_n 0.0194932f $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1084 N_A_1349_114#_c_1572_n N_VPWR_c_1833_n 3.72707e-19 $X=7.025 $Y=2.815
+ $X2=0 $Y2=0
cc_1085 N_A_1349_114#_c_1579_n A_1920_392# 0.00230006f $X=9.84 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_1086 N_A_1349_114#_M1033_g N_VGND_c_2157_n 0.00390708f $X=9.915 $Y=0.75 $X2=0
+ $Y2=0
cc_1087 N_A_1349_114#_M1033_g N_VGND_c_2160_n 0.00542671f $X=9.915 $Y=0.75 $X2=0
+ $Y2=0
cc_1088 N_A_1349_114#_c_1567_n A_1611_140# 0.0026403f $X=8.035 $Y=0.845
+ $X2=-0.19 $Y2=-0.245
cc_1089 N_A_1349_114#_c_1568_n A_1611_140# 9.34402e-19 $X=8.12 $Y=1.73 $X2=-0.19
+ $Y2=-0.245
cc_1090 N_A_1349_114#_M1033_g N_A_1818_76#_c_2312_n 0.0108598f $X=9.915 $Y=0.75
+ $X2=0 $Y2=0
cc_1091 N_RESET_B_M1011_g N_VPWR_c_1827_n 0.00377165f $X=10.91 $Y=2.16 $X2=0
+ $Y2=0
cc_1092 N_RESET_B_M1011_g N_VPWR_c_1812_n 0.00493777f $X=10.91 $Y=2.16 $X2=0
+ $Y2=0
cc_1093 N_RESET_B_M1008_g N_VGND_c_2157_n 5.97925e-19 $X=10.94 $Y=0.955 $X2=0
+ $Y2=0
cc_1094 N_A_2412_410#_M1037_g N_VPWR_c_1818_n 0.00464648f $X=12.945 $Y=2.4 $X2=0
+ $Y2=0
cc_1095 N_A_2412_410#_c_1758_n N_VPWR_c_1818_n 0.00557956f $X=12.855 $Y=1.42
+ $X2=0 $Y2=0
cc_1096 N_A_2412_410#_c_1761_n N_VPWR_c_1818_n 0.0440876f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1097 N_A_2412_410#_c_1762_n N_VPWR_c_1818_n 0.016421f $X=12.67 $Y=1.42 $X2=0
+ $Y2=0
cc_1098 N_A_2412_410#_c_1761_n N_VPWR_c_1828_n 0.00854762f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1099 N_A_2412_410#_M1037_g N_VPWR_c_1829_n 0.005209f $X=12.945 $Y=2.4 $X2=0
+ $Y2=0
cc_1100 N_A_2412_410#_M1037_g N_VPWR_c_1812_n 0.00991105f $X=12.945 $Y=2.4 $X2=0
+ $Y2=0
cc_1101 N_A_2412_410#_c_1761_n N_VPWR_c_1812_n 0.00873555f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1102 N_A_2412_410#_c_1760_n N_Q_N_c_2097_n 0.0657174f $X=12.25 $Y=0.58 $X2=0
+ $Y2=0
cc_1103 N_A_2412_410#_c_1761_n N_Q_N_c_2099_n 0.0999719f $X=12.195 $Y=2.195
+ $X2=0 $Y2=0
cc_1104 N_A_2412_410#_c_1763_n N_Q_N_c_2099_n 0.0240258f $X=12.235 $Y=1.42 $X2=0
+ $Y2=0
cc_1105 N_A_2412_410#_M1037_g Q 0.0261178f $X=12.945 $Y=2.4 $X2=0 $Y2=0
cc_1106 N_A_2412_410#_M1009_g Q 0.0190895f $X=12.96 $Y=0.74 $X2=0 $Y2=0
cc_1107 N_A_2412_410#_c_1759_n Q 0.0121736f $X=12.945 $Y=1.42 $X2=0 $Y2=0
cc_1108 N_A_2412_410#_c_1760_n Q 0.0118818f $X=12.25 $Y=0.58 $X2=0 $Y2=0
cc_1109 N_A_2412_410#_c_1761_n Q 0.00657613f $X=12.195 $Y=2.195 $X2=0 $Y2=0
cc_1110 N_A_2412_410#_c_1762_n Q 0.026211f $X=12.67 $Y=1.42 $X2=0 $Y2=0
cc_1111 N_A_2412_410#_M1009_g N_VGND_c_2152_n 0.00330721f $X=12.96 $Y=0.74 $X2=0
+ $Y2=0
cc_1112 N_A_2412_410#_c_1758_n N_VGND_c_2152_n 0.0048385f $X=12.855 $Y=1.42
+ $X2=0 $Y2=0
cc_1113 N_A_2412_410#_c_1760_n N_VGND_c_2152_n 0.00252997f $X=12.25 $Y=0.58
+ $X2=0 $Y2=0
cc_1114 N_A_2412_410#_c_1762_n N_VGND_c_2152_n 0.00977708f $X=12.67 $Y=1.42
+ $X2=0 $Y2=0
cc_1115 N_A_2412_410#_c_1760_n N_VGND_c_2158_n 0.011066f $X=12.25 $Y=0.58 $X2=0
+ $Y2=0
cc_1116 N_A_2412_410#_M1009_g N_VGND_c_2159_n 0.00428607f $X=12.96 $Y=0.74 $X2=0
+ $Y2=0
cc_1117 N_A_2412_410#_M1009_g N_VGND_c_2160_n 0.00806216f $X=12.96 $Y=0.74 $X2=0
+ $Y2=0
cc_1118 N_A_2412_410#_c_1760_n N_VGND_c_2160_n 0.00915947f $X=12.25 $Y=0.58
+ $X2=0 $Y2=0
cc_1119 N_VPWR_c_1817_n Q_N 0.0122422f $X=11.21 $Y=2.805 $X2=0 $Y2=0
cc_1120 N_VPWR_c_1818_n Q_N 0.00227672f $X=12.72 $Y=1.985 $X2=0 $Y2=0
cc_1121 N_VPWR_c_1828_n Q_N 0.0155281f $X=12.555 $Y=3.33 $X2=0 $Y2=0
cc_1122 N_VPWR_c_1812_n Q_N 0.0128528f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1123 N_VPWR_c_1818_n Q 0.0396567f $X=12.72 $Y=1.985 $X2=0 $Y2=0
cc_1124 N_VPWR_c_1829_n Q 0.0147721f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1125 N_VPWR_c_1812_n Q 0.0121589f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1126 N_A_311_119#_c_1985_n N_VGND_M1014_d 0.00783807f $X=2.58 $Y=0.925 $X2=0
+ $Y2=0
cc_1127 N_A_311_119#_c_1985_n N_VGND_c_2148_n 0.0287269f $X=2.58 $Y=0.925 $X2=0
+ $Y2=0
cc_1128 N_A_311_119#_c_1969_n N_VGND_c_2148_n 0.0155564f $X=2.665 $Y=0.84 $X2=0
+ $Y2=0
cc_1129 N_A_311_119#_c_1970_n N_VGND_c_2148_n 0.0151473f $X=2.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1130 N_A_311_119#_c_1975_n N_VGND_c_2148_n 0.00409119f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1131 N_A_311_119#_c_1975_n N_VGND_c_2154_n 0.00626553f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1132 N_A_311_119#_c_1970_n N_VGND_c_2155_n 0.0115893f $X=2.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1133 N_A_311_119#_c_1971_n N_VGND_c_2155_n 0.0115893f $X=3.975 $Y=0.435 $X2=0
+ $Y2=0
cc_1134 N_A_311_119#_c_1977_n N_VGND_c_2155_n 0.0801396f $X=3.46 $Y=0.435 $X2=0
+ $Y2=0
cc_1135 N_A_311_119#_c_1985_n N_VGND_c_2160_n 0.0111714f $X=2.58 $Y=0.925 $X2=0
+ $Y2=0
cc_1136 N_A_311_119#_c_1970_n N_VGND_c_2160_n 0.00583135f $X=2.75 $Y=0.34 $X2=0
+ $Y2=0
cc_1137 N_A_311_119#_c_1971_n N_VGND_c_2160_n 0.00583135f $X=3.975 $Y=0.435
+ $X2=0 $Y2=0
cc_1138 N_A_311_119#_c_1975_n N_VGND_c_2160_n 0.00761936f $X=1.7 $Y=0.79 $X2=0
+ $Y2=0
cc_1139 N_A_311_119#_c_1977_n N_VGND_c_2160_n 0.0413441f $X=3.46 $Y=0.435 $X2=0
+ $Y2=0
cc_1140 N_A_311_119#_c_1985_n A_523_119# 0.00260391f $X=2.58 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_1141 N_A_311_119#_c_1969_n A_523_119# 0.00211902f $X=2.665 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_1142 N_A_311_119#_c_1978_n N_A_867_119#_M1020_s 0.00382131f $X=4.39 $Y=1.08
+ $X2=-0.19 $Y2=-0.245
cc_1143 N_A_311_119#_c_1971_n N_A_867_119#_c_2279_n 0.0167755f $X=3.975 $Y=0.435
+ $X2=0 $Y2=0
cc_1144 N_A_311_119#_c_1973_n N_A_867_119#_c_2279_n 0.0166121f $X=4.06 $Y=0.995
+ $X2=0 $Y2=0
cc_1145 N_A_311_119#_c_1978_n N_A_867_119#_c_2279_n 0.0121158f $X=4.39 $Y=1.08
+ $X2=0 $Y2=0
cc_1146 N_A_311_119#_c_1971_n N_A_867_119#_c_2281_n 0.0159286f $X=3.975 $Y=0.435
+ $X2=0 $Y2=0
cc_1147 N_Q_N_c_2097_n N_VGND_c_2151_n 0.00159581f $X=11.72 $Y=0.57 $X2=0 $Y2=0
cc_1148 N_Q_N_c_2097_n N_VGND_c_2158_n 0.0133729f $X=11.72 $Y=0.57 $X2=0 $Y2=0
cc_1149 N_Q_N_c_2097_n N_VGND_c_2160_n 0.0131093f $X=11.72 $Y=0.57 $X2=0 $Y2=0
cc_1150 Q N_VGND_c_2152_n 0.0176449f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1151 Q N_VGND_c_2159_n 0.0147721f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1152 Q N_VGND_c_2160_n 0.0121589f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1153 N_VGND_c_2149_n N_A_867_119#_c_2280_n 0.0150385f $X=5.98 $Y=0.87 $X2=0
+ $Y2=0
cc_1154 N_VGND_c_2155_n N_A_867_119#_c_2280_n 0.0655844f $X=5.815 $Y=0 $X2=0
+ $Y2=0
cc_1155 N_VGND_c_2160_n N_A_867_119#_c_2280_n 0.0338323f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1156 N_VGND_c_2155_n N_A_867_119#_c_2281_n 0.0222128f $X=5.815 $Y=0 $X2=0
+ $Y2=0
cc_1157 N_VGND_c_2160_n N_A_867_119#_c_2281_n 0.0112618f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1158 N_VGND_c_2149_n N_A_867_119#_c_2282_n 0.030044f $X=5.98 $Y=0.87 $X2=0
+ $Y2=0
cc_1159 N_VGND_c_2160_n N_A_1818_76#_M1033_d 0.00252807f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1160 N_VGND_c_2150_n N_A_1818_76#_c_2311_n 0.0113368f $X=8.8 $Y=0.56 $X2=0
+ $Y2=0
cc_1161 N_VGND_c_2157_n N_A_1818_76#_c_2311_n 0.0174569f $X=11.055 $Y=0 $X2=0
+ $Y2=0
cc_1162 N_VGND_c_2160_n N_A_1818_76#_c_2311_n 0.00963343f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1163 N_VGND_c_2157_n N_A_1818_76#_c_2312_n 0.0661462f $X=11.055 $Y=0 $X2=0
+ $Y2=0
cc_1164 N_VGND_c_2160_n N_A_1818_76#_c_2312_n 0.039116f $X=13.2 $Y=0 $X2=0 $Y2=0

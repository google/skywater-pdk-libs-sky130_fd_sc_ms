* File: sky130_fd_sc_ms__bufinv_16.pex.spice
* Created: Wed Sep  2 12:00:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__BUFINV_16%A 3 7 11 15 19 23 25 26 27 41 43
c67 19 0 5.24737e-20 $X=1.41 $Y=2.4
r68 42 43 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.415 $Y2=1.515
r69 40 42 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.265 $Y=1.515
+ $X2=1.41 $Y2=1.515
r70 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r71 38 40 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=0.985 $Y=1.515
+ $X2=1.265 $Y2=1.515
r72 37 38 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.985 $Y2=1.515
r73 35 37 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.96 $Y2=1.515
r74 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r75 33 35 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.515
+ $X2=0.585 $Y2=1.515
r76 31 33 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.51 $Y2=1.515
r77 27 41 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r78 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r79 26 36 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r80 25 36 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r81 21 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.35
+ $X2=1.415 $Y2=1.515
r82 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.415 $Y=1.35
+ $X2=1.415 $Y2=0.74
r83 17 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.68
+ $X2=1.41 $Y2=1.515
r84 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.41 $Y=1.68
+ $X2=1.41 $Y2=2.4
r85 13 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=1.515
r86 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=0.74
r87 9 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=1.515
r88 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.96 $Y=1.68 $X2=0.96
+ $Y2=2.4
r89 5 33 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.68
+ $X2=0.51 $Y2=1.515
r90 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.51 $Y=1.68 $X2=0.51
+ $Y2=2.4
r91 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r92 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__BUFINV_16%A_27_74# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 53 57 61 63 66 68 70 72 73 74 78 82 84 86 89 95 101 102 103 119
c207 15 0 1.71373e-19 $X=1.845 $Y=0.74
r208 118 119 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.68 $Y=1.465
+ $X2=3.77 $Y2=1.465
r209 117 118 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.635 $Y=1.465
+ $X2=3.68 $Y2=1.465
r210 114 115 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.135 $Y=1.465
+ $X2=3.23 $Y2=1.465
r211 113 114 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.78 $Y=1.465
+ $X2=3.135 $Y2=1.465
r212 112 113 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=1.465
+ $X2=2.78 $Y2=1.465
r213 111 112 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.33 $Y=1.465
+ $X2=2.705 $Y2=1.465
r214 110 111 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.275 $Y=1.465
+ $X2=2.33 $Y2=1.465
r215 106 108 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.845 $Y=1.465
+ $X2=1.86 $Y2=1.465
r216 96 117 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.295 $Y=1.465
+ $X2=3.635 $Y2=1.465
r217 96 115 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.295 $Y=1.465
+ $X2=3.23 $Y2=1.465
r218 95 96 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.295
+ $Y=1.465 $X2=3.295 $Y2=1.465
r219 93 110 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.935 $Y=1.465
+ $X2=2.275 $Y2=1.465
r220 93 108 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.465
+ $X2=1.86 $Y2=1.465
r221 92 95 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=1.935 $Y=1.465
+ $X2=3.295 $Y2=1.465
r222 92 93 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.935
+ $Y=1.465 $X2=1.935 $Y2=1.465
r223 90 103 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.465
+ $X2=1.685 $Y2=1.095
r224 90 92 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=1.465
+ $X2=1.935 $Y2=1.465
r225 88 90 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.63
+ $X2=1.685 $Y2=1.465
r226 88 89 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.685 $Y=1.63
+ $X2=1.685 $Y2=1.95
r227 87 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=2.035
+ $X2=1.185 $Y2=2.035
r228 86 89 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=1.685 $Y2=1.95
r229 86 87 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=1.35 $Y2=2.035
r230 85 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.095
+ $X2=1.2 $Y2=1.095
r231 84 103 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=1.095
+ $X2=1.685 $Y2=1.095
r232 84 85 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.6 $Y=1.095
+ $X2=1.285 $Y2=1.095
r233 80 102 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.01 $X2=1.2
+ $Y2=1.095
r234 80 82 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.2 $Y=1.01
+ $X2=1.2 $Y2=0.515
r235 76 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r236 76 78 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r237 75 99 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=2.035
+ $X2=0.285 $Y2=2.035
r238 74 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.185 $Y2=2.035
r239 74 75 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.45 $Y2=2.035
r240 72 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.2 $Y2=1.095
r241 72 73 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.365 $Y2=1.095
r242 68 99 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.035
r243 68 70 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.815
r244 64 73 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r245 64 66 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r246 59 63 18.8402 $w=1.65e-07 $l=8.66025e-08 $layer=POLY_cond $X=4.13 $Y=1.45
+ $X2=4.105 $Y2=1.375
r247 59 61 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=4.13 $Y=1.45
+ $X2=4.13 $Y2=2.4
r248 55 63 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.065 $Y=1.3
+ $X2=4.105 $Y2=1.375
r249 55 57 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.065 $Y=1.3
+ $X2=4.065 $Y2=0.74
r250 53 63 6.66866 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=3.99 $Y=1.375
+ $X2=4.105 $Y2=1.375
r251 53 119 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.99 $Y=1.375
+ $X2=3.77 $Y2=1.375
r252 49 118 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.63
+ $X2=3.68 $Y2=1.465
r253 49 51 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.68 $Y=1.63
+ $X2=3.68 $Y2=2.4
r254 45 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=1.3
+ $X2=3.635 $Y2=1.465
r255 45 47 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.635 $Y=1.3
+ $X2=3.635 $Y2=0.74
r256 41 115 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.63
+ $X2=3.23 $Y2=1.465
r257 41 43 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.23 $Y=1.63
+ $X2=3.23 $Y2=2.4
r258 37 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.135 $Y=1.3
+ $X2=3.135 $Y2=1.465
r259 37 39 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.135 $Y=1.3
+ $X2=3.135 $Y2=0.74
r260 33 113 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.63
+ $X2=2.78 $Y2=1.465
r261 33 35 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.78 $Y=1.63
+ $X2=2.78 $Y2=2.4
r262 29 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.3
+ $X2=2.705 $Y2=1.465
r263 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.705 $Y=1.3
+ $X2=2.705 $Y2=0.74
r264 25 111 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.63
+ $X2=2.33 $Y2=1.465
r265 25 27 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.33 $Y=1.63
+ $X2=2.33 $Y2=2.4
r266 21 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.3
+ $X2=2.275 $Y2=1.465
r267 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.275 $Y=1.3
+ $X2=2.275 $Y2=0.74
r268 17 108 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.63
+ $X2=1.86 $Y2=1.465
r269 17 19 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.86 $Y=1.63
+ $X2=1.86 $Y2=2.4
r270 13 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.3
+ $X2=1.845 $Y2=1.465
r271 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.845 $Y=1.3
+ $X2=1.845 $Y2=0.74
r272 4 101 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.115
r273 4 78 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.815
r274 3 99 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r275 3 70 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r276 2 82 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.37 $X2=1.2 $Y2=0.515
r277 1 66 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFINV_16%A_384_74# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 155 157 158 159 160 163 167 171 173 177 179 181 185 186 210 220
+ 227 234 241 248 255 262 266
c468 160 0 5.24737e-20 $X=2.27 $Y=1.885
c469 158 0 1.71373e-19 $X=2.145 $Y=1.045
r470 265 266 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=11.435 $Y=1.465
+ $X2=11.48 $Y2=1.465
r471 264 265 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=11.005 $Y=1.465
+ $X2=11.435 $Y2=1.465
r472 263 264 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=10.99 $Y=1.465
+ $X2=11.005 $Y2=1.465
r473 261 263 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=10.71 $Y=1.465
+ $X2=10.99 $Y2=1.465
r474 261 262 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.71
+ $Y=1.465 $X2=10.71 $Y2=1.465
r475 259 261 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=10.53 $Y=1.465
+ $X2=10.71 $Y2=1.465
r476 258 259 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=10.505 $Y=1.465
+ $X2=10.53 $Y2=1.465
r477 257 258 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=10.08 $Y=1.465
+ $X2=10.505 $Y2=1.465
r478 256 257 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=10.075 $Y=1.465
+ $X2=10.08 $Y2=1.465
r479 254 256 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=9.78 $Y=1.465
+ $X2=10.075 $Y2=1.465
r480 254 255 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.465 $X2=9.78 $Y2=1.465
r481 252 254 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=9.58 $Y=1.465
+ $X2=9.78 $Y2=1.465
r482 251 252 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=9.575 $Y=1.465
+ $X2=9.58 $Y2=1.465
r483 250 251 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=9.145 $Y=1.465
+ $X2=9.575 $Y2=1.465
r484 249 250 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.13 $Y=1.465
+ $X2=9.145 $Y2=1.465
r485 247 249 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=8.85 $Y=1.465
+ $X2=9.13 $Y2=1.465
r486 247 248 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.85
+ $Y=1.465 $X2=8.85 $Y2=1.465
r487 245 247 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=8.645 $Y=1.465
+ $X2=8.85 $Y2=1.465
r488 244 245 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.63 $Y=1.465
+ $X2=8.645 $Y2=1.465
r489 243 244 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.215 $Y=1.465
+ $X2=8.63 $Y2=1.465
r490 242 243 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.18 $Y=1.465
+ $X2=8.215 $Y2=1.465
r491 240 242 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=7.925 $Y=1.465
+ $X2=8.18 $Y2=1.465
r492 240 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.925
+ $Y=1.465 $X2=7.925 $Y2=1.465
r493 238 240 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=7.73 $Y=1.465
+ $X2=7.925 $Y2=1.465
r494 237 238 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.715 $Y=1.465
+ $X2=7.73 $Y2=1.465
r495 236 237 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.285 $Y=1.465
+ $X2=7.715 $Y2=1.465
r496 235 236 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.28 $Y=1.465
+ $X2=7.285 $Y2=1.465
r497 233 235 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=7.005 $Y=1.465
+ $X2=7.28 $Y2=1.465
r498 233 234 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.005
+ $Y=1.465 $X2=7.005 $Y2=1.465
r499 231 233 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.83 $Y=1.465
+ $X2=7.005 $Y2=1.465
r500 230 231 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.785 $Y=1.465
+ $X2=6.83 $Y2=1.465
r501 229 230 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=6.38 $Y=1.465
+ $X2=6.785 $Y2=1.465
r502 228 229 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.355 $Y=1.465
+ $X2=6.38 $Y2=1.465
r503 226 228 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=6.065 $Y=1.465
+ $X2=6.355 $Y2=1.465
r504 226 227 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.465 $X2=6.065 $Y2=1.465
r505 224 226 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.465
+ $X2=6.065 $Y2=1.465
r506 223 224 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.855 $Y=1.465
+ $X2=5.93 $Y2=1.465
r507 222 223 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.48 $Y=1.465
+ $X2=5.855 $Y2=1.465
r508 221 222 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=5.425 $Y=1.465
+ $X2=5.48 $Y2=1.465
r509 219 221 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.175 $Y=1.465
+ $X2=5.425 $Y2=1.465
r510 219 220 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.465 $X2=5.175 $Y2=1.465
r511 217 219 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.03 $Y=1.465
+ $X2=5.175 $Y2=1.465
r512 216 217 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.995 $Y=1.465
+ $X2=5.03 $Y2=1.465
r513 215 216 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=4.58 $Y=1.465
+ $X2=4.995 $Y2=1.465
r514 213 215 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.565 $Y=1.465
+ $X2=4.58 $Y2=1.465
r515 211 262 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=10.71 $Y=1.665
+ $X2=10.71 $Y2=1.465
r516 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.71 $Y=1.665
+ $X2=10.71 $Y2=1.665
r517 208 255 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=9.78 $Y=1.665
+ $X2=9.78 $Y2=1.465
r518 207 210 0.5999 $w=2.3e-07 $l=9.35e-07 $layer=MET1_cond $X=9.775 $Y=1.665
+ $X2=10.71 $Y2=1.665
r519 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.775 $Y=1.665
+ $X2=9.775 $Y2=1.665
r520 205 248 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=8.85 $Y=1.665
+ $X2=8.85 $Y2=1.465
r521 204 207 0.593484 $w=2.3e-07 $l=9.25e-07 $layer=MET1_cond $X=8.85 $Y=1.665
+ $X2=9.775 $Y2=1.665
r522 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.85 $Y=1.665
+ $X2=8.85 $Y2=1.665
r523 202 241 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.925 $Y=1.665
+ $X2=7.925 $Y2=1.465
r524 201 204 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=7.92 $Y=1.665
+ $X2=8.85 $Y2=1.665
r525 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r526 199 234 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.005 $Y=1.665
+ $X2=7.005 $Y2=1.465
r527 198 201 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=7.005 $Y=1.665
+ $X2=7.92 $Y2=1.665
r528 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.005 $Y=1.665
+ $X2=7.005 $Y2=1.665
r529 196 227 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.065 $Y=1.665
+ $X2=6.065 $Y2=1.465
r530 195 198 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=6.065 $Y=1.665
+ $X2=7.005 $Y2=1.665
r531 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.065 $Y=1.665
+ $X2=6.065 $Y2=1.665
r532 193 220 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=5.17 $Y=1.665
+ $X2=5.17 $Y2=1.465
r533 192 195 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=5.175 $Y=1.665
+ $X2=6.065 $Y2=1.665
r534 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.665
+ $X2=5.175 $Y2=1.665
r535 189 298 5.77204 $w=4.65e-07 $l=2.2e-07 $layer=LI1_cond $X=4.06 $Y=1.665
+ $X2=4.06 $Y2=1.885
r536 188 192 0.554988 $w=2.3e-07 $l=8.65e-07 $layer=MET1_cond $X=4.31 $Y=1.665
+ $X2=5.175 $Y2=1.665
r537 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.31 $Y=1.665
+ $X2=4.31 $Y2=1.665
r538 181 183 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.905 $Y=1.985
+ $X2=3.905 $Y2=2.815
r539 179 298 3.27514 $w=4.65e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.905 $Y=1.97
+ $X2=4.06 $Y2=1.885
r540 179 181 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.905 $Y=1.97
+ $X2=3.905 $Y2=1.985
r541 175 177 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.81 $Y=0.96
+ $X2=3.81 $Y2=0.515
r542 174 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=1.885
+ $X2=3.005 $Y2=1.885
r543 173 298 6.7035 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=3.74 $Y=1.885
+ $X2=4.06 $Y2=1.885
r544 173 174 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.74 $Y=1.885
+ $X2=3.17 $Y2=1.885
r545 172 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.005 $Y=1.045
+ $X2=2.88 $Y2=1.045
r546 171 189 16.2667 $w=4.65e-07 $l=7.8543e-07 $layer=LI1_cond $X=3.685 $Y=1.045
+ $X2=4.06 $Y2=1.665
r547 171 175 4.82172 $w=4.65e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685
+ $Y=1.045 $X2=3.81 $Y2=0.96
r548 171 172 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.685 $Y=1.045
+ $X2=3.005 $Y2=1.045
r549 167 169 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.005 $Y=1.985
+ $X2=3.005 $Y2=2.815
r550 165 186 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=1.97
+ $X2=3.005 $Y2=1.885
r551 165 167 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.005 $Y=1.97
+ $X2=3.005 $Y2=1.985
r552 161 185 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.96
+ $X2=2.88 $Y2=1.045
r553 161 163 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.88 $Y=0.96
+ $X2=2.88 $Y2=0.515
r554 159 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=1.885
+ $X2=3.005 $Y2=1.885
r555 159 160 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.84 $Y=1.885
+ $X2=2.27 $Y2=1.885
r556 157 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=1.045
+ $X2=2.88 $Y2=1.045
r557 157 158 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.755 $Y=1.045
+ $X2=2.145 $Y2=1.045
r558 153 158 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=0.96
+ $X2=2.145 $Y2=1.045
r559 153 155 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.06 $Y=0.96
+ $X2=2.06 $Y2=0.515
r560 149 151 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.105 $Y=1.985
+ $X2=2.105 $Y2=2.815
r561 147 160 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.105 $Y=1.97
+ $X2=2.27 $Y2=1.885
r562 147 149 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.105 $Y=1.97
+ $X2=2.105 $Y2=1.985
r563 143 266 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.48 $Y=1.63
+ $X2=11.48 $Y2=1.465
r564 143 145 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.48 $Y=1.63
+ $X2=11.48 $Y2=2.4
r565 139 265 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.435 $Y=1.3
+ $X2=11.435 $Y2=1.465
r566 139 141 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.435 $Y=1.3
+ $X2=11.435 $Y2=0.74
r567 135 264 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.005 $Y=1.3
+ $X2=11.005 $Y2=1.465
r568 135 137 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.005 $Y=1.3
+ $X2=11.005 $Y2=0.74
r569 131 263 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.99 $Y=1.63
+ $X2=10.99 $Y2=1.465
r570 131 133 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.99 $Y=1.63
+ $X2=10.99 $Y2=2.4
r571 127 259 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.53 $Y=1.63
+ $X2=10.53 $Y2=1.465
r572 127 129 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.53 $Y=1.63
+ $X2=10.53 $Y2=2.4
r573 123 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.505 $Y=1.3
+ $X2=10.505 $Y2=1.465
r574 123 125 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.505 $Y=1.3
+ $X2=10.505 $Y2=0.74
r575 119 256 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.075 $Y=1.3
+ $X2=10.075 $Y2=1.465
r576 119 121 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.075 $Y=1.3
+ $X2=10.075 $Y2=0.74
r577 115 257 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.08 $Y=1.63
+ $X2=10.08 $Y2=1.465
r578 115 117 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.08 $Y=1.63
+ $X2=10.08 $Y2=2.4
r579 111 251 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.575 $Y=1.3
+ $X2=9.575 $Y2=1.465
r580 111 113 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.575 $Y=1.3
+ $X2=9.575 $Y2=0.74
r581 107 252 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.58 $Y=1.63
+ $X2=9.58 $Y2=1.465
r582 107 109 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=9.58 $Y=1.63
+ $X2=9.58 $Y2=2.4
r583 103 250 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.145 $Y=1.3
+ $X2=9.145 $Y2=1.465
r584 103 105 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.145 $Y=1.3
+ $X2=9.145 $Y2=0.74
r585 99 249 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.13 $Y=1.63
+ $X2=9.13 $Y2=1.465
r586 99 101 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=9.13 $Y=1.63
+ $X2=9.13 $Y2=2.4
r587 95 245 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.3
+ $X2=8.645 $Y2=1.465
r588 95 97 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.645 $Y=1.3
+ $X2=8.645 $Y2=0.74
r589 91 244 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.63
+ $X2=8.63 $Y2=1.465
r590 91 93 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.63 $Y=1.63
+ $X2=8.63 $Y2=2.4
r591 87 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=1.3
+ $X2=8.215 $Y2=1.465
r592 87 89 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.215 $Y=1.3
+ $X2=8.215 $Y2=0.74
r593 83 242 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.18 $Y=1.63
+ $X2=8.18 $Y2=1.465
r594 83 85 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.18 $Y=1.63
+ $X2=8.18 $Y2=2.4
r595 79 238 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.73 $Y=1.63
+ $X2=7.73 $Y2=1.465
r596 79 81 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.73 $Y=1.63
+ $X2=7.73 $Y2=2.4
r597 75 237 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.715 $Y=1.3
+ $X2=7.715 $Y2=1.465
r598 75 77 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.715 $Y=1.3
+ $X2=7.715 $Y2=0.74
r599 71 236 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.285 $Y=1.3
+ $X2=7.285 $Y2=1.465
r600 71 73 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.285 $Y=1.3
+ $X2=7.285 $Y2=0.74
r601 67 235 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.28 $Y=1.63
+ $X2=7.28 $Y2=1.465
r602 67 69 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.28 $Y=1.63
+ $X2=7.28 $Y2=2.4
r603 63 231 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.83 $Y=1.63
+ $X2=6.83 $Y2=1.465
r604 63 65 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.83 $Y=1.63
+ $X2=6.83 $Y2=2.4
r605 59 230 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.785 $Y=1.3
+ $X2=6.785 $Y2=1.465
r606 59 61 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.785 $Y=1.3
+ $X2=6.785 $Y2=0.74
r607 55 229 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=1.63
+ $X2=6.38 $Y2=1.465
r608 55 57 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.38 $Y=1.63
+ $X2=6.38 $Y2=2.4
r609 51 228 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.355 $Y=1.3
+ $X2=6.355 $Y2=1.465
r610 51 53 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.355 $Y=1.3
+ $X2=6.355 $Y2=0.74
r611 47 224 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.93 $Y=1.63
+ $X2=5.93 $Y2=1.465
r612 47 49 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.93 $Y=1.63
+ $X2=5.93 $Y2=2.4
r613 43 223 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.855 $Y=1.3
+ $X2=5.855 $Y2=1.465
r614 43 45 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.855 $Y=1.3
+ $X2=5.855 $Y2=0.74
r615 39 222 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.48 $Y=1.63
+ $X2=5.48 $Y2=1.465
r616 39 41 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.48 $Y=1.63
+ $X2=5.48 $Y2=2.4
r617 35 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.425 $Y=1.3
+ $X2=5.425 $Y2=1.465
r618 35 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.425 $Y=1.3
+ $X2=5.425 $Y2=0.74
r619 31 217 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.03 $Y=1.63
+ $X2=5.03 $Y2=1.465
r620 31 33 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.03 $Y=1.63
+ $X2=5.03 $Y2=2.4
r621 27 216 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.995 $Y=1.3
+ $X2=4.995 $Y2=1.465
r622 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.995 $Y=1.3
+ $X2=4.995 $Y2=0.74
r623 23 215 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.58 $Y=1.63
+ $X2=4.58 $Y2=1.465
r624 23 25 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.58 $Y=1.63
+ $X2=4.58 $Y2=2.4
r625 19 213 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.3
+ $X2=4.565 $Y2=1.465
r626 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.565 $Y=1.3
+ $X2=4.565 $Y2=0.74
r627 6 183 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=1.84 $X2=3.905 $Y2=2.815
r628 6 181 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=1.84 $X2=3.905 $Y2=1.985
r629 5 169 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.84 $X2=3.005 $Y2=2.815
r630 5 167 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.84 $X2=3.005 $Y2=1.985
r631 4 151 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.105 $Y2=2.815
r632 4 149 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.105 $Y2=1.985
r633 3 177 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.37 $X2=3.85 $Y2=0.515
r634 2 163 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.78
+ $Y=0.37 $X2=2.92 $Y2=0.515
r635 1 155 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.92
+ $Y=0.37 $X2=2.06 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 44 48
+ 52 56 60 66 72 78 82 86 92 98 104 108 110 115 116 118 119 121 122 124 125 127
+ 128 130 131 132 133 134 158 163 168 173 179 182 185 188 191 195
r222 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r223 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r224 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r225 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r226 182 183 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r227 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r228 177 195 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r229 177 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r230 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r231 174 191 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=10.885 $Y=3.33
+ $X2=10.777 $Y2=3.33
r232 174 176 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.885 $Y=3.33
+ $X2=11.28 $Y2=3.33
r233 173 194 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.62 $Y=3.33
+ $X2=11.81 $Y2=3.33
r234 173 176 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.62 $Y=3.33
+ $X2=11.28 $Y2=3.33
r235 172 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r236 172 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r237 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r238 169 188 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=9.955 $Y=3.33
+ $X2=9.837 $Y2=3.33
r239 169 171 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.955 $Y=3.33
+ $X2=10.32 $Y2=3.33
r240 168 191 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=10.67 $Y=3.33
+ $X2=10.777 $Y2=3.33
r241 168 171 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.67 $Y=3.33
+ $X2=10.32 $Y2=3.33
r242 167 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r243 167 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r244 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r245 164 185 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.995 $Y=3.33
+ $X2=8.882 $Y2=3.33
r246 164 166 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.995 $Y=3.33
+ $X2=9.36 $Y2=3.33
r247 163 188 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=9.72 $Y=3.33
+ $X2=9.837 $Y2=3.33
r248 163 166 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.72 $Y=3.33
+ $X2=9.36 $Y2=3.33
r249 162 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r250 162 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r251 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r252 159 182 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=7.955 $Y2=3.33
r253 159 161 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r254 158 185 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=8.77 $Y=3.33
+ $X2=8.882 $Y2=3.33
r255 158 161 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.77 $Y=3.33
+ $X2=8.4 $Y2=3.33
r256 157 183 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r258 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r259 148 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r260 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r261 145 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r262 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r263 142 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r264 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r265 139 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r266 139 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r267 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r268 136 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.735 $Y2=3.33
r269 136 138 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r270 134 157 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r271 134 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r272 134 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r273 132 156 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=6.96 $Y2=3.33
r274 132 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=7.055 $Y2=3.33
r275 130 153 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.07 $Y=3.33 $X2=6
+ $Y2=3.33
r276 130 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=6.155 $Y2=3.33
r277 129 156 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r278 129 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.155 $Y2=3.33
r279 127 150 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.04 $Y2=3.33
r280 127 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.255 $Y2=3.33
r281 126 153 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.34 $Y=3.33
+ $X2=6 $Y2=3.33
r282 126 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=3.33
+ $X2=5.255 $Y2=3.33
r283 124 147 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=3.33
+ $X2=4.08 $Y2=3.33
r284 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=3.33
+ $X2=4.355 $Y2=3.33
r285 123 150 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=5.04 $Y2=3.33
r286 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.355 $Y2=3.33
r287 121 144 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.12 $Y2=3.33
r288 121 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.455 $Y2=3.33
r289 120 147 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=4.08 $Y2=3.33
r290 120 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=3.455 $Y2=3.33
r291 118 141 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.16 $Y2=3.33
r292 118 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.555 $Y2=3.33
r293 117 144 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r294 117 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.555 $Y2=3.33
r295 115 138 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.2 $Y2=3.33
r296 115 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.635 $Y2=3.33
r297 114 141 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r298 114 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.635 $Y2=3.33
r299 110 113 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.745 $Y=1.985
+ $X2=11.745 $Y2=2.815
r300 108 194 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=11.745 $Y=3.245
+ $X2=11.81 $Y2=3.33
r301 108 113 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.745 $Y=3.245
+ $X2=11.745 $Y2=2.815
r302 104 107 39.1295 $w=2.13e-07 $l=7.3e-07 $layer=LI1_cond $X=10.777 $Y=2.085
+ $X2=10.777 $Y2=2.815
r303 102 191 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.777 $Y=3.245
+ $X2=10.777 $Y2=3.33
r304 102 107 23.0489 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=10.777 $Y=3.245
+ $X2=10.777 $Y2=2.815
r305 98 101 35.7993 $w=2.33e-07 $l=7.3e-07 $layer=LI1_cond $X=9.837 $Y=2.085
+ $X2=9.837 $Y2=2.815
r306 96 188 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=9.837 $Y=3.245
+ $X2=9.837 $Y2=3.33
r307 96 101 21.0873 $w=2.33e-07 $l=4.3e-07 $layer=LI1_cond $X=9.837 $Y=3.245
+ $X2=9.837 $Y2=2.815
r308 92 95 37.3904 $w=2.23e-07 $l=7.3e-07 $layer=LI1_cond $X=8.882 $Y=2.085
+ $X2=8.882 $Y2=2.815
r309 90 185 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.882 $Y=3.245
+ $X2=8.882 $Y2=3.33
r310 90 95 22.0245 $w=2.23e-07 $l=4.3e-07 $layer=LI1_cond $X=8.882 $Y=3.245
+ $X2=8.882 $Y2=2.815
r311 86 89 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.955 $Y=2.085
+ $X2=7.955 $Y2=2.815
r312 84 182 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=3.245
+ $X2=7.955 $Y2=3.33
r313 84 89 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.955 $Y=3.245
+ $X2=7.955 $Y2=2.815
r314 83 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=3.33
+ $X2=7.055 $Y2=3.33
r315 82 182 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=3.33
+ $X2=7.955 $Y2=3.33
r316 82 83 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.87 $Y=3.33
+ $X2=7.14 $Y2=3.33
r317 78 81 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.055 $Y=2.085
+ $X2=7.055 $Y2=2.815
r318 76 133 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=3.245
+ $X2=7.055 $Y2=3.33
r319 76 81 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.055 $Y=3.245
+ $X2=7.055 $Y2=2.815
r320 72 75 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.155 $Y=2.085
+ $X2=6.155 $Y2=2.815
r321 70 131 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=3.33
r322 70 75 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=2.815
r323 66 69 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.255 $Y=2.085
+ $X2=5.255 $Y2=2.815
r324 64 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.255 $Y=3.245
+ $X2=5.255 $Y2=3.33
r325 64 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.255 $Y=3.245
+ $X2=5.255 $Y2=2.815
r326 60 63 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.355 $Y=2.085
+ $X2=4.355 $Y2=2.815
r327 58 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=3.245
+ $X2=4.355 $Y2=3.33
r328 58 63 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.355 $Y=3.245
+ $X2=4.355 $Y2=2.815
r329 54 122 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=3.245
+ $X2=3.455 $Y2=3.33
r330 54 56 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.455 $Y=3.245
+ $X2=3.455 $Y2=2.305
r331 50 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=3.245
+ $X2=2.555 $Y2=3.33
r332 50 52 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.555 $Y=3.245
+ $X2=2.555 $Y2=2.305
r333 46 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=3.33
r334 46 48 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=2.455
r335 42 179 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r336 42 44 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.455
r337 13 113 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.705 $Y2=2.815
r338 13 110 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.705 $Y2=1.985
r339 12 107 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.755 $Y2=2.815
r340 12 104 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.755 $Y2=2.085
r341 11 101 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.67
+ $Y=1.84 $X2=9.805 $Y2=2.815
r342 11 98 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=9.67
+ $Y=1.84 $X2=9.805 $Y2=2.085
r343 10 95 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.84 $X2=8.855 $Y2=2.815
r344 10 92 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.84 $X2=8.855 $Y2=2.085
r345 9 89 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.82
+ $Y=1.84 $X2=7.955 $Y2=2.815
r346 9 86 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=7.82
+ $Y=1.84 $X2=7.955 $Y2=2.085
r347 8 81 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.84 $X2=7.055 $Y2=2.815
r348 8 78 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=1.84 $X2=7.055 $Y2=2.085
r349 7 75 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.02
+ $Y=1.84 $X2=6.155 $Y2=2.815
r350 7 72 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=6.02
+ $Y=1.84 $X2=6.155 $Y2=2.085
r351 6 69 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.12
+ $Y=1.84 $X2=5.255 $Y2=2.815
r352 6 66 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=5.12
+ $Y=1.84 $X2=5.255 $Y2=2.085
r353 5 63 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.84 $X2=4.355 $Y2=2.815
r354 5 60 400 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.84 $X2=4.355 $Y2=2.085
r355 4 56 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=3.32
+ $Y=1.84 $X2=3.455 $Y2=2.305
r356 3 52 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=2.42
+ $Y=1.84 $X2=2.555 $Y2=2.305
r357 2 48 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=2.455
r358 1 44 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__BUFINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 55 59 63 67 69 71 75 77 79 83 87 91 95 100 105 110 115 118 121 127 133 139
+ 145 146 151
r254 160 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.355 $Y=2.035
+ $X2=9.355 $Y2=2.035
r255 158 162 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=8.405 $Y=2.035
+ $X2=9.355 $Y2=2.035
r256 156 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.405 $Y=2.035
+ $X2=8.405 $Y2=2.035
r257 151 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.505 $Y=2.035
+ $X2=7.505 $Y2=2.035
r258 151 152 3.7572 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=2.005
+ $X2=7.505 $Y2=1.92
r259 145 148 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=11.255 $Y=2.035
+ $X2=11.255 $Y2=2.815
r260 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.255 $Y=2.035
+ $X2=11.255 $Y2=2.035
r261 140 146 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=10.305 $Y=2.035
+ $X2=11.255 $Y2=2.035
r262 140 162 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=10.305 $Y=2.035
+ $X2=9.355 $Y2=2.035
r263 139 142 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=10.305 $Y=2.035
+ $X2=10.305 $Y2=2.815
r264 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.305 $Y=2.035
+ $X2=10.305 $Y2=2.035
r265 134 154 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=6.605 $Y=2.035
+ $X2=7.505 $Y2=2.035
r266 133 136 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=6.605 $Y=2.035
+ $X2=6.605 $Y2=2.815
r267 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.605 $Y=2.035
+ $X2=6.605 $Y2=2.035
r268 128 134 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=5.705 $Y=2.035
+ $X2=6.605 $Y2=2.035
r269 127 130 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.705 $Y=2.035
+ $X2=5.705 $Y2=2.815
r270 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.705 $Y=2.035
+ $X2=5.705 $Y2=2.035
r271 122 128 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=4.815 $Y=2.035
+ $X2=5.705 $Y2=2.035
r272 121 124 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=4.805 $Y=2.035
+ $X2=4.805 $Y2=2.815
r273 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.815 $Y=2.035
+ $X2=4.815 $Y2=2.035
r274 118 158 0.240602 $w=2.3e-07 $l=3.75e-07 $layer=MET1_cond $X=8.03 $Y=2.035
+ $X2=8.405 $Y2=2.035
r275 118 154 0.336842 $w=2.3e-07 $l=5.25e-07 $layer=MET1_cond $X=8.03 $Y=2.035
+ $X2=7.505 $Y2=2.035
r276 117 145 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.255 $Y=2.02
+ $X2=11.255 $Y2=2.035
r277 115 117 1.23521 $w=3.63e-07 $l=3.5e-08 $layer=LI1_cond $X=11.237 $Y=1.985
+ $X2=11.237 $Y2=2.02
r278 115 116 6.28701 $w=3.63e-07 $l=1.95e-07 $layer=LI1_cond $X=11.237 $Y=1.985
+ $X2=11.237 $Y2=1.79
r279 112 139 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=10.305 $Y=2.02
+ $X2=10.305 $Y2=2.035
r280 110 112 0.501062 $w=3.43e-07 $l=1.5e-08 $layer=LI1_cond $X=10.297 $Y=2.005
+ $X2=10.297 $Y2=2.02
r281 110 111 3.73305 $w=3.43e-07 $l=8.5e-08 $layer=LI1_cond $X=10.297 $Y=2.005
+ $X2=10.297 $Y2=1.92
r282 107 133 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.605 $Y2=2.035
r283 105 107 0.545053 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=6.595 $Y=2.005
+ $X2=6.595 $Y2=2.02
r284 105 106 4.0474 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=2.005
+ $X2=6.595 $Y2=1.92
r285 102 127 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.705 $Y=2.02
+ $X2=5.705 $Y2=2.035
r286 100 102 0.581203 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.69 $Y=2.005
+ $X2=5.69 $Y2=2.02
r287 100 101 4.57587 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=5.69 $Y=2.005
+ $X2=5.69 $Y2=1.92
r288 97 121 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.805 $Y=2.02
+ $X2=4.805 $Y2=2.035
r289 95 97 0.561516 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=4.792 $Y=2.005
+ $X2=4.792 $Y2=2.02
r290 95 96 3.78181 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.792 $Y=2.005
+ $X2=4.792 $Y2=1.92
r291 91 116 44.5262 $w=3.28e-07 $l=1.275e-06 $layer=LI1_cond $X=11.22 $Y=0.515
+ $X2=11.22 $Y2=1.79
r292 87 111 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=10.25 $Y=0.515
+ $X2=10.25 $Y2=1.92
r293 81 160 3.13751 $w=3.28e-07 $l=8.06226e-08 $layer=LI1_cond $X=9.32 $Y=1.92
+ $X2=9.355 $Y2=1.985
r294 81 83 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=9.32 $Y=1.92
+ $X2=9.32 $Y2=0.515
r295 77 160 7.39394 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=9.355 $Y=2.185
+ $X2=9.355 $Y2=1.985
r296 77 79 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=9.355 $Y=2.185
+ $X2=9.355 $Y2=2.815
r297 73 156 3.09497 $w=3.2e-07 $l=7.2111e-08 $layer=LI1_cond $X=8.39 $Y=1.92
+ $X2=8.405 $Y2=1.985
r298 73 75 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=8.39 $Y=1.92
+ $X2=8.39 $Y2=0.515
r299 69 156 7.39394 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=8.405 $Y=2.185
+ $X2=8.405 $Y2=1.985
r300 69 71 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=8.405 $Y=2.185
+ $X2=8.405 $Y2=2.815
r301 65 151 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.505 $Y=2.085
+ $X2=7.505 $Y2=2.005
r302 65 67 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.505 $Y=2.085
+ $X2=7.505 $Y2=2.815
r303 63 152 66.0891 $w=2.43e-07 $l=1.405e-06 $layer=LI1_cond $X=7.462 $Y=0.515
+ $X2=7.462 $Y2=1.92
r304 59 106 68.9014 $w=2.33e-07 $l=1.405e-06 $layer=LI1_cond $X=6.537 $Y=0.515
+ $X2=6.537 $Y2=1.92
r305 55 101 75.3108 $w=2.13e-07 $l=1.405e-06 $layer=LI1_cond $X=5.617 $Y=0.515
+ $X2=5.617 $Y2=1.92
r306 51 96 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=4.74 $Y=0.515
+ $X2=4.74 $Y2=1.92
r307 16 148 400 $w=1.7e-07 $l=1.05889e-06 $layer=licon1_PDIFF $count=1 $X=11.08
+ $Y=1.84 $X2=11.255 $Y2=2.815
r308 16 115 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.08
+ $Y=1.84 $X2=11.255 $Y2=1.985
r309 15 142 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=2.815
r310 15 110 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=2.005
r311 14 160 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.84 $X2=9.355 $Y2=1.985
r312 14 79 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.22
+ $Y=1.84 $X2=9.355 $Y2=2.815
r313 13 156 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.84 $X2=8.405 $Y2=1.985
r314 13 71 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.84 $X2=8.405 $Y2=2.815
r315 12 151 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=1.84 $X2=7.505 $Y2=2.005
r316 12 67 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=1.84 $X2=7.505 $Y2=2.815
r317 11 136 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.47
+ $Y=1.84 $X2=6.605 $Y2=2.815
r318 11 105 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=6.47
+ $Y=1.84 $X2=6.605 $Y2=2.005
r319 10 130 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.84 $X2=5.705 $Y2=2.815
r320 10 100 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.84 $X2=5.705 $Y2=2.005
r321 9 124 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.84 $X2=4.805 $Y2=2.815
r322 9 95 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.84 $X2=4.805 $Y2=2.005
r323 8 91 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.08
+ $Y=0.37 $X2=11.22 $Y2=0.515
r324 7 87 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.15
+ $Y=0.37 $X2=10.29 $Y2=0.515
r325 6 83 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.22
+ $Y=0.37 $X2=9.36 $Y2=0.515
r326 5 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.29
+ $Y=0.37 $X2=8.43 $Y2=0.515
r327 4 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.36
+ $Y=0.37 $X2=7.5 $Y2=0.515
r328 3 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.43
+ $Y=0.37 $X2=6.57 $Y2=0.515
r329 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.5
+ $Y=0.37 $X2=5.64 $Y2=0.515
r330 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.64
+ $Y=0.37 $X2=4.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFINV_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 42 46
+ 50 54 58 62 66 70 74 78 82 86 88 90 93 94 96 97 99 100 102 103 104 106 111 129
+ 133 138 143 148 153 158 164 167 170 173 176 179 182 185 189
r214 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r215 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r216 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r217 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r218 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r219 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r220 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r221 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r222 162 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r223 162 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r224 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r225 159 185 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.885 $Y=0
+ $X2=10.72 $Y2=0
r226 159 161 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.885 $Y=0
+ $X2=11.28 $Y2=0
r227 158 188 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.555 $Y=0
+ $X2=11.777 $Y2=0
r228 158 161 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.555 $Y=0
+ $X2=11.28 $Y2=0
r229 157 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r230 157 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r231 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r232 154 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.955 $Y=0
+ $X2=9.79 $Y2=0
r233 154 156 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.955 $Y=0
+ $X2=10.32 $Y2=0
r234 153 185 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.555 $Y=0
+ $X2=10.72 $Y2=0
r235 153 156 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=10.555 $Y=0
+ $X2=10.32 $Y2=0
r236 152 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r237 152 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r238 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r239 149 179 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=8.86 $Y2=0
r240 149 151 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=9.36 $Y2=0
r241 148 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.625 $Y=0
+ $X2=9.79 $Y2=0
r242 148 151 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.625 $Y=0
+ $X2=9.36 $Y2=0
r243 147 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r244 147 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r245 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r246 144 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=0
+ $X2=7.93 $Y2=0
r247 144 146 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.095 $Y=0
+ $X2=8.4 $Y2=0
r248 143 179 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=0
+ $X2=8.86 $Y2=0
r249 143 146 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.695 $Y=0
+ $X2=8.4 $Y2=0
r250 142 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r251 142 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r252 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r253 139 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=0 $X2=7
+ $Y2=0
r254 139 141 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=7.44 $Y2=0
r255 138 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.93 $Y2=0
r256 138 141 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.44 $Y2=0
r257 137 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r258 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r259 134 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=0
+ $X2=6.07 $Y2=0
r260 134 136 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.235 $Y=0
+ $X2=6.48 $Y2=0
r261 133 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=0 $X2=7
+ $Y2=0
r262 133 136 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=0
+ $X2=6.48 $Y2=0
r263 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r264 129 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.07 $Y2=0
r265 129 131 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=5.52 $Y2=0
r266 128 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r267 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r268 125 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r269 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r270 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r271 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r272 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.12 $Y2=0
r273 119 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r274 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r275 116 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=1.63 $Y2=0
r276 116 118 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=2.16 $Y2=0
r277 115 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=1.68 $Y2=0
r278 115 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=0.72 $Y2=0
r279 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r280 112 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r281 112 114 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=1.2 $Y2=0
r282 111 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.63 $Y2=0
r283 111 114 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.2 $Y2=0
r284 109 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r285 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r286 106 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r287 106 108 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r288 104 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r289 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r290 104 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r291 102 127 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.04 $Y2=0
r292 102 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.17 $Y2=0
r293 101 131 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.52 $Y2=0
r294 101 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.17 $Y2=0
r295 99 124 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=4.08 $Y2=0
r296 99 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=4.28 $Y2=0
r297 98 127 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.445 $Y=0
+ $X2=5.04 $Y2=0
r298 98 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0
+ $X2=4.28 $Y2=0
r299 96 121 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.12 $Y2=0
r300 96 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.35
+ $Y2=0
r301 95 124 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=4.08 $Y2=0
r302 95 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.35
+ $Y2=0
r303 93 118 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.16 $Y2=0
r304 93 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.45
+ $Y2=0
r305 92 121 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.575 $Y=0
+ $X2=3.12 $Y2=0
r306 92 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.45
+ $Y2=0
r307 88 188 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.72 $Y=0.085
+ $X2=11.777 $Y2=0
r308 88 90 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.72 $Y=0.085
+ $X2=11.72 $Y2=0.515
r309 84 185 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.72 $Y=0.085
+ $X2=10.72 $Y2=0
r310 84 86 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.72 $Y=0.085
+ $X2=10.72 $Y2=0.515
r311 80 182 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=0.085
+ $X2=9.79 $Y2=0
r312 80 82 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.79 $Y=0.085
+ $X2=9.79 $Y2=0.515
r313 76 179 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=0.085
+ $X2=8.86 $Y2=0
r314 76 78 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.86 $Y=0.085
+ $X2=8.86 $Y2=0.515
r315 72 176 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r316 72 74 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.515
r317 68 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.085 $X2=7
+ $Y2=0
r318 68 70 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7 $Y=0.085 $X2=7
+ $Y2=0.515
r319 64 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0
r320 64 66 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0.515
r321 60 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.085
+ $X2=5.17 $Y2=0
r322 60 62 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.17 $Y=0.085
+ $X2=5.17 $Y2=0.515
r323 56 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0
r324 56 58 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0.515
r325 52 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r326 52 54 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.625
r327 48 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0
r328 48 50 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.625
r329 44 167 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0
r330 44 46 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0.675
r331 40 164 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r332 40 42 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.675
r333 13 90 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=11.51
+ $Y=0.37 $X2=11.72 $Y2=0.515
r334 12 86 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.58
+ $Y=0.37 $X2=10.72 $Y2=0.515
r335 11 82 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.65
+ $Y=0.37 $X2=9.79 $Y2=0.515
r336 10 78 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.37 $X2=8.86 $Y2=0.515
r337 9 74 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
r338 8 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.86
+ $Y=0.37 $X2=7 $Y2=0.515
r339 7 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.93
+ $Y=0.37 $X2=6.07 $Y2=0.515
r340 6 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.07
+ $Y=0.37 $X2=5.21 $Y2=0.515
r341 5 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
r342 4 54 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.37 $X2=3.35 $Y2=0.625
r343 3 50 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.37 $X2=2.49 $Y2=0.625
r344 2 46 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.37 $X2=1.63 $Y2=0.675
r345 1 42 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4_4 A B C D VGND VNB VPB VPWR X
M1000 a_83_264# D a_965_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=5.9e+11p ps=5.18e+06u
M1001 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=2.2402e+12p pd=1.413e+07u as=6.549e+11p ps=4.73e+06u
M1002 a_965_392# D a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_499_392# C a_965_392# VPB pshort w=1e+06u l=180000u
+  ad=9.3e+11p pd=7.86e+06u as=0p ps=0u
M1004 a_83_264# B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1005 X a_83_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=1.1996e+12p ps=1.092e+07u
M1006 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_264# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND D a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_591_392# B a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1015 a_83_264# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_591_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_591_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_499_392# B a_591_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_965_392# C a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

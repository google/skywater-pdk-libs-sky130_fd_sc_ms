* File: sky130_fd_sc_ms__o2bb2ai_2.spice
* Created: Wed Sep  2 12:24:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2bb2ai_2.pex.spice"
.subckt sky130_fd_sc_ms__o2bb2ai_2  VNB VPB A1_N A2_N B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1007 N_A_134_74#_M1007_d N_A1_N_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_136_387#_M1008_d N_A2_N_M1008_g N_A_134_74#_M1007_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1136 AS=0.0896 PD=0.995 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_136_387#_M1008_d N_A2_N_M1019_g N_A_134_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1136 AS=0.0896 PD=0.995 PS=0.92 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1012 N_A_134_74#_M1019_s N_A1_N_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_Y_M1000_d N_A_136_387#_M1000_g N_A_518_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1000_d N_A_136_387#_M1006_g N_A_518_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1147 PD=1.02 PS=1.05 NRD=0 NRS=4.86 M=1 R=4.93333
+ SA=75000.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1010 N_A_518_74#_M1006_s N_B1_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1010_s N_B2_M1002_g N_A_518_74#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1221 PD=1.09 PS=1.07 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75001.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_B2_M1015_g N_A_518_74#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1221 PD=1.035 PS=1.07 NRD=0.804 NRS=4.044 M=1 R=4.93333
+ SA=75002.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1017 N_A_518_74#_M1017_d N_B1_M1017_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.10915 PD=2.05 PS=1.035 NRD=0 NRS=1.62 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_136_387#_M1001_d N_A1_N_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.3675 PD=1.11 PS=2.83 NRD=0 NRS=89.6941 M=1 R=4.66667
+ SA=90000.3 SB=90004.4 A=0.1512 P=2.04 MULT=1
MM1003 N_VPWR_M1003_d N_A2_N_M1003_g N_A_136_387#_M1001_d VPB PSHORT L=0.18
+ W=0.84 AD=0.220325 AS=0.1134 PD=1.525 PS=1.11 NRD=48.5999 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90004 A=0.1512 P=2.04 MULT=1
MM1018 N_VPWR_M1003_d N_A2_N_M1018_g N_A_136_387#_M1018_s VPB PSHORT L=0.18
+ W=0.84 AD=0.220325 AS=0.159712 PD=1.525 PS=1.3 NRD=48.5999 NRS=1.1623 M=1
+ R=4.66667 SA=90001.3 SB=90003.4 A=0.1512 P=2.04 MULT=1
MM1014 N_A_136_387#_M1018_s N_A1_N_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18
+ W=0.84 AD=0.159712 AS=0.2196 PD=1.3 PS=1.40143 NRD=18.7544 NRS=55.1009 M=1
+ R=4.66667 SA=90001.7 SB=90003.2 A=0.1512 P=2.04 MULT=1
MM1011 N_Y_M1011_d N_A_136_387#_M1011_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.2928 PD=1.405 PS=1.86857 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.8
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1016 N_Y_M1011_d N_A_136_387#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.2016 PD=1.405 PS=1.48 NRD=1.7533 NRS=5.2599 M=1 R=6.22222
+ SA=90002.3 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1004 N_A_799_368#_M1004_d N_B1_M1004_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90002.8
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_799_368#_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1005_d N_B2_M1009_g N_A_799_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1013 N_A_799_368#_M1009_s N_B1_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
c_59 VNB 0 1.39855e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__o2bb2ai_2.pxi.spice"
*
.ends
*
*

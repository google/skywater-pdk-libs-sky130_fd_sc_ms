* File: sky130_fd_sc_ms__a41oi_1.pxi.spice
* Created: Fri Aug 28 17:09:51 2020
* 
x_PM_SKY130_FD_SC_MS__A41OI_1%B1 N_B1_M1003_g N_B1_M1007_g B1 N_B1_c_55_n
+ N_B1_c_56_n PM_SKY130_FD_SC_MS__A41OI_1%B1
x_PM_SKY130_FD_SC_MS__A41OI_1%A4 N_A4_M1002_g N_A4_M1005_g A4 N_A4_c_80_n
+ N_A4_c_81_n PM_SKY130_FD_SC_MS__A41OI_1%A4
x_PM_SKY130_FD_SC_MS__A41OI_1%A3 N_A3_M1006_g N_A3_M1009_g A3 N_A3_c_118_n
+ N_A3_c_119_n PM_SKY130_FD_SC_MS__A41OI_1%A3
x_PM_SKY130_FD_SC_MS__A41OI_1%A2 N_A2_M1008_g N_A2_M1000_g A2 N_A2_c_154_n
+ PM_SKY130_FD_SC_MS__A41OI_1%A2
x_PM_SKY130_FD_SC_MS__A41OI_1%A1 N_A1_M1001_g N_A1_M1004_g A1 N_A1_c_189_n
+ N_A1_c_190_n PM_SKY130_FD_SC_MS__A41OI_1%A1
x_PM_SKY130_FD_SC_MS__A41OI_1%Y N_Y_M1007_s N_Y_M1001_d N_Y_M1003_s N_Y_c_214_n
+ N_Y_c_219_n N_Y_c_215_n N_Y_c_216_n N_Y_c_217_n N_Y_c_220_n Y
+ PM_SKY130_FD_SC_MS__A41OI_1%Y
x_PM_SKY130_FD_SC_MS__A41OI_1%A_119_368# N_A_119_368#_M1003_d
+ N_A_119_368#_M1009_d N_A_119_368#_M1004_d N_A_119_368#_c_272_n
+ N_A_119_368#_c_274_n N_A_119_368#_c_268_n N_A_119_368#_c_269_n
+ N_A_119_368#_c_270_n PM_SKY130_FD_SC_MS__A41OI_1%A_119_368#
x_PM_SKY130_FD_SC_MS__A41OI_1%VPWR N_VPWR_M1002_d N_VPWR_M1000_d N_VPWR_c_308_n
+ VPWR N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_307_n
+ N_VPWR_c_313_n N_VPWR_c_314_n PM_SKY130_FD_SC_MS__A41OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A41OI_1%VGND N_VGND_M1007_d VGND N_VGND_c_344_n
+ N_VGND_c_345_n N_VGND_c_346_n PM_SKY130_FD_SC_MS__A41OI_1%VGND
cc_1 VNB N_B1_M1003_g 0.001973f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_B1_M1007_g 0.0333332f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_B1_c_55_n 0.00430714f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_B1_c_56_n 0.0604259f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_5 VNB N_A4_M1005_g 0.0271041f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_A4_c_80_n 0.00234054f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_7 VNB N_A4_c_81_n 0.0365182f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_8 VNB N_A3_M1006_g 0.0260165f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_9 VNB N_A3_c_118_n 0.0250766f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_A3_c_119_n 0.00452292f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_11 VNB N_A2_M1008_g 0.0284012f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB A2 0.00682758f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A2_c_154_n 0.0225947f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_14 VNB N_A1_M1001_g 0.031841f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_15 VNB N_A1_M1004_g 0.00188935f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_A1_c_189_n 0.0594419f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_17 VNB N_A1_c_190_n 0.0051843f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_18 VNB N_Y_c_214_n 0.0258829f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_19 VNB N_Y_c_215_n 0.0345375f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_20 VNB N_Y_c_216_n 0.0102107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_217_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.0120831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_307_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_344_n 0.0412642f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_VGND_c_345_n 0.0662801f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_26 VNB N_VGND_c_346_n 0.240368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_B1_M1003_g 0.0304184f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_28 VPB N_B1_c_55_n 0.00761464f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_29 VPB N_A4_M1002_g 0.0252853f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_30 VPB N_A4_c_80_n 0.00304716f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_31 VPB N_A4_c_81_n 0.0100288f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_32 VPB N_A3_M1009_g 0.0234408f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_33 VPB N_A3_c_118_n 0.00554261f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_34 VPB N_A3_c_119_n 0.003565f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_35 VPB N_A2_M1000_g 0.0224065f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_36 VPB A2 0.00526504f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_37 VPB N_A2_c_154_n 0.00545222f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_38 VPB N_A1_M1004_g 0.0309152f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_39 VPB N_A1_c_190_n 0.00761845f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_40 VPB N_Y_c_219_n 0.0353375f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_41 VPB N_Y_c_220_n 0.00719835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB Y 0.00351957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_119_368#_c_268_n 0.0142315f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_44 VPB N_A_119_368#_c_269_n 0.0288011f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_45 VPB N_A_119_368#_c_270_n 0.00275743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_308_n 0.00911553f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_47 VPB N_VPWR_c_309_n 0.0325002f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_48 VPB N_VPWR_c_310_n 0.0195071f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_49 VPB N_VPWR_c_311_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_307_n 0.0664811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_313_n 0.02216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_314_n 0.00651392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 N_B1_M1003_g N_A4_M1002_g 0.0170275f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_54 N_B1_M1007_g N_A4_M1005_g 0.0105574f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_55 N_B1_c_56_n N_A4_M1005_g 5.70607e-19 $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_56 N_B1_c_56_n N_A4_c_81_n 0.0170275f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_57 N_B1_M1007_g N_Y_c_214_n 0.0175621f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_58 N_B1_M1003_g N_Y_c_219_n 0.0123623f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_59 N_B1_M1007_g N_Y_c_216_n 0.0179726f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_60 N_B1_c_55_n N_Y_c_216_n 0.0247471f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_61 N_B1_c_56_n N_Y_c_216_n 0.00318727f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_62 N_B1_M1003_g N_Y_c_220_n 0.0186536f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_63 N_B1_c_55_n N_Y_c_220_n 0.0235439f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_64 N_B1_c_56_n N_Y_c_220_n 0.00136987f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_65 N_B1_M1007_g Y 0.00516025f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_66 N_B1_c_55_n Y 0.0368805f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_67 N_B1_c_56_n Y 0.00710565f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_68 N_B1_M1003_g N_A_119_368#_c_270_n 4.37331e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_69 N_B1_M1003_g N_VPWR_c_309_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_70 N_B1_M1003_g N_VPWR_c_307_n 0.00987672f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_71 N_B1_M1007_g N_VGND_c_344_n 0.00847491f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_72 N_B1_M1007_g N_VGND_c_346_n 0.00826401f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_73 N_A4_M1005_g N_A3_M1006_g 0.0399236f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A4_M1002_g N_A3_M1009_g 0.0133163f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_75 N_A4_c_80_n N_A3_M1009_g 3.01966e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A4_c_80_n N_A3_c_118_n 3.50935e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A4_c_81_n N_A3_c_118_n 0.0399236f $X=1.31 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A4_M1002_g N_A3_c_119_n 2.81338e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A4_c_80_n N_A3_c_119_n 0.0279517f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A4_c_81_n N_A3_c_119_n 0.00235304f $X=1.31 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A4_M1002_g N_Y_c_219_n 4.66361e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_82 N_A4_M1005_g N_Y_c_215_n 0.0171807f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A4_c_80_n N_Y_c_215_n 0.0204317f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A4_c_81_n N_Y_c_215_n 0.00510052f $X=1.31 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A4_M1002_g N_Y_c_220_n 0.00172065f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A4_M1005_g Y 0.00420733f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A4_c_80_n Y 0.0330364f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A4_c_81_n Y 0.00788563f $X=1.31 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A4_c_80_n N_A_119_368#_c_272_n 0.00491597f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_90 N_A4_c_81_n N_A_119_368#_c_272_n 0.00237233f $X=1.31 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A4_M1002_g N_A_119_368#_c_274_n 0.0180822f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A4_c_80_n N_A_119_368#_c_274_n 0.0156111f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_93 N_A4_c_81_n N_A_119_368#_c_274_n 9.02288e-19 $X=1.31 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A4_M1002_g N_A_119_368#_c_270_n 0.0085296f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A4_M1002_g N_VPWR_c_309_n 0.005209f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A4_M1002_g N_VPWR_c_307_n 0.00984912f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A4_M1002_g N_VPWR_c_313_n 0.00594853f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A4_M1005_g N_VGND_c_344_n 0.0118628f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A4_M1005_g N_VGND_c_345_n 0.00384553f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A4_M1005_g N_VGND_c_346_n 0.0075725f $X=1.31 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A3_M1006_g N_A2_M1008_g 0.0373965f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A3_M1009_g N_A2_M1000_g 0.0483083f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A3_c_119_n N_A2_M1000_g 3.75669e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A3_M1009_g A2 3.94809e-19 $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A3_c_118_n A2 0.00121024f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A3_c_119_n A2 0.0266982f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A3_c_118_n N_A2_c_154_n 0.017626f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A3_c_119_n N_A2_c_154_n 4.19879e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A3_M1006_g N_Y_c_215_n 0.0157189f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A3_c_118_n N_Y_c_215_n 0.00118184f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A3_c_119_n N_Y_c_215_n 0.024303f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A3_M1009_g N_A_119_368#_c_272_n 0.0225404f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A3_c_118_n N_A_119_368#_c_272_n 6.18717e-19 $X=1.79 $Y=1.515 $X2=0
+ $Y2=0
cc_114 N_A3_c_119_n N_A_119_368#_c_272_n 0.0282494f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A3_M1009_g N_A_119_368#_c_274_n 0.00362263f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A3_M1009_g N_VPWR_c_310_n 0.00460063f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A3_M1009_g N_VPWR_c_307_n 0.00904028f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A3_M1009_g N_VPWR_c_313_n 0.0181977f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A3_M1006_g N_VGND_c_344_n 0.00217763f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A3_M1006_g N_VGND_c_345_n 0.00461464f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A3_M1006_g N_VGND_c_346_n 0.0091028f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A2_M1008_g N_A1_M1001_g 0.0342424f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A2_M1000_g N_A1_M1004_g 0.0305753f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_124 A2 N_A1_c_189_n 0.00402425f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_c_154_n N_A1_c_189_n 0.0174186f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A2_M1008_g N_A1_c_190_n 2.13129e-19 $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_127 A2 N_A1_c_190_n 0.0354768f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A2_c_154_n N_A1_c_190_n 2.22391e-19 $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A2_M1008_g N_Y_c_215_n 0.0166695f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_130 A2 N_Y_c_215_n 0.0358367f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A2_c_154_n N_Y_c_215_n 0.004053f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A2_M1008_g N_Y_c_217_n 0.00278148f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_M1000_g N_A_119_368#_c_272_n 0.0218071f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_134 A2 N_A_119_368#_c_272_n 0.0409631f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A2_c_154_n N_A_119_368#_c_272_n 6.86384e-19 $X=2.36 $Y=1.515 $X2=0
+ $Y2=0
cc_136 N_A2_M1000_g N_A_119_368#_c_269_n 8.08672e-19 $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A2_M1000_g N_VPWR_c_308_n 0.00298851f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A2_M1000_g N_VPWR_c_310_n 0.00553757f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A2_M1000_g N_VPWR_c_307_n 0.0108916f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A2_M1000_g N_VPWR_c_313_n 0.00187567f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A2_M1008_g N_VGND_c_345_n 0.00461464f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A2_M1008_g N_VGND_c_346_n 0.00911823f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1001_g N_Y_c_215_n 0.0176533f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_c_189_n N_Y_c_215_n 0.00285738f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_145 N_A1_c_190_n N_Y_c_215_n 0.025569f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_146 N_A1_M1001_g N_Y_c_217_n 0.0142362f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A1_M1004_g N_A_119_368#_c_272_n 0.0240294f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_A_119_368#_c_268_n 0.00173708f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A1_c_189_n N_A_119_368#_c_268_n 0.00152648f $X=3.09 $Y=1.465 $X2=0
+ $Y2=0
cc_150 N_A1_c_190_n N_A_119_368#_c_268_n 0.0258519f $X=3.09 $Y=1.465 $X2=0 $Y2=0
cc_151 N_A1_M1004_g N_A_119_368#_c_269_n 0.0101825f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A1_M1004_g N_VPWR_c_308_n 0.00433115f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A1_M1004_g N_VPWR_c_311_n 0.005209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A1_M1004_g N_VPWR_c_307_n 0.00986397f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A1_M1001_g N_VGND_c_345_n 0.00434272f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A1_M1001_g N_VGND_c_346_n 0.00826262f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_157 N_Y_c_220_n N_A_119_368#_M1003_d 0.00471875f $X=0.72 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_158 Y N_A_119_368#_M1003_d 0.00211162f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_159 N_Y_c_220_n N_A_119_368#_c_274_n 0.0148699f $X=0.72 $Y=1.95 $X2=0 $Y2=0
cc_160 N_Y_c_219_n N_A_119_368#_c_270_n 0.0203021f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_161 N_Y_c_219_n N_VPWR_c_309_n 0.014549f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_162 N_Y_c_219_n N_VPWR_c_307_n 0.0119743f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_163 N_Y_c_215_n N_VGND_M1007_d 0.00637083f $X=2.89 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_164 N_Y_c_216_n N_VGND_M1007_d 0.0034772f $X=0.835 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_165 N_Y_c_214_n N_VGND_c_344_n 0.0277067f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_166 N_Y_c_216_n N_VGND_c_344_n 0.0321701f $X=0.835 $Y=1.045 $X2=0 $Y2=0
cc_167 N_Y_c_217_n N_VGND_c_345_n 0.0145639f $X=3.055 $Y=0.515 $X2=0 $Y2=0
cc_168 N_Y_c_214_n N_VGND_c_346_n 0.0119539f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_169 N_Y_c_217_n N_VGND_c_346_n 0.0119984f $X=3.055 $Y=0.515 $X2=0 $Y2=0
cc_170 N_Y_c_215_n A_277_74# 0.0048076f $X=2.89 $Y=1.045 $X2=-0.19 $Y2=-0.245
cc_171 N_Y_c_215_n A_355_74# 0.0121704f $X=2.89 $Y=1.045 $X2=-0.19 $Y2=-0.245
cc_172 N_Y_c_215_n A_469_74# 0.0121704f $X=2.89 $Y=1.045 $X2=-0.19 $Y2=-0.245
cc_173 N_A_119_368#_c_272_n N_VPWR_M1002_d 0.0208909f $X=2.915 $Y=2.12 $X2=-0.19
+ $Y2=1.66
cc_174 N_A_119_368#_c_274_n N_VPWR_M1002_d 0.00649923f $X=1.275 $Y=2.12
+ $X2=-0.19 $Y2=1.66
cc_175 N_A_119_368#_c_272_n N_VPWR_M1000_d 0.00599175f $X=2.915 $Y=2.12 $X2=0
+ $Y2=0
cc_176 N_A_119_368#_c_272_n N_VPWR_c_308_n 0.0227014f $X=2.915 $Y=2.12 $X2=0
+ $Y2=0
cc_177 N_A_119_368#_c_269_n N_VPWR_c_308_n 0.0203057f $X=3.08 $Y=2.815 $X2=0
+ $Y2=0
cc_178 N_A_119_368#_c_270_n N_VPWR_c_309_n 0.0145644f $X=0.78 $Y=2.375 $X2=0
+ $Y2=0
cc_179 N_A_119_368#_c_269_n N_VPWR_c_311_n 0.014549f $X=3.08 $Y=2.815 $X2=0
+ $Y2=0
cc_180 N_A_119_368#_c_269_n N_VPWR_c_307_n 0.0119743f $X=3.08 $Y=2.815 $X2=0
+ $Y2=0
cc_181 N_A_119_368#_c_270_n N_VPWR_c_307_n 0.0119803f $X=0.78 $Y=2.375 $X2=0
+ $Y2=0
cc_182 N_A_119_368#_c_272_n N_VPWR_c_313_n 0.0326655f $X=2.915 $Y=2.12 $X2=0
+ $Y2=0
cc_183 N_A_119_368#_c_274_n N_VPWR_c_313_n 0.0108583f $X=1.275 $Y=2.12 $X2=0
+ $Y2=0
cc_184 N_A_119_368#_c_270_n N_VPWR_c_313_n 0.0197993f $X=0.78 $Y=2.375 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__a221o_2.spice
* Created: Wed Sep  2 11:52:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a221o_2.pex.spice"
.subckt sky130_fd_sc_ms__a221o_2  VNB VPB A2 A1 B1 B2 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 N_X_M1002_d N_A_89_260#_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1003 N_X_M1002_d N_A_89_260#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.17575 PD=1.02 PS=1.215 NRD=0 NRS=15.396 M=1 R=4.93333
+ SA=75000.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1007 A_337_74# N_A2_M1007_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.17575 PD=0.95 PS=1.215 NRD=8.1 NRS=16.212 M=1 R=4.93333 SA=75001.2
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1001 N_A_89_260#_M1001_d N_A1_M1001_g A_337_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.3034 AS=0.0777 PD=1.56 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1008 A_603_74# N_B1_M1008_g N_A_89_260#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.3034 PD=0.95 PS=1.56 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_B2_M1009_g A_603_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0777 PD=1.13 PS=0.95 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002.9 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1010 N_A_89_260#_M1010_d N_C1_M1010_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75003.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1011_d N_A_89_260#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1011_d N_A_89_260#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.193464 PD=1.39 PS=1.53736 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001 A=0.2016 P=2.6 MULT=1
MM1013 N_A_319_392#_M1013_d N_A2_M1013_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.172736 PD=1.27 PS=1.37264 NRD=0 NRS=11.8003 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_319_392#_M1013_d VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_319_392#_M1004_d N_B1_M1004_g N_A_515_392#_M1004_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_A_515_392#_M1005_d N_B2_M1005_g N_A_319_392#_M1004_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_A_89_260#_M1006_d N_C1_M1006_g N_A_515_392#_M1005_d VPB PSHORT L=0.18
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__a221o_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a22oi_4.pex.spice
* Created: Fri Aug 28 17:03:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A22OI_4%B2 1 3 6 10 14 18 22 26 30 32 33 34 49 50
c81 49 0 1.11174e-19 $X=1.79 $Y=1.515
c82 26 0 8.01953e-20 $X=1.87 $Y=0.74
r83 48 50 11.4762 $w=3.36e-07 $l=8e-08 $layer=POLY_cond $X=1.79 $Y=1.56 $X2=1.87
+ $Y2=1.56
r84 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=1.515 $X2=1.79 $Y2=1.515
r85 41 43 34.4286 $w=3.36e-07 $l=2.4e-07 $layer=POLY_cond $X=0.77 $Y=1.56
+ $X2=1.01 $Y2=1.56
r86 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.77
+ $Y=1.515 $X2=0.77 $Y2=1.515
r87 39 41 27.256 $w=3.36e-07 $l=1.9e-07 $layer=POLY_cond $X=0.58 $Y=1.56
+ $X2=0.77 $Y2=1.56
r88 38 39 0.717262 $w=3.36e-07 $l=5e-09 $layer=POLY_cond $X=0.575 $Y=1.56
+ $X2=0.58 $Y2=1.56
r89 34 49 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.79 $Y2=1.565
r90 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r91 33 42 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.77 $Y2=1.565
r92 32 42 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.77
+ $Y2=1.565
r93 28 50 7.88988 $w=3.36e-07 $l=5.5e-08 $layer=POLY_cond $X=1.925 $Y=1.56
+ $X2=1.87 $Y2=1.56
r94 28 30 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.925 $Y=1.68
+ $X2=1.925 $Y2=2.4
r95 24 50 21.6522 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.56
r96 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.74
r97 20 48 45.1875 $w=3.36e-07 $l=3.15e-07 $layer=POLY_cond $X=1.475 $Y=1.56
+ $X2=1.79 $Y2=1.56
r98 20 45 5.02083 $w=3.36e-07 $l=3.5e-08 $layer=POLY_cond $X=1.475 $Y=1.56
+ $X2=1.44 $Y2=1.56
r99 20 22 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.475 $Y=1.68
+ $X2=1.475 $Y2=2.4
r100 16 45 21.6522 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.44 $Y=1.35
+ $X2=1.44 $Y2=1.56
r101 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.44 $Y=1.35
+ $X2=1.44 $Y2=0.74
r102 12 45 59.5327 $w=3.36e-07 $l=4.15e-07 $layer=POLY_cond $X=1.025 $Y=1.56
+ $X2=1.44 $Y2=1.56
r103 12 43 2.15179 $w=3.36e-07 $l=1.5e-08 $layer=POLY_cond $X=1.025 $Y=1.56
+ $X2=1.01 $Y2=1.56
r104 12 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.025 $Y=1.68
+ $X2=1.025 $Y2=2.4
r105 8 43 21.6522 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.01 $Y=1.35
+ $X2=1.01 $Y2=1.56
r106 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.01 $Y=1.35
+ $X2=1.01 $Y2=0.74
r107 4 39 21.6522 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.58 $Y=1.35
+ $X2=0.58 $Y2=1.56
r108 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.58 $Y=1.35 $X2=0.58
+ $Y2=0.74
r109 1 38 17.3521 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.575 $Y=1.77
+ $X2=0.575 $Y2=1.56
r110 1 3 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.575 $Y=1.77 $X2=0.575
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%B1 3 7 11 15 19 23 27 31 33 34 49
c93 7 0 1.11174e-19 $X=2.375 $Y=2.4
c94 3 0 1.9142e-19 $X=2.3 $Y=0.74
r95 49 50 18.3814 $w=3.54e-07 $l=1.35e-07 $layer=POLY_cond $X=3.59 $Y=1.5
+ $X2=3.725 $Y2=1.5
r96 48 49 42.8898 $w=3.54e-07 $l=3.15e-07 $layer=POLY_cond $X=3.275 $Y=1.5
+ $X2=3.59 $Y2=1.5
r97 47 48 15.6582 $w=3.54e-07 $l=1.15e-07 $layer=POLY_cond $X=3.16 $Y=1.5
+ $X2=3.275 $Y2=1.5
r98 45 47 6.80791 $w=3.54e-07 $l=5e-08 $layer=POLY_cond $X=3.11 $Y=1.5 $X2=3.16
+ $Y2=1.5
r99 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.515 $X2=3.11 $Y2=1.515
r100 43 45 38.8051 $w=3.54e-07 $l=2.85e-07 $layer=POLY_cond $X=2.825 $Y=1.5
+ $X2=3.11 $Y2=1.5
r101 42 43 12.935 $w=3.54e-07 $l=9.5e-08 $layer=POLY_cond $X=2.73 $Y=1.5
+ $X2=2.825 $Y2=1.5
r102 40 42 40.8475 $w=3.54e-07 $l=3e-07 $layer=POLY_cond $X=2.43 $Y=1.5 $X2=2.73
+ $Y2=1.5
r103 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.515 $X2=2.43 $Y2=1.515
r104 38 40 7.4887 $w=3.54e-07 $l=5.5e-08 $layer=POLY_cond $X=2.375 $Y=1.5
+ $X2=2.43 $Y2=1.5
r105 37 38 10.2119 $w=3.54e-07 $l=7.5e-08 $layer=POLY_cond $X=2.3 $Y=1.5
+ $X2=2.375 $Y2=1.5
r106 34 46 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.11 $Y2=1.565
r107 33 46 12.5965 $w=4.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.11 $Y2=1.565
r108 33 41 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.43 $Y2=1.565
r109 29 50 18.5736 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=3.725 $Y=1.68
+ $X2=3.725 $Y2=1.5
r110 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.725 $Y=1.68
+ $X2=3.725 $Y2=2.4
r111 25 49 22.9014 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.59 $Y=1.32
+ $X2=3.59 $Y2=1.5
r112 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.59 $Y=1.32
+ $X2=3.59 $Y2=0.74
r113 21 48 18.5736 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=3.275 $Y=1.68
+ $X2=3.275 $Y2=1.5
r114 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.275 $Y=1.68
+ $X2=3.275 $Y2=2.4
r115 17 47 22.9014 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.16 $Y=1.32
+ $X2=3.16 $Y2=1.5
r116 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.16 $Y=1.32
+ $X2=3.16 $Y2=0.74
r117 13 43 18.5736 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.825 $Y=1.68
+ $X2=2.825 $Y2=1.5
r118 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.825 $Y=1.68
+ $X2=2.825 $Y2=2.4
r119 9 42 22.9014 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.73 $Y=1.32
+ $X2=2.73 $Y2=1.5
r120 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.73 $Y=1.32
+ $X2=2.73 $Y2=0.74
r121 5 38 18.5736 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.375 $Y=1.68
+ $X2=2.375 $Y2=1.5
r122 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.375 $Y=1.68
+ $X2=2.375 $Y2=2.4
r123 1 37 22.9014 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.3 $Y=1.32 $X2=2.3
+ $Y2=1.5
r124 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.3 $Y=1.32 $X2=2.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%A1 3 5 6 9 13 17 21 25 29 33 35 36 37 52
c89 52 0 7.9229e-20 $X=5.755 $Y=1.515
c90 37 0 1.97869e-19 $X=5.52 $Y=1.665
c91 13 0 1.96393e-19 $X=4.625 $Y=2.4
c92 5 0 9.70149e-20 $X=4.465 $Y=1.575
r93 52 53 11.0213 $w=3.28e-07 $l=7.5e-08 $layer=POLY_cond $X=5.755 $Y=1.515
+ $X2=5.83 $Y2=1.515
r94 50 52 50.6982 $w=3.28e-07 $l=3.45e-07 $layer=POLY_cond $X=5.41 $Y=1.515
+ $X2=5.755 $Y2=1.515
r95 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.41
+ $Y=1.515 $X2=5.41 $Y2=1.515
r96 48 50 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=5.4 $Y=1.515 $X2=5.41
+ $Y2=1.515
r97 47 48 47.7591 $w=3.28e-07 $l=3.25e-07 $layer=POLY_cond $X=5.075 $Y=1.515
+ $X2=5.4 $Y2=1.515
r98 46 51 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.07 $Y=1.565
+ $X2=5.41 $Y2=1.565
r99 45 47 0.734756 $w=3.28e-07 $l=5e-09 $layer=POLY_cond $X=5.07 $Y=1.515
+ $X2=5.075 $Y2=1.515
r100 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.07
+ $Y=1.515 $X2=5.07 $Y2=1.515
r101 43 45 14.6951 $w=3.28e-07 $l=1e-07 $layer=POLY_cond $X=4.97 $Y=1.515
+ $X2=5.07 $Y2=1.515
r102 42 43 50.6982 $w=3.28e-07 $l=3.45e-07 $layer=POLY_cond $X=4.625 $Y=1.515
+ $X2=4.97 $Y2=1.515
r103 41 42 12.4909 $w=3.28e-07 $l=8.5e-08 $layer=POLY_cond $X=4.54 $Y=1.515
+ $X2=4.625 $Y2=1.515
r104 37 51 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.41 $Y2=1.565
r105 36 46 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.07 $Y2=1.565
r106 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r107 31 53 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=1.35
+ $X2=5.83 $Y2=1.515
r108 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.83 $Y=1.35
+ $X2=5.83 $Y2=0.74
r109 27 52 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=1.68
+ $X2=5.755 $Y2=1.515
r110 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.755 $Y=1.68
+ $X2=5.755 $Y2=2.4
r111 23 48 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=1.35
+ $X2=5.4 $Y2=1.515
r112 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.4 $Y=1.35 $X2=5.4
+ $Y2=0.74
r113 19 47 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.075 $Y=1.68
+ $X2=5.075 $Y2=1.515
r114 19 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.075 $Y=1.68
+ $X2=5.075 $Y2=2.4
r115 15 43 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.35
+ $X2=4.97 $Y2=1.515
r116 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.97 $Y=1.35
+ $X2=4.97 $Y2=0.74
r117 11 42 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.625 $Y=1.68
+ $X2=4.625 $Y2=1.515
r118 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.625 $Y=1.68
+ $X2=4.625 $Y2=2.4
r119 7 41 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=1.35
+ $X2=4.54 $Y2=1.515
r120 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.54 $Y=1.35 $X2=4.54
+ $Y2=0.74
r121 5 41 25.362 $w=3.28e-07 $l=1.00623e-07 $layer=POLY_cond $X=4.465 $Y=1.575
+ $X2=4.54 $Y2=1.515
r122 5 6 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.465 $Y=1.575
+ $X2=4.265 $Y2=1.575
r123 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.175 $Y=1.65
+ $X2=4.265 $Y2=1.575
r124 1 3 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.175 $Y=1.65
+ $X2=4.175 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%A2 3 7 11 15 19 23 27 31 33 34 35 51 53
c79 53 0 1.97869e-19 $X=7.555 $Y=1.515
c80 7 0 2.04552e-19 $X=6.26 $Y=0.74
r81 52 53 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.55 $Y=1.515
+ $X2=7.555 $Y2=1.515
r82 50 52 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.3 $Y=1.515
+ $X2=7.55 $Y2=1.515
r83 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.3
+ $Y=1.515 $X2=7.3 $Y2=1.515
r84 48 50 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.12 $Y=1.515 $X2=7.3
+ $Y2=1.515
r85 47 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.105 $Y=1.515
+ $X2=7.12 $Y2=1.515
r86 46 47 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=6.69 $Y=1.515
+ $X2=7.105 $Y2=1.515
r87 45 46 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.655 $Y=1.515
+ $X2=6.69 $Y2=1.515
r88 43 45 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=6.28 $Y=1.515
+ $X2=6.655 $Y2=1.515
r89 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.28
+ $Y=1.515 $X2=6.28 $Y2=1.515
r90 41 43 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.26 $Y=1.515 $X2=6.28
+ $Y2=1.515
r91 39 41 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.205 $Y=1.515
+ $X2=6.26 $Y2=1.515
r92 35 51 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.3 $Y2=1.565
r93 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r94 34 44 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.565 $X2=6.28
+ $Y2=1.565
r95 33 44 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=6.28
+ $Y2=1.565
r96 29 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.55 $Y=1.35
+ $X2=7.55 $Y2=1.515
r97 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.55 $Y=1.35
+ $X2=7.55 $Y2=0.74
r98 25 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.555 $Y=1.68
+ $X2=7.555 $Y2=1.515
r99 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.555 $Y=1.68
+ $X2=7.555 $Y2=2.4
r100 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.12 $Y=1.35
+ $X2=7.12 $Y2=1.515
r101 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.12 $Y=1.35
+ $X2=7.12 $Y2=0.74
r102 17 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=1.68
+ $X2=7.105 $Y2=1.515
r103 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.105 $Y=1.68
+ $X2=7.105 $Y2=2.4
r104 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.35
+ $X2=6.69 $Y2=1.515
r105 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.69 $Y=1.35
+ $X2=6.69 $Y2=0.74
r106 9 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.655 $Y=1.68
+ $X2=6.655 $Y2=1.515
r107 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.655 $Y=1.68
+ $X2=6.655 $Y2=2.4
r108 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.26 $Y=1.35
+ $X2=6.26 $Y2=1.515
r109 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.26 $Y=1.35 $X2=6.26
+ $Y2=0.74
r110 1 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.68
+ $X2=6.205 $Y2=1.515
r111 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.205 $Y=1.68
+ $X2=6.205 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%A_45_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40
+ 44 46 50 52 54 57 58 62 64 68 70 74 76 78 80 82 83 84 88 90 92
c138 90 0 7.9229e-20 $X=5.98 $Y=2.035
c139 62 0 1.96393e-19 $X=4.85 $Y=2.415
r140 78 94 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=7.82 $Y=2.12 $X2=7.82
+ $Y2=1.97
r141 78 80 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=7.82 $Y=2.12
+ $X2=7.82 $Y2=2.4
r142 77 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=2.035
+ $X2=6.88 $Y2=2.035
r143 76 94 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=7.695 $Y=2.035
+ $X2=7.82 $Y2=1.97
r144 76 77 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.695 $Y=2.035
+ $X2=6.965 $Y2=2.035
r145 72 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.88 $Y=2.12
+ $X2=6.88 $Y2=2.035
r146 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.88 $Y=2.12
+ $X2=6.88 $Y2=2.465
r147 71 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=2.035
+ $X2=5.94 $Y2=2.035
r148 70 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.035
+ $X2=6.88 $Y2=2.035
r149 70 71 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.795 $Y=2.035
+ $X2=6.065 $Y2=2.035
r150 66 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.035
r151 66 68 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.465
r152 65 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.015 $Y=2.035
+ $X2=4.89 $Y2=2.035
r153 64 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.815 $Y=2.035
+ $X2=5.94 $Y2=2.035
r154 64 65 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.815 $Y=2.035
+ $X2=5.015 $Y2=2.035
r155 60 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.89 $Y=2.12
+ $X2=4.89 $Y2=2.035
r156 60 62 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.89 $Y=2.12
+ $X2=4.89 $Y2=2.415
r157 59 86 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.035 $Y=2.035
+ $X2=3.91 $Y2=1.97
r158 58 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.765 $Y=2.035
+ $X2=4.89 $Y2=2.035
r159 58 59 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.765 $Y=2.035
+ $X2=4.035 $Y2=2.035
r160 55 57 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=3.91 $Y=2.905
+ $X2=3.91 $Y2=2.4
r161 54 86 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.91 $Y=2.12 $X2=3.91
+ $Y2=1.97
r162 54 57 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.91 $Y=2.12
+ $X2=3.91 $Y2=2.4
r163 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=2.99
+ $X2=3.05 $Y2=2.99
r164 52 55 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.785 $Y=2.99
+ $X2=3.91 $Y2=2.905
r165 52 53 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.785 $Y=2.99
+ $X2=3.215 $Y2=2.99
r166 48 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.99
r167 48 50 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.375
r168 47 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=2.99
+ $X2=2.15 $Y2=2.99
r169 46 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=2.99
+ $X2=3.05 $Y2=2.99
r170 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.885 $Y=2.99
+ $X2=2.315 $Y2=2.99
r171 42 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.99
r172 42 44 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.375
r173 41 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=2.99
+ $X2=1.25 $Y2=2.99
r174 40 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=2.15 $Y2=2.99
r175 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=1.415 $Y2=2.99
r176 36 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.905
+ $X2=1.25 $Y2=2.99
r177 36 38 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=1.25 $Y=2.905
+ $X2=1.25 $Y2=2.375
r178 34 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.25 $Y2=2.99
r179 34 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.435 $Y2=2.99
r180 30 33 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.31 $Y=1.985
+ $X2=0.31 $Y2=2.815
r181 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.31 $Y=2.905
+ $X2=0.435 $Y2=2.99
r182 28 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.31 $Y=2.905
+ $X2=0.31 $Y2=2.815
r183 9 94 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.645
+ $Y=1.84 $X2=7.78 $Y2=1.985
r184 9 80 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=7.645
+ $Y=1.84 $X2=7.78 $Y2=2.4
r185 8 92 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.88 $Y2=2.035
r186 8 74 300 $w=1.7e-07 $l=6.89202e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.84 $X2=6.88 $Y2=2.465
r187 7 90 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.98 $Y2=2.035
r188 7 68 300 $w=1.7e-07 $l=6.89202e-07 $layer=licon1_PDIFF $count=2 $X=5.845
+ $Y=1.84 $X2=5.98 $Y2=2.465
r189 6 88 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=1.84 $X2=4.85 $Y2=2.035
r190 6 62 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=4.715
+ $Y=1.84 $X2=4.85 $Y2=2.415
r191 5 86 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.815
+ $Y=1.84 $X2=3.95 $Y2=1.985
r192 5 57 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=3.815
+ $Y=1.84 $X2=3.95 $Y2=2.4
r193 4 50 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.915
+ $Y=1.84 $X2=3.05 $Y2=2.375
r194 3 44 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.84 $X2=2.15 $Y2=2.375
r195 2 38 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=1.115
+ $Y=1.84 $X2=1.25 $Y2=2.375
r196 1 33 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.35 $Y2=2.815
r197 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.35 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%Y 1 2 3 4 5 6 7 8 25 27 29 33 35 39 43 45 46
+ 47 52 54 60 62 64 66 67 69 70
c99 67 0 9.70149e-20 $X=5.45 $Y=0.95
c100 66 0 4.29123e-20 $X=5.615 $Y=0.95
c101 46 0 8.01953e-20 $X=2.68 $Y=1.095
r102 74 75 2.90031 $w=6.52e-07 $l=1.55e-07 $layer=LI1_cond $X=3.375 $Y=1.145
+ $X2=3.53 $Y2=1.145
r103 69 70 8.9816 $w=6.52e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.145
+ $X2=4.08 $Y2=1.145
r104 69 75 1.30982 $w=6.52e-07 $l=7e-08 $layer=LI1_cond $X=3.6 $Y=1.145 $X2=3.53
+ $Y2=1.145
r105 66 67 5.88189 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.615 $Y=0.95
+ $X2=5.45 $Y2=0.95
r106 56 67 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=4.755 $Y=0.99
+ $X2=5.45 $Y2=0.99
r107 54 70 6.20325 $w=6.52e-07 $l=2.04573e-07 $layer=LI1_cond $X=4.195 $Y=0.99
+ $X2=4.08 $Y2=1.145
r108 54 56 23.0489 $w=2.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.195 $Y=0.99
+ $X2=4.755 $Y2=0.99
r109 52 64 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.53 $Y=1.95
+ $X2=3.515 $Y2=2.035
r110 51 75 8.85584 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=3.53 $Y=1.52
+ $X2=3.53 $Y2=1.145
r111 51 52 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.53 $Y=1.52
+ $X2=3.53 $Y2=1.95
r112 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=2.035
+ $X2=2.6 $Y2=2.035
r113 47 64 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.415 $Y=2.035
+ $X2=3.515 $Y2=2.035
r114 47 48 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.415 $Y=2.035
+ $X2=2.685 $Y2=2.035
r115 45 74 10.7048 $w=6.52e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.375 $Y2=1.145
r116 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=2.68 $Y2=1.095
r117 41 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=2.12 $X2=2.6
+ $Y2=2.035
r118 41 43 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.6 $Y=2.12 $X2=2.6
+ $Y2=2.57
r119 37 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.68 $Y2=1.095
r120 37 39 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.515 $Y2=0.76
r121 36 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.7 $Y2=2.035
r122 35 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=2.6 $Y2=2.035
r123 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=1.785 $Y2=2.035
r124 31 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.12 $X2=1.7
+ $Y2=2.035
r125 31 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.7 $Y=2.12 $X2=1.7
+ $Y2=2.57
r126 30 58 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=2.035
+ $X2=0.76 $Y2=2.035
r127 29 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=1.7 $Y2=2.035
r128 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=0.885 $Y2=2.035
r129 25 58 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.12
+ $X2=0.76 $Y2=2.035
r130 25 27 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.76 $Y=2.12
+ $X2=0.76 $Y2=2.57
r131 8 64 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=3.365
+ $Y=1.84 $X2=3.5 $Y2=2.115
r132 7 62 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=2.035
r133 7 43 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.84 $X2=2.6 $Y2=2.57
r134 6 60 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.84 $X2=1.7 $Y2=2.035
r135 6 33 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.84 $X2=1.7 $Y2=2.57
r136 5 58 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.84 $X2=0.8 $Y2=2.035
r137 5 27 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.84 $X2=0.8 $Y2=2.57
r138 4 66 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.475
+ $Y=0.37 $X2=5.615 $Y2=0.95
r139 3 56 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.37 $X2=4.755 $Y2=0.95
r140 2 74 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.37 $X2=3.375 $Y2=0.91
r141 1 39 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.37 $X2=2.515 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 44
+ 48 58 59 62 65
r100 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r103 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 56 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 53 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.43 $Y2=3.33
r107 53 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r109 52 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r110 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r111 49 62 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.415 $Y2=3.33
r112 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=6 $Y2=3.33
r113 48 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6.43 $Y2=3.33
r114 48 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6 $Y2=3.33
r115 47 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r116 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 44 62 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.415 $Y2=3.33
r118 44 46 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 38 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r120 38 39 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r121 35 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 35 39 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=0.24 $Y2=3.33
r123 35 42 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 33 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.165 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=3.33
+ $X2=7.33 $Y2=3.33
r126 32 58 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.495 $Y=3.33
+ $X2=7.92 $Y2=3.33
r127 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.495 $Y=3.33
+ $X2=7.33 $Y2=3.33
r128 30 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.4 $Y2=3.33
r130 29 46 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.565 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=3.33
+ $X2=4.4 $Y2=3.33
r132 25 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=3.245
+ $X2=7.33 $Y2=3.33
r133 25 27 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.33 $Y=3.245
+ $X2=7.33 $Y2=2.375
r134 21 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=3.33
r135 21 23 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=2.375
r136 17 62 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=3.245
+ $X2=5.415 $Y2=3.33
r137 17 19 22.6215 $w=4.58e-07 $l=8.7e-07 $layer=LI1_cond $X=5.415 $Y=3.245
+ $X2=5.415 $Y2=2.375
r138 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=3.245 $X2=4.4
+ $Y2=3.33
r139 13 15 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=4.4 $Y=3.245
+ $X2=4.4 $Y2=2.375
r140 4 27 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=7.195
+ $Y=1.84 $X2=7.33 $Y2=2.375
r141 3 23 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.375
r142 2 19 300 $w=1.7e-07 $l=6.48055e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.84 $X2=5.415 $Y2=2.375
r143 1 15 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=4.265
+ $Y=1.84 $X2=4.4 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%A_48_74# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 39
r66 34 43 10.9604 $w=1.68e-07 $l=1.68e-07 $layer=LI1_cond $X=2.945 $Y=0.427
+ $X2=2.945 $Y2=0.595
r67 34 39 5.67594 $w=1.68e-07 $l=8.7e-08 $layer=LI1_cond $X=2.945 $Y=0.427
+ $X2=2.945 $Y2=0.34
r68 34 36 25.8882 $w=3.43e-07 $l=7.75e-07 $layer=LI1_cond $X=3.03 $Y=0.427
+ $X2=3.805 $Y2=0.427
r69 32 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.34
+ $X2=2.945 $Y2=0.34
r70 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.86 $Y=0.34 $X2=2.17
+ $Y2=0.34
r71 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.085 $Y=1.01
+ $X2=2.085 $Y2=0.515
r72 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=0.425
+ $X2=2.17 $Y2=0.34
r73 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.085 $Y=0.425
+ $X2=2.085 $Y2=0.515
r74 27 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.31 $Y=1.095
+ $X2=1.185 $Y2=1.095
r75 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2 $Y=1.095
+ $X2=2.085 $Y2=1.01
r76 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2 $Y=1.095 $X2=1.31
+ $Y2=1.095
r77 22 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.01
+ $X2=1.185 $Y2=1.095
r78 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.185 $Y=1.01
+ $X2=1.185 $Y2=0.515
r79 20 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.06 $Y=1.095
+ $X2=1.185 $Y2=1.095
r80 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.06 $Y=1.095
+ $X2=0.45 $Y2=1.095
r81 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.325 $Y=1.01
+ $X2=0.45 $Y2=1.095
r82 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.325 $Y=1.01
+ $X2=0.325 $Y2=0.515
r83 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.37 $X2=3.805 $Y2=0.515
r84 4 43 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.37 $X2=2.945 $Y2=0.595
r85 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.37 $X2=2.085 $Y2=0.515
r86 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.37 $X2=1.225 $Y2=0.515
r87 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.24
+ $Y=0.37 $X2=0.365 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 42 58 59 62 65
c94 19 0 1.9142e-19 $X=1.655 $Y=0.675
r95 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r96 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r98 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r99 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r100 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r101 52 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r102 50 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r103 49 52 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r104 49 50 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r105 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.655
+ $Y2=0
r106 47 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=2.16
+ $Y2=0
r107 46 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r108 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r110 43 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.755
+ $Y2=0
r111 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r112 42 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.655
+ $Y2=0
r113 42 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.2
+ $Y2=0
r114 40 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r115 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r116 37 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.755
+ $Y2=0
r117 37 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r118 35 53 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r119 35 50 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.16 $Y2=0
r120 33 55 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=6.96
+ $Y2=0
r121 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.295
+ $Y2=0
r122 32 58 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.92
+ $Y2=0
r123 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.295
+ $Y2=0
r124 30 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.31 $Y=0 $X2=6
+ $Y2=0
r125 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.31 $Y=0 $X2=6.435
+ $Y2=0
r126 29 55 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.96
+ $Y2=0
r127 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.435
+ $Y2=0
r128 25 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0
r129 25 27 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0.595
r130 21 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0
r131 21 23 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0.595
r132 17 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0
r133 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0.675
r134 13 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r135 13 15 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.675
r136 4 27 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.37 $X2=7.335 $Y2=0.595
r137 3 23 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.37 $X2=6.475 $Y2=0.595
r138 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.37 $X2=1.655 $Y2=0.675
r139 1 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.655
+ $Y=0.37 $X2=0.795 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_4%A_840_74# 1 2 3 4 5 16 20 24 25 28 30 34 39
+ 42
c62 20 0 1.6164e-19 $X=6.045 $Y=0.6
r63 37 39 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0.515
+ $X2=4.49 $Y2=0.515
r64 32 34 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.765 $Y=1.01
+ $X2=7.765 $Y2=0.515
r65 31 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.99 $Y=1.095
+ $X2=6.865 $Y2=1.095
r66 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.6 $Y=1.095
+ $X2=7.765 $Y2=1.01
r67 30 31 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.6 $Y=1.095
+ $X2=6.99 $Y2=1.095
r68 26 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=1.01
+ $X2=6.865 $Y2=1.095
r69 26 28 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=6.865 $Y=1.01
+ $X2=6.865 $Y2=0.515
r70 24 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.74 $Y=1.095
+ $X2=6.865 $Y2=1.095
r71 24 25 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.74 $Y=1.095
+ $X2=6.13 $Y2=1.095
r72 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.045 $Y=1.01
+ $X2=6.13 $Y2=1.095
r73 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.045 $Y=1.01
+ $X2=6.045 $Y2=0.965
r74 20 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.045 $Y=0.6
+ $X2=6.045 $Y2=0.475
r75 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.045 $Y=0.6
+ $X2=6.045 $Y2=0.965
r76 19 39 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.185 $Y=0.475
+ $X2=4.49 $Y2=0.475
r77 16 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=0.475
+ $X2=6.045 $Y2=0.475
r78 16 19 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=5.96 $Y=0.475
+ $X2=5.185 $Y2=0.475
r79 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.625
+ $Y=0.37 $X2=7.765 $Y2=0.515
r80 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.37 $X2=6.905 $Y2=0.515
r81 3 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.515
r82 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.965
r83 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.37 $X2=5.185 $Y2=0.515
r84 1 37 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.37 $X2=4.325 $Y2=0.515
.ends


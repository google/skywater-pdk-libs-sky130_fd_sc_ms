* NGSPICE file created from sky130_fd_sc_ms__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR D a_27_112# VPB pshort w=840000u l=180000u
+  ad=2.6463e+12p pd=2.068e+07u as=2.352e+11p ps=2.24e+06u
M1001 VPWR a_230_74# a_363_82# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1002 VGND a_230_74# a_363_82# VNB nlowvt w=740000u l=150000u
+  ad=1.8561e+12p pd=1.54e+07u as=2.109e+11p ps=2.05e+06u
M1003 a_773_124# a_230_74# a_641_80# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.692e+11p ps=2.3e+06u
M1004 a_569_80# a_27_112# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 Q_N a_1449_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1006 VGND a_821_98# a_1449_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1007 VPWR a_821_98# a_760_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1008 VPWR a_1449_368# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND RESET_B a_1049_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1010 a_569_392# a_27_112# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1011 Q_N a_1449_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1012 VPWR a_821_98# a_1449_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1013 a_230_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_641_80# a_230_74# a_569_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=0p ps=0u
M1015 VGND D a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1016 a_1049_74# a_641_80# a_821_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_230_74# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.772e+11p pd=2.34e+06u as=0p ps=0u
M1018 VGND a_821_98# a_773_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1449_368# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_760_508# a_363_82# a_641_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q a_821_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1022 VPWR a_821_98# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_641_80# a_363_82# a_569_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_821_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1025 VGND a_821_98# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR RESET_B a_821_98# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=2.88e+06u
M1027 a_821_98# a_641_80# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__maj3_2.pex.spice
* Created: Fri Aug 28 17:38:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MAJ3_2%A_87_264# 1 2 3 4 15 19 23 27 29 32 33 35 39
+ 41 43 46 47 53 55
r134 63 64 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.945 $Y=1.485
+ $X2=0.975 $Y2=1.485
r135 62 63 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.525 $Y=1.485
+ $X2=0.945 $Y2=1.485
r136 60 62 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.515 $Y=1.485
+ $X2=0.525 $Y2=1.485
r137 55 57 1.38244 $w=7.06e-07 $l=8e-08 $layer=LI1_cond $X=2.375 $Y=2.035
+ $X2=2.375 $Y2=2.115
r138 52 53 10.9648 $w=7.23e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0.712
+ $X2=2.76 $Y2=0.712
r139 49 52 8.99121 $w=7.23e-07 $l=5.45e-07 $layer=LI1_cond $X=2.05 $Y=0.712
+ $X2=2.595 $Y2=0.712
r140 47 64 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.06 $Y=1.485
+ $X2=0.975 $Y2=1.485
r141 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.485 $X2=1.06 $Y2=1.485
r142 41 59 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.52 $Y=2.12 $X2=4.52
+ $Y2=1.97
r143 41 43 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=4.52 $Y=2.12
+ $X2=4.52 $Y2=2.695
r144 37 39 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.495 $Y=0.905
+ $X2=4.495 $Y2=0.515
r145 36 55 9.37777 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=2.785 $Y=2.035
+ $X2=2.375 $Y2=2.035
r146 35 59 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=4.355 $Y=2.035
+ $X2=4.52 $Y2=1.97
r147 35 36 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=4.355 $Y=2.035
+ $X2=2.785 $Y2=2.035
r148 33 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.33 $Y=0.99
+ $X2=4.495 $Y2=0.905
r149 33 53 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=4.33 $Y=0.99
+ $X2=2.76 $Y2=0.99
r150 31 49 9.55322 $w=1.7e-07 $l=3.63e-07 $layer=LI1_cond $X=2.05 $Y=1.075
+ $X2=2.05 $Y2=0.712
r151 31 32 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.05 $Y=1.075
+ $X2=2.05 $Y2=1.78
r152 30 46 17.2342 $w=2.69e-07 $l=4.61302e-07 $layer=LI1_cond $X=1.255 $Y=1.865
+ $X2=1.075 $Y2=1.485
r153 29 55 2.93768 $w=7.06e-07 $l=4.87647e-07 $layer=LI1_cond $X=1.965 $Y=1.865
+ $X2=2.375 $Y2=2.035
r154 29 32 9.67802 $w=7.06e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.965 $Y=1.865
+ $X2=2.05 $Y2=1.78
r155 29 30 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.965 $Y=1.865
+ $X2=1.255 $Y2=1.865
r156 25 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.65
+ $X2=0.975 $Y2=1.485
r157 25 27 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.975 $Y=1.65
+ $X2=0.975 $Y2=2.4
r158 21 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.32
+ $X2=0.945 $Y2=1.485
r159 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.945 $Y=1.32
+ $X2=0.945 $Y2=0.74
r160 17 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.32
+ $X2=0.515 $Y2=1.485
r161 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.515 $Y=1.32
+ $X2=0.515 $Y2=0.74
r162 13 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.65
+ $X2=0.525 $Y2=1.485
r163 13 15 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.525 $Y=1.65
+ $X2=0.525 $Y2=2.4
r164 4 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=1.985
r165 4 43 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.695
r166 3 57 300 $w=1.7e-07 $l=4.4238e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=1.735 $X2=2.62 $Y2=2.115
r167 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.37 $X2=4.495 $Y2=0.515
r168 1 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.455
+ $Y=0.37 $X2=2.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_2%B 3 7 11 15 17 24 25
r45 23 25 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.81 $Y=1.41
+ $X2=2.845 $Y2=1.41
r46 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.81
+ $Y=1.41 $X2=2.81 $Y2=1.41
r47 21 23 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.81 $Y2=1.41
r48 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.38 $Y=1.41
+ $X2=2.395 $Y2=1.41
r49 17 24 4.55224 $w=6.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.41
r50 13 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.575
+ $X2=2.845 $Y2=1.41
r51 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.845 $Y=1.575
+ $X2=2.845 $Y2=2.235
r52 9 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.245
+ $X2=2.81 $Y2=1.41
r53 9 11 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.81 $Y=1.245
+ $X2=2.81 $Y2=0.74
r54 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.575
+ $X2=2.395 $Y2=1.41
r55 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.395 $Y=1.575
+ $X2=2.395 $Y2=2.235
r56 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.245
+ $X2=2.38 $Y2=1.41
r57 1 3 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.38 $Y=1.245
+ $X2=2.38 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_2%C 3 7 11 15 19 20 22 25 26
r62 26 34 1.31569 $w=4.98e-07 $l=5.5e-08 $layer=LI1_cond $X=3.465 $Y=1.41
+ $X2=3.465 $Y2=1.465
r63 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.575
r64 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.245
r65 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.41 $X2=3.38 $Y2=1.41
r66 22 34 4.78431 $w=4.98e-07 $l=2e-07 $layer=LI1_cond $X=3.465 $Y=1.665
+ $X2=3.465 $Y2=1.465
r67 20 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.465
+ $X2=4.37 $Y2=1.63
r68 20 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.465
+ $X2=4.37 $Y2=1.3
r69 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=1.465 $X2=4.37 $Y2=1.465
r70 17 34 3.16914 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=3.715 $Y=1.465
+ $X2=3.465 $Y2=1.465
r71 17 19 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.715 $Y=1.465
+ $X2=4.37 $Y2=1.465
r72 15 31 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=4.295 $Y=2.34
+ $X2=4.295 $Y2=1.63
r73 11 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.28 $Y=0.74
+ $X2=4.28 $Y2=1.3
r74 7 28 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.305 $Y=2.235
+ $X2=3.305 $Y2=1.575
r75 3 27 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.29 $Y=0.74
+ $X2=3.29 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_2%A 4 5 7 8 9 10 13 16 18 19 21
r70 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.385 $X2=1.63 $Y2=1.385
r71 21 25 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.63 $Y=1.295 $X2=1.63
+ $Y2=1.385
r72 18 24 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.8 $Y=1.385
+ $X2=1.63 $Y2=1.385
r73 18 19 3.90195 $w=3.3e-07 $l=1.32e-07 $layer=POLY_cond $X=1.8 $Y=1.385
+ $X2=1.932 $Y2=1.385
r74 16 20 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.89 $Y=0.74
+ $X2=3.89 $Y2=1.615
r75 11 13 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=3.875 $Y=3.075
+ $X2=3.875 $Y2=2.34
r76 10 20 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.875 $Y=1.705
+ $X2=3.875 $Y2=1.615
r77 10 13 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=3.875 $Y=1.705
+ $X2=3.875 $Y2=2.34
r78 8 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.785 $Y=3.15
+ $X2=3.875 $Y2=3.075
r79 8 9 925.543 $w=1.5e-07 $l=1.805e-06 $layer=POLY_cond $X=3.785 $Y=3.15
+ $X2=1.98 $Y2=3.15
r80 5 19 34.7346 $w=1.65e-07 $l=1.9182e-07 $layer=POLY_cond $X=1.99 $Y=1.22
+ $X2=1.932 $Y2=1.385
r81 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.99 $Y=1.22 $X2=1.99
+ $Y2=0.74
r82 2 9 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.89 $Y=3.075
+ $X2=1.98 $Y2=3.15
r83 2 4 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=1.89 $Y=3.075
+ $X2=1.89 $Y2=2.34
r84 1 19 34.7346 $w=1.65e-07 $l=1.84811e-07 $layer=POLY_cond $X=1.89 $Y=1.55
+ $X2=1.932 $Y2=1.385
r85 1 4 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.89 $Y=1.55 $X2=1.89
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_2%VPWR 1 2 3 10 12 18 24 26 28 33 43 44 50 53
r48 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 44 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r53 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.65 $Y2=3.33
r54 41 43 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=4.56 $Y2=3.33
r55 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r59 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 34 50 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=1.78 $Y=3.33
+ $X2=1.432 $Y2=3.33
r61 34 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 33 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.65 $Y2=3.33
r63 33 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 32 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 29 47 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.192 $Y2=3.33
r68 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 28 50 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.432 $Y2=3.33
r70 28 31 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 26 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 22 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=3.245
+ $X2=3.65 $Y2=3.33
r74 22 24 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.65 $Y=3.245
+ $X2=3.65 $Y2=2.375
r75 18 21 9.03512 $w=6.93e-07 $l=5.25e-07 $layer=LI1_cond $X=1.432 $Y=2.285
+ $X2=1.432 $Y2=2.81
r76 16 50 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.432 $Y=3.245
+ $X2=1.432 $Y2=3.33
r77 16 21 7.48625 $w=6.93e-07 $l=4.35e-07 $layer=LI1_cond $X=1.432 $Y=3.245
+ $X2=1.432 $Y2=2.81
r78 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.26 $Y=1.985
+ $X2=0.26 $Y2=2.815
r79 10 47 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.192 $Y2=3.33
r80 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.815
r81 3 24 300 $w=1.7e-07 $l=7.56836e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=1.735 $X2=3.65 $Y2=2.375
r82 2 21 300 $w=1.7e-07 $l=1.03764e-06 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=1.84 $X2=1.205 $Y2=2.81
r83 2 18 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=1.84 $X2=1.205 $Y2=2.285
r84 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.3 $Y2=2.815
r85 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.3 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_2%X 1 2 9 13 14 15 16 23 32
r31 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.735 $Y=2 $X2=0.735
+ $Y2=2.035
r32 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.735 $Y=2.405
+ $X2=0.735 $Y2=2.775
r33 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.735 $Y=1.975
+ $X2=0.735 $Y2=2
r34 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.735 $Y=1.975
+ $X2=0.735 $Y2=1.82
r35 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.735 $Y=2.06
+ $X2=0.735 $Y2=2.405
r36 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.735 $Y=2.06
+ $X2=0.735 $Y2=2.035
r37 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.64 $Y=1.13 $X2=0.64
+ $Y2=1.82
r38 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.725 $Y=0.96
+ $X2=0.725 $Y2=1.13
r39 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=0.725 $Y=0.96
+ $X2=0.725 $Y2=0.515
r40 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.84 $X2=0.75 $Y2=1.985
r41 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.84 $X2=0.75 $Y2=2.815
r42 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 51
r50 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 47 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r52 46 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 40 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r56 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r57 37 51 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.59
+ $Y2=0
r58 37 39 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r59 36 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r60 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r63 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r64 30 46 13.8654 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.435
+ $Y2=0
r65 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=2.16
+ $Y2=0
r66 29 51 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.59
+ $Y2=0
r67 29 35 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.34 $Y=0 $X2=3.12
+ $Y2=0
r68 28 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r69 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r70 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 25 43 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r72 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.72
+ $Y2=0
r73 24 46 13.8654 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.435
+ $Y2=0
r74 24 27 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.72
+ $Y2=0
r75 22 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r76 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r77 18 51 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=0.085 $X2=3.59
+ $Y2=0
r78 18 20 11.4824 $w=4.98e-07 $l=4.8e-07 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0.565
r79 14 46 2.92113 $w=7.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0.085
+ $X2=1.435 $Y2=0
r80 14 16 6.97712 $w=7.18e-07 $l=4.2e-07 $layer=LI1_cond $X=1.435 $Y=0.085
+ $X2=1.435 $Y2=0.505
r81 10 43 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.192 $Y2=0
r82 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.515
r83 3 20 182 $w=1.7e-07 $l=3.07409e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.37 $X2=3.59 $Y2=0.565
r84 2 16 45.5 $w=1.7e-07 $l=7.54487e-07 $layer=licon1_NDIFF $count=4 $X=1.02
+ $Y=0.37 $X2=1.71 $Y2=0.505
r85 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__ebufn_4.pex.spice
* Created: Wed Sep  2 12:07:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EBUFN_4%A 3 7 9 12
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.465
+ $X2=0.515 $Y2=1.63
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.465
+ $X2=0.515 $Y2=1.3
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.465 $X2=0.515 $Y2=1.465
r38 9 13 5.10825 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.515 $Y2=1.54
r39 7 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.535 $Y=0.74
+ $X2=0.535 $Y2=1.3
r40 3 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%TE_B 3 5 6 8 9 11 13 14 16 18 19 21 23 24 26
+ 28 29 30 31 32 33 36 38
c119 26 0 6.07806e-20 $X=3.46 $Y=1.725
c120 21 0 1.01045e-19 $X=3.01 $Y=1.725
c121 19 0 1.6749e-19 $X=2.92 $Y=1.65
c122 16 0 1.60162e-19 $X=2.56 $Y=1.725
c123 14 0 1.23507e-19 $X=2.47 $Y=1.65
r124 36 38 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.385
+ $X2=1.065 $Y2=1.22
r125 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.385 $X2=1.075 $Y2=1.385
r126 33 37 3.89339 $w=3.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=1.075 $Y2=1.365
r127 26 28 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.46 $Y=1.725
+ $X2=3.46 $Y2=2.4
r128 25 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.1 $Y=1.65 $X2=3.01
+ $Y2=1.65
r129 24 26 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.37 $Y=1.65
+ $X2=3.46 $Y2=1.725
r130 24 25 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.37 $Y=1.65
+ $X2=3.1 $Y2=1.65
r131 21 32 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.01 $Y=1.725
+ $X2=3.01 $Y2=1.65
r132 21 23 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.01 $Y=1.725
+ $X2=3.01 $Y2=2.4
r133 20 31 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.65 $Y=1.65 $X2=2.56
+ $Y2=1.65
r134 19 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.92 $Y=1.65 $X2=3.01
+ $Y2=1.65
r135 19 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.92 $Y=1.65
+ $X2=2.65 $Y2=1.65
r136 16 31 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.725
+ $X2=2.56 $Y2=1.65
r137 16 18 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.56 $Y=1.725
+ $X2=2.56 $Y2=2.4
r138 15 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.2 $Y=1.65 $X2=2.11
+ $Y2=1.65
r139 14 31 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.47 $Y=1.65 $X2=2.56
+ $Y2=1.65
r140 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.47 $Y=1.65
+ $X2=2.2 $Y2=1.65
r141 11 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.11 $Y=1.725
+ $X2=2.11 $Y2=1.65
r142 11 13 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.11 $Y=1.725
+ $X2=2.11 $Y2=2.4
r143 10 29 13.6393 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.24 $Y=1.65
+ $X2=1.065 $Y2=1.65
r144 9 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.02 $Y=1.65 $X2=2.11
+ $Y2=1.65
r145 9 10 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.02 $Y=1.65
+ $X2=1.24 $Y2=1.65
r146 6 29 12.4285 $w=2.65e-07 $l=1.16619e-07 $layer=POLY_cond $X=0.98 $Y=1.725
+ $X2=1.065 $Y2=1.65
r147 6 8 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=0.98 $Y=1.725
+ $X2=0.98 $Y2=2.4
r148 5 29 12.4285 $w=2.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.065 $Y=1.575
+ $X2=1.065 $Y2=1.65
r149 4 36 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=1.065 $Y=1.395
+ $X2=1.065 $Y2=1.385
r150 4 5 29.6765 $w=3.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.065 $Y=1.395
+ $X2=1.065 $Y2=1.575
r151 3 38 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.965 $Y=0.74
+ $X2=0.965 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%A_208_74# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 28 29 30 33 36 38 48 49
c107 24 0 2.0941e-19 $X=3.535 $Y=1.185
c108 22 0 1.06758e-19 $X=3.46 $Y=1.26
c109 19 0 1.27021e-19 $X=3.105 $Y=1.185
c110 14 0 8.52094e-20 $X=2.675 $Y=1.185
r111 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=0.465 $X2=1.615 $Y2=0.465
r112 45 48 7.32809 $w=7.08e-07 $l=4.35e-07 $layer=LI1_cond $X=1.18 $Y=0.655
+ $X2=1.615 $Y2=0.655
r113 39 49 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=1.615 $Y=1.145
+ $X2=1.615 $Y2=0.465
r114 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.615
+ $Y=1.145 $X2=1.615 $Y2=1.145
r115 36 38 20.708 $w=3.18e-07 $l=5.75e-07 $layer=LI1_cond $X=1.615 $Y=1.72
+ $X2=1.615 $Y2=1.145
r116 35 48 5.42292 $w=3.2e-07 $l=3.55e-07 $layer=LI1_cond $X=1.615 $Y=1.01
+ $X2=1.615 $Y2=0.655
r117 35 38 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=1.615 $Y=1.01
+ $X2=1.615 $Y2=1.145
r118 31 36 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.165 $Y=1.805
+ $X2=1.615 $Y2=1.805
r119 31 33 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.165 $Y=1.89
+ $X2=1.165 $Y2=2.02
r120 27 39 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.615 $Y=1.185
+ $X2=1.615 $Y2=1.145
r121 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.535 $Y=1.185
+ $X2=3.535 $Y2=0.74
r122 23 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=1.26
+ $X2=3.105 $Y2=1.26
r123 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.46 $Y=1.26
+ $X2=3.535 $Y2=1.185
r124 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.46 $Y=1.26
+ $X2=3.18 $Y2=1.26
r125 19 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=1.185
+ $X2=3.105 $Y2=1.26
r126 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.105 $Y=1.185
+ $X2=3.105 $Y2=0.74
r127 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.75 $Y=1.26
+ $X2=2.675 $Y2=1.26
r128 17 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.03 $Y=1.26
+ $X2=3.105 $Y2=1.26
r129 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.03 $Y=1.26
+ $X2=2.75 $Y2=1.26
r130 14 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=1.185
+ $X2=2.675 $Y2=1.26
r131 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.675 $Y=1.185
+ $X2=2.675 $Y2=0.74
r132 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.32 $Y=1.26
+ $X2=2.245 $Y2=1.26
r133 12 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.6 $Y=1.26
+ $X2=2.675 $Y2=1.26
r134 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.6 $Y=1.26
+ $X2=2.32 $Y2=1.26
r135 9 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.245 $Y=1.185
+ $X2=2.245 $Y2=1.26
r136 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.245 $Y=1.185
+ $X2=2.245 $Y2=0.74
r137 8 27 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.78 $Y=1.26
+ $X2=1.615 $Y2=1.185
r138 7 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.17 $Y=1.26
+ $X2=2.245 $Y2=1.26
r139 7 8 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.17 $Y=1.26 $X2=1.78
+ $Y2=1.26
r140 2 33 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.84 $X2=1.205 $Y2=2.02
r141 1 45 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.04
+ $Y=0.37 $X2=1.18 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%A_27_368# 1 2 9 13 17 21 25 29 33 37 41 45
+ 48 51 53 56 57 58 60 62 65 68 71 72 73 74 85
c167 65 0 1.06758e-19 $X=3.985 $Y=1.485
c168 9 0 1.71649e-19 $X=3.91 $Y=2.4
r169 84 85 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.26 $Y=1.485
+ $X2=5.275 $Y2=1.485
r170 83 84 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=4.825 $Y=1.485
+ $X2=5.26 $Y2=1.485
r171 82 83 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.81 $Y=1.485
+ $X2=4.825 $Y2=1.485
r172 79 80 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.36 $Y=1.485
+ $X2=4.395 $Y2=1.485
r173 75 77 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.91 $Y=1.485
+ $X2=3.965 $Y2=1.485
r174 71 72 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.17 $Y=1.13
+ $X2=0.17 $Y2=1.95
r175 69 82 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.665 $Y=1.485
+ $X2=4.81 $Y2=1.485
r176 69 80 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.665 $Y=1.485
+ $X2=4.395 $Y2=1.485
r177 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.665
+ $Y=1.485 $X2=4.665 $Y2=1.485
r178 66 79 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.985 $Y=1.485
+ $X2=4.36 $Y2=1.485
r179 66 77 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.985 $Y=1.485
+ $X2=3.965 $Y2=1.485
r180 65 74 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=1.485
+ $X2=3.82 $Y2=1.485
r181 65 68 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.985 $Y=1.485
+ $X2=4.665 $Y2=1.485
r182 65 66 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.985
+ $Y=1.485 $X2=3.985 $Y2=1.485
r183 62 74 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.53 $Y=1.565
+ $X2=3.82 $Y2=1.565
r184 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=1.65
+ $X2=2.53 $Y2=1.565
r185 59 60 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.445 $Y=1.65
+ $X2=2.445 $Y2=2.06
r186 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=2.145
+ $X2=2.445 $Y2=2.06
r187 57 58 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.36 $Y=2.145
+ $X2=1.63 $Y2=2.145
r188 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.545 $Y=2.23
+ $X2=1.63 $Y2=2.145
r189 55 56 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.545 $Y=2.23
+ $X2=1.545 $Y2=2.39
r190 54 73 3.18746 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=2.475
+ $X2=0.225 $Y2=2.475
r191 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=2.475
+ $X2=1.545 $Y2=2.39
r192 53 54 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=1.46 $Y=2.475
+ $X2=0.365 $Y2=2.475
r193 49 73 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=2.56
+ $X2=0.225 $Y2=2.475
r194 49 51 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=2.56
+ $X2=0.225 $Y2=2.815
r195 46 73 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=2.39
+ $X2=0.225 $Y2=2.475
r196 46 48 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=0.225 $Y=2.39
+ $X2=0.225 $Y2=2.115
r197 45 72 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=2.09
+ $X2=0.225 $Y2=1.95
r198 45 48 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.225 $Y=2.09
+ $X2=0.225 $Y2=2.115
r199 39 71 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.245 $Y=0.97
+ $X2=0.245 $Y2=1.13
r200 39 41 16.3863 $w=3.18e-07 $l=4.55e-07 $layer=LI1_cond $X=0.245 $Y=0.97
+ $X2=0.245 $Y2=0.515
r201 35 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.32
+ $X2=5.275 $Y2=1.485
r202 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.275 $Y=1.32
+ $X2=5.275 $Y2=0.74
r203 31 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.26 $Y=1.65
+ $X2=5.26 $Y2=1.485
r204 31 33 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.26 $Y=1.65
+ $X2=5.26 $Y2=2.4
r205 27 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=1.32
+ $X2=4.825 $Y2=1.485
r206 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.825 $Y=1.32
+ $X2=4.825 $Y2=0.74
r207 23 82 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.65
+ $X2=4.81 $Y2=1.485
r208 23 25 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.81 $Y=1.65
+ $X2=4.81 $Y2=2.4
r209 19 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.32
+ $X2=4.395 $Y2=1.485
r210 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.395 $Y=1.32
+ $X2=4.395 $Y2=0.74
r211 15 79 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.65
+ $X2=4.36 $Y2=1.485
r212 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.36 $Y=1.65
+ $X2=4.36 $Y2=2.4
r213 11 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.32
+ $X2=3.965 $Y2=1.485
r214 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.965 $Y=1.32
+ $X2=3.965 $Y2=0.74
r215 7 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=1.65
+ $X2=3.91 $Y2=1.485
r216 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.91 $Y=1.65 $X2=3.91
+ $Y2=2.4
r217 2 51 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r218 2 48 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r219 1 41 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.175
+ $Y=0.37 $X2=0.32 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%VPWR 1 2 3 12 16 18 22 24 25 26 28 45 46 49
+ 52
r70 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 43 46 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 43 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 42 45 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r76 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r77 40 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.32 $Y=3.33
+ $X2=3.195 $Y2=3.33
r78 40 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.32 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r81 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r83 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r84 33 49 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=0.742 $Y2=3.33
r85 33 35 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=1.2
+ $Y2=3.33
r86 31 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 28 49 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.742 $Y2=3.33
r89 28 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 26 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r91 26 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 24 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.17 $Y=3.33 $X2=2.16
+ $Y2=3.33
r93 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=3.33
+ $X2=2.335 $Y2=3.33
r94 20 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=3.245
+ $X2=3.195 $Y2=3.33
r95 20 22 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=3.195 $Y=3.245
+ $X2=3.195 $Y2=2.325
r96 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=3.33
+ $X2=2.335 $Y2=3.33
r97 18 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=3.195 $Y2=3.33
r98 18 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.07 $Y=3.33 $X2=2.5
+ $Y2=3.33
r99 14 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=3.245
+ $X2=2.335 $Y2=3.33
r100 14 16 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.335 $Y=3.245
+ $X2=2.335 $Y2=2.825
r101 10 49 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=3.33
r102 10 12 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=0.742 $Y=3.245
+ $X2=0.742 $Y2=2.815
r103 3 22 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=3.1
+ $Y=1.84 $X2=3.235 $Y2=2.325
r104 2 16 600 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=1.84 $X2=2.335 $Y2=2.825
r105 1 12 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.74 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%A_348_368# 1 2 3 4 5 16 18 22 24 26 29 30 31
+ 34 36 40 46 53
c65 31 0 1.01045e-19 $X=3.77 $Y=2.99
c66 26 0 1.71649e-19 $X=3.645 $Y=1.99
c67 18 0 1.60162e-19 $X=2.785 $Y=1.99
c68 16 0 1.23507e-19 $X=2.7 $Y=2.485
r69 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.525 $Y=1.985
+ $X2=5.525 $Y2=2.815
r70 38 43 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.525 $Y=2.905
+ $X2=5.525 $Y2=2.815
r71 37 53 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.7 $Y=2.99
+ $X2=4.585 $Y2=2.99
r72 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.4 $Y=2.99
+ $X2=5.525 $Y2=2.905
r73 36 37 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.4 $Y=2.99 $X2=4.7
+ $Y2=2.99
r74 32 53 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=2.905
+ $X2=4.585 $Y2=2.99
r75 32 34 29.0616 $w=2.28e-07 $l=5.8e-07 $layer=LI1_cond $X=4.585 $Y=2.905
+ $X2=4.585 $Y2=2.325
r76 30 53 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.47 $Y=2.99
+ $X2=4.585 $Y2=2.99
r77 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.47 $Y=2.99 $X2=3.77
+ $Y2=2.99
r78 27 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.645 $Y=2.905
+ $X2=3.77 $Y2=2.99
r79 27 29 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.645 $Y=2.905
+ $X2=3.645 $Y2=2.815
r80 26 52 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=1.99
+ $X2=3.645 $Y2=1.905
r81 26 29 38.0306 $w=2.48e-07 $l=8.25e-07 $layer=LI1_cond $X=3.645 $Y=1.99
+ $X2=3.645 $Y2=2.815
r82 25 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.905
+ $X2=2.785 $Y2=1.905
r83 24 52 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.52 $Y=1.905
+ $X2=3.645 $Y2=1.905
r84 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.52 $Y=1.905
+ $X2=2.87 $Y2=1.905
r85 20 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=2.57
+ $X2=2.785 $Y2=2.485
r86 20 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.785 $Y=2.57
+ $X2=2.785 $Y2=2.815
r87 19 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=2.4
+ $X2=2.785 $Y2=2.485
r88 18 49 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.99
+ $X2=2.785 $Y2=1.905
r89 18 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.785 $Y=1.99
+ $X2=2.785 $Y2=2.4
r90 17 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=2.485
+ $X2=1.885 $Y2=2.485
r91 16 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=2.485
+ $X2=2.785 $Y2=2.485
r92 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.7 $Y=2.485
+ $X2=1.97 $Y2=2.485
r93 5 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.84 $X2=5.485 $Y2=2.815
r94 5 40 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.84 $X2=5.485 $Y2=1.985
r95 4 34 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=4.45
+ $Y=1.84 $X2=4.585 $Y2=2.325
r96 3 52 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.84 $X2=3.685 $Y2=1.985
r97 3 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.84 $X2=3.685 $Y2=2.815
r98 2 49 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.65
+ $Y=1.84 $X2=2.785 $Y2=1.985
r99 2 22 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.84 $X2=2.785 $Y2=2.815
r100 1 46 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.84 $X2=1.885 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%Z 1 2 3 4 13 15 19 21 23 24 27 30 33 34 35
+ 41
c67 24 0 6.7572e-20 $X=4.345 $Y=1.065
c68 19 0 1.41838e-19 $X=4.18 $Y=0.82
c69 13 0 6.07806e-20 $X=4.135 $Y=1.99
r70 39 41 1.54806 $w=3.33e-07 $l=4.5e-08 $layer=LI1_cond $X=5.037 $Y=1.99
+ $X2=5.037 $Y2=2.035
r71 35 46 8.42831 $w=3.33e-07 $l=2.45e-07 $layer=LI1_cond $X=5.037 $Y=2.405
+ $X2=5.037 $Y2=2.65
r72 34 39 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=5.037 $Y=1.905
+ $X2=5.037 $Y2=1.99
r73 34 35 12.0404 $w=3.33e-07 $l=3.5e-07 $layer=LI1_cond $X=5.037 $Y=2.055
+ $X2=5.037 $Y2=2.405
r74 34 41 0.688026 $w=3.33e-07 $l=2e-08 $layer=LI1_cond $X=5.037 $Y=2.055
+ $X2=5.037 $Y2=2.035
r75 30 34 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=5.12 $Y=1.82
+ $X2=5.037 $Y2=1.905
r76 29 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.12 $Y=1.15
+ $X2=5.04 $Y2=1.065
r77 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.12 $Y=1.15
+ $X2=5.12 $Y2=1.82
r78 25 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0.98 $X2=5.04
+ $Y2=1.065
r79 25 27 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=0.98 $X2=5.04
+ $Y2=0.86
r80 23 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=1.065
+ $X2=5.04 $Y2=1.065
r81 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.875 $Y=1.065
+ $X2=4.345 $Y2=1.065
r82 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=1.905
+ $X2=4.135 $Y2=1.905
r83 21 34 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.87 $Y=1.905
+ $X2=5.037 $Y2=1.905
r84 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.87 $Y=1.905
+ $X2=4.3 $Y2=1.905
r85 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.18 $Y=0.98
+ $X2=4.345 $Y2=1.065
r86 17 19 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.18 $Y=0.98 $X2=4.18
+ $Y2=0.82
r87 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=1.99
+ $X2=4.135 $Y2=1.905
r88 13 15 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=4.135 $Y=1.99
+ $X2=4.135 $Y2=2.65
r89 4 34 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=4.9
+ $Y=1.84 $X2=5.035 $Y2=1.97
r90 4 46 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=4.9 $Y=1.84
+ $X2=5.035 $Y2=2.65
r91 3 32 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=4 $Y=1.84
+ $X2=4.135 $Y2=1.97
r92 3 15 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=4 $Y=1.84
+ $X2=4.135 $Y2=2.65
r93 2 27 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=4.9
+ $Y=0.37 $X2=5.04 $Y2=0.86
r94 1 19 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.37 $X2=4.18 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%VGND 1 2 3 12 16 20 23 24 26 27 28 30 49 50
+ 53
r72 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r73 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r74 47 50 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=5.52
+ $Y2=0
r75 46 49 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.52
+ $Y2=0
r76 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r77 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r78 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r79 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r80 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r81 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r82 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r83 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r84 35 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r85 35 37 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r86 33 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r87 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r88 30 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r89 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r90 28 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.12
+ $Y2=0
r91 28 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r92 26 43 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.12
+ $Y2=0
r93 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.28
+ $Y2=0
r94 25 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.6
+ $Y2=0
r95 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.28
+ $Y2=0
r96 23 40 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.16
+ $Y2=0
r97 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.46
+ $Y2=0
r98 22 43 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=3.12
+ $Y2=0
r99 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.46
+ $Y2=0
r100 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0
r101 18 20 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0.645
r102 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r103 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.515
r104 10 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r105 10 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.495
r106 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.37 $X2=3.32 $Y2=0.645
r107 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.32
+ $Y=0.37 $X2=2.46 $Y2=0.515
r108 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.61
+ $Y=0.37 $X2=0.75 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__EBUFN_4%A_378_74# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 42 44 47
c81 44 0 2.52699e-19 $X=2.89 $Y=1.065
c82 33 0 1.27021e-19 $X=3.835 $Y=0.34
r83 44 45 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.89 $Y=1.065
+ $X2=2.89 $Y2=1.225
r84 40 42 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.53 $Y=0.425 $X2=5.53
+ $Y2=0.515
r85 39 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=0.34
+ $X2=4.61 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.405 $Y=0.34
+ $X2=5.53 $Y2=0.425
r87 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.405 $Y=0.34
+ $X2=4.695 $Y2=0.34
r88 34 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=0.425
+ $X2=4.61 $Y2=0.34
r89 34 36 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.61 $Y=0.425
+ $X2=4.61 $Y2=0.58
r90 32 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=0.34
+ $X2=4.61 $Y2=0.34
r91 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.525 $Y=0.34
+ $X2=3.835 $Y2=0.34
r92 29 31 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=3.71 $Y=0.98
+ $X2=3.71 $Y2=0.515
r93 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.71 $Y=0.425
+ $X2=3.835 $Y2=0.34
r94 28 31 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.71 $Y=0.425 $X2=3.71
+ $Y2=0.515
r95 27 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=1.065
+ $X2=2.89 $Y2=1.065
r96 26 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.585 $Y=1.065
+ $X2=3.71 $Y2=0.98
r97 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.585 $Y=1.065
+ $X2=2.975 $Y2=1.065
r98 22 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=0.98
+ $X2=2.89 $Y2=1.065
r99 22 24 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.89 $Y=0.98
+ $X2=2.89 $Y2=0.515
r100 20 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=1.225
+ $X2=2.89 $Y2=1.225
r101 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.805 $Y=1.225
+ $X2=2.115 $Y2=1.225
r102 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.03 $Y=1.14
+ $X2=2.115 $Y2=1.225
r103 16 18 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.03 $Y=1.14
+ $X2=2.03 $Y2=0.515
r104 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.35
+ $Y=0.37 $X2=5.49 $Y2=0.515
r105 4 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.47
+ $Y=0.37 $X2=4.61 $Y2=0.58
r106 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.61
+ $Y=0.37 $X2=3.75 $Y2=0.515
r107 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.75
+ $Y=0.37 $X2=2.89 $Y2=0.515
r108 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.89
+ $Y=0.37 $X2=2.03 $Y2=0.515
.ends


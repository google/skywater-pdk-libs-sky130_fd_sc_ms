* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ms__sedfxbp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
*.PININFO CLK:I D:I DE:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I Q:O
*.PININFO Q_N:O
MI14 net86 M1 VPB pshort m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI637 clkpos clkneg VPB pshort m=1 w=1.12 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI13 S0 clkneg VPB pshort m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI651 db clkpos VPB pshort m=1 w=0.42 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI645 Q S0 VPB pshort m=1 w=1.12 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net122 M1 VPB pshort m=1 w=0.42 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI638 clkneg CLK VPB pshort m=1 w=1.12 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI643 net114 q1 VPB pshort m=1 w=0.42 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI639 M1 M0 VPB pshort m=1 w=0.84 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI644 S0 clkpos VPB pshort m=1 w=0.42 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q_N q1 VPB pshort m=1 w=1.12 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI659 M0 clkneg VPB pshort m=1 w=0.42 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI17 q1 S0 VPB pshort m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net131 deneg VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI47 net138 sceneg VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI46 VPWR SCD VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI31 net143 D VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI42 net143 SCE VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI40 net158 q1 VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI36 deneg DE VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI38 VPWR DE VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI44 sceneg SCE VPB pshort m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI634 M1 M0 VNB nlowvt m=1 w=0.64 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkpos clkneg VNB nlowvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg CLK VNB nlowvt m=1 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI661 Q_N q1 VNB nlowvt m=1 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI641 net186 q1 VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI642 S0 clkneg VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI648 db clkneg VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI646 Q S0 VNB nlowvt m=1 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net199 M1 VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI657 M0 clkpos VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI43 net143 sceneg VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI18 q1 S0 VNB nlowvt m=1 w=0.64 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI45 sceneg SCE VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI32 net143 D VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI16 net223 M1 VNB nlowvt m=1 w=0.64 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI15 S0 clkpos VNB nlowvt m=1 w=0.64 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI41 net231 q1 VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI39 VGND deneg VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI37 deneg DE VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net218 DE VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI49 net247 SCE VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI48 VGND SCD VNB nlowvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ms__sedfxbp_1

* File: sky130_fd_sc_ms__nand2_8.spice
* Created: Fri Aug 28 17:42:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand2_8.pex.spice"
.subckt sky130_fd_sc_ms__nand2_8  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_B_M1000_g N_A_27_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1000_d N_B_M1001_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75006.5 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1002_d N_B_M1010_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75006.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.222 AS=0.1036 PD=1.34 PS=1.02 NRD=25.944 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75005.6 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1011_d N_B_M1012_g N_A_27_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.222 AS=0.1184 PD=1.34 PS=1.06 NRD=25.944 NRS=3.24 M=1 R=4.93333
+ SA=75002.7 SB=75004.9 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_B_M1017_g N_A_27_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75003.1
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1017_d N_B_M1018_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1018_s N_A_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1004_d N_A_M1004_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.4
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1004_d N_A_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.9
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1008 N_A_27_74#_M1008_d N_A_M1008_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_27_74#_M1008_d N_A_M1013_g N_Y_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.7
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_A_M1014_g N_Y_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2368 AS=0.1036 PD=1.38 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.1
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1014_d N_A_M1019_g N_Y_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2368 AS=0.1036 PD=1.38 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.9
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_A_27_74#_M1023_d N_A_M1023_g N_Y_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19805 AS=0.1036 PD=2.07 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1016_d N_B_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12 AD=0.1792
+ AS=1.4784 PD=1.44 PS=4.88 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.2 SB=90002.9
+ A=0.2016 P=2.6 MULT=1
MM1020 N_Y_M1016_d N_B_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12 AD=0.1792
+ AS=0.8736 PD=1.44 PS=2.68 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.7 SB=90002.4
+ A=0.2016 P=2.6 MULT=1
MM1021 N_Y_M1021_d N_B_M1021_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.8736 PD=1.39 PS=2.68 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.5 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1022 N_Y_M1021_d N_B_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.9 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.3696
+ AS=0.1792 PD=2.9 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90002
+ A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_Y_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.364
+ AS=0.1792 PD=1.77 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7 SB=90001.5
+ A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1007_d N_A_M1009_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12 AD=0.364
+ AS=0.1512 PD=1.77 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12 AD=0.308
+ AS=0.1512 PD=2.79 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__nand2_8.pxi.spice"
*
.ends
*
*

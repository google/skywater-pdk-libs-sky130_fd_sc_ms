* File: sky130_fd_sc_ms__or3_1.pxi.spice
* Created: Wed Sep  2 12:28:11 2020
* 
x_PM_SKY130_FD_SC_MS__OR3_1%C N_C_c_51_n N_C_M1000_g N_C_M1007_g C N_C_c_53_n
+ PM_SKY130_FD_SC_MS__OR3_1%C
x_PM_SKY130_FD_SC_MS__OR3_1%B N_B_M1002_g N_B_M1003_g B N_B_c_80_n
+ PM_SKY130_FD_SC_MS__OR3_1%B
x_PM_SKY130_FD_SC_MS__OR3_1%A N_A_M1006_g N_A_M1001_g A N_A_c_112_n N_A_c_113_n
+ PM_SKY130_FD_SC_MS__OR3_1%A
x_PM_SKY130_FD_SC_MS__OR3_1%A_27_74# N_A_27_74#_M1007_s N_A_27_74#_M1003_d
+ N_A_27_74#_M1000_s N_A_27_74#_M1004_g N_A_27_74#_M1005_g N_A_27_74#_c_149_n
+ N_A_27_74#_c_150_n N_A_27_74#_c_163_n N_A_27_74#_c_151_n N_A_27_74#_c_152_n
+ N_A_27_74#_c_153_n N_A_27_74#_c_159_n N_A_27_74#_c_154_n N_A_27_74#_c_155_n
+ N_A_27_74#_c_156_n PM_SKY130_FD_SC_MS__OR3_1%A_27_74#
x_PM_SKY130_FD_SC_MS__OR3_1%VPWR N_VPWR_M1006_d N_VPWR_c_237_n VPWR
+ N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_236_n N_VPWR_c_241_n
+ PM_SKY130_FD_SC_MS__OR3_1%VPWR
x_PM_SKY130_FD_SC_MS__OR3_1%X N_X_M1005_d N_X_M1004_d N_X_c_266_n N_X_c_267_n
+ N_X_c_263_n X X X PM_SKY130_FD_SC_MS__OR3_1%X
x_PM_SKY130_FD_SC_MS__OR3_1%VGND N_VGND_M1007_d N_VGND_M1001_d N_VGND_c_287_n
+ N_VGND_c_288_n VGND N_VGND_c_289_n N_VGND_c_290_n N_VGND_c_291_n
+ N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n PM_SKY130_FD_SC_MS__OR3_1%VGND
cc_1 VNB N_C_c_51_n 0.0279743f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.77
cc_2 VNB N_C_M1007_g 0.0444924f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_3 VNB N_C_c_53_n 0.0153111f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_4 VNB N_B_M1003_g 0.0402646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB B 0.00552308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B_c_80_n 0.0228865f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_7 VNB N_A_M1001_g 0.0411168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_112_n 0.00231998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_113_n 0.0363227f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_10 VNB N_A_27_74#_M1004_g 0.00187093f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.515
cc_11 VNB N_A_27_74#_M1005_g 0.0287882f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_12 VNB N_A_27_74#_c_149_n 0.0277943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_150_n 0.00992268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_151_n 0.00979143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_152_n 0.00746217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_153_n 4.2489e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_154_n 0.0157854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_155_n 0.0109349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_156_n 0.0336134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_236_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_263_n 0.0247379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB X 0.0267037f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.565
cc_23 VNB X 0.0139384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_287_n 0.00651905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_288_n 0.00981015f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_26 VNB N_VGND_c_289_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_290_n 0.028973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_291_n 0.0190372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_292_n 0.186353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_293_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_294_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_C_c_51_n 0.0345756f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.77
cc_33 VPB N_C_c_53_n 0.00745261f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_34 VPB N_B_M1002_g 0.0212032f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_35 VPB B 0.00437076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_B_c_80_n 0.00547205f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_37 VPB N_A_M1006_g 0.0244947f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_38 VPB N_A_c_112_n 0.00297478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_c_113_n 0.0103796f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.565
cc_40 VPB N_A_27_74#_M1004_g 0.031627f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.515
cc_41 VPB N_A_27_74#_c_153_n 0.00334823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_27_74#_c_159_n 0.0388119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_237_n 0.0142325f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_44 VPB N_VPWR_c_238_n 0.0496025f $X=-0.19 $Y=1.66 $X2=0.417 $Y2=1.515
cc_45 VPB N_VPWR_c_239_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_236_n 0.0860025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_241_n 0.0143983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_X_c_266_n 0.0101022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_X_c_267_n 0.0417369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_X_c_263_n 0.00756894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 N_C_c_51_n N_B_M1002_g 0.0720051f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_52 N_C_M1007_g N_B_M1003_g 0.0293272f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_53 N_C_c_51_n B 7.49167e-19 $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_54 N_C_c_53_n B 0.0238235f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_55 N_C_c_51_n N_B_c_80_n 0.0160621f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_56 N_C_c_53_n N_B_c_80_n 4.21721e-19 $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_57 N_C_M1007_g N_A_27_74#_c_149_n 0.00712316f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_58 N_C_c_51_n N_A_27_74#_c_150_n 0.00291196f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_59 N_C_c_53_n N_A_27_74#_c_150_n 0.0211058f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_60 N_C_c_51_n N_A_27_74#_c_163_n 0.0133533f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_61 N_C_c_53_n N_A_27_74#_c_163_n 0.00908651f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_62 N_C_c_51_n N_A_27_74#_c_159_n 0.0201358f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_63 N_C_c_53_n N_A_27_74#_c_159_n 0.025494f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_64 N_C_c_51_n N_A_27_74#_c_154_n 0.00198478f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_65 N_C_M1007_g N_A_27_74#_c_154_n 0.0160891f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_66 N_C_c_53_n N_A_27_74#_c_154_n 0.0151257f $X=0.405 $Y=1.515 $X2=0 $Y2=0
cc_67 N_C_M1007_g N_A_27_74#_c_155_n 8.67149e-19 $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_68 N_C_c_51_n N_VPWR_c_238_n 0.00567889f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_69 N_C_c_51_n N_VPWR_c_236_n 0.00610055f $X=0.505 $Y=1.77 $X2=0 $Y2=0
cc_70 N_C_M1007_g N_VGND_c_287_n 0.0130729f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_71 N_C_M1007_g N_VGND_c_289_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_72 N_C_M1007_g N_VGND_c_292_n 0.00761198f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_73 N_B_M1002_g N_A_M1006_g 0.0434391f $X=0.925 $Y=2.34 $X2=0 $Y2=0
cc_74 N_B_M1003_g N_A_M1001_g 0.0120173f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_75 B N_A_c_112_n 0.0350348f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_76 N_B_c_80_n N_A_c_112_n 2.7993e-19 $X=1 $Y=1.515 $X2=0 $Y2=0
cc_77 B N_A_c_113_n 0.00340053f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_78 N_B_c_80_n N_A_c_113_n 0.0176805f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B_M1002_g N_A_27_74#_c_163_n 0.0175218f $X=0.925 $Y=2.34 $X2=0 $Y2=0
cc_80 B N_A_27_74#_c_163_n 0.0349587f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_81 N_B_c_80_n N_A_27_74#_c_163_n 7.11116e-19 $X=1 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B_M1002_g N_A_27_74#_c_159_n 0.00355274f $X=0.925 $Y=2.34 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_A_27_74#_c_154_n 0.0114826f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_84 B N_A_27_74#_c_154_n 0.0392242f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_85 N_B_c_80_n N_A_27_74#_c_154_n 0.00224064f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B_M1003_g N_A_27_74#_c_155_n 0.0163295f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_87 N_B_c_80_n N_A_27_74#_c_155_n 0.00221201f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B_M1002_g N_VPWR_c_237_n 0.00306046f $X=0.925 $Y=2.34 $X2=0 $Y2=0
cc_89 N_B_M1002_g N_VPWR_c_238_n 0.0059286f $X=0.925 $Y=2.34 $X2=0 $Y2=0
cc_90 N_B_M1002_g N_VPWR_c_236_n 0.00610055f $X=0.925 $Y=2.34 $X2=0 $Y2=0
cc_91 N_B_M1003_g N_VGND_c_287_n 0.00593102f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_92 N_B_M1003_g N_VGND_c_290_n 0.00435437f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_VGND_c_292_n 0.0082237f $X=0.995 $Y=0.645 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_A_27_74#_M1004_g 0.00635048f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_95 N_A_c_113_n N_A_27_74#_M1004_g 0.00116328f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_M1001_g N_A_27_74#_M1005_g 0.0220159f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_97 N_A_M1006_g N_A_27_74#_c_163_n 0.0206941f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_98 N_A_c_112_n N_A_27_74#_c_163_n 0.0235064f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A_c_113_n N_A_27_74#_c_163_n 0.00378607f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_M1001_g N_A_27_74#_c_151_n 0.0135443f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_101 N_A_M1001_g N_A_27_74#_c_152_n 0.00572869f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_102 N_A_c_112_n N_A_27_74#_c_152_n 0.0156671f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A_M1006_g N_A_27_74#_c_153_n 0.00304023f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_104 N_A_c_112_n N_A_27_74#_c_153_n 0.00827244f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A_c_113_n N_A_27_74#_c_153_n 4.33638e-19 $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A_M1001_g N_A_27_74#_c_155_n 0.0162445f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_107 N_A_c_112_n N_A_27_74#_c_155_n 0.0273553f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_c_113_n N_A_27_74#_c_155_n 0.0058749f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A_M1001_g N_A_27_74#_c_156_n 0.0177468f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_110 N_A_c_112_n N_A_27_74#_c_156_n 3.03321e-19 $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A_M1006_g N_VPWR_c_237_n 0.0190349f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_112 N_A_M1006_g N_VPWR_c_238_n 0.00492916f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_113 N_A_M1006_g N_VPWR_c_236_n 0.00511769f $X=1.495 $Y=2.34 $X2=0 $Y2=0
cc_114 N_A_M1001_g X 7.18714e-19 $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_VGND_c_288_n 0.00642087f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_116 N_A_M1001_g N_VGND_c_290_n 0.00435437f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_117 N_A_M1001_g N_VGND_c_292_n 0.0082291f $X=1.81 $Y=0.645 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_163_n A_119_368# 0.0096152f $X=2.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_27_74#_c_163_n A_203_368# 0.0144757f $X=2.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_27_74#_c_163_n N_VPWR_M1006_d 0.0206763f $X=2.09 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_27_74#_c_153_n N_VPWR_M1006_d 0.00251301f $X=2.175 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_27_74#_M1004_g N_VPWR_c_237_n 0.0193868f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_163_n N_VPWR_c_237_n 0.0509764f $X=2.09 $Y=2.035 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_152_n N_VPWR_c_237_n 0.00103513f $X=2.175 $Y=1.63 $X2=0
+ $Y2=0
cc_125 N_A_27_74#_c_156_n N_VPWR_c_237_n 3.65473e-19 $X=2.29 $Y=1.465 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_c_159_n N_VPWR_c_238_n 0.00975961f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_127 N_A_27_74#_M1004_g N_VPWR_c_239_n 0.00460063f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_27_74#_M1004_g N_VPWR_c_236_n 0.00912296f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_159_n N_VPWR_c_236_n 0.0111753f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_130 N_A_27_74#_M1004_g N_X_c_266_n 0.00196268f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A_27_74#_c_153_n N_X_c_266_n 0.00111918f $X=2.175 $Y=1.95 $X2=0 $Y2=0
cc_132 N_A_27_74#_M1005_g N_X_c_263_n 0.0025312f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_27_74#_c_152_n N_X_c_263_n 0.0304389f $X=2.175 $Y=1.63 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_153_n N_X_c_263_n 0.0061697f $X=2.175 $Y=1.95 $X2=0 $Y2=0
cc_135 N_A_27_74#_c_156_n N_X_c_263_n 0.0106236f $X=2.29 $Y=1.465 $X2=0 $Y2=0
cc_136 N_A_27_74#_M1005_g X 0.00941145f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_27_74#_c_155_n X 0.0050994f $X=1.76 $Y=0.817 $X2=0 $Y2=0
cc_138 N_A_27_74#_M1005_g X 0.0032303f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_27_74#_c_152_n X 0.00740597f $X=2.175 $Y=1.63 $X2=0 $Y2=0
cc_140 N_A_27_74#_c_156_n X 4.83855e-19 $X=2.29 $Y=1.465 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_151_n N_VGND_M1001_d 5.19034e-19 $X=2.09 $Y=1.095 $X2=0
+ $Y2=0
cc_142 N_A_27_74#_c_152_n N_VGND_M1001_d 0.00275048f $X=2.175 $Y=1.63 $X2=0
+ $Y2=0
cc_143 N_A_27_74#_c_149_n N_VGND_c_287_n 0.017215f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_144 N_A_27_74#_c_154_n N_VGND_c_287_n 0.0211984f $X=1.045 $Y=0.817 $X2=0
+ $Y2=0
cc_145 N_A_27_74#_M1005_g N_VGND_c_288_n 0.00604382f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_27_74#_c_151_n N_VGND_c_288_n 0.0111634f $X=2.09 $Y=1.095 $X2=0 $Y2=0
cc_147 N_A_27_74#_c_152_n N_VGND_c_288_n 0.0126115f $X=2.175 $Y=1.63 $X2=0 $Y2=0
cc_148 N_A_27_74#_c_156_n N_VGND_c_288_n 5.51659e-19 $X=2.29 $Y=1.465 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_c_149_n N_VGND_c_289_n 0.011066f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_150 N_A_27_74#_c_155_n N_VGND_c_290_n 0.0198465f $X=1.76 $Y=0.817 $X2=0 $Y2=0
cc_151 N_A_27_74#_M1005_g N_VGND_c_291_n 0.00434272f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_27_74#_M1005_g N_VGND_c_292_n 0.00824987f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_27_74#_c_149_n N_VGND_c_292_n 0.00915947f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_154 N_A_27_74#_c_155_n N_VGND_c_292_n 0.0243841f $X=1.76 $Y=0.817 $X2=0 $Y2=0
cc_155 N_VPWR_c_237_n N_X_c_267_n 0.0260873f $X=2.15 $Y=2.375 $X2=0 $Y2=0
cc_156 N_VPWR_c_239_n N_X_c_267_n 0.0124046f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_c_236_n N_X_c_267_n 0.0102675f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_158 X N_VGND_c_288_n 0.0183192f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_159 X N_VGND_c_291_n 0.0161257f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_160 X N_VGND_c_292_n 0.013291f $X=2.555 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__xor2_1.spice
* Created: Fri Aug 28 18:18:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xor2_1.pex.spice"
.subckt sky130_fd_sc_ms__xor2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1008 N_A_194_125#_M1008_d N_A_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.177375 AS=0.33275 PD=1.195 PS=2.31 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.5
+ SB=75002.6 A=0.0825 P=1.4 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_194_125#_M1008_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.107506 AS=0.177375 PD=0.937984 PS=1.195 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75001.3 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1004 A_455_87# N_A_M1004_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.144644 PD=0.98 PS=1.26202 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_B_M1005_g A_455_87# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75001.8 SB=75000.9
+ A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_194_125#_M1009_g N_X_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2997 AS=0.1554 PD=2.29 PS=1.16 NRD=0 NRS=22.692 M=1 R=4.93333 SA=75002.4
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 A_161_392# N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90000.6
+ A=0.18 P=2.36 MULT=1
MM1001 N_A_194_125#_M1001_d N_B_M1001_g A_161_392# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90000.2
+ A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_355_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2184 AS=0.3584 PD=1.51 PS=2.88 NRD=10.5395 NRS=6.1464 M=1 R=6.22222
+ SA=90000.2 SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1006 N_A_355_368#_M1006_d N_B_M1006_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2184 PD=1.44 PS=1.51 NRD=7.8997 NRS=8.7862 M=1 R=6.22222
+ SA=90000.8 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1007_d N_A_194_125#_M1007_g N_A_355_368#_M1006_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3696 AS=0.1792 PD=2.9 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90001.3 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__xor2_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o311ai_4.pxi.spice
* Created: Wed Sep  2 12:25:22 2020
* 
x_PM_SKY130_FD_SC_MS__O311AI_4%C1 N_C1_M1010_g N_C1_c_149_n N_C1_M1005_g
+ N_C1_c_150_n N_C1_M1019_g N_C1_M1021_g N_C1_c_152_n N_C1_M1020_g N_C1_c_153_n
+ N_C1_c_154_n N_C1_c_155_n N_C1_M1032_g C1 C1 N_C1_c_156_n
+ PM_SKY130_FD_SC_MS__O311AI_4%C1
x_PM_SKY130_FD_SC_MS__O311AI_4%B1 N_B1_c_224_n N_B1_M1022_g N_B1_c_216_n
+ N_B1_c_217_n N_B1_c_227_n N_B1_M1023_g N_B1_M1003_g N_B1_M1016_g N_B1_M1017_g
+ N_B1_M1031_g B1 B1 B1 B1 N_B1_c_223_n PM_SKY130_FD_SC_MS__O311AI_4%B1
x_PM_SKY130_FD_SC_MS__O311AI_4%A3 N_A3_M1000_g N_A3_M1011_g N_A3_M1012_g
+ N_A3_M1013_g N_A3_M1025_g N_A3_M1027_g N_A3_M1034_g N_A3_M1035_g A3 A3
+ N_A3_c_289_n N_A3_c_283_n N_A3_c_291_n N_A3_c_284_n A3
+ PM_SKY130_FD_SC_MS__O311AI_4%A3
x_PM_SKY130_FD_SC_MS__O311AI_4%A2 N_A2_M1024_g N_A2_M1004_g N_A2_M1026_g
+ N_A2_M1006_g N_A2_M1028_g N_A2_c_379_n N_A2_M1018_g N_A2_M1030_g N_A2_c_381_n
+ N_A2_M1029_g A2 A2 N_A2_c_387_n N_A2_c_382_n PM_SKY130_FD_SC_MS__O311AI_4%A2
x_PM_SKY130_FD_SC_MS__O311AI_4%A1 N_A1_M1001_g N_A1_c_471_n N_A1_c_472_n
+ N_A1_M1002_g N_A1_M1008_g N_A1_M1009_g N_A1_M1014_g N_A1_c_474_n N_A1_M1007_g
+ N_A1_M1033_g N_A1_c_475_n N_A1_M1015_g A1 A1 A1 N_A1_c_483_n N_A1_c_476_n
+ PM_SKY130_FD_SC_MS__O311AI_4%A1
x_PM_SKY130_FD_SC_MS__O311AI_4%VPWR N_VPWR_M1010_s N_VPWR_M1021_s N_VPWR_M1023_s
+ N_VPWR_M1008_s N_VPWR_M1009_s N_VPWR_M1033_s N_VPWR_c_553_n N_VPWR_c_554_n
+ N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n
+ N_VPWR_c_560_n N_VPWR_c_561_n VPWR N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n
+ N_VPWR_c_552_n PM_SKY130_FD_SC_MS__O311AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O311AI_4%Y N_Y_M1005_d N_Y_M1020_d N_Y_M1010_d N_Y_M1022_d
+ N_Y_M1000_d N_Y_M1025_d N_Y_c_673_n N_Y_c_667_n N_Y_c_678_n N_Y_c_664_n
+ N_Y_c_668_n N_Y_c_669_n N_Y_c_723_n N_Y_c_725_n N_Y_c_730_n N_Y_c_685_n
+ N_Y_c_690_n N_Y_c_670_n N_Y_c_671_n N_Y_c_737_n Y Y N_Y_c_665_n Y
+ PM_SKY130_FD_SC_MS__O311AI_4%Y
x_PM_SKY130_FD_SC_MS__O311AI_4%A_841_368# N_A_841_368#_M1000_s
+ N_A_841_368#_M1012_s N_A_841_368#_M1034_s N_A_841_368#_M1026_s
+ N_A_841_368#_M1030_s N_A_841_368#_c_800_n N_A_841_368#_c_801_n
+ N_A_841_368#_c_802_n N_A_841_368#_c_815_n N_A_841_368#_c_803_n
+ N_A_841_368#_c_819_n N_A_841_368#_c_804_n N_A_841_368#_c_869_p
+ N_A_841_368#_c_805_n N_A_841_368#_c_806_n N_A_841_368#_c_807_n
+ N_A_841_368#_c_808_n N_A_841_368#_c_809_n
+ PM_SKY130_FD_SC_MS__O311AI_4%A_841_368#
x_PM_SKY130_FD_SC_MS__O311AI_4%A_1353_368# N_A_1353_368#_M1024_d
+ N_A_1353_368#_M1028_d N_A_1353_368#_M1008_d N_A_1353_368#_M1014_d
+ N_A_1353_368#_c_877_n N_A_1353_368#_c_881_n N_A_1353_368#_c_874_n
+ N_A_1353_368#_c_875_n N_A_1353_368#_c_895_n N_A_1353_368#_c_899_n
+ N_A_1353_368#_c_876_n N_A_1353_368#_c_884_n N_A_1353_368#_c_888_n
+ N_A_1353_368#_c_904_n PM_SKY130_FD_SC_MS__O311AI_4%A_1353_368#
x_PM_SKY130_FD_SC_MS__O311AI_4%A_27_74# N_A_27_74#_M1005_s N_A_27_74#_M1019_s
+ N_A_27_74#_M1032_s N_A_27_74#_M1016_s N_A_27_74#_M1031_s N_A_27_74#_c_929_n
+ N_A_27_74#_c_930_n N_A_27_74#_c_931_n N_A_27_74#_c_954_n N_A_27_74#_c_932_n
+ PM_SKY130_FD_SC_MS__O311AI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O311AI_4%A_459_74# N_A_459_74#_M1003_d N_A_459_74#_M1017_d
+ N_A_459_74#_M1011_s N_A_459_74#_M1027_s N_A_459_74#_M1004_s
+ N_A_459_74#_M1018_s N_A_459_74#_M1001_s N_A_459_74#_M1007_s
+ N_A_459_74#_c_969_n N_A_459_74#_c_970_n N_A_459_74#_c_971_n
+ N_A_459_74#_c_972_n N_A_459_74#_c_973_n N_A_459_74#_c_997_n
+ N_A_459_74#_c_974_n N_A_459_74#_c_1002_n N_A_459_74#_c_975_n
+ N_A_459_74#_c_976_n N_A_459_74#_c_977_n N_A_459_74#_c_978_n
+ N_A_459_74#_c_979_n N_A_459_74#_c_980_n N_A_459_74#_c_981_n
+ N_A_459_74#_c_982_n N_A_459_74#_c_1004_n N_A_459_74#_c_1005_n
+ N_A_459_74#_c_983_n N_A_459_74#_c_984_n N_A_459_74#_c_1045_n
+ PM_SKY130_FD_SC_MS__O311AI_4%A_459_74#
x_PM_SKY130_FD_SC_MS__O311AI_4%VGND N_VGND_M1011_d N_VGND_M1013_d N_VGND_M1035_d
+ N_VGND_M1006_d N_VGND_M1029_d N_VGND_M1002_d N_VGND_M1015_d N_VGND_c_1118_n
+ N_VGND_c_1119_n N_VGND_c_1120_n N_VGND_c_1121_n N_VGND_c_1122_n
+ N_VGND_c_1123_n N_VGND_c_1124_n VGND N_VGND_c_1125_n N_VGND_c_1126_n
+ N_VGND_c_1127_n N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n
+ N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n
+ N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n
+ PM_SKY130_FD_SC_MS__O311AI_4%VGND
cc_1 VNB N_C1_M1010_g 0.00196751f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_C1_c_149_n 0.0204707f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_3 VNB N_C1_c_150_n 0.0152712f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_4 VNB N_C1_M1021_g 0.00173962f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=2.4
cc_5 VNB N_C1_c_152_n 0.0149102f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_6 VNB N_C1_c_153_n 0.0223569f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.26
cc_7 VNB N_C1_c_154_n 0.112274f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.26
cc_8 VNB N_C1_c_155_n 0.0147616f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.185
cc_9 VNB N_C1_c_156_n 0.0156012f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_10 VNB N_B1_c_216_n 0.00879774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_217_n 0.00674136f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_12 VNB N_B1_M1003_g 0.023123f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.63
cc_13 VNB N_B1_M1016_g 0.0221713f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_14 VNB N_B1_M1017_g 0.0223226f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.26
cc_15 VNB N_B1_M1031_g 0.0304926f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB B1 0.0110294f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_17 VNB N_B1_c_223_n 0.0824487f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.54
cc_18 VNB N_A3_M1011_g 0.0287422f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_19 VNB N_A3_M1013_g 0.0244469f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_20 VNB N_A3_M1027_g 0.0244287f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A3_M1035_g 0.0247143f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.407
cc_22 VNB N_A3_c_283_n 0.094389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A3_c_284_n 0.0023959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_M1004_g 0.0258894f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_A2_M1006_g 0.0230723f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_26 VNB N_A2_c_379_n 0.016486f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=0.74
cc_27 VNB N_A2_M1030_g 0.00108962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_c_381_n 0.0161012f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_29 VNB N_A2_c_382_n 0.100719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_M1001_g 0.0315883f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_31 VNB N_A1_c_471_n 0.00596486f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_32 VNB N_A1_c_472_n 0.00495433f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_33 VNB N_A1_M1002_g 0.0316257f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_34 VNB N_A1_c_474_n 0.0189372f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_A1_c_475_n 0.0198259f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.407
cc_36 VNB N_A1_c_476_n 0.118955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_552_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_664_n 0.0471346f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_39 VNB N_Y_c_665_n 0.00164207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB Y 0.00406123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_929_n 0.012589f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=0.74
cc_42 VNB N_A_27_74#_c_930_n 0.0218403f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.26
cc_43 VNB N_A_27_74#_c_931_n 0.00963967f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.185
cc_44 VNB N_A_27_74#_c_932_n 0.00205354f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.407
cc_45 VNB N_A_459_74#_c_969_n 0.0207409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_459_74#_c_970_n 0.00525772f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.407
cc_47 VNB N_A_459_74#_c_971_n 0.00638704f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.407
cc_48 VNB N_A_459_74#_c_972_n 0.00387414f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.465
cc_49 VNB N_A_459_74#_c_973_n 0.00206045f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_50 VNB N_A_459_74#_c_974_n 0.00239415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_459_74#_c_975_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_459_74#_c_976_n 0.00672511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_459_74#_c_977_n 0.00181921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_459_74#_c_978_n 0.012969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_459_74#_c_979_n 0.00206647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_459_74#_c_980_n 0.00159982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_459_74#_c_981_n 0.0106354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_459_74#_c_982_n 0.00220643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_459_74#_c_983_n 0.00190558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_459_74#_c_984_n 0.0010144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1118_n 0.0105224f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_62 VNB N_VGND_c_1119_n 0.00794664f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_63 VNB N_VGND_c_1120_n 0.00801909f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.407
cc_64 VNB N_VGND_c_1121_n 0.00512538f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.407
cc_65 VNB N_VGND_c_1122_n 0.00647008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1123_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_67 VNB N_VGND_c_1124_n 0.0505272f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=1.54
cc_68 VNB N_VGND_c_1125_n 0.109865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1126_n 0.0159624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1127_n 0.0180412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1128_n 0.0166074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1129_n 0.0189911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1130_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1131_n 0.00613127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1132_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1133_n 0.00651315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1134_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1135_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1136_n 0.0172515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1137_n 0.0262931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1138_n 0.564514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VPB N_C1_M1010_g 0.0290335f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_83 VPB N_C1_M1021_g 0.0246651f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=2.4
cc_84 VPB N_C1_c_156_n 0.0164782f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.465
cc_85 VPB N_B1_c_224_n 0.0196927f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_86 VPB N_B1_c_216_n 0.00378507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_B1_c_217_n 0.00263664f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_88 VPB N_B1_c_227_n 0.0216538f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_89 VPB B1 0.0220548f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.465
cc_90 VPB N_B1_c_223_n 0.0517997f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.54
cc_91 VPB N_A3_M1000_g 0.0256846f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_92 VPB N_A3_M1012_g 0.0216932f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=1.63
cc_93 VPB N_A3_M1025_g 0.0222345f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.26
cc_94 VPB N_A3_M1034_g 0.0221222f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.407
cc_95 VPB N_A3_c_289_n 0.00417977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A3_c_283_n 0.0207182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A3_c_291_n 0.00402652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A2_M1024_g 0.0199866f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_99 VPB N_A2_M1026_g 0.0213141f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=1.63
cc_100 VPB N_A2_M1028_g 0.0211471f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.26
cc_101 VPB N_A2_M1030_g 0.0286155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A2_c_387_n 0.00701871f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.54
cc_103 VPB N_A2_c_382_n 0.0126329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A1_c_471_n 0.00794688f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_105 VPB N_A1_c_472_n 0.00495506f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_106 VPB N_A1_M1008_g 0.0272532f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=2.4
cc_107 VPB N_A1_M1009_g 0.0198927f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=0.74
cc_108 VPB N_A1_M1014_g 0.0198946f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=0.74
cc_109 VPB N_A1_M1033_g 0.0263926f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.465
cc_110 VPB N_A1_c_483_n 0.00851772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A1_c_476_n 0.0140247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_553_n 0.0119967f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.26
cc_113 VPB N_VPWR_c_554_n 0.0487491f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=0.74
cc_114 VPB N_VPWR_c_555_n 0.00565803f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.407
cc_115 VPB N_VPWR_c_556_n 0.0113936f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.407
cc_116 VPB N_VPWR_c_557_n 0.00271781f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.465
cc_117 VPB N_VPWR_c_558_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.36 $Y2=1.185
cc_118 VPB N_VPWR_c_559_n 0.0639253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_560_n 0.0223565f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.54
cc_120 VPB N_VPWR_c_561_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_562_n 0.113124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_563_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_564_n 0.0182909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_565_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_566_n 0.0614384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_567_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_568_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_552_n 0.109272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_Y_c_667_n 0.00330473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_Y_c_668_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.407
cc_131 VPB N_Y_c_669_n 0.0148222f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.465
cc_132 VPB N_Y_c_670_n 0.00281502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_Y_c_671_n 0.00258192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB Y 0.00137865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_841_368#_c_800_n 0.00748204f $X=-0.19 $Y=1.66 $X2=1.715 $Y2=1.26
cc_136 VPB N_A_841_368#_c_801_n 0.00241371f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.185
cc_137 VPB N_A_841_368#_c_802_n 0.00466382f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=0.74
cc_138 VPB N_A_841_368#_c_803_n 0.00358353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_841_368#_c_804_n 0.00241371f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.407
cc_140 VPB N_A_841_368#_c_805_n 0.00618927f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_141 VPB N_A_841_368#_c_806_n 0.00524903f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_142 VPB N_A_841_368#_c_807_n 0.0023295f $X=-0.19 $Y=1.66 $X2=1.075 $Y2=1.54
cc_143 VPB N_A_841_368#_c_808_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_841_368#_c_809_n 0.00244483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1353_368#_c_874_n 0.0132311f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=0.74
cc_146 VPB N_A_1353_368#_c_875_n 0.00233077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1353_368#_c_876_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=1.407
cc_148 N_C1_M1021_g N_B1_c_224_n 0.0161135f $X=1.18 $Y=2.4 $X2=-0.19 $Y2=-0.245
cc_149 N_C1_c_153_n N_B1_c_217_n 0.0169735f $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_150 N_C1_c_154_n N_B1_c_217_n 0.0161135f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_151 N_C1_c_156_n N_B1_c_217_n 0.00133236f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_152 N_C1_c_155_n N_B1_M1003_g 0.0324285f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_153 N_C1_M1010_g N_VPWR_c_554_n 0.02101f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_154 N_C1_M1021_g N_VPWR_c_554_n 7.08416e-19 $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_155 N_C1_c_154_n N_VPWR_c_554_n 8.88842e-19 $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_156 N_C1_c_156_n N_VPWR_c_554_n 0.0256434f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_157 N_C1_M1010_g N_VPWR_c_555_n 5.89761e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_158 N_C1_M1021_g N_VPWR_c_555_n 0.0128732f $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_159 N_C1_M1010_g N_VPWR_c_560_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_160 N_C1_M1021_g N_VPWR_c_560_n 0.00460063f $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_161 N_C1_M1010_g N_VPWR_c_552_n 0.00910426f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_162 N_C1_M1021_g N_VPWR_c_552_n 0.00910426f $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_163 N_C1_M1010_g N_Y_c_673_n 0.00191215f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_164 N_C1_c_154_n N_Y_c_673_n 0.00142304f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_165 N_C1_c_156_n N_Y_c_673_n 0.027751f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_166 N_C1_M1010_g N_Y_c_667_n 0.00891715f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_167 N_C1_M1021_g N_Y_c_667_n 2.18333e-19 $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_168 N_C1_M1021_g N_Y_c_678_n 0.0153755f $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_169 N_C1_c_153_n N_Y_c_678_n 5.45325e-19 $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_170 N_C1_c_154_n N_Y_c_678_n 0.00681504f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_171 N_C1_c_156_n N_Y_c_678_n 0.0118912f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_172 N_C1_c_153_n N_Y_c_664_n 0.00350562f $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_173 N_C1_c_155_n N_Y_c_664_n 0.00520798f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_174 N_C1_M1021_g N_Y_c_668_n 6.27806e-19 $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_175 N_C1_c_149_n N_Y_c_685_n 0.00429752f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_176 N_C1_c_150_n N_Y_c_685_n 0.0128945f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_177 N_C1_c_152_n N_Y_c_685_n 0.0147571f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_178 N_C1_c_154_n N_Y_c_685_n 0.00593628f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_179 N_C1_c_156_n N_Y_c_685_n 0.0419281f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_180 N_C1_c_150_n N_Y_c_690_n 4.05917e-19 $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_181 N_C1_c_152_n N_Y_c_690_n 0.0036256f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_182 N_C1_c_153_n N_Y_c_690_n 0.0130927f $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_183 N_C1_c_154_n N_Y_c_690_n 0.00507672f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_184 N_C1_c_155_n N_Y_c_690_n 0.00632997f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_185 N_C1_M1021_g N_Y_c_670_n 6.08944e-19 $X=1.18 $Y=2.4 $X2=0 $Y2=0
cc_186 N_C1_c_153_n N_Y_c_670_n 7.60047e-19 $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_187 N_C1_c_149_n N_A_27_74#_c_930_n 0.00194058f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_188 N_C1_c_154_n N_A_27_74#_c_930_n 0.00381029f $X=1.435 $Y=1.26 $X2=0 $Y2=0
cc_189 N_C1_c_156_n N_A_27_74#_c_930_n 0.0211412f $X=1.075 $Y=1.465 $X2=0 $Y2=0
cc_190 N_C1_c_149_n N_A_27_74#_c_931_n 0.0144205f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_191 N_C1_c_150_n N_A_27_74#_c_931_n 0.0102631f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_192 N_C1_c_152_n N_A_27_74#_c_931_n 0.0101492f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_193 N_C1_c_153_n N_A_27_74#_c_931_n 3.14401e-19 $X=1.715 $Y=1.26 $X2=0 $Y2=0
cc_194 N_C1_c_155_n N_A_27_74#_c_931_n 0.0121821f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_195 N_C1_c_155_n N_A_459_74#_c_969_n 2.00992e-19 $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_196 N_C1_c_149_n N_VGND_c_1125_n 0.00291649f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_197 N_C1_c_150_n N_VGND_c_1125_n 0.00291649f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_198 N_C1_c_152_n N_VGND_c_1125_n 0.00291649f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_199 N_C1_c_155_n N_VGND_c_1125_n 0.00291649f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_200 N_C1_c_149_n N_VGND_c_1138_n 0.00362829f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_201 N_C1_c_150_n N_VGND_c_1138_n 0.00359171f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_202 N_C1_c_152_n N_VGND_c_1138_n 0.00359121f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_203 N_C1_c_155_n N_VGND_c_1138_n 0.00359219f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_204 B1 N_A3_c_283_n 0.00689953f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_205 B1 N_A3_c_284_n 0.0124194f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B1_c_224_n N_VPWR_c_555_n 0.00194871f $X=1.68 $Y=1.725 $X2=0 $Y2=0
cc_207 N_B1_c_224_n N_VPWR_c_565_n 0.005209f $X=1.68 $Y=1.725 $X2=0 $Y2=0
cc_208 N_B1_c_227_n N_VPWR_c_565_n 0.005209f $X=2.13 $Y=1.725 $X2=0 $Y2=0
cc_209 N_B1_c_227_n N_VPWR_c_566_n 0.00419671f $X=2.13 $Y=1.725 $X2=0 $Y2=0
cc_210 N_B1_c_224_n N_VPWR_c_552_n 0.0098216f $X=1.68 $Y=1.725 $X2=0 $Y2=0
cc_211 N_B1_c_227_n N_VPWR_c_552_n 0.00986704f $X=2.13 $Y=1.725 $X2=0 $Y2=0
cc_212 N_B1_c_224_n N_Y_c_678_n 0.0139775f $X=1.68 $Y=1.725 $X2=0 $Y2=0
cc_213 N_B1_c_216_n N_Y_c_664_n 0.00807475f $X=2.04 $Y=1.65 $X2=0 $Y2=0
cc_214 N_B1_M1003_g N_Y_c_664_n 0.013432f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B1_M1016_g N_Y_c_664_n 0.0104926f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B1_M1017_g N_Y_c_664_n 0.0105534f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B1_M1031_g N_Y_c_664_n 0.0125939f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_218 B1 N_Y_c_664_n 0.147849f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B1_c_223_n N_Y_c_664_n 0.00784304f $X=3.43 $Y=1.515 $X2=0 $Y2=0
cc_220 N_B1_c_224_n N_Y_c_668_n 0.0124012f $X=1.68 $Y=1.725 $X2=0 $Y2=0
cc_221 N_B1_c_227_n N_Y_c_668_n 0.0166663f $X=2.13 $Y=1.725 $X2=0 $Y2=0
cc_222 N_B1_c_227_n N_Y_c_669_n 0.0177271f $X=2.13 $Y=1.725 $X2=0 $Y2=0
cc_223 B1 N_Y_c_669_n 0.151962f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 N_B1_c_223_n N_Y_c_669_n 0.00805248f $X=3.43 $Y=1.515 $X2=0 $Y2=0
cc_225 N_B1_c_217_n N_Y_c_690_n 7.37935e-19 $X=1.77 $Y=1.65 $X2=0 $Y2=0
cc_226 N_B1_M1003_g N_Y_c_690_n 9.07448e-19 $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B1_c_224_n N_Y_c_670_n 0.00382687f $X=1.68 $Y=1.725 $X2=0 $Y2=0
cc_228 N_B1_c_216_n N_Y_c_670_n 0.00254734f $X=2.04 $Y=1.65 $X2=0 $Y2=0
cc_229 N_B1_c_227_n N_Y_c_670_n 0.00705031f $X=2.13 $Y=1.725 $X2=0 $Y2=0
cc_230 N_B1_M1003_g N_A_27_74#_c_931_n 4.56461e-19 $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B1_M1003_g N_A_27_74#_c_932_n 0.0106751f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B1_M1016_g N_A_27_74#_c_932_n 0.00838518f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B1_M1017_g N_A_27_74#_c_932_n 0.00849254f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B1_M1031_g N_A_27_74#_c_932_n 0.00849254f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B1_M1003_g N_A_459_74#_c_969_n 0.00375385f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B1_M1016_g N_A_459_74#_c_969_n 0.0103107f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B1_M1017_g N_A_459_74#_c_969_n 0.0103245f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_M1031_g N_A_459_74#_c_969_n 0.0131979f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_M1031_g N_A_459_74#_c_970_n 0.00284982f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1003_g N_VGND_c_1125_n 0.00329872f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B1_M1016_g N_VGND_c_1125_n 0.00288916f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B1_M1017_g N_VGND_c_1125_n 0.00288916f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_243 N_B1_M1031_g N_VGND_c_1125_n 0.00288916f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B1_M1003_g N_VGND_c_1138_n 0.00428036f $X=2.22 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B1_M1016_g N_VGND_c_1138_n 0.0035719f $X=2.65 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B1_M1017_g N_VGND_c_1138_n 0.0035729f $X=3.08 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B1_M1031_g N_VGND_c_1138_n 0.00362289f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A3_M1034_g N_A2_M1024_g 0.0238523f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A3_M1035_g N_A2_M1004_g 0.0234798f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A3_c_289_n N_A2_c_382_n 2.5456e-19 $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_251 N_A3_c_283_n N_A2_c_382_n 0.0238523f $X=6.24 $Y=1.515 $X2=0 $Y2=0
cc_252 N_A3_M1000_g N_VPWR_c_562_n 0.00333896f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A3_M1012_g N_VPWR_c_562_n 0.00333926f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A3_M1025_g N_VPWR_c_562_n 0.00333916f $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A3_M1034_g N_VPWR_c_562_n 0.00333896f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A3_M1000_g N_VPWR_c_566_n 0.0023861f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A3_M1000_g N_VPWR_c_552_n 0.00428307f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A3_M1012_g N_VPWR_c_552_n 0.00423847f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A3_M1025_g N_VPWR_c_552_n 0.00424916f $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A3_M1034_g N_VPWR_c_552_n 0.00424355f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A3_M1011_g N_Y_c_664_n 0.0125331f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A3_M1013_g N_Y_c_664_n 0.011293f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A3_M1027_g N_Y_c_664_n 0.0112465f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A3_M1035_g N_Y_c_664_n 0.0144061f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A3_c_283_n N_Y_c_664_n 0.0195424f $X=6.24 $Y=1.515 $X2=0 $Y2=0
cc_266 N_A3_c_284_n N_Y_c_664_n 0.125235f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_267 N_A3_M1000_g N_Y_c_669_n 0.0169965f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_268 N_A3_c_284_n N_Y_c_669_n 0.00639096f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_269 N_A3_M1012_g N_Y_c_723_n 0.00898357f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A3_M1025_g N_Y_c_723_n 4.54754e-19 $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A3_M1012_g N_Y_c_725_n 0.0141209f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A3_M1025_g N_Y_c_725_n 0.0152718f $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A3_c_283_n N_Y_c_725_n 8.63305e-19 $X=6.24 $Y=1.515 $X2=0 $Y2=0
cc_274 N_A3_c_291_n N_Y_c_725_n 0.0344934f $X=5.535 $Y=1.605 $X2=0 $Y2=0
cc_275 N_A3_c_284_n N_Y_c_725_n 0.00678134f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_276 N_A3_M1034_g N_Y_c_730_n 0.0208039f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A3_c_289_n N_Y_c_730_n 0.0115976f $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_278 N_A3_M1000_g N_Y_c_671_n 5.59553e-19 $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A3_M1012_g N_Y_c_671_n 0.00375725f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_280 N_A3_M1025_g N_Y_c_671_n 6.0418e-19 $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A3_c_283_n N_Y_c_671_n 0.00397658f $X=6.24 $Y=1.515 $X2=0 $Y2=0
cc_282 N_A3_c_284_n N_Y_c_671_n 0.0257279f $X=5.185 $Y=1.605 $X2=0 $Y2=0
cc_283 N_A3_M1034_g N_Y_c_737_n 0.00906877f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A3_c_289_n N_Y_c_737_n 0.0261729f $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_285 N_A3_c_283_n N_Y_c_737_n 0.00146526f $X=6.24 $Y=1.515 $X2=0 $Y2=0
cc_286 N_A3_M1035_g Y 0.00958083f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A3_c_289_n Y 0.0283828f $X=6.03 $Y=1.515 $X2=0 $Y2=0
cc_288 N_A3_M1000_g N_A_841_368#_c_800_n 0.00895541f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A3_M1012_g N_A_841_368#_c_800_n 2.72638e-19 $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A3_M1000_g N_A_841_368#_c_801_n 0.0119307f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A3_M1012_g N_A_841_368#_c_801_n 0.01459f $X=5.075 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A3_M1000_g N_A_841_368#_c_802_n 0.00291744f $X=4.575 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A3_M1025_g N_A_841_368#_c_815_n 0.00802203f $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A3_M1034_g N_A_841_368#_c_815_n 7.99633e-19 $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_295 N_A3_M1025_g N_A_841_368#_c_803_n 0.0138388f $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A3_M1034_g N_A_841_368#_c_803_n 0.012538f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A3_M1025_g N_A_841_368#_c_819_n 7.9395e-19 $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A3_M1034_g N_A_841_368#_c_819_n 0.0102581f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A3_M1025_g N_A_841_368#_c_807_n 0.00179757f $X=5.595 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A3_M1034_g N_A_841_368#_c_808_n 0.001916f $X=6.225 $Y=2.4 $X2=0 $Y2=0
cc_301 N_A3_M1011_g N_A_459_74#_c_969_n 5.29638e-19 $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A3_M1011_g N_A_459_74#_c_970_n 0.00284982f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A3_M1011_g N_A_459_74#_c_971_n 0.0128625f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A3_M1011_g N_A_459_74#_c_973_n 4.39567e-19 $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A3_M1013_g N_A_459_74#_c_973_n 0.00688453f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A3_M1027_g N_A_459_74#_c_973_n 8.14332e-19 $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A3_M1013_g N_A_459_74#_c_997_n 0.0095689f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A3_M1027_g N_A_459_74#_c_997_n 0.0095689f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A3_M1013_g N_A_459_74#_c_974_n 8.11586e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A3_M1027_g N_A_459_74#_c_974_n 0.00724443f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A3_M1035_g N_A_459_74#_c_974_n 0.0072728f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A3_M1035_g N_A_459_74#_c_1002_n 0.00947961f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A3_M1035_g N_A_459_74#_c_975_n 8.13633e-19 $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A3_M1013_g N_A_459_74#_c_1004_n 0.00181289f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A3_M1027_g N_A_459_74#_c_1005_n 0.00181289f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A3_M1035_g N_A_459_74#_c_1005_n 0.00181289f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A3_M1035_g N_A_459_74#_c_983_n 9.18816e-19 $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A3_M1011_g N_VGND_c_1118_n 0.0078527f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A3_M1013_g N_VGND_c_1118_n 4.46147e-19 $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A3_M1013_g N_VGND_c_1119_n 0.00320743f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A3_M1027_g N_VGND_c_1119_n 0.00465809f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A3_M1035_g N_VGND_c_1120_n 0.00471422f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A3_M1011_g N_VGND_c_1126_n 0.00281141f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A3_M1013_g N_VGND_c_1126_n 0.00331438f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A3_M1027_g N_VGND_c_1127_n 0.00331438f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A3_M1035_g N_VGND_c_1127_n 0.00331438f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A3_M1011_g N_VGND_c_1138_n 0.00365066f $X=4.79 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A3_M1013_g N_VGND_c_1138_n 0.00427695f $X=5.22 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A3_M1027_g N_VGND_c_1138_n 0.00427695f $X=5.81 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A3_M1035_g N_VGND_c_1138_n 0.00427774f $X=6.24 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A2_c_381_n N_A1_M1001_g 0.0181944f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_332 N_A2_c_382_n N_A1_M1001_g 0.00761232f $X=8.175 $Y=1.44 $X2=0 $Y2=0
cc_333 N_A2_M1030_g N_A1_c_472_n 0.00761232f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_334 N_A2_M1030_g N_VPWR_c_556_n 0.00191284f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A2_M1024_g N_VPWR_c_562_n 0.00333896f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A2_M1026_g N_VPWR_c_562_n 0.00333926f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_337 N_A2_M1028_g N_VPWR_c_562_n 0.00333926f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_338 N_A2_M1030_g N_VPWR_c_562_n 0.00333896f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_339 N_A2_M1024_g N_VPWR_c_552_n 0.00423284f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_340 N_A2_M1026_g N_VPWR_c_552_n 0.00424108f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_341 N_A2_M1028_g N_VPWR_c_552_n 0.00423619f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_342 N_A2_M1030_g N_VPWR_c_552_n 0.00427818f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A2_M1024_g N_Y_c_730_n 0.00383501f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_344 N_A2_M1004_g N_Y_c_665_n 0.00324583f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A2_M1024_g Y 0.00672158f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_346 N_A2_M1004_g Y 0.00210281f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A2_M1026_g Y 7.70243e-19 $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A2_c_387_n Y 0.0332185f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_349 N_A2_c_382_n Y 0.00788086f $X=8.175 $Y=1.44 $X2=0 $Y2=0
cc_350 N_A2_M1024_g N_A_841_368#_c_819_n 0.00965153f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A2_M1026_g N_A_841_368#_c_819_n 5.88728e-19 $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A2_M1024_g N_A_841_368#_c_804_n 0.0119307f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_353 N_A2_M1026_g N_A_841_368#_c_804_n 0.0146917f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_354 N_A2_M1028_g N_A_841_368#_c_805_n 0.0143955f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_355 N_A2_M1030_g N_A_841_368#_c_805_n 0.014552f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_356 N_A2_M1028_g N_A_841_368#_c_806_n 5.70966e-19 $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A2_M1030_g N_A_841_368#_c_806_n 0.00851312f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_358 N_A2_M1024_g N_A_841_368#_c_808_n 0.001916f $X=6.675 $Y=2.4 $X2=0 $Y2=0
cc_359 N_A2_M1026_g N_A_1353_368#_c_877_n 0.0134861f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A2_M1028_g N_A_1353_368#_c_877_n 0.013761f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A2_c_387_n N_A_1353_368#_c_877_n 0.0464562f $X=7.61 $Y=1.515 $X2=0
+ $Y2=0
cc_362 N_A2_c_382_n N_A_1353_368#_c_877_n 0.00103042f $X=8.175 $Y=1.44 $X2=0
+ $Y2=0
cc_363 N_A2_M1026_g N_A_1353_368#_c_881_n 4.56234e-19 $X=7.175 $Y=2.4 $X2=0
+ $Y2=0
cc_364 N_A2_M1028_g N_A_1353_368#_c_881_n 0.00975709f $X=7.725 $Y=2.4 $X2=0
+ $Y2=0
cc_365 N_A2_M1030_g N_A_1353_368#_c_874_n 0.019644f $X=8.175 $Y=2.4 $X2=0 $Y2=0
cc_366 N_A2_M1026_g N_A_1353_368#_c_884_n 0.0106569f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_367 N_A2_M1028_g N_A_1353_368#_c_884_n 5.48326e-19 $X=7.725 $Y=2.4 $X2=0
+ $Y2=0
cc_368 N_A2_c_387_n N_A_1353_368#_c_884_n 0.0246996f $X=7.61 $Y=1.515 $X2=0
+ $Y2=0
cc_369 N_A2_c_382_n N_A_1353_368#_c_884_n 8.53086e-19 $X=8.175 $Y=1.44 $X2=0
+ $Y2=0
cc_370 N_A2_M1028_g N_A_1353_368#_c_888_n 0.00260767f $X=7.725 $Y=2.4 $X2=0
+ $Y2=0
cc_371 N_A2_c_382_n N_A_1353_368#_c_888_n 0.00281866f $X=8.175 $Y=1.44 $X2=0
+ $Y2=0
cc_372 N_A2_M1004_g N_A_459_74#_c_974_n 8.06429e-19 $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A2_M1004_g N_A_459_74#_c_1002_n 0.0114917f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A2_c_387_n N_A_459_74#_c_1002_n 0.00430774f $X=7.61 $Y=1.515 $X2=0
+ $Y2=0
cc_375 N_A2_c_382_n N_A_459_74#_c_1002_n 0.00466587f $X=8.175 $Y=1.44 $X2=0
+ $Y2=0
cc_376 N_A2_M1004_g N_A_459_74#_c_975_n 0.00661943f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A2_M1006_g N_A_459_74#_c_975_n 3.97481e-19 $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A2_M1006_g N_A_459_74#_c_976_n 0.0127949f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A2_c_379_n N_A_459_74#_c_976_n 0.0159019f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_380 N_A2_c_387_n N_A_459_74#_c_976_n 0.0477395f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_381 N_A2_c_382_n N_A_459_74#_c_976_n 0.00509226f $X=8.175 $Y=1.44 $X2=0 $Y2=0
cc_382 N_A2_c_379_n N_A_459_74#_c_977_n 0.00814722f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_383 N_A2_c_381_n N_A_459_74#_c_977_n 0.00156085f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_384 N_A2_c_382_n N_A_459_74#_c_978_n 0.0184133f $X=8.175 $Y=1.44 $X2=0 $Y2=0
cc_385 N_A2_c_381_n N_A_459_74#_c_979_n 2.1934e-19 $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_386 N_A2_c_381_n N_A_459_74#_c_980_n 6.00311e-19 $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_387 N_A2_M1004_g N_A_459_74#_c_983_n 0.00668147f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A2_c_387_n N_A_459_74#_c_983_n 0.0211953f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_389 N_A2_c_382_n N_A_459_74#_c_983_n 0.00272398f $X=8.175 $Y=1.44 $X2=0 $Y2=0
cc_390 N_A2_M1006_g N_A_459_74#_c_984_n 5.55763e-19 $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A2_c_379_n N_A_459_74#_c_984_n 7.16428e-19 $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_392 N_A2_c_387_n N_A_459_74#_c_984_n 0.00906486f $X=7.61 $Y=1.515 $X2=0 $Y2=0
cc_393 N_A2_c_382_n N_A_459_74#_c_984_n 0.0182807f $X=8.175 $Y=1.44 $X2=0 $Y2=0
cc_394 N_A2_M1004_g N_VGND_c_1120_n 0.00325376f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_395 N_A2_M1004_g N_VGND_c_1121_n 5.16425e-19 $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A2_M1006_g N_VGND_c_1121_n 0.0103635f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A2_c_379_n N_VGND_c_1121_n 0.00243974f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_398 N_A2_c_379_n N_VGND_c_1122_n 5.07467e-19 $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_399 N_A2_c_381_n N_VGND_c_1122_n 0.0130384f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_400 N_A2_M1004_g N_VGND_c_1128_n 0.00331438f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A2_M1006_g N_VGND_c_1128_n 0.00383152f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_402 N_A2_c_379_n N_VGND_c_1129_n 0.00461464f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_403 N_A2_c_381_n N_VGND_c_1129_n 0.00383152f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_404 N_A2_M1004_g N_VGND_c_1138_n 0.00427774f $X=6.84 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A2_M1006_g N_VGND_c_1138_n 0.0075754f $X=7.27 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A2_c_379_n N_VGND_c_1138_n 0.00908525f $X=7.74 $Y=1.2 $X2=0 $Y2=0
cc_407 N_A2_c_381_n N_VGND_c_1138_n 0.00758242f $X=8.245 $Y=1.2 $X2=0 $Y2=0
cc_408 N_A1_M1008_g N_VPWR_c_556_n 0.0131746f $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_409 N_A1_M1009_g N_VPWR_c_556_n 4.99668e-19 $X=9.635 $Y=2.4 $X2=0 $Y2=0
cc_410 N_A1_M1008_g N_VPWR_c_557_n 4.99668e-19 $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A1_M1009_g N_VPWR_c_557_n 0.0119877f $X=9.635 $Y=2.4 $X2=0 $Y2=0
cc_412 N_A1_M1014_g N_VPWR_c_557_n 0.0121164f $X=10.085 $Y=2.4 $X2=0 $Y2=0
cc_413 N_A1_M1033_g N_VPWR_c_557_n 5.18631e-19 $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A1_M1033_g N_VPWR_c_559_n 0.00551672f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_415 N_A1_M1008_g N_VPWR_c_563_n 0.00460063f $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_416 N_A1_M1009_g N_VPWR_c_563_n 0.00460063f $X=9.635 $Y=2.4 $X2=0 $Y2=0
cc_417 N_A1_M1014_g N_VPWR_c_564_n 0.00460063f $X=10.085 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A1_M1033_g N_VPWR_c_564_n 0.005209f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A1_M1008_g N_VPWR_c_552_n 0.00908554f $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_420 N_A1_M1009_g N_VPWR_c_552_n 0.00908554f $X=9.635 $Y=2.4 $X2=0 $Y2=0
cc_421 N_A1_M1014_g N_VPWR_c_552_n 0.00908554f $X=10.085 $Y=2.4 $X2=0 $Y2=0
cc_422 N_A1_M1033_g N_VPWR_c_552_n 0.00986008f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_423 N_A1_M1008_g N_A_841_368#_c_805_n 6.08298e-19 $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_424 N_A1_M1008_g N_A_841_368#_c_806_n 0.00102674f $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_425 N_A1_c_472_n N_A_1353_368#_c_874_n 0.0128386f $X=8.75 $Y=1.605 $X2=0
+ $Y2=0
cc_426 N_A1_M1008_g N_A_1353_368#_c_874_n 0.0199043f $X=9.185 $Y=2.4 $X2=0 $Y2=0
cc_427 N_A1_c_483_n N_A_1353_368#_c_874_n 0.00895228f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_428 N_A1_M1008_g N_A_1353_368#_c_875_n 2.89602e-19 $X=9.185 $Y=2.4 $X2=0
+ $Y2=0
cc_429 N_A1_M1009_g N_A_1353_368#_c_875_n 2.89602e-19 $X=9.635 $Y=2.4 $X2=0
+ $Y2=0
cc_430 N_A1_M1009_g N_A_1353_368#_c_895_n 0.0152674f $X=9.635 $Y=2.4 $X2=0 $Y2=0
cc_431 N_A1_M1014_g N_A_1353_368#_c_895_n 0.0152674f $X=10.085 $Y=2.4 $X2=0
+ $Y2=0
cc_432 N_A1_c_483_n N_A_1353_368#_c_895_n 0.045745f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_433 N_A1_c_476_n N_A_1353_368#_c_895_n 4.96975e-19 $X=10.535 $Y=1.44 $X2=0
+ $Y2=0
cc_434 N_A1_M1033_g N_A_1353_368#_c_899_n 0.00401886f $X=10.535 $Y=2.4 $X2=0
+ $Y2=0
cc_435 N_A1_c_483_n N_A_1353_368#_c_899_n 0.0174453f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_436 N_A1_c_476_n N_A_1353_368#_c_899_n 5.51705e-19 $X=10.535 $Y=1.44 $X2=0
+ $Y2=0
cc_437 N_A1_M1014_g N_A_1353_368#_c_876_n 2.92425e-19 $X=10.085 $Y=2.4 $X2=0
+ $Y2=0
cc_438 N_A1_M1033_g N_A_1353_368#_c_876_n 0.011127f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_439 N_A1_c_483_n N_A_1353_368#_c_904_n 0.0170101f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_440 N_A1_c_476_n N_A_1353_368#_c_904_n 5.54777e-19 $X=10.535 $Y=1.44 $X2=0
+ $Y2=0
cc_441 N_A1_M1001_g N_A_459_74#_c_978_n 0.0142591f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_442 N_A1_c_471_n N_A_459_74#_c_978_n 0.00285025f $X=9.03 $Y=1.605 $X2=0 $Y2=0
cc_443 N_A1_M1002_g N_A_459_74#_c_978_n 0.0028354f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_444 N_A1_c_483_n N_A_459_74#_c_978_n 0.00974864f $X=10.35 $Y=1.515 $X2=0
+ $Y2=0
cc_445 N_A1_M1001_g N_A_459_74#_c_979_n 0.00725305f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_446 N_A1_M1002_g N_A_459_74#_c_979_n 3.97173e-19 $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_447 N_A1_M1001_g N_A_459_74#_c_980_n 0.00467801f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_448 N_A1_M1002_g N_A_459_74#_c_980_n 0.00432461f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_449 N_A1_M1002_g N_A_459_74#_c_981_n 0.0185175f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_450 N_A1_c_474_n N_A_459_74#_c_981_n 0.0150704f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_451 N_A1_c_483_n N_A_459_74#_c_981_n 0.0802473f $X=10.35 $Y=1.515 $X2=0 $Y2=0
cc_452 N_A1_c_476_n N_A_459_74#_c_981_n 0.0196647f $X=10.535 $Y=1.44 $X2=0 $Y2=0
cc_453 N_A1_c_474_n N_A_459_74#_c_982_n 0.0120086f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_454 N_A1_c_475_n N_A_459_74#_c_982_n 4.13268e-19 $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_455 N_A1_M1001_g N_A_459_74#_c_984_n 3.35826e-19 $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A1_M1001_g N_A_459_74#_c_1045_n 0.00199342f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_457 N_A1_M1001_g N_VGND_c_1122_n 0.0019818f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A1_c_474_n N_VGND_c_1124_n 6.05373e-19 $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_459 N_A1_c_475_n N_VGND_c_1124_n 0.0160519f $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_460 N_A1_c_476_n N_VGND_c_1124_n 2.29254e-19 $X=10.535 $Y=1.44 $X2=0 $Y2=0
cc_461 N_A1_c_474_n N_VGND_c_1130_n 0.00451267f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_462 N_A1_c_475_n N_VGND_c_1130_n 0.00383152f $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_463 N_A1_M1001_g N_VGND_c_1136_n 0.00434272f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_464 N_A1_M1002_g N_VGND_c_1136_n 0.00383152f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_465 N_A1_M1001_g N_VGND_c_1137_n 5.00706e-19 $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_466 N_A1_M1002_g N_VGND_c_1137_n 0.0120529f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A1_c_474_n N_VGND_c_1137_n 0.00510378f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_468 N_A1_M1001_g N_VGND_c_1138_n 0.00820382f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A1_M1002_g N_VGND_c_1138_n 0.00752925f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A1_c_474_n N_VGND_c_1138_n 0.00879879f $X=10.1 $Y=1.2 $X2=0 $Y2=0
cc_471 N_A1_c_475_n N_VGND_c_1138_n 0.00757689f $X=10.545 $Y=1.2 $X2=0 $Y2=0
cc_472 N_VPWR_c_554_n N_Y_c_673_n 0.00919206f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_473 N_VPWR_c_554_n N_Y_c_667_n 0.0437611f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_474 N_VPWR_c_555_n N_Y_c_667_n 0.0266809f $X=1.405 $Y=2.455 $X2=0 $Y2=0
cc_475 N_VPWR_c_560_n N_Y_c_667_n 0.0146357f $X=1.24 $Y=3.33 $X2=0 $Y2=0
cc_476 N_VPWR_c_552_n N_Y_c_667_n 0.0121141f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_M1021_s N_Y_c_678_n 0.00568561f $X=1.27 $Y=1.84 $X2=0 $Y2=0
cc_478 N_VPWR_c_555_n N_Y_c_678_n 0.0189268f $X=1.405 $Y=2.455 $X2=0 $Y2=0
cc_479 N_VPWR_c_555_n N_Y_c_668_n 0.0266809f $X=1.405 $Y=2.455 $X2=0 $Y2=0
cc_480 N_VPWR_c_565_n N_Y_c_668_n 0.0144623f $X=2.24 $Y=2.852 $X2=0 $Y2=0
cc_481 N_VPWR_c_566_n N_Y_c_668_n 0.0268614f $X=3.905 $Y=2.852 $X2=0 $Y2=0
cc_482 N_VPWR_c_552_n N_Y_c_668_n 0.0118344f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_M1023_s N_Y_c_669_n 0.045746f $X=2.22 $Y=1.84 $X2=0 $Y2=0
cc_484 N_VPWR_c_566_n N_Y_c_669_n 0.131886f $X=3.905 $Y=2.852 $X2=0 $Y2=0
cc_485 N_VPWR_c_566_n N_A_841_368#_c_800_n 0.0383127f $X=3.905 $Y=2.852 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_562_n N_A_841_368#_c_801_n 0.0421443f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_552_n N_A_841_368#_c_801_n 0.0236813f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_562_n N_A_841_368#_c_802_n 0.0235512f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_566_n N_A_841_368#_c_802_n 0.0112248f $X=3.905 $Y=2.852 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_552_n N_A_841_368#_c_802_n 0.0126924f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_562_n N_A_841_368#_c_803_n 0.0486181f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_552_n N_A_841_368#_c_803_n 0.0274872f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_562_n N_A_841_368#_c_804_n 0.0421443f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_552_n N_A_841_368#_c_804_n 0.0236813f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_556_n N_A_841_368#_c_805_n 0.0121616f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_562_n N_A_841_368#_c_805_n 0.0624745f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_552_n N_A_841_368#_c_805_n 0.0344938f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_556_n N_A_841_368#_c_806_n 0.0387318f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_562_n N_A_841_368#_c_807_n 0.0236215f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_552_n N_A_841_368#_c_807_n 0.0127839f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_562_n N_A_841_368#_c_808_n 0.0234458f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_552_n N_A_841_368#_c_808_n 0.0125551f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_562_n N_A_841_368#_c_809_n 0.0236566f $X=8.795 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_552_n N_A_841_368#_c_809_n 0.0128296f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_M1008_s N_A_1353_368#_c_874_n 0.00650996f $X=8.815 $Y=1.84 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_556_n N_A_1353_368#_c_874_n 0.0212273f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_556_n N_A_1353_368#_c_875_n 0.025138f $X=8.96 $Y=2.415 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_557_n N_A_1353_368#_c_875_n 0.025138f $X=9.86 $Y=2.415 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_563_n N_A_1353_368#_c_875_n 0.0101736f $X=9.695 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_552_n N_A_1353_368#_c_875_n 0.0084208f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_511 N_VPWR_M1009_s N_A_1353_368#_c_895_n 0.00320006f $X=9.725 $Y=1.84 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_557_n N_A_1353_368#_c_895_n 0.0164816f $X=9.86 $Y=2.415 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_557_n N_A_1353_368#_c_876_n 0.0251606f $X=9.86 $Y=2.415 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_559_n N_A_1353_368#_c_876_n 0.0273089f $X=10.76 $Y=1.985 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_564_n N_A_1353_368#_c_876_n 0.0123179f $X=10.675 $Y=3.33 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_552_n N_A_1353_368#_c_876_n 0.0101276f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_517 N_Y_c_669_n N_A_841_368#_M1000_s 0.0118091f $X=4.685 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_518 N_Y_c_725_n N_A_841_368#_M1012_s 0.00449621f $X=5.685 $Y=2.035 $X2=0
+ $Y2=0
cc_519 N_Y_c_730_n N_A_841_368#_M1034_s 0.00172633f $X=6.365 $Y=2.035 $X2=0
+ $Y2=0
cc_520 N_Y_c_669_n N_A_841_368#_c_800_n 0.0219147f $X=4.685 $Y=2.035 $X2=0 $Y2=0
cc_521 N_Y_M1000_d N_A_841_368#_c_801_n 0.00218982f $X=4.665 $Y=1.84 $X2=0 $Y2=0
cc_522 N_Y_c_723_n N_A_841_368#_c_801_n 0.0177084f $X=4.85 $Y=2.31 $X2=0 $Y2=0
cc_523 N_Y_c_725_n N_A_841_368#_c_815_n 0.0190305f $X=5.685 $Y=2.035 $X2=0 $Y2=0
cc_524 N_Y_c_737_n N_A_841_368#_c_815_n 0.032507f $X=5.85 $Y=2.115 $X2=0 $Y2=0
cc_525 N_Y_M1025_d N_A_841_368#_c_803_n 0.00560237f $X=5.685 $Y=1.84 $X2=0 $Y2=0
cc_526 N_Y_c_737_n N_A_841_368#_c_803_n 0.0207027f $X=5.85 $Y=2.115 $X2=0 $Y2=0
cc_527 N_Y_c_730_n N_A_841_368#_c_819_n 0.0169941f $X=6.365 $Y=2.035 $X2=0 $Y2=0
cc_528 N_Y_c_737_n N_A_841_368#_c_819_n 0.0242292f $X=5.85 $Y=2.115 $X2=0 $Y2=0
cc_529 N_Y_c_685_n N_A_27_74#_M1019_s 0.00342755f $X=1.41 $Y=1.015 $X2=0 $Y2=0
cc_530 N_Y_c_664_n N_A_27_74#_M1032_s 0.00176461f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_531 N_Y_c_664_n N_A_27_74#_M1016_s 0.00176891f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_532 N_Y_c_664_n N_A_27_74#_M1031_s 0.00213024f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_533 N_Y_M1005_d N_A_27_74#_c_931_n 0.00174304f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_534 N_Y_M1020_d N_A_27_74#_c_931_n 0.00169393f $X=1.435 $Y=0.37 $X2=0 $Y2=0
cc_535 N_Y_c_664_n N_A_27_74#_c_931_n 0.0036578f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_536 N_Y_c_685_n N_A_27_74#_c_931_n 0.0633287f $X=1.41 $Y=1.015 $X2=0 $Y2=0
cc_537 N_Y_c_664_n N_A_27_74#_c_954_n 0.0133131f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_538 N_Y_c_664_n N_A_27_74#_c_932_n 0.0955773f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_539 N_Y_c_664_n N_A_459_74#_M1003_d 0.00176891f $X=6.365 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_540 N_Y_c_664_n N_A_459_74#_M1017_d 0.00187547f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_541 N_Y_c_664_n N_A_459_74#_M1011_s 0.00176461f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_542 N_Y_c_664_n N_A_459_74#_M1027_s 0.00176461f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_543 N_Y_c_664_n N_A_459_74#_c_969_n 0.0061464f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_544 N_Y_c_664_n N_A_459_74#_c_971_n 0.0410903f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_545 N_Y_c_664_n N_A_459_74#_c_972_n 0.0141908f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_546 N_Y_c_664_n N_A_459_74#_c_997_n 0.0405558f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_547 N_Y_c_664_n N_A_459_74#_c_1002_n 0.00843866f $X=6.365 $Y=1.175 $X2=0
+ $Y2=0
cc_548 N_Y_c_665_n N_A_459_74#_c_1002_n 0.018143f $X=6.48 $Y=1.26 $X2=0 $Y2=0
cc_549 N_Y_c_664_n N_A_459_74#_c_1004_n 0.0151907f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_550 N_Y_c_664_n N_A_459_74#_c_1005_n 0.0170682f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_551 N_Y_c_665_n N_A_459_74#_c_983_n 0.00490592f $X=6.48 $Y=1.26 $X2=0 $Y2=0
cc_552 N_Y_c_664_n N_VGND_M1011_d 0.00213024f $X=6.365 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_553 N_Y_c_664_n N_VGND_M1013_d 0.00355802f $X=6.365 $Y=1.175 $X2=0 $Y2=0
cc_554 N_Y_c_665_n N_VGND_M1035_d 0.002798f $X=6.48 $Y=1.26 $X2=0 $Y2=0
cc_555 N_A_841_368#_c_804_n N_A_1353_368#_M1024_d 0.00218982f $X=7.285 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_556 N_A_841_368#_c_805_n N_A_1353_368#_M1028_d 0.00165831f $X=8.235 $Y=2.99
+ $X2=0 $Y2=0
cc_557 N_A_841_368#_M1026_s N_A_1353_368#_c_877_n 0.00516882f $X=7.265 $Y=1.84
+ $X2=0 $Y2=0
cc_558 N_A_841_368#_c_869_p N_A_1353_368#_c_877_n 0.0208278f $X=7.45 $Y=2.455
+ $X2=0 $Y2=0
cc_559 N_A_841_368#_c_805_n N_A_1353_368#_c_881_n 0.0139027f $X=8.235 $Y=2.99
+ $X2=0 $Y2=0
cc_560 N_A_841_368#_M1030_s N_A_1353_368#_c_874_n 0.00749925f $X=8.265 $Y=1.84
+ $X2=0 $Y2=0
cc_561 N_A_841_368#_c_806_n N_A_1353_368#_c_874_n 0.0212273f $X=8.4 $Y=2.415
+ $X2=0 $Y2=0
cc_562 N_A_841_368#_c_804_n N_A_1353_368#_c_884_n 0.0177084f $X=7.285 $Y=2.99
+ $X2=0 $Y2=0
cc_563 N_A_1353_368#_c_874_n N_A_459_74#_c_978_n 0.0296093f $X=9.295 $Y=2.05
+ $X2=0 $Y2=0
cc_564 N_A_1353_368#_c_874_n N_A_459_74#_c_984_n 0.00130388f $X=9.295 $Y=2.05
+ $X2=0 $Y2=0
cc_565 N_A_1353_368#_c_888_n N_A_459_74#_c_984_n 0.00385768f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_566 N_A_27_74#_c_932_n N_A_459_74#_M1003_d 0.00335829f $X=3.735 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_567 N_A_27_74#_c_932_n N_A_459_74#_M1017_d 0.003555f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_568 N_A_27_74#_M1016_s N_A_459_74#_c_969_n 0.00179007f $X=2.725 $Y=0.37 $X2=0
+ $Y2=0
cc_569 N_A_27_74#_M1031_s N_A_459_74#_c_969_n 0.002891f $X=3.595 $Y=0.37 $X2=0
+ $Y2=0
cc_570 N_A_27_74#_c_931_n N_A_459_74#_c_969_n 0.0101071f $X=1.92 $Y=0.475 $X2=0
+ $Y2=0
cc_571 N_A_27_74#_c_932_n N_A_459_74#_c_969_n 0.0865605f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_572 N_A_27_74#_c_932_n N_A_459_74#_c_972_n 0.015741f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_573 N_A_27_74#_c_929_n N_VGND_c_1125_n 0.0111552f $X=0.24 $Y=0.6 $X2=0 $Y2=0
cc_574 N_A_27_74#_c_931_n N_VGND_c_1125_n 0.0702753f $X=1.92 $Y=0.475 $X2=0
+ $Y2=0
cc_575 N_A_27_74#_c_932_n N_VGND_c_1125_n 0.00197884f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_576 N_A_27_74#_c_929_n N_VGND_c_1138_n 0.00923333f $X=0.24 $Y=0.6 $X2=0 $Y2=0
cc_577 N_A_27_74#_c_931_n N_VGND_c_1138_n 0.0589522f $X=1.92 $Y=0.475 $X2=0
+ $Y2=0
cc_578 N_A_27_74#_c_932_n N_VGND_c_1138_n 0.00654682f $X=3.735 $Y=0.835 $X2=0
+ $Y2=0
cc_579 N_A_459_74#_c_971_n N_VGND_M1011_d 0.00447087f $X=4.92 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_580 N_A_459_74#_c_997_n N_VGND_M1013_d 0.00724158f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_581 N_A_459_74#_c_1002_n N_VGND_M1035_d 0.00831277f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_582 N_A_459_74#_c_976_n N_VGND_M1006_d 0.0022694f $X=7.945 $Y=1.095 $X2=0
+ $Y2=0
cc_583 N_A_459_74#_c_981_n N_VGND_M1002_d 0.0117895f $X=10.165 $Y=1.045 $X2=0
+ $Y2=0
cc_584 N_A_459_74#_c_969_n N_VGND_c_1118_n 0.0221151f $X=4.07 $Y=0.455 $X2=0
+ $Y2=0
cc_585 N_A_459_74#_c_971_n N_VGND_c_1118_n 0.0212697f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_586 N_A_459_74#_c_973_n N_VGND_c_1118_n 0.00897147f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_587 N_A_459_74#_c_973_n N_VGND_c_1119_n 0.00865936f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_588 N_A_459_74#_c_997_n N_VGND_c_1119_n 0.0256608f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_589 N_A_459_74#_c_974_n N_VGND_c_1119_n 0.00900273f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_590 N_A_459_74#_c_974_n N_VGND_c_1120_n 0.00900616f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_591 N_A_459_74#_c_1002_n N_VGND_c_1120_n 0.0264479f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_592 N_A_459_74#_c_975_n N_VGND_c_1120_n 0.0086628f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_593 N_A_459_74#_c_975_n N_VGND_c_1121_n 0.0177526f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_594 N_A_459_74#_c_976_n N_VGND_c_1121_n 0.017402f $X=7.945 $Y=1.095 $X2=0
+ $Y2=0
cc_595 N_A_459_74#_c_977_n N_VGND_c_1121_n 0.0120634f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_596 N_A_459_74#_c_977_n N_VGND_c_1122_n 0.0281649f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_597 N_A_459_74#_c_978_n N_VGND_c_1122_n 0.0207473f $X=8.725 $Y=1.385 $X2=0
+ $Y2=0
cc_598 N_A_459_74#_c_979_n N_VGND_c_1122_n 0.0216462f $X=8.89 $Y=0.515 $X2=0
+ $Y2=0
cc_599 N_A_459_74#_c_1045_n N_VGND_c_1122_n 0.00756924f $X=8.85 $Y=1.045 $X2=0
+ $Y2=0
cc_600 N_A_459_74#_c_981_n N_VGND_c_1124_n 0.00697079f $X=10.165 $Y=1.045 $X2=0
+ $Y2=0
cc_601 N_A_459_74#_c_982_n N_VGND_c_1124_n 0.0225912f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
cc_602 N_A_459_74#_c_969_n N_VGND_c_1125_n 0.0878111f $X=4.07 $Y=0.455 $X2=0
+ $Y2=0
cc_603 N_A_459_74#_c_971_n N_VGND_c_1125_n 0.0024506f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_604 N_A_459_74#_c_971_n N_VGND_c_1126_n 0.00197156f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_605 N_A_459_74#_c_973_n N_VGND_c_1126_n 0.0108551f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_606 N_A_459_74#_c_997_n N_VGND_c_1126_n 0.00197156f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_607 N_A_459_74#_c_997_n N_VGND_c_1127_n 0.00197156f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_608 N_A_459_74#_c_974_n N_VGND_c_1127_n 0.0143093f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_609 N_A_459_74#_c_1002_n N_VGND_c_1127_n 0.00197156f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_610 N_A_459_74#_c_1002_n N_VGND_c_1128_n 0.00197695f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_611 N_A_459_74#_c_975_n N_VGND_c_1128_n 0.0109942f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_612 N_A_459_74#_c_977_n N_VGND_c_1129_n 0.00749631f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_613 N_A_459_74#_c_982_n N_VGND_c_1130_n 0.0110391f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
cc_614 N_A_459_74#_c_979_n N_VGND_c_1136_n 0.0109942f $X=8.89 $Y=0.515 $X2=0
+ $Y2=0
cc_615 N_A_459_74#_c_979_n N_VGND_c_1137_n 0.01839f $X=8.89 $Y=0.515 $X2=0 $Y2=0
cc_616 N_A_459_74#_c_981_n N_VGND_c_1137_n 0.0610657f $X=10.165 $Y=1.045 $X2=0
+ $Y2=0
cc_617 N_A_459_74#_c_982_n N_VGND_c_1137_n 0.0167469f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0
cc_618 N_A_459_74#_c_969_n N_VGND_c_1138_n 0.0692687f $X=4.07 $Y=0.455 $X2=0
+ $Y2=0
cc_619 N_A_459_74#_c_971_n N_VGND_c_1138_n 0.00976958f $X=4.92 $Y=0.835 $X2=0
+ $Y2=0
cc_620 N_A_459_74#_c_973_n N_VGND_c_1138_n 0.00898945f $X=5.005 $Y=0.635 $X2=0
+ $Y2=0
cc_621 N_A_459_74#_c_997_n N_VGND_c_1138_n 0.00943478f $X=5.86 $Y=0.835 $X2=0
+ $Y2=0
cc_622 N_A_459_74#_c_974_n N_VGND_c_1138_n 0.0118109f $X=6.025 $Y=0.635 $X2=0
+ $Y2=0
cc_623 N_A_459_74#_c_1002_n N_VGND_c_1138_n 0.00947592f $X=6.89 $Y=0.835 $X2=0
+ $Y2=0
cc_624 N_A_459_74#_c_975_n N_VGND_c_1138_n 0.00904371f $X=7.055 $Y=0.515 $X2=0
+ $Y2=0
cc_625 N_A_459_74#_c_977_n N_VGND_c_1138_n 0.0062048f $X=8.03 $Y=0.515 $X2=0
+ $Y2=0
cc_626 N_A_459_74#_c_979_n N_VGND_c_1138_n 0.00904371f $X=8.89 $Y=0.515 $X2=0
+ $Y2=0
cc_627 N_A_459_74#_c_982_n N_VGND_c_1138_n 0.00911606f $X=10.33 $Y=0.515 $X2=0
+ $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__buf_16 A VGND VNB VPB VPWR X
X0 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X25 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X33 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X41 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

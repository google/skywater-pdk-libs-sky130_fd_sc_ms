* NGSPICE file created from sky130_fd_sc_ms__or2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__or2b_2 A B_N VGND VNB VPB VPWR X
M1000 a_187_48# a_27_368# a_473_368# VPB pshort w=1e+06u l=180000u
+  ad=4e+11p pd=2.8e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR B_N a_27_368# VPB pshort w=840000u l=180000u
+  ad=8.002e+11p pd=5.97e+06u as=2.352e+11p ps=2.24e+06u
M1002 VGND B_N a_27_368# VNB nlowvt w=550000u l=150000u
+  ad=9.5555e+11p pd=7.08e+06u as=1.5675e+11p ps=1.67e+06u
M1003 a_187_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=2.208e+11p pd=1.97e+06u as=0p ps=0u
M1004 X a_187_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 VGND a_187_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_473_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_27_368# a_187_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_187_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=5.432e+11p ps=3.21e+06u
M1009 X a_187_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


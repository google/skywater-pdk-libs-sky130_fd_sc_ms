* File: sky130_fd_sc_ms__ebufn_2.spice
* Created: Fri Aug 28 17:31:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__ebufn_2.pex.spice"
.subckt sky130_fd_sc_ms__ebufn_2  VNB VPB TE_B A Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1008 N_Z_M1008_d N_A_84_48#_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 N_Z_M1008_d N_A_84_48#_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.15355 PD=1.02 PS=1.155 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_283_48#_M1002_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.15355 PD=1.025 PS=1.155 NRD=0.804 NRS=10.536 M=1
+ R=4.93333 SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1002_d N_A_283_48#_M1003_g N_A_27_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.2109 PD=1.025 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_TE_B_M1011_g N_A_283_48#_M1011_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_84_48#_M1000_d N_A_M1000_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_33_368#_M1005_d N_A_84_48#_M1005_g N_Z_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.2 SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1007 N_A_33_368#_M1007_d N_A_84_48#_M1007_g N_Z_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_TE_B_M1004_g N_A_33_368#_M1007_d VPB PSHORT L=0.18
+ W=1.12 AD=0.27395 AS=0.1792 PD=1.75 PS=1.44 NRD=33.3324 NRS=0 M=1 R=6.22222
+ SA=90001.2 SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1004_d N_TE_B_M1006_g N_A_33_368#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.27395 AS=0.3136 PD=1.75 PS=2.8 NRD=33.3324 NRS=0 M=1 R=6.22222
+ SA=90001.8 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1001_d N_TE_B_M1001_g N_A_283_48#_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.235 AS=0.28 PD=1.47 PS=2.56 NRD=13.7703 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1010 N_A_84_48#_M1010_d N_A_M1010_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.235 PD=2.56 PS=1.47 NRD=0 NRS=23.6203 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__ebufn_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand4b_4.pxi.spice
* Created: Wed Sep  2 12:14:44 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4B_4%A_N N_A_N_M1023_g N_A_N_c_123_n N_A_N_M1018_g
+ N_A_N_c_120_n N_A_N_c_125_n N_A_N_M1022_g A_N A_N N_A_N_c_122_n
+ PM_SKY130_FD_SC_MS__NAND4B_4%A_N
x_PM_SKY130_FD_SC_MS__NAND4B_4%A_27_158# N_A_27_158#_M1023_s N_A_27_158#_M1018_d
+ N_A_27_158#_c_162_n N_A_27_158#_M1005_g N_A_27_158#_c_163_n
+ N_A_27_158#_c_164_n N_A_27_158#_c_165_n N_A_27_158#_M1011_g
+ N_A_27_158#_M1002_g N_A_27_158#_c_166_n N_A_27_158#_M1024_g
+ N_A_27_158#_c_167_n N_A_27_158#_M1025_g N_A_27_158#_c_174_n
+ N_A_27_158#_M1004_g N_A_27_158#_c_168_n N_A_27_158#_c_169_n
+ N_A_27_158#_c_175_n N_A_27_158#_c_170_n N_A_27_158#_c_171_n
+ N_A_27_158#_c_196_n N_A_27_158#_c_172_n PM_SKY130_FD_SC_MS__NAND4B_4%A_27_158#
x_PM_SKY130_FD_SC_MS__NAND4B_4%B N_B_M1003_g N_B_M1009_g N_B_M1019_g N_B_M1016_g
+ N_B_M1021_g N_B_M1020_g B N_B_c_267_n N_B_c_264_n
+ PM_SKY130_FD_SC_MS__NAND4B_4%B
x_PM_SKY130_FD_SC_MS__NAND4B_4%C N_C_M1000_g N_C_M1008_g N_C_M1012_g N_C_M1013_g
+ N_C_M1017_g N_C_M1026_g C C C C C C N_C_c_330_n PM_SKY130_FD_SC_MS__NAND4B_4%C
x_PM_SKY130_FD_SC_MS__NAND4B_4%D N_D_M1001_g N_D_c_394_n N_D_c_395_n N_D_M1007_g
+ N_D_M1014_g N_D_M1006_g N_D_M1010_g N_D_M1015_g N_D_c_401_n D D D N_D_c_403_n
+ N_D_c_404_n PM_SKY130_FD_SC_MS__NAND4B_4%D
x_PM_SKY130_FD_SC_MS__NAND4B_4%VPWR N_VPWR_M1018_s N_VPWR_M1022_s N_VPWR_M1004_s
+ N_VPWR_M1020_s N_VPWR_M1017_d N_VPWR_M1010_s N_VPWR_c_464_n N_VPWR_c_465_n
+ N_VPWR_c_466_n N_VPWR_c_467_n VPWR N_VPWR_c_468_n N_VPWR_c_469_n
+ N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n
+ N_VPWR_c_475_n N_VPWR_c_476_n N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_463_n
+ PM_SKY130_FD_SC_MS__NAND4B_4%VPWR
x_PM_SKY130_FD_SC_MS__NAND4B_4%Y N_Y_M1005_s N_Y_M1024_s N_Y_M1002_d N_Y_M1016_d
+ N_Y_M1012_s N_Y_M1006_d N_Y_c_544_n N_Y_c_561_n N_Y_c_548_n N_Y_c_545_n
+ N_Y_c_549_n N_Y_c_583_n N_Y_c_550_n N_Y_c_602_n N_Y_c_612_n N_Y_c_551_n
+ N_Y_c_568_n N_Y_c_573_n N_Y_c_552_n N_Y_c_604_n Y N_Y_c_546_n Y
+ PM_SKY130_FD_SC_MS__NAND4B_4%Y
x_PM_SKY130_FD_SC_MS__NAND4B_4%VGND N_VGND_M1023_d N_VGND_M1001_d N_VGND_M1014_d
+ N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n VGND N_VGND_c_658_n
+ N_VGND_c_659_n N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n
+ N_VGND_c_664_n N_VGND_c_665_n PM_SKY130_FD_SC_MS__NAND4B_4%VGND
x_PM_SKY130_FD_SC_MS__NAND4B_4%A_225_74# N_A_225_74#_M1005_d N_A_225_74#_M1011_d
+ N_A_225_74#_M1025_d N_A_225_74#_M1009_d N_A_225_74#_M1021_d
+ N_A_225_74#_c_746_n N_A_225_74#_c_755_n N_A_225_74#_c_747_n
+ N_A_225_74#_c_781_n N_A_225_74#_c_748_n N_A_225_74#_c_749_n
+ N_A_225_74#_c_750_n PM_SKY130_FD_SC_MS__NAND4B_4%A_225_74#
x_PM_SKY130_FD_SC_MS__NAND4B_4%A_656_74# N_A_656_74#_M1003_s N_A_656_74#_M1019_s
+ N_A_656_74#_M1000_d N_A_656_74#_M1013_d N_A_656_74#_c_802_n
+ N_A_656_74#_c_803_n N_A_656_74#_c_804_n N_A_656_74#_c_805_n
+ PM_SKY130_FD_SC_MS__NAND4B_4%A_656_74#
x_PM_SKY130_FD_SC_MS__NAND4B_4%A_1025_158# N_A_1025_158#_M1000_s
+ N_A_1025_158#_M1008_s N_A_1025_158#_M1026_s N_A_1025_158#_M1007_s
+ N_A_1025_158#_M1015_s N_A_1025_158#_c_847_n N_A_1025_158#_c_848_n
+ N_A_1025_158#_c_849_n N_A_1025_158#_c_850_n N_A_1025_158#_c_851_n
+ N_A_1025_158#_c_852_n N_A_1025_158#_c_853_n N_A_1025_158#_c_854_n
+ N_A_1025_158#_c_855_n N_A_1025_158#_c_856_n N_A_1025_158#_c_857_n
+ PM_SKY130_FD_SC_MS__NAND4B_4%A_1025_158#
cc_1 VNB N_A_N_M1023_g 0.0333164f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_N_c_120_n 0.0169027f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.65
cc_3 VNB A_N 0.0150716f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_N_c_122_n 0.0690338f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.512
cc_5 VNB N_A_27_158#_c_162_n 0.0165976f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.26
cc_6 VNB N_A_27_158#_c_163_n 0.0132022f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.725
cc_7 VNB N_A_27_158#_c_164_n 0.00931297f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.26
cc_8 VNB N_A_27_158#_c_165_n 0.0142122f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.26
cc_9 VNB N_A_27_158#_c_166_n 0.0140099f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.512
cc_10 VNB N_A_27_158#_c_167_n 0.0138142f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.512
cc_11 VNB N_A_27_158#_c_168_n 0.0153016f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_12 VNB N_A_27_158#_c_169_n 0.00671405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_158#_c_170_n 0.00780183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_158#_c_171_n 0.0169482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_158#_c_172_n 0.0723198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1003_g 0.0226992f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_17 VNB N_B_M1009_g 0.022168f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.26
cc_18 VNB N_B_M1019_g 0.022142f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.26
cc_19 VNB N_B_M1021_g 0.0286524f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.512
cc_20 VNB N_B_c_264_n 0.0859529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_M1000_g 0.0332392f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_22 VNB N_C_M1008_g 0.0230318f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.26
cc_23 VNB N_C_M1013_g 0.0230618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_M1026_g 0.0237321f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.512
cc_25 VNB C 0.0205651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C_c_330_n 0.0699767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_D_M1001_g 0.0205853f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_28 VNB N_D_c_394_n 0.0146865f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.725
cc_29 VNB N_D_c_395_n 0.00900825f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.26
cc_30 VNB N_D_M1007_g 0.0203441f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.65
cc_31 VNB N_D_M1014_g 0.021724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_D_M1006_g 0.00178153f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.512
cc_33 VNB N_D_M1010_g 0.00178153f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.512
cc_34 VNB N_D_M1015_g 0.0310968f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.54
cc_35 VNB N_D_c_401_n 0.00735939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB D 0.0169158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_D_c_403_n 0.0149615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_D_c_404_n 0.0766171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_463_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_544_n 0.0055499f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.512
cc_41 VNB N_Y_c_545_n 0.0186163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_546_n 0.0055714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB Y 0.00320909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_655_n 0.00863836f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.26
cc_45 VNB N_VGND_c_656_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_657_n 0.00617711f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.465
cc_47 VNB N_VGND_c_658_n 0.0193283f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_48 VNB N_VGND_c_659_n 0.154047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_660_n 0.0150174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_661_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_662_n 0.486338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_663_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_664_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_665_n 0.00702348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_225_74#_c_746_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_225_74#_c_747_n 0.00523745f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.512
cc_57 VNB N_A_225_74#_c_748_n 0.00250726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_225_74#_c_749_n 0.00795952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_225_74#_c_750_n 0.00161948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_656_74#_c_802_n 0.0263677f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_61 VNB N_A_656_74#_c_803_n 0.00264577f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.512
cc_62 VNB N_A_656_74#_c_804_n 0.0019256f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.465
cc_63 VNB N_A_656_74#_c_805_n 0.00243302f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.512
cc_64 VNB N_A_1025_158#_c_847_n 0.00248004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1025_158#_c_848_n 0.00187418f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=1.512
cc_66 VNB N_A_1025_158#_c_849_n 0.0044611f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_67 VNB N_A_1025_158#_c_850_n 0.00195975f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_68 VNB N_A_1025_158#_c_851_n 0.0123218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1025_158#_c_852_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1025_158#_c_853_n 0.00802292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1025_158#_c_854_n 0.00189026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1025_158#_c_855_n 0.00348098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1025_158#_c_856_n 0.00207621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1025_158#_c_857_n 0.00255592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VPB N_A_N_c_123_n 0.0207886f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.725
cc_76 VPB N_A_N_c_120_n 0.00702868f $X=-0.19 $Y=1.66 $X2=1.305 $Y2=1.65
cc_77 VPB N_A_N_c_125_n 0.0192165f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.725
cc_78 VPB A_N 0.0231175f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_79 VPB N_A_N_c_122_n 0.0280141f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.512
cc_80 VPB N_A_27_158#_M1002_g 0.027319f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.512
cc_81 VPB N_A_27_158#_c_174_n 0.0225058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_27_158#_c_175_n 0.0035517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_27_158#_c_170_n 0.00492307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_27_158#_c_172_n 0.0231513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_B_M1016_g 0.0249274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_B_M1020_g 0.0257075f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.512
cc_87 VPB N_B_c_267_n 0.0112877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_B_c_264_n 0.0326459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_C_M1012_g 0.0287155f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.26
cc_90 VPB N_C_M1017_g 0.028744f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.512
cc_91 VPB C 0.0265354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_C_c_330_n 0.0302347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_D_M1006_g 0.026917f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.512
cc_94 VPB N_D_M1010_g 0.0261603f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.512
cc_95 VPB D 0.0165945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_464_n 0.0652448f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.465
cc_97 VPB N_VPWR_c_465_n 0.0169263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_466_n 0.0128241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_467_n 0.0118994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_468_n 0.0182134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_469_n 0.0208961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_470_n 0.0160859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_471_n 0.0178937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_472_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_473_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_474_n 0.0259773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_475_n 0.0383574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_476_n 0.0319815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_477_n 0.0252488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_478_n 0.034283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_463_n 0.0985303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_Y_c_548_n 0.00598444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_Y_c_549_n 0.00224521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_Y_c_550_n 0.00574731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_Y_c_551_n 0.00239158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_Y_c_552_n 0.0017422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB Y 0.00171176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 N_A_N_c_120_n N_A_27_158#_c_164_n 0.00415792f $X=1.305 $Y=1.65 $X2=0
+ $Y2=0
cc_119 N_A_N_c_122_n N_A_27_158#_c_164_n 0.00104584f $X=1.035 $Y=1.512 $X2=0
+ $Y2=0
cc_120 N_A_N_c_125_n N_A_27_158#_M1002_g 0.0111617f $X=1.395 $Y=1.725 $X2=0
+ $Y2=0
cc_121 N_A_N_M1023_g N_A_27_158#_c_168_n 0.0132267f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_122 A_N N_A_27_158#_c_168_n 0.0297062f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A_N_c_122_n N_A_27_158#_c_168_n 0.0132438f $X=1.035 $Y=1.512 $X2=0
+ $Y2=0
cc_124 N_A_N_M1023_g N_A_27_158#_c_169_n 0.00473994f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_125 A_N N_A_27_158#_c_169_n 0.0102955f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A_N_c_122_n N_A_27_158#_c_169_n 0.00507609f $X=1.035 $Y=1.512 $X2=0
+ $Y2=0
cc_127 N_A_N_c_123_n N_A_27_158#_c_175_n 0.0208586f $X=0.945 $Y=1.725 $X2=0
+ $Y2=0
cc_128 N_A_N_c_120_n N_A_27_158#_c_175_n 0.00417844f $X=1.305 $Y=1.65 $X2=0
+ $Y2=0
cc_129 N_A_N_c_125_n N_A_27_158#_c_175_n 0.0167379f $X=1.395 $Y=1.725 $X2=0
+ $Y2=0
cc_130 A_N N_A_27_158#_c_175_n 0.00809884f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A_N_c_122_n N_A_27_158#_c_175_n 7.38215e-19 $X=1.035 $Y=1.512 $X2=0
+ $Y2=0
cc_132 N_A_N_c_120_n N_A_27_158#_c_170_n 0.011598f $X=1.305 $Y=1.65 $X2=0 $Y2=0
cc_133 N_A_N_M1023_g N_A_27_158#_c_171_n 0.0104346f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_134 A_N N_A_27_158#_c_171_n 0.0263292f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A_N_c_122_n N_A_27_158#_c_171_n 0.00613351f $X=1.035 $Y=1.512 $X2=0
+ $Y2=0
cc_136 N_A_N_c_120_n N_A_27_158#_c_196_n 0.00990809f $X=1.305 $Y=1.65 $X2=0
+ $Y2=0
cc_137 A_N N_A_27_158#_c_196_n 0.0212325f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A_N_c_122_n N_A_27_158#_c_196_n 0.0079642f $X=1.035 $Y=1.512 $X2=0
+ $Y2=0
cc_139 N_A_N_c_120_n N_A_27_158#_c_172_n 0.0111617f $X=1.305 $Y=1.65 $X2=0 $Y2=0
cc_140 N_A_N_c_123_n N_VPWR_c_464_n 0.00600499f $X=0.945 $Y=1.725 $X2=0 $Y2=0
cc_141 A_N N_VPWR_c_464_n 0.0276508f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A_N_c_122_n N_VPWR_c_464_n 0.00213732f $X=1.035 $Y=1.512 $X2=0 $Y2=0
cc_143 N_A_N_c_125_n N_VPWR_c_465_n 0.00776524f $X=1.395 $Y=1.725 $X2=0 $Y2=0
cc_144 N_A_N_c_123_n N_VPWR_c_469_n 0.00465228f $X=0.945 $Y=1.725 $X2=0 $Y2=0
cc_145 N_A_N_c_125_n N_VPWR_c_469_n 0.00465228f $X=1.395 $Y=1.725 $X2=0 $Y2=0
cc_146 N_A_N_c_123_n N_VPWR_c_463_n 0.00555093f $X=0.945 $Y=1.725 $X2=0 $Y2=0
cc_147 N_A_N_c_125_n N_VPWR_c_463_n 0.00555093f $X=1.395 $Y=1.725 $X2=0 $Y2=0
cc_148 N_A_N_M1023_g N_VGND_c_655_n 0.0191059f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_N_M1023_g N_VGND_c_658_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_N_M1023_g N_VGND_c_662_n 0.00687202f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_N_M1023_g N_A_225_74#_c_749_n 8.50533e-19 $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_27_158#_c_167_n N_B_M1003_g 0.0245946f $X=2.775 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_27_158#_c_170_n N_B_c_267_n 0.0139961f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_27_158#_c_172_n N_B_c_267_n 0.00413082f $X=2.775 $Y=1.477 $X2=0 $Y2=0
cc_155 N_A_27_158#_c_170_n N_B_c_264_n 0.00111951f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A_27_158#_c_172_n N_B_c_264_n 0.0245946f $X=2.775 $Y=1.477 $X2=0 $Y2=0
cc_157 N_A_27_158#_c_175_n N_VPWR_c_464_n 0.0289323f $X=1.17 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_27_158#_M1002_g N_VPWR_c_465_n 0.0221499f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_27_158#_c_175_n N_VPWR_c_465_n 0.0281499f $X=1.17 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_27_158#_c_170_n N_VPWR_c_465_n 0.02503f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A_27_158#_c_175_n N_VPWR_c_469_n 0.00657675f $X=1.17 $Y=1.985 $X2=0
+ $Y2=0
cc_162 N_A_27_158#_M1002_g N_VPWR_c_474_n 0.00460063f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_27_158#_c_174_n N_VPWR_c_474_n 0.00460063f $X=2.79 $Y=1.77 $X2=0
+ $Y2=0
cc_164 N_A_27_158#_c_174_n N_VPWR_c_475_n 0.0188265f $X=2.79 $Y=1.77 $X2=0 $Y2=0
cc_165 N_A_27_158#_M1002_g N_VPWR_c_463_n 0.00911461f $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_27_158#_c_174_n N_VPWR_c_463_n 0.00906823f $X=2.79 $Y=1.77 $X2=0
+ $Y2=0
cc_167 N_A_27_158#_c_175_n N_VPWR_c_463_n 0.00992028f $X=1.17 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_27_158#_c_162_n N_Y_c_544_n 0.00678753f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_27_158#_c_163_n N_Y_c_544_n 0.00241988f $X=1.84 $Y=1.26 $X2=0 $Y2=0
cc_170 N_A_27_158#_c_165_n N_Y_c_544_n 0.0127999f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_171 N_A_27_158#_c_166_n N_Y_c_544_n 0.012572f $X=2.345 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A_27_158#_c_168_n N_Y_c_544_n 0.0130492f $X=1.005 $Y=1.045 $X2=0 $Y2=0
cc_173 N_A_27_158#_c_170_n N_Y_c_544_n 0.0427778f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A_27_158#_c_172_n N_Y_c_544_n 0.00308687f $X=2.775 $Y=1.477 $X2=0 $Y2=0
cc_175 N_A_27_158#_c_170_n N_Y_c_561_n 0.0481643f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A_27_158#_c_172_n N_Y_c_561_n 0.013283f $X=2.775 $Y=1.477 $X2=0 $Y2=0
cc_177 N_A_27_158#_M1002_g N_Y_c_548_n 4.5815e-19 $X=1.93 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A_27_158#_c_174_n N_Y_c_548_n 4.57751e-19 $X=2.79 $Y=1.77 $X2=0 $Y2=0
cc_179 N_A_27_158#_c_167_n N_Y_c_545_n 0.00620792f $X=2.775 $Y=1.185 $X2=0 $Y2=0
cc_180 N_A_27_158#_c_170_n N_Y_c_545_n 0.0087312f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A_27_158#_c_172_n N_Y_c_545_n 0.00465633f $X=2.775 $Y=1.477 $X2=0 $Y2=0
cc_182 N_A_27_158#_c_165_n N_Y_c_568_n 0.00118267f $X=1.915 $Y=1.185 $X2=0 $Y2=0
cc_183 N_A_27_158#_c_166_n N_Y_c_568_n 0.00934096f $X=2.345 $Y=1.185 $X2=0 $Y2=0
cc_184 N_A_27_158#_c_167_n N_Y_c_568_n 0.00968259f $X=2.775 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A_27_158#_c_170_n N_Y_c_568_n 0.0256206f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A_27_158#_c_172_n N_Y_c_568_n 0.0131921f $X=2.775 $Y=1.477 $X2=0 $Y2=0
cc_187 N_A_27_158#_c_174_n N_Y_c_573_n 0.0174211f $X=2.79 $Y=1.77 $X2=0 $Y2=0
cc_188 N_A_27_158#_c_170_n N_Y_c_573_n 0.00579184f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A_27_158#_c_168_n N_VGND_M1023_d 0.00350363f $X=1.005 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_190 N_A_27_158#_c_162_n N_VGND_c_655_n 0.00117816f $X=1.485 $Y=1.185 $X2=0
+ $Y2=0
cc_191 N_A_27_158#_c_168_n N_VGND_c_655_n 0.0126491f $X=1.005 $Y=1.045 $X2=0
+ $Y2=0
cc_192 N_A_27_158#_c_162_n N_VGND_c_659_n 0.00279469f $X=1.485 $Y=1.185 $X2=0
+ $Y2=0
cc_193 N_A_27_158#_c_165_n N_VGND_c_659_n 0.00278247f $X=1.915 $Y=1.185 $X2=0
+ $Y2=0
cc_194 N_A_27_158#_c_166_n N_VGND_c_659_n 0.00278271f $X=2.345 $Y=1.185 $X2=0
+ $Y2=0
cc_195 N_A_27_158#_c_167_n N_VGND_c_659_n 0.00278271f $X=2.775 $Y=1.185 $X2=0
+ $Y2=0
cc_196 N_A_27_158#_c_162_n N_VGND_c_662_n 0.00357517f $X=1.485 $Y=1.185 $X2=0
+ $Y2=0
cc_197 N_A_27_158#_c_165_n N_VGND_c_662_n 0.00353427f $X=1.915 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_A_27_158#_c_166_n N_VGND_c_662_n 0.00353428f $X=2.345 $Y=1.185 $X2=0
+ $Y2=0
cc_199 N_A_27_158#_c_167_n N_VGND_c_662_n 0.00353526f $X=2.775 $Y=1.185 $X2=0
+ $Y2=0
cc_200 N_A_27_158#_c_171_n N_VGND_c_662_n 0.0127184f $X=0.28 $Y=0.95 $X2=0 $Y2=0
cc_201 N_A_27_158#_c_168_n N_A_225_74#_M1005_d 0.00511261f $X=1.005 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_202 N_A_27_158#_c_162_n N_A_225_74#_c_746_n 0.0101479f $X=1.485 $Y=1.185
+ $X2=0 $Y2=0
cc_203 N_A_27_158#_c_165_n N_A_225_74#_c_746_n 0.00750248f $X=1.915 $Y=1.185
+ $X2=0 $Y2=0
cc_204 N_A_27_158#_c_162_n N_A_225_74#_c_755_n 8.39771e-19 $X=1.485 $Y=1.185
+ $X2=0 $Y2=0
cc_205 N_A_27_158#_c_165_n N_A_225_74#_c_755_n 0.00528291f $X=1.915 $Y=1.185
+ $X2=0 $Y2=0
cc_206 N_A_27_158#_c_166_n N_A_225_74#_c_747_n 0.00966901f $X=2.345 $Y=1.185
+ $X2=0 $Y2=0
cc_207 N_A_27_158#_c_167_n N_A_225_74#_c_747_n 0.0105758f $X=2.775 $Y=1.185
+ $X2=0 $Y2=0
cc_208 N_A_27_158#_c_162_n N_A_225_74#_c_749_n 0.00937192f $X=1.485 $Y=1.185
+ $X2=0 $Y2=0
cc_209 N_A_27_158#_c_165_n N_A_225_74#_c_749_n 9.20446e-19 $X=1.915 $Y=1.185
+ $X2=0 $Y2=0
cc_210 N_A_27_158#_c_168_n N_A_225_74#_c_749_n 0.0152408f $X=1.005 $Y=1.045
+ $X2=0 $Y2=0
cc_211 N_A_27_158#_c_165_n N_A_225_74#_c_750_n 0.00187501f $X=1.915 $Y=1.185
+ $X2=0 $Y2=0
cc_212 N_B_c_264_n C 0.00700821f $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_213 N_B_c_264_n N_C_c_330_n 0.00425553f $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_214 N_B_M1016_g N_VPWR_c_470_n 0.00460063f $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_215 N_B_M1020_g N_VPWR_c_470_n 0.00461464f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_216 N_B_M1016_g N_VPWR_c_475_n 0.0153729f $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_217 N_B_M1020_g N_VPWR_c_475_n 5.15764e-19 $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_218 N_B_M1016_g N_VPWR_c_476_n 5.05806e-19 $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_219 N_B_M1020_g N_VPWR_c_476_n 0.0151413f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_220 N_B_M1016_g N_VPWR_c_463_n 0.00903917f $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B_M1020_g N_VPWR_c_463_n 0.00908554f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B_M1003_g N_Y_c_545_n 0.0104262f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B_M1009_g N_Y_c_545_n 0.0104864f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_224 N_B_M1019_g N_Y_c_545_n 0.0104262f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B_M1021_g N_Y_c_545_n 0.00328941f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B_c_267_n N_Y_c_545_n 0.0748019f $X=3.295 $Y=1.515 $X2=0 $Y2=0
cc_227 N_B_c_264_n N_Y_c_545_n 0.00922038f $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_228 N_B_M1016_g N_Y_c_549_n 3.75297e-19 $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B_M1020_g N_Y_c_549_n 3.80419e-19 $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_230 N_B_M1020_g N_Y_c_583_n 0.0148668f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_231 N_B_M1003_g N_Y_c_568_n 0.00100316f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B_M1016_g N_Y_c_573_n 0.0168449f $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_233 N_B_c_267_n N_Y_c_573_n 0.0780115f $X=3.295 $Y=1.515 $X2=0 $Y2=0
cc_234 N_B_c_264_n N_Y_c_573_n 0.00536498f $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_235 N_B_M1016_g N_Y_c_552_n 0.00853921f $X=4.25 $Y=2.4 $X2=0 $Y2=0
cc_236 N_B_M1020_g N_Y_c_552_n 0.0105426f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_237 N_B_c_264_n N_Y_c_552_n 8.76085e-19 $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_238 N_B_M1021_g N_Y_c_546_n 0.0065941f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B_M1019_g Y 5.28058e-19 $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B_M1021_g Y 0.00366525f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B_M1020_g Y 0.0052722f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_242 N_B_c_267_n Y 0.0179388f $X=3.295 $Y=1.515 $X2=0 $Y2=0
cc_243 N_B_c_264_n Y 0.0229886f $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B_M1003_g N_VGND_c_659_n 0.00329872f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B_M1009_g N_VGND_c_659_n 0.00288916f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B_M1019_g N_VGND_c_659_n 0.00288916f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B_M1021_g N_VGND_c_659_n 0.00288916f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B_M1003_g N_VGND_c_662_n 0.00428036f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B_M1009_g N_VGND_c_662_n 0.0035719f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B_M1019_g N_VGND_c_662_n 0.0035719f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B_M1021_g N_VGND_c_662_n 0.00362189f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B_M1003_g N_A_225_74#_c_747_n 0.00295514f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B_M1003_g N_A_225_74#_c_748_n 0.0106614f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B_M1009_g N_A_225_74#_c_748_n 0.00838518f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B_M1019_g N_A_225_74#_c_748_n 0.00841805f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B_M1021_g N_A_225_74#_c_748_n 0.00842664f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B_c_264_n N_A_225_74#_c_748_n 0.00397412f $X=4.495 $Y=1.515 $X2=0 $Y2=0
cc_258 N_B_M1003_g N_A_656_74#_c_802_n 0.00357851f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_259 N_B_M1009_g N_A_656_74#_c_802_n 0.0103107f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B_M1019_g N_A_656_74#_c_802_n 0.0103107f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B_M1021_g N_A_656_74#_c_802_n 0.013323f $X=4.495 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B_M1021_g N_A_1025_158#_c_853_n 0.00326063f $X=4.495 $Y=0.74 $X2=0
+ $Y2=0
cc_263 N_C_M1026_g N_D_M1001_g 0.0119435f $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_264 C N_D_c_394_n 0.0128675f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_265 C N_D_c_395_n 0.00806403f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_266 N_C_c_330_n N_D_c_395_n 0.0119435f $X=6.79 $Y=1.515 $X2=0 $Y2=0
cc_267 C D 0.0296351f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_268 C N_D_c_404_n 0.00166444f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_269 N_C_M1012_g N_VPWR_c_476_n 0.0187634f $X=5.945 $Y=2.4 $X2=0 $Y2=0
cc_270 N_C_M1012_g N_VPWR_c_477_n 0.00461464f $X=5.945 $Y=2.4 $X2=0 $Y2=0
cc_271 N_C_M1017_g N_VPWR_c_477_n 0.00460063f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_272 N_C_M1017_g N_VPWR_c_478_n 0.0187373f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_273 N_C_M1012_g N_VPWR_c_463_n 0.00911317f $X=5.945 $Y=2.4 $X2=0 $Y2=0
cc_274 N_C_M1017_g N_VPWR_c_463_n 0.0090668f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_275 N_C_M1012_g N_Y_c_583_n 0.0163793f $X=5.945 $Y=2.4 $X2=0 $Y2=0
cc_276 C N_Y_c_583_n 0.0864049f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_277 N_C_c_330_n N_Y_c_583_n 0.00229929f $X=6.79 $Y=1.515 $X2=0 $Y2=0
cc_278 N_C_M1012_g N_Y_c_550_n 3.07561e-19 $X=5.945 $Y=2.4 $X2=0 $Y2=0
cc_279 N_C_M1017_g N_Y_c_550_n 3.08235e-19 $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_280 N_C_M1017_g N_Y_c_602_n 0.0163499f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_281 C N_Y_c_602_n 0.0670722f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_282 C N_Y_c_604_n 0.0499482f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_283 N_C_c_330_n N_Y_c_604_n 0.00287383f $X=6.79 $Y=1.515 $X2=0 $Y2=0
cc_284 C Y 0.0263965f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_285 N_C_M1026_g N_VGND_c_656_n 6.33938e-19 $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_286 N_C_M1000_g N_VGND_c_659_n 0.00288893f $X=5.485 $Y=0.74 $X2=0 $Y2=0
cc_287 N_C_M1008_g N_VGND_c_659_n 0.00288916f $X=5.915 $Y=0.74 $X2=0 $Y2=0
cc_288 N_C_M1013_g N_VGND_c_659_n 0.00290044f $X=6.345 $Y=0.74 $X2=0 $Y2=0
cc_289 N_C_M1026_g N_VGND_c_659_n 0.00451103f $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_290 N_C_M1000_g N_VGND_c_662_n 0.00362175f $X=5.485 $Y=0.74 $X2=0 $Y2=0
cc_291 N_C_M1008_g N_VGND_c_662_n 0.0035719f $X=5.915 $Y=0.74 $X2=0 $Y2=0
cc_292 N_C_M1013_g N_VGND_c_662_n 0.00356391f $X=6.345 $Y=0.74 $X2=0 $Y2=0
cc_293 N_C_M1026_g N_VGND_c_662_n 0.00876431f $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_294 N_C_M1000_g N_A_225_74#_c_748_n 3.60088e-19 $X=5.485 $Y=0.74 $X2=0 $Y2=0
cc_295 N_C_M1000_g N_A_656_74#_c_802_n 0.0124709f $X=5.485 $Y=0.74 $X2=0 $Y2=0
cc_296 N_C_M1008_g N_A_656_74#_c_803_n 0.011702f $X=5.915 $Y=0.74 $X2=0 $Y2=0
cc_297 N_C_M1013_g N_A_656_74#_c_803_n 0.0118633f $X=6.345 $Y=0.74 $X2=0 $Y2=0
cc_298 N_C_M1000_g N_A_656_74#_c_804_n 0.00270258f $X=5.485 $Y=0.74 $X2=0 $Y2=0
cc_299 N_C_M1008_g N_A_656_74#_c_805_n 7.20203e-19 $X=5.915 $Y=0.74 $X2=0 $Y2=0
cc_300 N_C_M1013_g N_A_656_74#_c_805_n 0.00731775f $X=6.345 $Y=0.74 $X2=0 $Y2=0
cc_301 N_C_M1026_g N_A_656_74#_c_805_n 0.00676657f $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_302 N_C_M1000_g N_A_1025_158#_c_847_n 0.00911542f $X=5.485 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_C_M1008_g N_A_1025_158#_c_847_n 0.00915993f $X=5.915 $Y=0.74 $X2=0
+ $Y2=0
cc_304 C N_A_1025_158#_c_847_n 0.0325459f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_305 N_C_c_330_n N_A_1025_158#_c_847_n 0.0021687f $X=6.79 $Y=1.515 $X2=0 $Y2=0
cc_306 N_C_M1026_g N_A_1025_158#_c_848_n 3.34174e-19 $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_307 C N_A_1025_158#_c_849_n 0.0237998f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_308 N_C_M1000_g N_A_1025_158#_c_853_n 0.00532122f $X=5.485 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_C_M1008_g N_A_1025_158#_c_853_n 6.3885e-19 $X=5.915 $Y=0.74 $X2=0 $Y2=0
cc_310 C N_A_1025_158#_c_853_n 0.0232973f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_311 N_C_M1000_g N_A_1025_158#_c_854_n 8.87619e-19 $X=5.485 $Y=0.74 $X2=0
+ $Y2=0
cc_312 N_C_M1008_g N_A_1025_158#_c_854_n 0.00638082f $X=5.915 $Y=0.74 $X2=0
+ $Y2=0
cc_313 C N_A_1025_158#_c_854_n 0.0203551f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_314 N_C_c_330_n N_A_1025_158#_c_854_n 0.00247032f $X=6.79 $Y=1.515 $X2=0
+ $Y2=0
cc_315 N_C_M1013_g N_A_1025_158#_c_855_n 0.00991537f $X=6.345 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_C_M1026_g N_A_1025_158#_c_855_n 0.0135723f $X=6.79 $Y=0.74 $X2=0 $Y2=0
cc_317 C N_A_1025_158#_c_855_n 0.0735753f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_318 N_C_c_330_n N_A_1025_158#_c_855_n 0.00269656f $X=6.79 $Y=1.515 $X2=0
+ $Y2=0
cc_319 N_D_M1010_g N_VPWR_c_467_n 0.00386341f $X=8.565 $Y=2.4 $X2=0 $Y2=0
cc_320 D N_VPWR_c_467_n 0.0231613f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_321 N_D_c_404_n N_VPWR_c_467_n 0.00145428f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_322 N_D_M1006_g N_VPWR_c_471_n 0.00460063f $X=8.095 $Y=2.4 $X2=0 $Y2=0
cc_323 N_D_M1010_g N_VPWR_c_471_n 0.005209f $X=8.565 $Y=2.4 $X2=0 $Y2=0
cc_324 N_D_M1006_g N_VPWR_c_478_n 0.0155248f $X=8.095 $Y=2.4 $X2=0 $Y2=0
cc_325 N_D_M1010_g N_VPWR_c_478_n 5.25645e-19 $X=8.565 $Y=2.4 $X2=0 $Y2=0
cc_326 N_D_M1006_g N_VPWR_c_463_n 0.00904118f $X=8.095 $Y=2.4 $X2=0 $Y2=0
cc_327 N_D_M1010_g N_VPWR_c_463_n 0.00985698f $X=8.565 $Y=2.4 $X2=0 $Y2=0
cc_328 N_D_c_394_n N_Y_c_602_n 0.00730719f $X=7.575 $Y=1.375 $X2=0 $Y2=0
cc_329 N_D_c_395_n N_Y_c_602_n 0.00141204f $X=7.295 $Y=1.375 $X2=0 $Y2=0
cc_330 N_D_M1006_g N_Y_c_602_n 0.0163499f $X=8.095 $Y=2.4 $X2=0 $Y2=0
cc_331 D N_Y_c_602_n 0.0285459f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_332 N_D_c_403_n N_Y_c_602_n 6.24251e-19 $X=8.005 $Y=1.465 $X2=0 $Y2=0
cc_333 N_D_M1010_g N_Y_c_612_n 0.00242423f $X=8.565 $Y=2.4 $X2=0 $Y2=0
cc_334 D N_Y_c_612_n 0.0218221f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_335 N_D_c_404_n N_Y_c_612_n 6.08557e-19 $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_336 N_D_M1010_g N_Y_c_551_n 0.0106141f $X=8.565 $Y=2.4 $X2=0 $Y2=0
cc_337 N_D_M1001_g N_VGND_c_656_n 0.00936142f $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_338 N_D_M1007_g N_VGND_c_656_n 0.00924442f $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_339 N_D_M1014_g N_VGND_c_656_n 4.47062e-19 $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_340 N_D_M1007_g N_VGND_c_657_n 4.46513e-19 $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_341 N_D_M1014_g N_VGND_c_657_n 0.0095322f $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_342 N_D_M1015_g N_VGND_c_657_n 0.0057749f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_343 N_D_M1001_g N_VGND_c_659_n 0.00383152f $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_344 N_D_M1007_g N_VGND_c_660_n 0.00383152f $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_345 N_D_M1014_g N_VGND_c_660_n 0.00383152f $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_346 N_D_M1015_g N_VGND_c_661_n 0.00434272f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_347 N_D_M1001_g N_VGND_c_662_n 0.00757637f $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_348 N_D_M1007_g N_VGND_c_662_n 0.0075754f $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_349 N_D_M1014_g N_VGND_c_662_n 0.0075754f $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_350 N_D_M1015_g N_VGND_c_662_n 0.00824755f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_351 N_D_M1001_g N_A_656_74#_c_805_n 2.08848e-19 $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_352 N_D_M1001_g N_A_1025_158#_c_848_n 3.33944e-19 $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_353 N_D_M1001_g N_A_1025_158#_c_849_n 0.010673f $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_354 N_D_c_394_n N_A_1025_158#_c_849_n 0.0019675f $X=7.575 $Y=1.375 $X2=0
+ $Y2=0
cc_355 N_D_M1007_g N_A_1025_158#_c_849_n 0.0164691f $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_356 N_D_M1007_g N_A_1025_158#_c_850_n 3.34629e-19 $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_357 N_D_M1014_g N_A_1025_158#_c_850_n 3.34629e-19 $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_358 N_D_M1014_g N_A_1025_158#_c_851_n 0.0131094f $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_359 N_D_M1015_g N_A_1025_158#_c_851_n 0.012892f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_360 D N_A_1025_158#_c_851_n 0.0826332f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_361 N_D_c_404_n N_A_1025_158#_c_851_n 0.0123393f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_362 N_D_M1014_g N_A_1025_158#_c_852_n 8.80469e-19 $X=8.08 $Y=0.74 $X2=0 $Y2=0
cc_363 N_D_M1015_g N_A_1025_158#_c_852_n 0.00983615f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_D_M1001_g N_A_1025_158#_c_856_n 0.00359034f $X=7.22 $Y=0.74 $X2=0 $Y2=0
cc_365 N_D_M1007_g N_A_1025_158#_c_856_n 2.36785e-19 $X=7.65 $Y=0.74 $X2=0 $Y2=0
cc_366 D N_A_1025_158#_c_857_n 0.0134174f $X=8.795 $Y=1.58 $X2=0 $Y2=0
cc_367 N_D_c_403_n N_A_1025_158#_c_857_n 0.00199624f $X=8.005 $Y=1.465 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_465_n N_Y_c_548_n 0.0316586f $X=1.705 $Y=2.015 $X2=0 $Y2=0
cc_369 N_VPWR_c_474_n N_Y_c_548_n 0.0275757f $X=2.85 $Y=2.852 $X2=0 $Y2=0
cc_370 N_VPWR_c_475_n N_Y_c_548_n 0.028554f $X=4.19 $Y=2.852 $X2=0 $Y2=0
cc_371 N_VPWR_c_463_n N_Y_c_548_n 0.0228248f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_372 N_VPWR_c_470_n N_Y_c_549_n 0.00972736f $X=4.76 $Y=3.33 $X2=0 $Y2=0
cc_373 N_VPWR_c_475_n N_Y_c_549_n 0.0284324f $X=4.19 $Y=2.852 $X2=0 $Y2=0
cc_374 N_VPWR_c_476_n N_Y_c_549_n 0.0296717f $X=4.925 $Y=2.375 $X2=0 $Y2=0
cc_375 N_VPWR_c_463_n N_Y_c_549_n 0.00805147f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_M1020_s N_Y_c_583_n 0.0281813f $X=4.79 $Y=1.84 $X2=0 $Y2=0
cc_377 N_VPWR_c_476_n N_Y_c_583_n 0.0817059f $X=4.925 $Y=2.375 $X2=0 $Y2=0
cc_378 N_VPWR_c_476_n N_Y_c_550_n 0.0284622f $X=4.925 $Y=2.375 $X2=0 $Y2=0
cc_379 N_VPWR_c_477_n N_Y_c_550_n 0.0264602f $X=6.835 $Y=2.852 $X2=0 $Y2=0
cc_380 N_VPWR_c_478_n N_Y_c_550_n 0.0292023f $X=8.035 $Y=2.852 $X2=0 $Y2=0
cc_381 N_VPWR_c_463_n N_Y_c_550_n 0.0219015f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPWR_M1017_d N_Y_c_602_n 0.0296509f $X=6.865 $Y=1.84 $X2=0 $Y2=0
cc_383 N_VPWR_c_478_n N_Y_c_602_n 0.0875729f $X=8.035 $Y=2.852 $X2=0 $Y2=0
cc_384 N_VPWR_c_467_n N_Y_c_551_n 0.0323712f $X=8.79 $Y=2.115 $X2=0 $Y2=0
cc_385 N_VPWR_c_471_n N_Y_c_551_n 0.0127641f $X=8.675 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_c_478_n N_Y_c_551_n 0.0284631f $X=8.035 $Y=2.852 $X2=0 $Y2=0
cc_387 N_VPWR_c_463_n N_Y_c_551_n 0.0104969f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_M1004_s N_Y_c_573_n 0.0368106f $X=2.88 $Y=1.84 $X2=0 $Y2=0
cc_389 N_VPWR_c_475_n N_Y_c_573_n 0.0989131f $X=4.19 $Y=2.852 $X2=0 $Y2=0
cc_390 N_Y_c_544_n N_A_225_74#_M1011_d 0.00178571f $X=2.395 $Y=1.005 $X2=0 $Y2=0
cc_391 N_Y_c_545_n N_A_225_74#_M1025_d 0.00176461f $X=4.445 $Y=1.175 $X2=0 $Y2=0
cc_392 N_Y_c_545_n N_A_225_74#_M1009_d 0.00176891f $X=4.445 $Y=1.175 $X2=0 $Y2=0
cc_393 N_Y_c_546_n N_A_225_74#_M1021_d 8.81272e-19 $X=4.56 $Y=1.26 $X2=0 $Y2=0
cc_394 N_Y_M1005_s N_A_225_74#_c_746_n 0.00285125f $X=1.56 $Y=0.37 $X2=0 $Y2=0
cc_395 N_Y_c_544_n N_A_225_74#_c_746_n 0.0106717f $X=2.395 $Y=1.005 $X2=0 $Y2=0
cc_396 N_Y_c_544_n N_A_225_74#_c_755_n 0.0152131f $X=2.395 $Y=1.005 $X2=0 $Y2=0
cc_397 N_Y_M1024_s N_A_225_74#_c_747_n 0.00176461f $X=2.42 $Y=0.37 $X2=0 $Y2=0
cc_398 N_Y_c_544_n N_A_225_74#_c_747_n 0.00391529f $X=2.395 $Y=1.005 $X2=0 $Y2=0
cc_399 N_Y_c_545_n N_A_225_74#_c_747_n 0.00271156f $X=4.445 $Y=1.175 $X2=0 $Y2=0
cc_400 N_Y_c_568_n N_A_225_74#_c_747_n 0.0160271f $X=2.56 $Y=0.86 $X2=0 $Y2=0
cc_401 N_Y_c_545_n N_A_225_74#_c_781_n 0.0134809f $X=4.445 $Y=1.175 $X2=0 $Y2=0
cc_402 N_Y_c_545_n N_A_225_74#_c_748_n 0.0682654f $X=4.445 $Y=1.175 $X2=0 $Y2=0
cc_403 N_Y_c_546_n N_A_225_74#_c_748_n 0.0133931f $X=4.56 $Y=1.26 $X2=0 $Y2=0
cc_404 N_Y_c_545_n N_A_656_74#_M1003_s 0.00176891f $X=4.445 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_405 N_Y_c_545_n N_A_656_74#_M1019_s 0.00176891f $X=4.445 $Y=1.175 $X2=0 $Y2=0
cc_406 N_Y_c_546_n N_A_1025_158#_c_853_n 0.00182029f $X=4.56 $Y=1.26 $X2=0 $Y2=0
cc_407 N_VGND_c_659_n N_A_225_74#_c_746_n 0.0333877f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_662_n N_A_225_74#_c_746_n 0.0187857f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_659_n N_A_225_74#_c_747_n 0.0556832f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_662_n N_A_225_74#_c_747_n 0.0311746f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_659_n N_A_225_74#_c_748_n 0.00197884f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_662_n N_A_225_74#_c_748_n 0.00653056f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_655_n N_A_225_74#_c_749_n 0.0232594f $X=0.71 $Y=0.515 $X2=0
+ $Y2=0
cc_414 N_VGND_c_659_n N_A_225_74#_c_749_n 0.0227371f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_662_n N_A_225_74#_c_749_n 0.0125119f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_659_n N_A_225_74#_c_750_n 0.0173119f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_662_n N_A_225_74#_c_750_n 0.00950667f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_659_n N_A_656_74#_c_802_n 0.100903f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_c_662_n N_A_656_74#_c_802_n 0.07974f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_659_n N_A_656_74#_c_803_n 0.0263582f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_662_n N_A_656_74#_c_803_n 0.0204706f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_659_n N_A_656_74#_c_804_n 0.0119499f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_662_n N_A_656_74#_c_804_n 0.00939712f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_656_n N_A_656_74#_c_805_n 5.76843e-19 $X=7.435 $Y=0.615 $X2=0
+ $Y2=0
cc_425 N_VGND_c_659_n N_A_656_74#_c_805_n 0.0154821f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_662_n N_A_656_74#_c_805_n 0.0119879f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_656_n N_A_1025_158#_c_848_n 0.0168557f $X=7.435 $Y=0.615 $X2=0
+ $Y2=0
cc_428 N_VGND_c_659_n N_A_1025_158#_c_848_n 0.00787994f $X=7.27 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_662_n N_A_1025_158#_c_848_n 0.00654995f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_M1001_d N_A_1025_158#_c_849_n 0.00180746f $X=7.295 $Y=0.37 $X2=0
+ $Y2=0
cc_431 N_VGND_c_656_n N_A_1025_158#_c_849_n 0.0163515f $X=7.435 $Y=0.615 $X2=0
+ $Y2=0
cc_432 N_VGND_c_656_n N_A_1025_158#_c_850_n 0.0168617f $X=7.435 $Y=0.615 $X2=0
+ $Y2=0
cc_433 N_VGND_c_657_n N_A_1025_158#_c_850_n 0.0171804f $X=8.315 $Y=0.615 $X2=0
+ $Y2=0
cc_434 N_VGND_c_660_n N_A_1025_158#_c_850_n 0.00838873f $X=8.13 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_662_n N_A_1025_158#_c_850_n 0.00694347f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_M1014_d N_A_1025_158#_c_851_n 0.00334827f $X=8.155 $Y=0.37 $X2=0
+ $Y2=0
cc_437 N_VGND_c_657_n N_A_1025_158#_c_851_n 0.0236105f $X=8.315 $Y=0.615 $X2=0
+ $Y2=0
cc_438 N_VGND_c_657_n N_A_1025_158#_c_852_n 0.0169405f $X=8.315 $Y=0.615 $X2=0
+ $Y2=0
cc_439 N_VGND_c_661_n N_A_1025_158#_c_852_n 0.0145639f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_662_n N_A_1025_158#_c_852_n 0.0119984f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_441 N_A_225_74#_c_748_n N_A_656_74#_M1003_s 0.00335829f $X=4.71 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_442 N_A_225_74#_c_748_n N_A_656_74#_M1019_s 0.00335829f $X=4.71 $Y=0.835
+ $X2=0 $Y2=0
cc_443 N_A_225_74#_M1009_d N_A_656_74#_c_802_n 0.00179007f $X=3.71 $Y=0.37 $X2=0
+ $Y2=0
cc_444 N_A_225_74#_M1021_d N_A_656_74#_c_802_n 0.002891f $X=4.57 $Y=0.37 $X2=0
+ $Y2=0
cc_445 N_A_225_74#_c_747_n N_A_656_74#_c_802_n 0.00550602f $X=2.905 $Y=0.34
+ $X2=0 $Y2=0
cc_446 N_A_225_74#_c_748_n N_A_656_74#_c_802_n 0.0858378f $X=4.71 $Y=0.835 $X2=0
+ $Y2=0
cc_447 N_A_225_74#_c_748_n N_A_1025_158#_c_853_n 0.0106593f $X=4.71 $Y=0.835
+ $X2=0 $Y2=0
cc_448 N_A_656_74#_c_802_n N_A_1025_158#_M1000_s 0.00298648f $X=5.535 $Y=0.455
+ $X2=-0.19 $Y2=-0.245
cc_449 N_A_656_74#_c_803_n N_A_1025_158#_M1008_s 0.00178994f $X=6.395 $Y=0.465
+ $X2=0 $Y2=0
cc_450 N_A_656_74#_M1000_d N_A_1025_158#_c_847_n 0.00209695f $X=5.56 $Y=0.37
+ $X2=0 $Y2=0
cc_451 N_A_656_74#_c_802_n N_A_1025_158#_c_847_n 0.00363923f $X=5.535 $Y=0.455
+ $X2=0 $Y2=0
cc_452 N_A_656_74#_c_803_n N_A_1025_158#_c_847_n 0.00479011f $X=6.395 $Y=0.465
+ $X2=0 $Y2=0
cc_453 N_A_656_74#_c_804_n N_A_1025_158#_c_847_n 0.010631f $X=5.795 $Y=0.465
+ $X2=0 $Y2=0
cc_454 N_A_656_74#_c_805_n N_A_1025_158#_c_848_n 0.0171277f $X=6.56 $Y=0.465
+ $X2=0 $Y2=0
cc_455 N_A_656_74#_c_802_n N_A_1025_158#_c_853_n 0.0189665f $X=5.535 $Y=0.455
+ $X2=0 $Y2=0
cc_456 N_A_656_74#_c_803_n N_A_1025_158#_c_854_n 0.0146773f $X=6.395 $Y=0.465
+ $X2=0 $Y2=0
cc_457 N_A_656_74#_M1013_d N_A_1025_158#_c_855_n 0.00192406f $X=6.42 $Y=0.37
+ $X2=0 $Y2=0
cc_458 N_A_656_74#_c_803_n N_A_1025_158#_c_855_n 0.00430203f $X=6.395 $Y=0.465
+ $X2=0 $Y2=0
cc_459 N_A_656_74#_c_805_n N_A_1025_158#_c_855_n 0.0168408f $X=6.56 $Y=0.465
+ $X2=0 $Y2=0

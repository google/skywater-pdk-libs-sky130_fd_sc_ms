* File: sky130_fd_sc_ms__and3_2.spice
* Created: Fri Aug 28 17:12:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and3_2.pex.spice"
.subckt sky130_fd_sc_ms__and3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_133_136# N_A_M1005_g N_A_41_384#_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=29.052 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1004 A_247_136# N_B_M1004_g A_133_136# VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1344 PD=0.88 PS=1.06 NRD=12.18 NRS=29.052 M=1 R=4.26667 SA=75000.8
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_C_M1003_g A_247_136# VNB NLOWVT L=0.15 W=0.64 AD=0.15789
+ AS=0.0768 PD=1.2429 PS=0.88 NRD=14.988 NRS=12.18 M=1 R=4.26667 SA=75001.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_X_M1000_d N_A_41_384#_M1000_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.18256 PD=1.06 PS=1.4371 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1000_d N_A_41_384#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.3552 PD=1.06 PS=2.44 NRD=6.48 NRS=27.564 M=1 R=4.93333
+ SA=75001.7 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_41_384#_M1006_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1638 AS=0.2352 PD=1.23 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1007 N_A_41_384#_M1007_d N_B_M1007_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1638 PD=1.11 PS=1.23 NRD=0 NRS=15.2281 M=1 R=4.66667 SA=90000.8
+ SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1008_d N_C_M1008_g N_A_41_384#_M1007_d VPB PSHORT L=0.18 W=0.84
+ AD=0.231257 AS=0.1134 PD=1.42286 PS=1.11 NRD=114.91 NRS=0 M=1 R=4.66667
+ SA=90001.2 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1001 N_X_M1001_d N_A_41_384#_M1001_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308343 PD=1.39 PS=1.89714 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.5 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1002 N_X_M1001_d N_A_41_384#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.392 PD=1.39 PS=2.94 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90002
+ SB=90000.3 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_56 VPB 0 1.15e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__and3_2.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dlrtp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dlrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.515000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.097600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.175000 1.800000 8.995000 1.970000 ;
        RECT 7.175000 1.970000 7.425000 2.980000 ;
        RECT 7.385000 0.365000 7.645000 0.880000 ;
        RECT 7.385000 0.880000 8.995000 1.130000 ;
        RECT 8.095000 1.970000 8.425000 2.980000 ;
        RECT 8.315000 0.365000 8.505000 0.880000 ;
        RECT 8.765000 1.130000 8.995000 1.800000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.494400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.120000 6.595000 1.450000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.262200 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.450000 1.290000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.120000 0.085000 ;
        RECT 0.680000  0.085000 1.010000 0.940000 ;
        RECT 2.335000  0.085000 2.665000 0.600000 ;
        RECT 4.190000  0.085000 4.440000 0.810000 ;
        RECT 5.965000  0.085000 6.295000 0.600000 ;
        RECT 6.955000  0.085000 7.215000 1.130000 ;
        RECT 7.815000  0.085000 8.145000 0.710000 ;
        RECT 8.675000  0.085000 9.005000 0.710000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.120000 3.415000 ;
        RECT 0.650000 2.710000 0.980000 3.245000 ;
        RECT 2.335000 2.710000 2.665000 3.245000 ;
        RECT 4.345000 2.650000 4.905000 3.245000 ;
        RECT 5.610000 1.960000 5.940000 3.245000 ;
        RECT 6.645000 1.960000 6.975000 3.245000 ;
        RECT 7.595000 2.140000 7.925000 3.245000 ;
        RECT 8.595000 2.140000 8.925000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.610000 0.445000 1.110000 ;
      RECT 0.115000 1.110000 0.855000 1.280000 ;
      RECT 0.115000 1.950000 0.855000 2.370000 ;
      RECT 0.115000 2.370000 2.665000 2.540000 ;
      RECT 0.115000 2.540000 0.445000 2.830000 ;
      RECT 0.685000 1.280000 0.855000 1.950000 ;
      RECT 1.185000 1.950000 1.630000 2.200000 ;
      RECT 1.240000 0.420000 1.630000 0.770000 ;
      RECT 1.240000 0.770000 3.005000 0.940000 ;
      RECT 1.240000 0.940000 1.630000 1.200000 ;
      RECT 1.460000 1.200000 1.630000 1.450000 ;
      RECT 1.460000 1.450000 1.900000 1.780000 ;
      RECT 1.460000 1.780000 1.630000 1.950000 ;
      RECT 1.800000 1.110000 3.340000 1.280000 ;
      RECT 1.800000 2.020000 2.240000 2.200000 ;
      RECT 2.070000 1.280000 2.240000 2.020000 ;
      RECT 2.495000 1.470000 2.785000 1.800000 ;
      RECT 2.495000 1.800000 2.665000 2.370000 ;
      RECT 2.835000 0.255000 4.020000 0.425000 ;
      RECT 2.835000 0.425000 3.005000 0.770000 ;
      RECT 2.845000 1.970000 3.125000 2.140000 ;
      RECT 2.845000 2.140000 3.015000 2.905000 ;
      RECT 2.845000 2.905000 3.985000 3.075000 ;
      RECT 2.955000 1.280000 3.340000 1.450000 ;
      RECT 2.955000 1.450000 3.125000 1.970000 ;
      RECT 3.175000 0.595000 3.680000 0.925000 ;
      RECT 3.185000 2.405000 3.465000 2.735000 ;
      RECT 3.295000 1.725000 5.020000 1.895000 ;
      RECT 3.295000 1.895000 3.465000 2.405000 ;
      RECT 3.510000 0.925000 3.680000 1.725000 ;
      RECT 3.655000 2.065000 3.985000 2.905000 ;
      RECT 3.850000 0.425000 4.020000 1.225000 ;
      RECT 3.850000 1.225000 4.150000 1.555000 ;
      RECT 4.195000 2.065000 5.440000 2.480000 ;
      RECT 4.670000 0.280000 5.785000 0.450000 ;
      RECT 4.670000 0.450000 5.000000 1.030000 ;
      RECT 4.720000 1.350000 5.020000 1.725000 ;
      RECT 5.110000 2.480000 5.440000 2.700000 ;
      RECT 5.180000 0.620000 5.360000 0.950000 ;
      RECT 5.190000 0.950000 5.360000 1.620000 ;
      RECT 5.190000 1.620000 8.595000 1.630000 ;
      RECT 5.190000 1.630000 6.935000 1.790000 ;
      RECT 5.190000 1.790000 5.440000 2.065000 ;
      RECT 5.535000 0.450000 5.785000 0.770000 ;
      RECT 5.535000 0.770000 6.725000 0.950000 ;
      RECT 6.110000 1.790000 6.440000 2.700000 ;
      RECT 6.465000 0.345000 6.725000 0.770000 ;
      RECT 6.765000 1.300000 8.595000 1.620000 ;
  END
END sky130_fd_sc_ms__dlrtp_4

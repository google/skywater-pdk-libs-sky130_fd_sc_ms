* File: sky130_fd_sc_ms__mux2i_1.pxi.spice
* Created: Wed Sep  2 12:11:59 2020
* 
x_PM_SKY130_FD_SC_MS__MUX2I_1%S N_S_M1009_g N_S_M1007_g N_S_c_70_n N_S_M1002_g
+ N_S_c_72_n N_S_M1008_g N_S_c_73_n N_S_c_79_n N_S_c_74_n S S N_S_c_76_n
+ PM_SKY130_FD_SC_MS__MUX2I_1%S
x_PM_SKY130_FD_SC_MS__MUX2I_1%A_114_74# N_A_114_74#_M1007_d N_A_114_74#_M1009_d
+ N_A_114_74#_M1003_g N_A_114_74#_M1001_g N_A_114_74#_c_130_n
+ N_A_114_74#_c_131_n N_A_114_74#_c_132_n N_A_114_74#_c_138_n
+ N_A_114_74#_c_133_n N_A_114_74#_c_134_n N_A_114_74#_c_135_n
+ N_A_114_74#_c_136_n PM_SKY130_FD_SC_MS__MUX2I_1%A_114_74#
x_PM_SKY130_FD_SC_MS__MUX2I_1%A0 N_A0_M1000_g N_A0_c_203_n N_A0_M1005_g A0
+ N_A0_c_201_n N_A0_c_202_n PM_SKY130_FD_SC_MS__MUX2I_1%A0
x_PM_SKY130_FD_SC_MS__MUX2I_1%A1 N_A1_c_235_n N_A1_M1004_g N_A1_M1006_g A1
+ N_A1_c_238_n PM_SKY130_FD_SC_MS__MUX2I_1%A1
x_PM_SKY130_FD_SC_MS__MUX2I_1%VPWR N_VPWR_M1009_s N_VPWR_M1002_d N_VPWR_c_258_n
+ N_VPWR_c_259_n N_VPWR_c_260_n VPWR N_VPWR_c_261_n N_VPWR_c_262_n
+ N_VPWR_c_257_n N_VPWR_c_264_n PM_SKY130_FD_SC_MS__MUX2I_1%VPWR
x_PM_SKY130_FD_SC_MS__MUX2I_1%A_223_368# N_A_223_368#_M1002_s
+ N_A_223_368#_M1005_s N_A_223_368#_c_293_n N_A_223_368#_c_294_n
+ N_A_223_368#_c_295_n N_A_223_368#_c_296_n
+ PM_SKY130_FD_SC_MS__MUX2I_1%A_223_368#
x_PM_SKY130_FD_SC_MS__MUX2I_1%A_402_368# N_A_402_368#_M1003_d
+ N_A_402_368#_M1006_d N_A_402_368#_c_323_n N_A_402_368#_c_324_n
+ N_A_402_368#_c_325_n N_A_402_368#_c_326_n
+ PM_SKY130_FD_SC_MS__MUX2I_1%A_402_368#
x_PM_SKY130_FD_SC_MS__MUX2I_1%Y N_Y_M1000_d N_Y_M1005_d N_Y_c_366_p N_Y_c_348_n
+ N_Y_c_350_n Y PM_SKY130_FD_SC_MS__MUX2I_1%Y
x_PM_SKY130_FD_SC_MS__MUX2I_1%VGND N_VGND_M1007_s N_VGND_M1008_d N_VGND_c_368_n
+ N_VGND_c_369_n N_VGND_c_370_n VGND N_VGND_c_371_n N_VGND_c_372_n
+ N_VGND_c_373_n N_VGND_c_374_n PM_SKY130_FD_SC_MS__MUX2I_1%VGND
x_PM_SKY130_FD_SC_MS__MUX2I_1%A_225_74# N_A_225_74#_M1008_s N_A_225_74#_M1004_d
+ N_A_225_74#_c_404_n N_A_225_74#_c_405_n N_A_225_74#_c_406_n
+ N_A_225_74#_c_415_n N_A_225_74#_c_407_n N_A_225_74#_c_408_n
+ N_A_225_74#_c_409_n PM_SKY130_FD_SC_MS__MUX2I_1%A_225_74#
cc_1 VNB N_S_M1007_g 0.0378713f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_S_c_70_n 0.0500851f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.26
cc_3 VNB N_S_M1002_g 0.020162f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_4 VNB N_S_c_72_n 0.0203248f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.185
cc_5 VNB N_S_c_73_n 0.0155613f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.26
cc_6 VNB N_S_c_74_n 0.00664804f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.26
cc_7 VNB S 0.0234095f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_S_c_76_n 0.0290861f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_9 VNB N_A_114_74#_M1001_g 0.0251947f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_10 VNB N_A_114_74#_c_130_n 0.00541105f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.335
cc_11 VNB N_A_114_74#_c_131_n 0.0201137f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.26
cc_12 VNB N_A_114_74#_c_132_n 0.00490111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_114_74#_c_133_n 0.00341769f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_14 VNB N_A_114_74#_c_134_n 0.00106462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_114_74#_c_135_n 0.00166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_114_74#_c_136_n 0.0269708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A0_M1000_g 0.0286315f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_18 VNB N_A0_c_201_n 0.04568f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_19 VNB N_A0_c_202_n 0.00549587f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_20 VNB N_A1_c_235_n 0.0257716f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.945
cc_21 VNB N_A1_M1006_g 0.00944997f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_22 VNB A1 0.00924341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_238_n 0.0633283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_257_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_25 VNB N_Y_c_348_n 0.0122596f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.26
cc_26 VNB N_VGND_c_368_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_27 VNB N_VGND_c_369_n 0.0325289f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.26
cc_28 VNB N_VGND_c_370_n 0.00969314f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_29 VNB N_VGND_c_371_n 0.034428f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_30 VNB N_VGND_c_372_n 0.0504776f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_31 VNB N_VGND_c_373_n 0.240757f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.35
cc_32 VNB N_VGND_c_374_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_225_74#_c_404_n 0.00874347f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.26
cc_34 VNB N_A_225_74#_c_405_n 0.0100806f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=1.335
cc_35 VNB N_A_225_74#_c_406_n 0.00386611f $X=-0.19 $Y=-0.245 $X2=1.47 $Y2=2.4
cc_36 VNB N_A_225_74#_c_407_n 0.0070932f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.185
cc_37 VNB N_A_225_74#_c_408_n 0.00124385f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_38 VNB N_A_225_74#_c_409_n 0.0279156f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.68
cc_39 VPB N_S_M1009_g 0.0323486f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_40 VPB N_S_M1002_g 0.0275322f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_41 VPB N_S_c_79_n 0.0298646f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.68
cc_42 VPB S 0.0120179f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB N_S_c_76_n 0.00170579f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_44 VPB N_A_114_74#_M1003_g 0.0250126f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.26
cc_45 VPB N_A_114_74#_c_138_n 0.0162142f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_46 VPB N_A_114_74#_c_133_n 0.00990288f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.295
cc_47 VPB N_A_114_74#_c_135_n 0.00163415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_114_74#_c_136_n 0.00576402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A0_c_203_n 0.0199904f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_50 VPB N_A0_c_201_n 0.0164255f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_51 VPB N_A0_c_202_n 0.0041961f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_52 VPB N_A1_M1006_g 0.0292517f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_53 VPB N_VPWR_c_258_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_54 VPB N_VPWR_c_259_n 0.0472706f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.26
cc_55 VPB N_VPWR_c_260_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_56 VPB N_VPWR_c_261_n 0.0326305f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.74
cc_57 VPB N_VPWR_c_262_n 0.0489477f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_58 VPB N_VPWR_c_257_n 0.073045f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.35
cc_59 VPB N_VPWR_c_264_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_223_368#_c_293_n 0.00521825f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_61 VPB N_A_223_368#_c_294_n 0.0098828f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.26
cc_62 VPB N_A_223_368#_c_295_n 0.0135882f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.335
cc_63 VPB N_A_223_368#_c_296_n 0.00737697f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.335
cc_64 VPB N_A_402_368#_c_323_n 0.00685898f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.26
cc_65 VPB N_A_402_368#_c_324_n 0.0239108f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=1.335
cc_66 VPB N_A_402_368#_c_325_n 0.0036732f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.4
cc_67 VPB N_A_402_368#_c_326_n 0.0442133f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=1.185
cc_68 VPB N_Y_c_348_n 0.00399281f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.26
cc_69 N_S_M1002_g N_A_114_74#_M1003_g 0.0351196f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_70 N_S_c_72_n N_A_114_74#_M1001_g 0.026721f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_71 N_S_M1007_g N_A_114_74#_c_130_n 0.00968387f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_72 N_S_c_70_n N_A_114_74#_c_130_n 0.0189538f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_73 N_S_M1002_g N_A_114_74#_c_130_n 3.49755e-19 $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_74 S N_A_114_74#_c_130_n 0.0123511f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_S_c_76_n N_A_114_74#_c_130_n 3.2525e-19 $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_76 N_S_c_70_n N_A_114_74#_c_131_n 0.0129614f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_77 N_S_M1002_g N_A_114_74#_c_131_n 0.0150924f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_78 N_S_M1007_g N_A_114_74#_c_132_n 0.009213f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_79 N_S_c_70_n N_A_114_74#_c_132_n 0.0020895f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_80 N_S_c_72_n N_A_114_74#_c_132_n 0.0015289f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_81 N_S_M1009_g N_A_114_74#_c_138_n 0.0167311f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_82 N_S_M1002_g N_A_114_74#_c_133_n 0.0076579f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_83 N_S_c_79_n N_A_114_74#_c_133_n 0.00885853f $X=0.395 $Y=1.68 $X2=0 $Y2=0
cc_84 S N_A_114_74#_c_133_n 0.0255963f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_S_c_76_n N_A_114_74#_c_133_n 0.00775954f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_86 S N_A_114_74#_c_134_n 0.0145892f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_S_c_76_n N_A_114_74#_c_134_n 0.00410432f $X=0.385 $Y=1.35 $X2=0 $Y2=0
cc_88 N_S_M1002_g N_A_114_74#_c_135_n 0.00116992f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_89 N_S_M1002_g N_A_114_74#_c_136_n 0.0183745f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_90 N_S_M1009_g N_VPWR_c_259_n 0.00870081f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_91 N_S_c_79_n N_VPWR_c_259_n 0.00100521f $X=0.395 $Y=1.68 $X2=0 $Y2=0
cc_92 S N_VPWR_c_259_n 0.0158723f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_S_M1002_g N_VPWR_c_260_n 0.0158618f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_94 N_S_M1009_g N_VPWR_c_261_n 0.005209f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_95 N_S_M1002_g N_VPWR_c_261_n 0.00460063f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_96 N_S_M1009_g N_VPWR_c_257_n 0.00991105f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_97 N_S_M1002_g N_VPWR_c_257_n 0.00913687f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_98 N_S_M1002_g N_A_223_368#_c_293_n 8.13654e-19 $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_99 N_S_M1009_g N_A_223_368#_c_294_n 0.00167358f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_100 N_S_M1002_g N_A_223_368#_c_294_n 0.00147311f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_101 N_S_M1002_g N_A_223_368#_c_295_n 0.0158466f $X=1.47 $Y=2.4 $X2=0 $Y2=0
cc_102 N_S_M1007_g N_VGND_c_369_n 0.00800579f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_103 N_S_c_73_n N_VGND_c_369_n 0.0010506f $X=0.395 $Y=1.26 $X2=0 $Y2=0
cc_104 S N_VGND_c_369_n 0.015437f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_105 N_S_c_72_n N_VGND_c_370_n 0.00622602f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_106 N_S_M1007_g N_VGND_c_371_n 0.0043544f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_107 N_S_c_72_n N_VGND_c_371_n 0.00434272f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_108 N_S_M1007_g N_VGND_c_373_n 0.00830065f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_109 N_S_c_72_n N_VGND_c_373_n 0.00826311f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_110 N_S_M1007_g N_A_225_74#_c_404_n 0.0024493f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_111 N_S_c_72_n N_A_225_74#_c_404_n 0.0103339f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_112 N_S_c_72_n N_A_225_74#_c_405_n 0.0117984f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_113 N_S_c_70_n N_A_225_74#_c_406_n 0.00554277f $X=1.38 $Y=1.26 $X2=0 $Y2=0
cc_114 N_S_c_72_n N_A_225_74#_c_406_n 0.00214722f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_115 N_S_c_72_n N_A_225_74#_c_415_n 5.97863e-19 $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_116 N_A_114_74#_M1001_g N_A0_M1000_g 0.0329672f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_114_74#_c_135_n N_A0_c_201_n 8.89634e-19 $X=1.965 $Y=1.435 $X2=0
+ $Y2=0
cc_118 N_A_114_74#_c_136_n N_A0_c_201_n 0.0378784f $X=1.965 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A_114_74#_M1003_g N_A0_c_202_n 0.00263235f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_114_74#_c_135_n N_A0_c_202_n 0.013347f $X=1.965 $Y=1.435 $X2=0 $Y2=0
cc_121 N_A_114_74#_c_136_n N_A0_c_202_n 0.00174711f $X=1.965 $Y=1.515 $X2=0
+ $Y2=0
cc_122 N_A_114_74#_c_138_n N_VPWR_c_259_n 0.0303778f $X=0.72 $Y=2.265 $X2=0
+ $Y2=0
cc_123 N_A_114_74#_M1003_g N_VPWR_c_260_n 0.0128546f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_114_74#_c_138_n N_VPWR_c_261_n 0.0147721f $X=0.72 $Y=2.265 $X2=0
+ $Y2=0
cc_125 N_A_114_74#_M1003_g N_VPWR_c_262_n 0.00460063f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_114_74#_M1003_g N_VPWR_c_257_n 0.00913687f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_114_74#_c_138_n N_VPWR_c_257_n 0.0121589f $X=0.72 $Y=2.265 $X2=0
+ $Y2=0
cc_128 N_A_114_74#_c_131_n N_A_223_368#_c_293_n 0.0142143f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_129 N_A_114_74#_c_133_n N_A_223_368#_c_293_n 0.0226777f $X=0.722 $Y=2.1 $X2=0
+ $Y2=0
cc_130 N_A_114_74#_c_138_n N_A_223_368#_c_294_n 0.0648589f $X=0.72 $Y=2.265
+ $X2=0 $Y2=0
cc_131 N_A_114_74#_M1003_g N_A_223_368#_c_295_n 0.0190473f $X=1.92 $Y=2.4 $X2=0
+ $Y2=0
cc_132 N_A_114_74#_c_131_n N_A_223_368#_c_295_n 0.0143565f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_133 N_A_114_74#_c_135_n N_A_223_368#_c_295_n 0.0143711f $X=1.965 $Y=1.435
+ $X2=0 $Y2=0
cc_134 N_A_114_74#_c_136_n N_A_223_368#_c_295_n 5.96025e-19 $X=1.965 $Y=1.515
+ $X2=0 $Y2=0
cc_135 N_A_114_74#_M1003_g N_A_223_368#_c_296_n 0.00489007f $X=1.92 $Y=2.4 $X2=0
+ $Y2=0
cc_136 N_A_114_74#_M1003_g N_A_402_368#_c_325_n 0.0028276f $X=1.92 $Y=2.4 $X2=0
+ $Y2=0
cc_137 N_A_114_74#_M1001_g N_Y_c_350_n 2.75206e-19 $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_114_74#_M1001_g N_VGND_c_370_n 0.00622568f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_114_74#_c_132_n N_VGND_c_371_n 0.0111177f $X=0.71 $Y=0.645 $X2=0
+ $Y2=0
cc_140 N_A_114_74#_M1001_g N_VGND_c_372_n 0.00433139f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_114_74#_M1001_g N_VGND_c_373_n 0.00817354f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_114_74#_c_132_n N_VGND_c_373_n 0.0120515f $X=0.71 $Y=0.645 $X2=0
+ $Y2=0
cc_143 N_A_114_74#_M1001_g N_A_225_74#_c_404_n 6.28869e-19 $X=2.055 $Y=0.74
+ $X2=0 $Y2=0
cc_144 N_A_114_74#_c_132_n N_A_225_74#_c_404_n 0.0424364f $X=0.71 $Y=0.645 $X2=0
+ $Y2=0
cc_145 N_A_114_74#_M1001_g N_A_225_74#_c_405_n 0.0136151f $X=2.055 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_114_74#_c_131_n N_A_225_74#_c_405_n 0.0265109f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_147 N_A_114_74#_c_135_n N_A_225_74#_c_405_n 0.0243844f $X=1.965 $Y=1.435
+ $X2=0 $Y2=0
cc_148 N_A_114_74#_c_136_n N_A_225_74#_c_405_n 0.00124773f $X=1.965 $Y=1.515
+ $X2=0 $Y2=0
cc_149 N_A_114_74#_c_130_n N_A_225_74#_c_406_n 0.0121698f $X=0.805 $Y=1.35 $X2=0
+ $Y2=0
cc_150 N_A_114_74#_c_131_n N_A_225_74#_c_406_n 0.0275396f $X=1.8 $Y=1.435 $X2=0
+ $Y2=0
cc_151 N_A_114_74#_M1001_g N_A_225_74#_c_415_n 0.00985062f $X=2.055 $Y=0.74
+ $X2=0 $Y2=0
cc_152 N_A_114_74#_M1001_g N_A_225_74#_c_408_n 0.00375375f $X=2.055 $Y=0.74
+ $X2=0 $Y2=0
cc_153 N_A0_M1000_g N_A1_c_235_n 0.0101019f $X=2.445 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A0_c_201_n N_A1_M1006_g 0.0335879f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A0_c_201_n N_A1_c_238_n 0.00888505f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A0_c_203_n N_VPWR_c_262_n 0.00333926f $X=2.895 $Y=1.77 $X2=0 $Y2=0
cc_157 N_A0_c_203_n N_VPWR_c_257_n 0.00427931f $X=2.895 $Y=1.77 $X2=0 $Y2=0
cc_158 N_A0_c_201_n N_A_223_368#_c_295_n 0.00415885f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A0_c_203_n N_A_223_368#_c_296_n 0.0114497f $X=2.895 $Y=1.77 $X2=0 $Y2=0
cc_160 N_A0_c_201_n N_A_223_368#_c_296_n 0.00228146f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A0_c_202_n N_A_223_368#_c_296_n 0.0246446f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A0_c_203_n N_A_402_368#_c_323_n 0.004848f $X=2.895 $Y=1.77 $X2=0 $Y2=0
cc_163 N_A0_c_203_n N_A_402_368#_c_324_n 0.0167923f $X=2.895 $Y=1.77 $X2=0 $Y2=0
cc_164 N_A0_c_203_n N_A_402_368#_c_326_n 0.0010052f $X=2.895 $Y=1.77 $X2=0 $Y2=0
cc_165 N_A0_M1000_g N_Y_c_348_n 0.00502765f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A0_c_201_n N_Y_c_348_n 0.00563212f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A0_c_202_n N_Y_c_348_n 0.0326257f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A0_M1000_g N_Y_c_350_n 0.00510039f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A0_c_201_n N_Y_c_350_n 0.00634965f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A0_c_202_n N_Y_c_350_n 0.015419f $X=2.7 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A0_M1000_g N_VGND_c_372_n 0.00291649f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A0_M1000_g N_VGND_c_373_n 0.00361693f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A0_M1000_g N_A_225_74#_c_405_n 0.00451515f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A0_M1000_g N_A_225_74#_c_415_n 0.00611057f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A0_M1000_g N_A_225_74#_c_407_n 0.0149352f $X=2.445 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_M1006_g N_VPWR_c_262_n 0.00333896f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A1_M1006_g N_VPWR_c_257_n 0.00426502f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A1_M1006_g N_A_402_368#_c_324_n 0.0145133f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A1_M1006_g N_A_402_368#_c_326_n 0.0156015f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_180 A1 N_A_402_368#_c_326_n 0.0190699f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A1_c_238_n N_A_402_368#_c_326_n 0.00216224f $X=3.56 $Y=1.385 $X2=0
+ $Y2=0
cc_182 N_A1_c_235_n N_Y_c_348_n 0.00708472f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_183 N_A1_M1006_g N_Y_c_348_n 0.00788008f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_184 A1 N_Y_c_348_n 0.0282043f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A1_c_235_n N_VGND_c_372_n 0.00291649f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_186 N_A1_c_235_n N_VGND_c_373_n 0.00365785f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_187 N_A1_c_235_n N_A_225_74#_c_407_n 0.0142787f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_188 A1 N_A_225_74#_c_409_n 0.0232175f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A1_c_238_n N_A_225_74#_c_409_n 0.00189183f $X=3.56 $Y=1.385 $X2=0 $Y2=0
cc_190 N_VPWR_c_260_n N_A_223_368#_c_294_n 0.0234083f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_261_n N_A_223_368#_c_294_n 0.011066f $X=1.53 $Y=3.33 $X2=0 $Y2=0
cc_192 N_VPWR_c_257_n N_A_223_368#_c_294_n 0.00915947f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_193 N_VPWR_M1002_d N_A_223_368#_c_295_n 0.00425857f $X=1.56 $Y=1.84 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_260_n N_A_223_368#_c_295_n 0.0170259f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_262_n N_A_402_368#_c_324_n 0.0930732f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_257_n N_A_402_368#_c_324_n 0.0523528f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_260_n N_A_402_368#_c_325_n 0.0103602f $X=1.695 $Y=2.455 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_262_n N_A_402_368#_c_325_n 0.0179217f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_257_n N_A_402_368#_c_325_n 0.00971942f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_200 N_A_223_368#_c_295_n N_A_402_368#_M1003_d 0.00893085f $X=2.505 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_201 N_A_223_368#_c_295_n N_A_402_368#_c_323_n 0.0198097f $X=2.505 $Y=2.035
+ $X2=0 $Y2=0
cc_202 N_A_223_368#_c_296_n N_A_402_368#_c_323_n 0.0329563f $X=2.67 $Y=2.115
+ $X2=0 $Y2=0
cc_203 N_A_223_368#_M1005_s N_A_402_368#_c_324_n 0.00246514f $X=2.54 $Y=1.84
+ $X2=0 $Y2=0
cc_204 N_A_223_368#_c_296_n N_A_402_368#_c_324_n 0.0205469f $X=2.67 $Y=2.115
+ $X2=0 $Y2=0
cc_205 N_A_402_368#_c_324_n N_Y_M1005_d 0.00165831f $X=3.405 $Y=2.99 $X2=0 $Y2=0
cc_206 N_A_402_368#_c_324_n N_Y_c_348_n 0.0118736f $X=3.405 $Y=2.99 $X2=0 $Y2=0
cc_207 N_A_402_368#_c_326_n N_Y_c_348_n 0.0334931f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_208 N_Y_c_350_n N_A_225_74#_c_405_n 0.00171692f $X=3.035 $Y=0.87 $X2=0 $Y2=0
cc_209 N_Y_c_350_n N_A_225_74#_c_415_n 0.0195323f $X=3.035 $Y=0.87 $X2=0 $Y2=0
cc_210 N_Y_M1000_d N_A_225_74#_c_407_n 0.00935673f $X=2.52 $Y=0.37 $X2=0 $Y2=0
cc_211 N_Y_c_366_p N_A_225_74#_c_407_n 0.00960383f $X=3.13 $Y=1.035 $X2=0 $Y2=0
cc_212 N_Y_c_350_n N_A_225_74#_c_407_n 0.032664f $X=3.035 $Y=0.87 $X2=0 $Y2=0
cc_213 N_VGND_c_370_n N_A_225_74#_c_404_n 0.0191765f $X=1.77 $Y=0.675 $X2=0
+ $Y2=0
cc_214 N_VGND_c_371_n N_A_225_74#_c_404_n 0.0145639f $X=1.605 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_373_n N_A_225_74#_c_404_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_M1008_d N_A_225_74#_c_405_n 0.00358162f $X=1.56 $Y=0.37 $X2=0
+ $Y2=0
cc_217 N_VGND_c_370_n N_A_225_74#_c_405_n 0.0248957f $X=1.77 $Y=0.675 $X2=0
+ $Y2=0
cc_218 N_VGND_c_372_n N_A_225_74#_c_407_n 0.044415f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_373_n N_A_225_74#_c_407_n 0.0381644f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_370_n N_A_225_74#_c_408_n 0.00795492f $X=1.77 $Y=0.675 $X2=0
+ $Y2=0
cc_221 N_VGND_c_372_n N_A_225_74#_c_408_n 0.00751083f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_373_n N_A_225_74#_c_408_n 0.00615808f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_372_n N_A_225_74#_c_409_n 0.0126895f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_373_n N_A_225_74#_c_409_n 0.0105154f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_A_225_74#_c_405_n A_426_74# 0.00122604f $X=2.105 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_225_74#_c_415_n A_426_74# 0.00479875f $X=2.19 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_225_74#_c_407_n A_426_74# 0.00141176f $X=3.395 $Y=0.435 $X2=-0.19
+ $Y2=-0.245

* File: sky130_fd_sc_ms__edfxbp_1.spice
* Created: Fri Aug 28 17:32:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__edfxbp_1.pex.spice"
.subckt sky130_fd_sc_ms__edfxbp_1  VNB VPB D DE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1032 A_145_74# N_D_M1032_g N_A_27_74#_M1032_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1848 PD=0.66 PS=1.72 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_DE_M1018_g A_145_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_DE_M1024_g N_A_161_446#_M1024_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.1281 PD=0.78 PS=1.45 NRD=19.992 NRS=2.856 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_527_74# N_A_161_446#_M1001_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=2.856 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_27_74#_M1002_d N_A_575_48#_M1002_g A_527_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_818_74#_M1025_d N_CLK_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.2109 PD=2.01 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1029 N_A_1008_74#_M1029_d N_A_818_74#_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1034 N_A_1198_97#_M1034_d N_A_818_74#_M1034_g N_A_27_74#_M1034_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1014 A_1334_97# N_A_1008_74#_M1014_g N_A_1198_97#_M1034_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08925 AS=0.1113 PD=0.845 PS=0.95 NRD=45 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_1419_71#_M1019_g A_1334_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109992 AS=0.08925 PD=0.92717 PS=0.845 NRD=0 NRS=45 M=1 R=2.8 SA=75001.4
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1015 N_A_1419_71#_M1015_d N_A_1198_97#_M1015_g N_VGND_M1019_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.167608 PD=1.85 PS=1.41283 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 A_1807_74# N_A_1419_71#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.2109 PD=0.95 PS=2.05 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1006 N_A_1879_74#_M1006_d N_A_1008_74#_M1006_g A_1807_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.477045 AS=0.0777 PD=2.97276 PS=0.95 NRD=14.592 NRS=8.1 M=1
+ R=4.93333 SA=75000.6 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1021 A_2227_118# N_A_818_74#_M1021_g N_A_1879_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.270755 PD=0.66 PS=1.68724 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_575_48#_M1010_g A_2227_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.114985 AS=0.0504 PD=0.907358 PS=0.66 NRD=45 NRS=18.564 M=1 R=2.8
+ SA=75002.7 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_575_48#_M1016_d N_A_1879_74#_M1016_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.175215 PD=1.85 PS=1.38264 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A_1879_74#_M1017_g N_Q_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2257 AS=0.2109 PD=1.35 PS=2.05 NRD=53.508 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1020 N_Q_N_M1020_d N_A_575_48#_M1020_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2257 PD=2.05 PS=1.35 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 A_119_508# N_D_M1027_g N_A_27_74#_M1027_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=23.443 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_161_446#_M1011_g A_119_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333 SA=90000.6
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_DE_M1008_g N_A_161_446#_M1008_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.3766 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1009 A_559_504# N_DE_M1009_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=0.42 AD=0.0441
+ AS=0.105 PD=0.63 PS=0.903396 NRD=23.443 NRS=0 M=1 R=2.33333 SA=90000.9
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1033 N_A_27_74#_M1033_d N_A_575_48#_M1033_g A_559_504# VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333
+ SA=90001.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1031 N_A_818_74#_M1031_d N_CLK_M1031_g N_VPWR_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1028 N_A_1008_74#_M1028_d N_A_818_74#_M1028_g N_VPWR_M1028_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_1198_97#_M1000_d N_A_1008_74#_M1000_g N_A_27_74#_M1000_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1997 PD=0.69 PS=1.89 NRD=0 NRS=39.8531 M=1
+ R=2.33333 SA=90000.3 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1007 A_1426_508# N_A_818_74#_M1007_g N_A_1198_97#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0693 AS=0.0567 PD=0.75 PS=0.69 NRD=51.5943 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1023 N_VPWR_M1023_d N_A_1419_71#_M1023_g A_1426_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.119317 AS=0.0693 PD=1.01 PS=0.75 NRD=107.444 NRS=51.5943 M=1 R=2.33333
+ SA=90001.2 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1005 N_A_1419_71#_M1005_d N_A_1198_97#_M1005_g N_VPWR_M1023_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.238633 PD=2.24 PS=2.02 NRD=0 NRS=53.7219 M=1
+ R=4.66667 SA=90001 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1012 A_2011_392# N_A_1419_71#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1035 N_A_1879_74#_M1035_d N_A_818_74#_M1035_g A_2011_392# VPB PSHORT L=0.18
+ W=1 AD=0.229718 AS=0.12 PD=1.95775 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1003 A_2209_443# N_A_1008_74#_M1003_g N_A_1879_74#_M1035_d VPB PSHORT L=0.18
+ W=0.42 AD=0.063 AS=0.0964817 PD=0.72 PS=0.822254 NRD=44.5417 NRS=53.9386 M=1
+ R=2.33333 SA=90001.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1022 N_VPWR_M1022_d N_A_575_48#_M1022_g A_2209_443# VPB PSHORT L=0.18 W=0.42
+ AD=0.139162 AS=0.063 PD=1.05 PS=0.72 NRD=0 NRS=44.5417 M=1 R=2.33333
+ SA=90001.7 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1013 N_A_575_48#_M1013_d N_A_1879_74#_M1013_g N_VPWR_M1022_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.331338 PD=2.56 PS=2.5 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_A_1879_74#_M1026_g N_Q_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1030 N_Q_N_M1030_d N_A_575_48#_M1030_g N_VPWR_M1026_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX36_noxref VNB VPB NWDIODE A=27.5178 P=33.33
*
.include "sky130_fd_sc_ms__edfxbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sdfbbn_2.pex.spice
* Created: Wed Sep  2 12:29:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%SCD 2 5 9 10 11 15 16 17 19
r31 19 21 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.97
+ $X2=0.407 $Y2=2.135
r32 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.97 $X2=0.385 $Y2=1.97
r33 15 17 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.29
+ $X2=0.407 $Y2=1.125
r34 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.29 $X2=0.385 $Y2=1.29
r35 11 20 8.27047 $w=4.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.97
r36 10 11 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r37 10 16 0.135582 $w=4.23e-07 $l=5e-09 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.29
r38 9 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.805
+ $X2=0.52 $Y2=1.125
r39 5 21 196.298 $w=1.8e-07 $l=5.05e-07 $layer=POLY_cond $X=0.505 $Y=2.64
+ $X2=0.505 $Y2=2.135
r40 2 19 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.948
+ $X2=0.407 $Y2=1.97
r41 1 15 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.312
+ $X2=0.407 $Y2=1.29
r42 1 2 94.3237 $w=3.75e-07 $l=6.36e-07 $layer=POLY_cond $X=0.407 $Y=1.312
+ $X2=0.407 $Y2=1.948
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%D 3 9 11 12 13 20
c58 13 0 1.16291e-19 $X=1.68 $Y=1.665
r59 18 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.65 $Y=1.625 $X2=1.74
+ $Y2=1.625
r60 15 18 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.42 $Y=1.625
+ $X2=1.65 $Y2=1.625
r61 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.625 $X2=1.65 $Y2=1.625
r62 11 12 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.375 $Y=2.035
+ $X2=1.375 $Y2=2.185
r63 7 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.46
+ $X2=1.74 $Y2=1.625
r64 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=1.74 $Y=1.46 $X2=1.74
+ $Y2=0.805
r65 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.79
+ $X2=1.42 $Y2=1.625
r66 5 11 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.42 $Y=1.79
+ $X2=1.42 $Y2=2.035
r67 3 12 176.863 $w=1.8e-07 $l=4.55e-07 $layer=POLY_cond $X=1.345 $Y=2.64
+ $X2=1.345 $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_341_410# 1 2 7 9 10 11 14 17 18 20 21 24
+ 28 32 34
c80 34 0 4.36151e-19 $X=3.067 $Y=1.645
c81 28 0 1.21362e-19 $X=3.025 $Y=0.815
c82 24 0 7.30946e-20 $X=2.77 $Y=1.645
c83 21 0 3.06618e-19 $X=2.94 $Y=1.645
c84 11 0 1.16291e-19 $X=1.885 $Y=2.125
r85 30 34 6.41553 $w=2.52e-07 $l=1.66493e-07 $layer=LI1_cond $X=3.07 $Y=1.81
+ $X2=3.067 $Y2=1.645
r86 30 32 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=3.07 $Y=1.81
+ $X2=3.07 $Y2=2.465
r87 26 34 6.41553 $w=2.52e-07 $l=1.65e-07 $layer=LI1_cond $X=3.067 $Y=1.48
+ $X2=3.067 $Y2=1.645
r88 26 28 30.0539 $w=2.53e-07 $l=6.65e-07 $layer=LI1_cond $X=3.067 $Y=1.48
+ $X2=3.067 $Y2=0.815
r89 24 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.77 $Y=1.645 $X2=2.77
+ $Y2=1.735
r90 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.645 $X2=2.77 $Y2=1.645
r91 21 34 0.398883 $w=3.3e-07 $l=1.27e-07 $layer=LI1_cond $X=2.94 $Y=1.645
+ $X2=3.067 $Y2=1.645
r92 21 23 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.94 $Y=1.645
+ $X2=2.77 $Y2=1.645
r93 19 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=1.735
+ $X2=2.13 $Y2=1.735
r94 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.605 $Y=1.735
+ $X2=2.77 $Y2=1.735
r95 18 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.605 $Y=1.735
+ $X2=2.205 $Y2=1.735
r96 16 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=1.735
r97 16 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=2.05
r98 12 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.66
+ $X2=2.13 $Y2=1.735
r99 12 14 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.13 $Y=1.66
+ $X2=2.13 $Y2=0.805
r100 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.055 $Y=2.125
+ $X2=2.13 $Y2=2.05
r101 10 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.055 $Y=2.125
+ $X2=1.885 $Y2=2.125
r102 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.795 $Y=2.2
+ $X2=1.885 $Y2=2.125
r103 7 9 117.822 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=1.795 $Y=2.2
+ $X2=1.795 $Y2=2.64
r104 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.32 $X2=3.03 $Y2=2.465
r105 1 28 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.595 $X2=3.025 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%SCE 4 7 9 10 11 13 17 18 19 20 21 23 26 27
+ 28 29 33 34
c100 20 0 3.4396e-19 $X=3.175 $Y=2.125
c101 18 0 1.53309e-19 $X=3.175 $Y=1.165
c102 7 0 2.32243e-19 $X=0.955 $Y=2.64
c103 4 0 1.01507e-19 $X=0.91 $Y=0.805
r104 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.97
+ $Y=1.29 $X2=0.97 $Y2=1.29
r105 28 29 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=1.295
+ $X2=1.06 $Y2=1.665
r106 28 34 0.117263 $w=5.08e-07 $l=5e-09 $layer=LI1_cond $X=1.06 $Y=1.295
+ $X2=1.06 $Y2=1.29
r107 26 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.97 $Y=1.63
+ $X2=0.97 $Y2=1.29
r108 26 27 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.63
+ $X2=0.97 $Y2=1.795
r109 25 33 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.125
+ $X2=0.97 $Y2=1.29
r110 22 23 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.25 $Y=1.24
+ $X2=3.25 $Y2=2.05
r111 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.175 $Y=2.125
+ $X2=3.25 $Y2=2.05
r112 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.175 $Y=2.125
+ $X2=2.895 $Y2=2.125
r113 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.175 $Y=1.165
+ $X2=3.25 $Y2=1.24
r114 18 19 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.175 $Y=1.165
+ $X2=2.885 $Y2=1.165
r115 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=1.09
+ $X2=2.885 $Y2=1.165
r116 15 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.81 $Y=1.09
+ $X2=2.81 $Y2=0.805
r117 14 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.81 $Y=0.255
+ $X2=2.81 $Y2=0.805
r118 11 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.805 $Y=2.2
+ $X2=2.895 $Y2=2.125
r119 11 13 117.822 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=2.805 $Y=2.2
+ $X2=2.805 $Y2=2.64
r120 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.735 $Y=0.18
+ $X2=2.81 $Y2=0.255
r121 9 10 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=2.735 $Y=0.18
+ $X2=0.985 $Y2=0.18
r122 7 27 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=0.955 $Y=2.64
+ $X2=0.955 $Y2=1.795
r123 4 25 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.91 $Y=0.805
+ $X2=0.91 $Y2=1.125
r124 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.985 $Y2=0.18
r125 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.91 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%CLK_N 3 6 8 11 12 13
c42 12 0 1.13063e-19 $X=3.73 $Y=1.515
c43 11 0 3.06916e-19 $X=3.73 $Y=1.515
r44 11 14 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.735 $Y=1.515
+ $X2=3.735 $Y2=1.68
r45 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.735 $Y=1.515
+ $X2=3.735 $Y2=1.35
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.515 $X2=3.73 $Y2=1.515
r47 8 12 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=1.515
r48 6 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.815 $Y=2.4
+ $X2=3.815 $Y2=1.68
r49 3 13 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.8 $Y=0.86 $X2=3.8
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_1007_366# 1 2 3 12 16 17 18 20 23 27 30
+ 32 33 34 36 38 41 43 47 51 55 56 58 60 63 64 65 69 71 76
c192 65 0 4.51061e-21 $X=9.07 $Y=2.035
c193 56 0 1.26757e-20 $X=5.2 $Y=1.995
c194 55 0 3.62521e-20 $X=5.2 $Y=1.995
c195 51 0 1.46444e-19 $X=9.78 $Y=1.745
c196 23 0 8.54043e-20 $X=9.435 $Y=0.9
c197 16 0 8.01569e-20 $X=5.775 $Y=1.195
r198 67 69 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=9.07 $Y=2.21
+ $X2=9.07 $Y2=2.265
r199 65 67 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=9.07 $Y=2.035
+ $X2=9.07 $Y2=2.21
r200 62 63 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.077 $Y=0.945
+ $X2=8.077 $Y2=1.115
r201 60 61 14.878 $w=2.46e-07 $l=3e-07 $layer=LI1_cond $X=7.66 $Y=2.9 $X2=7.96
+ $Y2=2.9
r202 56 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.995
+ $X2=5.2 $Y2=2.16
r203 56 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.995
+ $X2=5.2 $Y2=1.83
r204 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.995 $X2=5.2 $Y2=1.995
r205 52 76 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.78 $Y=1.745
+ $X2=9.855 $Y2=1.745
r206 52 73 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=9.78 $Y=1.745
+ $X2=9.435 $Y2=1.745
r207 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.745 $X2=9.78 $Y2=1.745
r208 49 51 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.78 $Y=1.95
+ $X2=9.78 $Y2=1.745
r209 48 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.235 $Y=2.035
+ $X2=9.07 $Y2=2.035
r210 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.615 $Y=2.035
+ $X2=9.78 $Y2=1.95
r211 47 48 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.615 $Y=2.035
+ $X2=9.235 $Y2=2.035
r212 44 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=2.21
+ $X2=7.96 $Y2=2.21
r213 43 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.905 $Y=2.21
+ $X2=9.07 $Y2=2.21
r214 43 44 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=8.905 $Y=2.21
+ $X2=8.045 $Y2=2.21
r215 41 62 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.86
+ $X2=8.115 $Y2=0.945
r216 38 61 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.96 $Y=2.73
+ $X2=7.96 $Y2=2.9
r217 37 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=2.295
+ $X2=7.96 $Y2=2.21
r218 37 38 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.96 $Y=2.295
+ $X2=7.96 $Y2=2.73
r219 36 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=2.125
+ $X2=7.96 $Y2=2.21
r220 36 63 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=7.96 $Y=2.125
+ $X2=7.96 $Y2=1.115
r221 34 58 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=7.072 $Y=2.902
+ $X2=6.9 $Y2=2.902
r222 33 60 1.26986 $w=3.45e-07 $l=7.93725e-09 $layer=LI1_cond $X=7.653 $Y=2.902
+ $X2=7.66 $Y2=2.9
r223 33 34 19.4078 $w=3.43e-07 $l=5.81e-07 $layer=LI1_cond $X=7.653 $Y=2.902
+ $X2=7.072 $Y2=2.902
r224 32 58 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.555 $Y=2.99
+ $X2=6.9 $Y2=2.99
r225 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.47 $Y=2.905
+ $X2=5.555 $Y2=2.99
r226 29 55 11.5986 $w=2.84e-07 $l=3.46627e-07 $layer=LI1_cond $X=5.47 $Y=2.18
+ $X2=5.2 $Y2=2.005
r227 29 30 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.47 $Y=2.18
+ $X2=5.47 $Y2=2.905
r228 25 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.855 $Y=1.91
+ $X2=9.855 $Y2=1.745
r229 25 27 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=9.855 $Y=1.91
+ $X2=9.855 $Y2=2.54
r230 21 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.435 $Y=1.58
+ $X2=9.435 $Y2=1.745
r231 21 23 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.435 $Y=1.58
+ $X2=9.435 $Y2=0.9
r232 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.85 $Y=1.12
+ $X2=5.85 $Y2=0.835
r233 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.775 $Y=1.195
+ $X2=5.85 $Y2=1.12
r234 16 17 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.775 $Y=1.195
+ $X2=5.355 $Y2=1.195
r235 14 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.28 $Y=1.27
+ $X2=5.355 $Y2=1.195
r236 14 71 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.28 $Y=1.27
+ $X2=5.28 $Y2=1.83
r237 12 72 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.275 $Y=2.53
+ $X2=5.275 $Y2=2.16
r238 3 69 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.935
+ $Y=2.12 $X2=9.07 $Y2=2.265
r239 2 60 300 $w=1.7e-07 $l=1.03049e-06 $layer=licon1_PDIFF $count=2 $X=6.92
+ $Y=2.12 $X2=7.66 $Y2=2.815
r240 1 41 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.625 $X2=8.115 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_871_368# 1 2 9 13 17 21 25 31 33 39 40 43
+ 44 45 47 48 49 51 52 58 59 62 70 77
c202 77 0 1.26757e-20 $X=5.855 $Y=1.265
c203 70 0 1.62439e-20 $X=10.32 $Y=1.59
c204 62 0 1.15277e-19 $X=5.76 $Y=1.675
c205 52 0 1.27085e-19 $X=6.145 $Y=1.295
c206 51 0 6.70526e-20 $X=10.175 $Y=1.295
c207 47 0 9.35685e-20 $X=6.66 $Y=1.69
c208 21 0 1.08678e-19 $X=11.16 $Y=0.62
r209 71 85 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=10.32 $Y=1.59
+ $X2=10.32 $Y2=1.43
r210 70 73 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.32 $Y=1.59
+ $X2=10.32 $Y2=1.755
r211 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.32
+ $Y=1.59 $X2=10.32 $Y2=1.59
r212 63 81 0.161011 $w=5.18e-07 $l=7e-09 $layer=LI1_cond $X=5.855 $Y=1.675
+ $X2=5.855 $Y2=1.682
r213 62 65 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.76 $Y=1.675
+ $X2=5.76 $Y2=1.84
r214 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.675 $X2=5.76 $Y2=1.675
r215 59 85 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.43
r216 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.295
r217 55 63 8.74057 $w=5.18e-07 $l=3.8e-07 $layer=LI1_cond $X=5.855 $Y=1.295
+ $X2=5.855 $Y2=1.675
r218 55 77 0.690045 $w=5.18e-07 $l=3e-08 $layer=LI1_cond $X=5.855 $Y=1.295
+ $X2=5.855 $Y2=1.265
r219 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=1.295 $X2=6
+ $Y2=1.295
r220 52 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=1.295
+ $X2=6 $Y2=1.295
r221 51 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=10.32 $Y2=1.295
r222 51 52 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=6.145 $Y2=1.295
r223 48 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.66 $Y=1.69
+ $X2=6.66 $Y2=1.525
r224 47 49 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.66 $Y=1.69
+ $X2=6.495 $Y2=1.69
r225 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.69 $X2=6.66 $Y2=1.69
r226 43 44 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.595 $Y=2.005
+ $X2=4.595 $Y2=1.84
r227 40 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.22 $Y=1.43
+ $X2=11.22 $Y2=1.265
r228 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.22
+ $Y=1.43 $X2=11.22 $Y2=1.43
r229 37 85 1.29116 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=1.43
+ $X2=10.32 $Y2=1.43
r230 37 39 28.2349 $w=2.98e-07 $l=7.35e-07 $layer=LI1_cond $X=10.485 $Y=1.43
+ $X2=11.22 $Y2=1.43
r231 36 81 3.68146 $w=3.15e-07 $l=2.6e-07 $layer=LI1_cond $X=6.115 $Y=1.682
+ $X2=5.855 $Y2=1.682
r232 36 49 13.9025 $w=3.13e-07 $l=3.8e-07 $layer=LI1_cond $X=6.115 $Y=1.682
+ $X2=6.495 $Y2=1.682
r233 34 45 2.11342 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.94 $Y=1.265
+ $X2=4.777 $Y2=1.265
r234 33 77 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=5.595 $Y=1.265
+ $X2=5.855 $Y2=1.265
r235 33 34 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.595 $Y=1.265
+ $X2=4.94 $Y2=1.265
r236 29 45 4.3182 $w=2.1e-07 $l=1.0225e-07 $layer=LI1_cond $X=4.815 $Y=1.18
+ $X2=4.777 $Y2=1.265
r237 29 31 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=4.815 $Y=1.18
+ $X2=4.815 $Y2=0.76
r238 27 45 4.3182 $w=2.1e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.7 $Y=1.35
+ $X2=4.777 $Y2=1.265
r239 27 44 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.7 $Y=1.35 $X2=4.7
+ $Y2=1.84
r240 23 43 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.595 $Y=2.03
+ $X2=4.595 $Y2=2.005
r241 23 25 23.807 $w=3.78e-07 $l=7.85e-07 $layer=LI1_cond $X=4.595 $Y=2.03
+ $X2=4.595 $Y2=2.815
r242 21 75 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=11.16 $Y=0.62
+ $X2=11.16 $Y2=1.265
r243 17 73 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=10.245 $Y=2.54
+ $X2=10.245 $Y2=1.755
r244 13 67 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.665 $Y=0.835
+ $X2=6.665 $Y2=1.525
r245 9 65 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.695 $Y=2.53
+ $X2=5.695 $Y2=1.84
r246 2 43 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=4.355
+ $Y=1.84 $X2=4.49 $Y2=2.005
r247 2 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.355
+ $Y=1.84 $X2=4.49 $Y2=2.815
r248 1 31 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=4.715
+ $Y=0.49 $X2=4.855 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_1157_464# 1 2 7 8 11 13 15 17 20 22 23 26
+ 28 29 33 34
c98 29 0 8.01569e-20 $X=6.615 $Y=1.27
c99 26 0 1.27085e-19 $X=6.45 $Y=0.835
c100 8 0 6.70526e-20 $X=7.365 $Y=1.36
r101 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.2
+ $Y=1.45 $X2=7.2 $Y2=1.45
r102 31 33 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=7.2 $Y=2.04 $X2=7.2
+ $Y2=1.45
r103 30 33 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.2 $Y=1.355
+ $X2=7.2 $Y2=1.45
r104 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.035 $Y=1.27
+ $X2=7.2 $Y2=1.355
r105 28 29 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.035 $Y=1.27
+ $X2=6.615 $Y2=1.27
r106 24 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.45 $Y=1.185
+ $X2=6.615 $Y2=1.27
r107 24 26 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.45 $Y=1.185
+ $X2=6.45 $Y2=0.835
r108 22 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.035 $Y=2.125
+ $X2=7.2 $Y2=2.04
r109 22 23 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=7.035 $Y=2.125
+ $X2=6.17 $Y2=2.125
r110 18 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.005 $Y=2.21
+ $X2=6.17 $Y2=2.125
r111 18 20 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.005 $Y=2.21
+ $X2=6.005 $Y2=2.515
r112 16 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.2 $Y=1.435
+ $X2=7.2 $Y2=1.45
r113 13 17 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.9 $Y=1.285
+ $X2=7.885 $Y2=1.36
r114 13 15 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.9 $Y=1.285
+ $X2=7.9 $Y2=0.9
r115 9 17 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.885 $Y=1.435
+ $X2=7.885 $Y2=1.36
r116 9 11 429.524 $w=1.8e-07 $l=1.105e-06 $layer=POLY_cond $X=7.885 $Y=1.435
+ $X2=7.885 $Y2=2.54
r117 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.365 $Y=1.36
+ $X2=7.2 $Y2=1.435
r118 7 17 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.795 $Y=1.36
+ $X2=7.885 $Y2=1.36
r119 7 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.795 $Y=1.36
+ $X2=7.365 $Y2=1.36
r120 2 20 600 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=2.32 $X2=6.005 $Y2=2.515
r121 1 26 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.625 $X2=6.45 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_1643_257# 1 2 9 13 16 20 22 23 24 27 30
+ 31 32 34 35 36 37 41 44 47 51 52 53 57 58 61 63 67 71
c201 71 0 1.11129e-19 $X=12.66 $Y=1.22
c202 58 0 1.91513e-19 $X=12.66 $Y=1.13
c203 57 0 1.28025e-19 $X=12.66 $Y=1.215
c204 32 0 7.74904e-20 $X=9.725 $Y=0.345
c205 24 0 4.51061e-21 $X=8.38 $Y=1.955
r206 64 67 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=13.69 $Y=2.17
+ $X2=13.91 $Y2=2.17
r207 61 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.66 $Y=1.385
+ $X2=12.66 $Y2=1.55
r208 61 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.66 $Y=1.385
+ $X2=12.66 $Y2=1.22
r209 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.66
+ $Y=1.385 $X2=12.66 $Y2=1.385
r210 57 60 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.66 $Y=1.215
+ $X2=12.66 $Y2=1.385
r211 57 58 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=12.66 $Y=1.215
+ $X2=12.66 $Y2=1.13
r212 53 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.98 $Y=0.685
+ $X2=11.98 $Y2=0.855
r213 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.38
+ $Y=1.45 $X2=8.38 $Y2=1.45
r214 45 63 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.775 $Y=1.17
+ $X2=13.69 $Y2=1.17
r215 45 47 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=13.775 $Y=1.17
+ $X2=13.985 $Y2=1.17
r216 44 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.69 $Y=2.005
+ $X2=13.69 $Y2=2.17
r217 43 63 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.69 $Y=1.335
+ $X2=13.69 $Y2=1.17
r218 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.69 $Y=1.335
+ $X2=13.69 $Y2=2.005
r219 42 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.825 $Y=1.215
+ $X2=12.66 $Y2=1.215
r220 41 63 3.70735 $w=2.5e-07 $l=1.05119e-07 $layer=LI1_cond $X=13.605 $Y=1.215
+ $X2=13.69 $Y2=1.17
r221 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.605 $Y=1.215
+ $X2=12.825 $Y2=1.215
r222 39 58 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.58 $Y=0.94
+ $X2=12.58 $Y2=1.13
r223 38 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.065 $Y=0.855
+ $X2=11.98 $Y2=0.855
r224 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.495 $Y=0.855
+ $X2=12.58 $Y2=0.94
r225 37 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.495 $Y=0.855
+ $X2=12.065 $Y2=0.855
r226 35 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.895 $Y=0.685
+ $X2=11.98 $Y2=0.685
r227 35 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.895 $Y=0.685
+ $X2=11.51 $Y2=0.685
r228 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.425 $Y=0.6
+ $X2=11.51 $Y2=0.685
r229 33 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.425 $Y=0.43
+ $X2=11.425 $Y2=0.6
r230 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.34 $Y=0.345
+ $X2=11.425 $Y2=0.43
r231 31 32 105.364 $w=1.68e-07 $l=1.615e-06 $layer=LI1_cond $X=11.34 $Y=0.345
+ $X2=9.725 $Y2=0.345
r232 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.64 $Y=0.43
+ $X2=9.725 $Y2=0.345
r233 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.64 $Y=0.43
+ $X2=9.64 $Y2=1.11
r234 28 51 10.5458 $w=2.95e-07 $l=3.41746e-07 $layer=LI1_cond $X=8.62 $Y=1.195
+ $X2=8.417 $Y2=1.45
r235 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.555 $Y=1.195
+ $X2=9.64 $Y2=1.11
r236 27 28 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=9.555 $Y=1.195 $X2=8.62
+ $Y2=1.195
r237 23 52 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.38 $Y=1.79
+ $X2=8.38 $Y2=1.45
r238 23 24 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.38 $Y=1.79
+ $X2=8.38 $Y2=1.955
r239 22 52 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.38 $Y=1.285
+ $X2=8.38 $Y2=1.45
r240 20 71 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.705 $Y=0.74
+ $X2=12.705 $Y2=1.22
r241 16 72 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=12.705 $Y=2.46
+ $X2=12.705 $Y2=1.55
r242 13 22 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.33 $Y=0.9
+ $X2=8.33 $Y2=1.285
r243 9 24 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=8.305 $Y=2.54
+ $X2=8.305 $Y2=1.955
r244 2 67 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.765
+ $Y=1.995 $X2=13.91 $Y2=2.17
r245 1 47 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=13.845
+ $Y=0.9 $X2=13.985 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%SET_B 3 7 11 15 16 17 20 22 25 30 31 32
c133 32 0 1.96837e-19 $X=12.12 $Y=1.22
c134 31 0 1.11129e-19 $X=12.12 $Y=1.385
c135 25 0 1.46444e-19 $X=8.955 $Y=1.615
c136 16 0 1.54515e-19 $X=12.095 $Y=1.665
r137 31 41 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=12.14 $Y=1.385
+ $X2=12.14 $Y2=1.665
r138 30 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.12 $Y=1.385
+ $X2=12.12 $Y2=1.55
r139 30 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.12 $Y=1.385
+ $X2=12.12 $Y2=1.22
r140 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.12
+ $Y=1.385 $X2=12.12 $Y2=1.385
r141 25 28 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.937 $Y=1.615
+ $X2=8.937 $Y2=1.78
r142 25 27 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.937 $Y=1.615
+ $X2=8.937 $Y2=1.45
r143 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.955
+ $Y=1.615 $X2=8.955 $Y2=1.615
r144 22 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=1.665
+ $X2=12.24 $Y2=1.665
r145 20 26 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=9.36 $Y=1.615
+ $X2=8.955 $Y2=1.615
r146 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r147 17 19 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.505 $Y=1.665
+ $X2=9.36 $Y2=1.665
r148 16 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=12.24 $Y2=1.665
r149 16 17 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=9.505 $Y2=1.665
r150 15 32 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.185 $Y=0.74
+ $X2=12.185 $Y2=1.22
r151 11 33 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=12.195 $Y=2.46
+ $X2=12.195 $Y2=1.55
r152 7 27 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.935 $Y=0.9
+ $X2=8.935 $Y2=1.45
r153 3 28 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=8.845 $Y=2.54
+ $X2=8.845 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_688_98# 1 2 9 14 15 16 20 23 24 29 30 31
+ 32 34 38 40 41 42 46 48 50 55 59 61 66
c176 66 0 1.16265e-19 $X=4.64 $Y=1.505
c177 32 0 1.32086e-19 $X=10.78 $Y=2.085
c178 20 0 9.35685e-20 $X=6.21 $Y=0.835
c179 9 0 1.13063e-19 $X=4.265 $Y=2.4
r180 60 66 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.28 $Y=1.505
+ $X2=4.64 $Y2=1.505
r181 60 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.28 $Y=1.505
+ $X2=4.265 $Y2=1.505
r182 59 62 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=1.505
+ $X2=4.255 $Y2=1.67
r183 59 61 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=1.505
+ $X2=4.255 $Y2=1.34
r184 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=1.505 $X2=4.28 $Y2=1.505
r185 55 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.15 $Y=1.95
+ $X2=4.15 $Y2=1.67
r186 52 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.15 $Y=1.17
+ $X2=4.15 $Y2=1.34
r187 51 57 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.675 $Y=2.035
+ $X2=3.55 $Y2=2.035
r188 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=2.035
+ $X2=4.15 $Y2=1.95
r189 50 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.065 $Y=2.035
+ $X2=3.675 $Y2=2.035
r190 46 57 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.12
+ $X2=3.55 $Y2=2.035
r191 46 48 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.55 $Y=2.12
+ $X2=3.55 $Y2=2.815
r192 42 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=1.085
+ $X2=4.15 $Y2=1.17
r193 42 44 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.065 $Y=1.085
+ $X2=3.585 $Y2=1.085
r194 39 40 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.227 $Y=2.095
+ $X2=6.227 $Y2=2.245
r195 36 41 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.77 $Y=1.185
+ $X2=10.77 $Y2=1.995
r196 32 41 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.78 $Y=2.085
+ $X2=10.78 $Y2=1.995
r197 32 34 258.492 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=10.78 $Y=2.085
+ $X2=10.78 $Y2=2.75
r198 30 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.695 $Y=1.11
+ $X2=10.77 $Y2=1.185
r199 30 31 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=10.695 $Y=1.11
+ $X2=9.985 $Y2=1.11
r200 27 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.91 $Y=1.035
+ $X2=9.985 $Y2=1.11
r201 27 29 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.91 $Y=1.035
+ $X2=9.91 $Y2=0.685
r202 26 29 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.91 $Y=0.255
+ $X2=9.91 $Y2=0.685
r203 25 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.285 $Y=0.18
+ $X2=6.21 $Y2=0.18
r204 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.835 $Y=0.18
+ $X2=9.91 $Y2=0.255
r205 24 25 1820.32 $w=1.5e-07 $l=3.55e-06 $layer=POLY_cond $X=9.835 $Y=0.18
+ $X2=6.285 $Y2=0.18
r206 23 40 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.23 $Y=2.64
+ $X2=6.23 $Y2=2.245
r207 20 39 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=6.21 $Y=0.835
+ $X2=6.21 $Y2=2.095
r208 17 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.21 $Y=0.255
+ $X2=6.21 $Y2=0.18
r209 17 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.21 $Y=0.255
+ $X2=6.21 $Y2=0.835
r210 15 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.135 $Y=0.18
+ $X2=6.21 $Y2=0.18
r211 15 16 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=6.135 $Y=0.18
+ $X2=4.715 $Y2=0.18
r212 12 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.64 $Y=1.34
+ $X2=4.64 $Y2=1.505
r213 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.64 $Y=1.34
+ $X2=4.64 $Y2=0.86
r214 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.64 $Y=0.255
+ $X2=4.715 $Y2=0.18
r215 11 14 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=4.64 $Y=0.255
+ $X2=4.64 $Y2=0.86
r216 7 63 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.67
+ $X2=4.265 $Y2=1.505
r217 7 9 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=4.265 $Y=1.67
+ $X2=4.265 $Y2=2.4
r218 2 57 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.59 $Y2=2.115
r219 2 48 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.59 $Y2=2.815
r220 1 44 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.49 $X2=3.585 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_2216_410# 1 2 3 12 14 16 18 20 25 29 33
+ 37 39 40 43 47 51 54 58 59 63 65 69 71 73 76 78 84 88 90 96 98 100 104
c213 51 0 7.20841e-20 $X=11.67 $Y=0.98
c214 20 0 2.75443e-20 $X=11.67 $Y=2.05
r215 97 104 10.142 $w=3.3e-07 $l=5.8e-08 $layer=POLY_cond $X=14.65 $Y=1.595
+ $X2=14.65 $Y2=1.537
r216 96 99 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.65 $Y=1.595
+ $X2=14.65 $Y2=1.76
r217 96 98 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.65 $Y=1.595
+ $X2=14.65 $Y2=1.43
r218 96 97 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.65
+ $Y=1.595 $X2=14.65 $Y2=1.595
r219 92 93 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=13.31 $Y=2.345
+ $X2=13.31 $Y2=2.59
r220 90 92 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=13.31 $Y=2.225
+ $X2=13.31 $Y2=2.345
r221 86 88 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=12.92 $Y=0.777
+ $X2=13.085 $Y2=0.777
r222 79 103 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.245 $Y=2.215
+ $X2=11.245 $Y2=2.38
r223 79 100 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.245 $Y=2.215
+ $X2=11.245 $Y2=2.125
r224 78 81 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=11.245 $Y=2.215
+ $X2=11.245 $Y2=2.345
r225 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.245
+ $Y=2.215 $X2=11.245 $Y2=2.215
r226 76 99 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=14.57 $Y=2.505
+ $X2=14.57 $Y2=1.76
r227 73 94 13.6427 $w=2.52e-07 $l=2.93581e-07 $layer=LI1_cond $X=14.57 $Y=1.005
+ $X2=14.487 $Y2=0.75
r228 73 98 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=14.57 $Y=1.005
+ $X2=14.57 $Y2=1.43
r229 72 93 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.435 $Y=2.59
+ $X2=13.31 $Y2=2.59
r230 71 76 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.485 $Y=2.59
+ $X2=14.57 $Y2=2.505
r231 71 72 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=14.485 $Y=2.59
+ $X2=13.435 $Y2=2.59
r232 67 93 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=13.31 $Y=2.675
+ $X2=13.31 $Y2=2.59
r233 67 69 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=13.31 $Y=2.675
+ $X2=13.31 $Y2=2.815
r234 65 94 3.04159 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=14.32 $Y=0.75
+ $X2=14.487 $Y2=0.75
r235 65 88 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=14.32 $Y=0.75
+ $X2=13.085 $Y2=0.75
r236 64 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=2.345
+ $X2=11.97 $Y2=2.345
r237 63 92 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.185 $Y=2.345
+ $X2=13.31 $Y2=2.345
r238 63 64 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=13.185 $Y=2.345
+ $X2=12.135 $Y2=2.345
r239 60 81 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.41 $Y=2.345
+ $X2=11.245 $Y2=2.345
r240 59 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.805 $Y=2.345
+ $X2=11.97 $Y2=2.345
r241 59 60 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.805 $Y=2.345
+ $X2=11.41 $Y2=2.345
r242 49 51 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=11.55 $Y=0.98
+ $X2=11.67 $Y2=0.98
r243 45 58 32.0891 $w=1.65e-07 $l=4.4379e-07 $layer=POLY_cond $X=16.76 $Y=1.74
+ $X2=16.645 $Y2=1.35
r244 45 47 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=16.76 $Y=1.74
+ $X2=16.76 $Y2=2.42
r245 41 58 32.0891 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=16.72 $Y=1.35
+ $X2=16.645 $Y2=1.35
r246 41 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.72 $Y=1.35
+ $X2=16.72 $Y2=0.79
r247 40 57 18.3011 $w=2.95e-07 $l=9e-08 $layer=POLY_cond $X=15.855 $Y=1.497
+ $X2=15.765 $Y2=1.497
r248 39 58 2.52421 $w=2.95e-07 $l=1.47e-07 $layer=POLY_cond $X=16.645 $Y=1.497
+ $X2=16.645 $Y2=1.35
r249 39 40 160.643 $w=2.95e-07 $l=7.9e-07 $layer=POLY_cond $X=16.645 $Y=1.497
+ $X2=15.855 $Y2=1.497
r250 35 57 14.3312 $w=1.8e-07 $l=1.48e-07 $layer=POLY_cond $X=15.765 $Y=1.645
+ $X2=15.765 $Y2=1.497
r251 35 37 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=15.765 $Y=1.645
+ $X2=15.765 $Y2=2.4
r252 31 57 21.3513 $w=2.95e-07 $l=1.05e-07 $layer=POLY_cond $X=15.66 $Y=1.497
+ $X2=15.765 $Y2=1.497
r253 31 55 70.1542 $w=2.95e-07 $l=3.45e-07 $layer=POLY_cond $X=15.66 $Y=1.497
+ $X2=15.315 $Y2=1.497
r254 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=15.66 $Y=1.35
+ $X2=15.66 $Y2=0.74
r255 27 55 14.3312 $w=1.8e-07 $l=1.48e-07 $layer=POLY_cond $X=15.315 $Y=1.645
+ $X2=15.315 $Y2=1.497
r256 27 29 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=15.315 $Y=1.645
+ $X2=15.315 $Y2=2.4
r257 23 55 17.2844 $w=2.95e-07 $l=8.5e-08 $layer=POLY_cond $X=15.23 $Y=1.497
+ $X2=15.315 $Y2=1.497
r258 23 54 19.7714 $w=2.95e-07 $l=7.5e-08 $layer=POLY_cond $X=15.23 $Y=1.497
+ $X2=15.155 $Y2=1.497
r259 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=15.23 $Y=1.35
+ $X2=15.23 $Y2=0.74
r260 22 104 12.8918 $w=2.15e-07 $l=1.65e-07 $layer=POLY_cond $X=14.815 $Y=1.537
+ $X2=14.65 $Y2=1.537
r261 22 54 101.481 $w=2.15e-07 $l=3.4e-07 $layer=POLY_cond $X=14.815 $Y=1.537
+ $X2=15.155 $Y2=1.537
r262 19 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.67 $Y=1.055
+ $X2=11.67 $Y2=0.98
r263 19 20 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=11.67 $Y=1.055
+ $X2=11.67 $Y2=2.05
r264 16 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.55 $Y=0.905
+ $X2=11.55 $Y2=0.98
r265 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.55 $Y=0.905
+ $X2=11.55 $Y2=0.62
r266 15 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.41 $Y=2.125
+ $X2=11.245 $Y2=2.125
r267 14 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.595 $Y=2.125
+ $X2=11.67 $Y2=2.05
r268 14 15 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=11.595 $Y=2.125
+ $X2=11.41 $Y2=2.125
r269 12 103 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=11.17 $Y=2.75
+ $X2=11.17 $Y2=2.38
r270 3 90 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=13.215
+ $Y=1.96 $X2=13.35 $Y2=2.225
r271 3 69 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=13.215
+ $Y=1.96 $X2=13.35 $Y2=2.815
r272 2 84 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=11.825
+ $Y=1.96 $X2=11.97 $Y2=2.425
r273 1 86 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=12.78
+ $Y=0.37 $X2=12.92 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_1997_82# 1 2 9 13 21 24 25 26 27 30 31 33
+ 38 41 45 47 52 53
c156 41 0 1.85877e-19 $X=10.945 $Y=0.685
c157 26 0 1.62439e-20 $X=10.91 $Y=1.835
r158 53 59 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.2 $Y=1.635
+ $X2=13.2 $Y2=1.8
r159 53 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.2 $Y=1.635
+ $X2=13.2 $Y2=1.47
r160 52 55 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=13.2 $Y=1.635
+ $X2=13.2 $Y2=1.805
r161 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.2
+ $Y=1.635 $X2=13.2 $Y2=1.635
r162 47 49 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=12.58 $Y=1.805
+ $X2=12.58 $Y2=2.005
r163 45 46 11.3956 $w=1.82e-07 $l=1.7e-07 $layer=LI1_cond $X=11.652 $Y=1.835
+ $X2=11.652 $Y2=2.005
r164 41 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.025 $Y=0.685
+ $X2=11.025 $Y2=1.025
r165 36 38 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.47 $Y=2.185
+ $X2=10.825 $Y2=2.185
r166 34 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.665 $Y=1.805
+ $X2=12.58 $Y2=1.805
r167 33 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.035 $Y=1.805
+ $X2=13.2 $Y2=1.805
r168 33 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.035 $Y=1.805
+ $X2=12.665 $Y2=1.805
r169 32 46 1.129 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=11.75 $Y=2.005
+ $X2=11.652 $Y2=2.005
r170 31 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.495 $Y=2.005
+ $X2=12.58 $Y2=2.005
r171 31 32 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=12.495 $Y=2.005
+ $X2=11.75 $Y2=2.005
r172 30 45 5.7679 $w=1.82e-07 $l=9.0802e-08 $layer=LI1_cond $X=11.64 $Y=1.75
+ $X2=11.652 $Y2=1.835
r173 29 30 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=11.64 $Y=1.11
+ $X2=11.64 $Y2=1.75
r174 28 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.11 $Y=1.025
+ $X2=11.025 $Y2=1.025
r175 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.555 $Y=1.025
+ $X2=11.64 $Y2=1.11
r176 27 28 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=11.555 $Y=1.025
+ $X2=11.11 $Y2=1.025
r177 25 45 1.129 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=11.555 $Y=1.835
+ $X2=11.652 $Y2=1.835
r178 25 26 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=11.555 $Y=1.835
+ $X2=10.91 $Y2=1.835
r179 24 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.825 $Y=2.1
+ $X2=10.825 $Y2=2.185
r180 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.825 $Y=1.92
+ $X2=10.91 $Y2=1.835
r181 23 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.825 $Y=1.92
+ $X2=10.825 $Y2=2.1
r182 21 36 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=10.47 $Y=2.815
+ $X2=10.47 $Y2=2.27
r183 17 41 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=10.125 $Y=0.725
+ $X2=10.94 $Y2=0.725
r184 13 58 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=13.135 $Y=0.74
+ $X2=13.135 $Y2=1.47
r185 9 59 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=13.125 $Y=2.46
+ $X2=13.125 $Y2=1.8
r186 2 36 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.335
+ $Y=2.12 $X2=10.47 $Y2=2.265
r187 2 21 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=10.335
+ $Y=2.12 $X2=10.47 $Y2=2.815
r188 1 41 91 $w=1.7e-07 $l=1.08885e-06 $layer=licon1_NDIFF $count=2 $X=9.985
+ $Y=0.41 $X2=10.945 $Y2=0.685
r189 1 17 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.985
+ $Y=0.41 $X2=10.125 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%RESET_B 3 7 9 12
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.11 $Y=1.67
+ $X2=14.11 $Y2=1.835
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.11 $Y=1.67
+ $X2=14.11 $Y2=1.505
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.11
+ $Y=1.67 $X2=14.11 $Y2=1.67
r39 7 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=14.2 $Y=1.11
+ $X2=14.2 $Y2=1.505
r40 3 15 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=14.135 $Y=2.315
+ $X2=14.135 $Y2=1.835
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_3272_94# 1 2 9 11 13 16 18 20 23 27 33 36
+ 42
c68 27 0 1.7776e-19 $X=16.535 $Y=2.065
r69 41 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=17.735 $Y=1.385
+ $X2=17.75 $Y2=1.385
r70 40 41 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=17.32 $Y=1.385
+ $X2=17.735 $Y2=1.385
r71 39 40 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=17.285 $Y=1.385
+ $X2=17.32 $Y2=1.385
r72 34 39 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=17.2 $Y=1.385
+ $X2=17.285 $Y2=1.385
r73 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.2
+ $Y=1.385 $X2=17.2 $Y2=1.385
r74 31 36 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=16.7 $Y=1.385
+ $X2=16.52 $Y2=1.385
r75 31 33 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=16.7 $Y=1.385 $X2=17.2
+ $Y2=1.385
r76 27 29 22.7287 $w=3.58e-07 $l=7.1e-07 $layer=LI1_cond $X=16.52 $Y=2.065
+ $X2=16.52 $Y2=2.775
r77 25 36 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=16.52 $Y=1.55
+ $X2=16.52 $Y2=1.385
r78 25 27 16.4863 $w=3.58e-07 $l=5.15e-07 $layer=LI1_cond $X=16.52 $Y=1.55
+ $X2=16.52 $Y2=2.065
r79 21 36 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=16.505 $Y=1.22
+ $X2=16.52 $Y2=1.385
r80 21 23 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=16.505 $Y=1.22
+ $X2=16.505 $Y2=0.645
r81 18 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.75 $Y=1.22
+ $X2=17.75 $Y2=1.385
r82 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.75 $Y=1.22
+ $X2=17.75 $Y2=0.74
r83 14 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=17.735 $Y=1.55
+ $X2=17.735 $Y2=1.385
r84 14 16 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=17.735 $Y=1.55
+ $X2=17.735 $Y2=2.4
r85 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.32 $Y=1.22
+ $X2=17.32 $Y2=1.385
r86 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.32 $Y=1.22
+ $X2=17.32 $Y2=0.74
r87 7 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=17.285 $Y=1.55
+ $X2=17.285 $Y2=1.385
r88 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=17.285 $Y=1.55
+ $X2=17.285 $Y2=2.4
r89 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=16.395
+ $Y=1.92 $X2=16.535 $Y2=2.775
r90 2 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=16.395
+ $Y=1.92 $X2=16.535 $Y2=2.065
r91 1 23 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=16.36
+ $Y=0.47 $X2=16.505 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_27_464# 1 2 9 12 13 14 17 20
r42 15 17 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.02 $Y=2.905
+ $X2=2.02 $Y2=2.465
r43 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.855 $Y=2.99
+ $X2=2.02 $Y2=2.905
r44 13 14 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.855 $Y=2.99
+ $X2=1.235 $Y2=2.99
r45 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.905
+ $X2=1.235 $Y2=2.99
r46 11 12 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.15 $Y=2.475
+ $X2=1.15 $Y2=2.905
r47 10 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.39
+ $X2=0.24 $Y2=2.39
r48 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.39
+ $X2=1.15 $Y2=2.475
r49 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.065 $Y=2.39 $X2=0.365
+ $Y2=2.39
r50 2 17 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.885
+ $Y=2.32 $X2=2.02 $Y2=2.465
r51 1 20 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 39 43 47 49
+ 53 57 61 65 69 73 77 83 87 89 94 95 97 98 100 101 102 104 109 117 122 131 150
+ 154 160 163 166 169 172 175 179 186 188 192
c209 47 0 1.16265e-19 $X=4.04 $Y=2.425
c210 43 0 7.30946e-20 $X=2.58 $Y=2.465
r211 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=3.33 $X2=18
+ $Y2=3.33
r212 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r213 185 186 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.005 $Y=3.13
+ $X2=15.17 $Y2=3.13
r214 183 185 0.167871 $w=5.68e-07 $l=8e-09 $layer=LI1_cond $X=14.997 $Y=3.13
+ $X2=15.005 $Y2=3.13
r215 181 183 7.49123 $w=5.68e-07 $l=3.57e-07 $layer=LI1_cond $X=14.64 $Y=3.13
+ $X2=14.997 $Y2=3.13
r216 181 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r217 178 181 4.09185 $w=5.68e-07 $l=1.95e-07 $layer=LI1_cond $X=14.445 $Y=3.13
+ $X2=14.64 $Y2=3.13
r218 178 179 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=14.445 $Y=3.13
+ $X2=14.28 $Y2=3.13
r219 175 176 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r220 172 173 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r221 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r222 167 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r223 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r224 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r225 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r226 158 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=18 $Y2=3.33
r227 158 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=17.04 $Y2=3.33
r228 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r229 155 188 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.225 $Y=3.33
+ $X2=17.06 $Y2=3.33
r230 155 157 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.225 $Y=3.33
+ $X2=17.52 $Y2=3.33
r231 154 191 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=17.875 $Y=3.33
+ $X2=18.057 $Y2=3.33
r232 154 157 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.875 $Y=3.33
+ $X2=17.52 $Y2=3.33
r233 153 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.04 $Y2=3.33
r234 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r235 150 188 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.895 $Y=3.33
+ $X2=17.06 $Y2=3.33
r236 150 152 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=16.895 $Y=3.33
+ $X2=16.56 $Y2=3.33
r237 149 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.56 $Y2=3.33
r238 149 182 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=14.64 $Y2=3.33
r239 148 186 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=15.6 $Y=3.33
+ $X2=15.17 $Y2=3.33
r240 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r241 145 182 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r242 144 179 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=14.16 $Y=3.33
+ $X2=14.28 $Y2=3.33
r243 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r244 142 145 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=14.16 $Y2=3.33
r245 141 144 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=14.16 $Y2=3.33
r246 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r247 138 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r248 138 176 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r249 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r250 135 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.56 $Y=3.33
+ $X2=11.395 $Y2=3.33
r251 135 137 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.56 $Y=3.33
+ $X2=12.24 $Y2=3.33
r252 134 176 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=11.28 $Y2=3.33
r253 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r254 131 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=11.395 $Y2=3.33
r255 131 133 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=9.84 $Y2=3.33
r256 130 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r257 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r258 127 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.53 $Y2=3.33
r259 127 129 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=9.36 $Y2=3.33
r260 126 173 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r261 126 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r262 125 126 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r263 123 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.215 $Y=3.33
+ $X2=5.09 $Y2=3.33
r264 123 125 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=3.33
+ $X2=5.52 $Y2=3.33
r265 122 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=8.53 $Y2=3.33
r266 122 125 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=5.52 $Y2=3.33
r267 121 167 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r268 121 164 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r269 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r270 118 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.58 $Y2=3.33
r271 118 120 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=3.6 $Y2=3.33
r272 117 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.04 $Y2=3.33
r273 117 120 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.6 $Y2=3.33
r274 116 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r275 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r276 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r277 113 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r278 112 115 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r279 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r280 110 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r281 110 112 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r282 109 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.58 $Y2=3.33
r283 109 115 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.16 $Y2=3.33
r284 107 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r285 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r286 104 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r287 104 106 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r288 102 130 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=9.36 $Y2=3.33
r289 102 173 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=8.4 $Y2=3.33
r290 100 148 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=15.825 $Y=3.33
+ $X2=15.6 $Y2=3.33
r291 100 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.825 $Y=3.33
+ $X2=15.99 $Y2=3.33
r292 99 152 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=16.56 $Y2=3.33
r293 99 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=15.99 $Y2=3.33
r294 97 137 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=12.305 $Y=3.33
+ $X2=12.24 $Y2=3.33
r295 97 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.305 $Y=3.33
+ $X2=12.47 $Y2=3.33
r296 96 141 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.72 $Y2=3.33
r297 96 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.47 $Y2=3.33
r298 94 129 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.36 $Y2=3.33
r299 94 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.63 $Y2=3.33
r300 93 133 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=9.795 $Y=3.33
+ $X2=9.84 $Y2=3.33
r301 93 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.795 $Y=3.33
+ $X2=9.63 $Y2=3.33
r302 89 92 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=18 $Y=1.985 $X2=18
+ $Y2=2.815
r303 87 191 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=18 $Y=3.245
+ $X2=18.057 $Y2=3.33
r304 87 92 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=18 $Y=3.245 $X2=18
+ $Y2=2.815
r305 83 86 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=17.06 $Y=2.045
+ $X2=17.06 $Y2=2.795
r306 81 188 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.06 $Y=3.245
+ $X2=17.06 $Y2=3.33
r307 81 86 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=17.06 $Y=3.245
+ $X2=17.06 $Y2=2.795
r308 77 80 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=15.99 $Y=2.115
+ $X2=15.99 $Y2=2.815
r309 75 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.99 $Y=3.245
+ $X2=15.99 $Y2=3.33
r310 75 80 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.99 $Y=3.245
+ $X2=15.99 $Y2=2.815
r311 71 183 3.68532 $w=3.45e-07 $l=2.85e-07 $layer=LI1_cond $X=14.997 $Y=2.845
+ $X2=14.997 $Y2=3.13
r312 71 73 23.2159 $w=3.43e-07 $l=6.95e-07 $layer=LI1_cond $X=14.997 $Y=2.845
+ $X2=14.997 $Y2=2.15
r313 67 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.47 $Y=3.245
+ $X2=12.47 $Y2=3.33
r314 67 69 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=12.47 $Y=3.245
+ $X2=12.47 $Y2=2.79
r315 63 175 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.395 $Y=3.245
+ $X2=11.395 $Y2=3.33
r316 63 65 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.395 $Y=3.245
+ $X2=11.395 $Y2=2.79
r317 59 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.63 $Y=3.245
+ $X2=9.63 $Y2=3.33
r318 59 61 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=9.63 $Y=3.245
+ $X2=9.63 $Y2=2.455
r319 55 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=3.245
+ $X2=8.53 $Y2=3.33
r320 55 57 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=8.53 $Y=3.245
+ $X2=8.53 $Y2=2.63
r321 51 169 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=3.245
+ $X2=5.09 $Y2=3.33
r322 51 53 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=5.09 $Y=3.245
+ $X2=5.09 $Y2=2.555
r323 50 166 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=3.33
+ $X2=4.04 $Y2=3.33
r324 49 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=5.09 $Y2=3.33
r325 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=4.205 $Y2=3.33
r326 45 166 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=3.33
r327 45 47 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.425
r328 41 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=3.245
+ $X2=2.58 $Y2=3.33
r329 41 43 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.58 $Y=3.245
+ $X2=2.58 $Y2=2.465
r330 37 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r331 37 39 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.81
r332 12 92 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=17.825
+ $Y=1.84 $X2=17.96 $Y2=2.815
r333 12 89 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=17.825
+ $Y=1.84 $X2=17.96 $Y2=1.985
r334 11 86 400 $w=1.7e-07 $l=9.74359e-07 $layer=licon1_PDIFF $count=1 $X=16.85
+ $Y=1.92 $X2=17.06 $Y2=2.795
r335 11 83 400 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=16.85
+ $Y=1.92 $X2=17.06 $Y2=2.045
r336 10 80 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=15.855
+ $Y=1.84 $X2=15.99 $Y2=2.815
r337 10 77 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=15.855
+ $Y=1.84 $X2=15.99 $Y2=2.115
r338 9 185 600 $w=1.7e-07 $l=1.34979e-06 $layer=licon1_PDIFF $count=1 $X=14.225
+ $Y=1.995 $X2=15.005 $Y2=3.01
r339 9 178 600 $w=1.7e-07 $l=1.11961e-06 $layer=licon1_PDIFF $count=1 $X=14.225
+ $Y=1.995 $X2=14.445 $Y2=3.01
r340 9 73 300 $w=1.7e-07 $l=8.53991e-07 $layer=licon1_PDIFF $count=2 $X=14.225
+ $Y=1.995 $X2=15.005 $Y2=2.15
r341 8 69 600 $w=1.7e-07 $l=9.17851e-07 $layer=licon1_PDIFF $count=1 $X=12.285
+ $Y=1.96 $X2=12.47 $Y2=2.79
r342 7 65 600 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=11.26
+ $Y=2.54 $X2=11.395 $Y2=2.79
r343 6 61 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=9.485
+ $Y=2.12 $X2=9.63 $Y2=2.455
r344 5 57 600 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=1 $X=8.395
+ $Y=2.12 $X2=8.53 $Y2=2.63
r345 4 53 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=2.32 $X2=5.05 $Y2=2.555
r346 3 47 300 $w=1.7e-07 $l=6.48999e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=2.425
r347 2 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.435
+ $Y=2.32 $X2=2.58 $Y2=2.465
r348 1 39 600 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.32 $X2=0.73 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_197_119# 1 2 3 4 15 17 19 20 23 24 25 26
+ 28 29 32 33 34 36 37 38 40 41 42 44 45 46 48 49 50 51 56 57 58 60 61 63 64 68
c222 48 0 1.91291e-19 $X=6.03 $Y=0.84
c223 45 0 7.90252e-20 $X=5.945 $Y=0.925
c224 26 0 1.01507e-19 $X=1.69 $Y=1.205
c225 17 0 8.61452e-20 $X=1.57 $Y=2.515
c226 15 0 1.46097e-19 $X=1.53 $Y=2.425
r227 66 68 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=2.557
+ $X2=6.67 $Y2=2.557
r228 59 60 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=7.62 $Y=1.015
+ $X2=7.62 $Y2=2.38
r229 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.535 $Y=0.93
+ $X2=7.62 $Y2=1.015
r230 57 58 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.535 $Y=0.93
+ $X2=7.115 $Y2=0.93
r231 54 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.95 $Y=0.845
+ $X2=7.115 $Y2=0.93
r232 54 56 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.95 $Y=0.845
+ $X2=6.95 $Y2=0.81
r233 53 56 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.95 $Y=0.435
+ $X2=6.95 $Y2=0.81
r234 51 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.535 $Y=2.465
+ $X2=7.62 $Y2=2.38
r235 51 68 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=7.535 $Y=2.465
+ $X2=6.67 $Y2=2.465
r236 49 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.785 $Y=0.35
+ $X2=6.95 $Y2=0.435
r237 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.785 $Y=0.35
+ $X2=6.115 $Y2=0.35
r238 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.03 $Y=0.435
+ $X2=6.115 $Y2=0.35
r239 47 48 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.03 $Y=0.435
+ $X2=6.03 $Y2=0.84
r240 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.945 $Y=0.925
+ $X2=6.03 $Y2=0.84
r241 45 46 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.945 $Y=0.925
+ $X2=5.28 $Y2=0.925
r242 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.195 $Y=0.84
+ $X2=5.28 $Y2=0.925
r243 43 44 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.195 $Y=0.425
+ $X2=5.195 $Y2=0.84
r244 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.11 $Y=0.34
+ $X2=5.195 $Y2=0.425
r245 41 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.11 $Y=0.34
+ $X2=4.52 $Y2=0.34
r246 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.52 $Y2=0.34
r247 39 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.435 $Y2=0.66
r248 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.745
+ $X2=4.435 $Y2=0.66
r249 37 38 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=4.35 $Y=0.745
+ $X2=3.535 $Y2=0.745
r250 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.45 $Y=0.66
+ $X2=3.535 $Y2=0.745
r251 35 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.66
r252 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=3.45 $Y2=0.425
r253 33 34 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=2.77 $Y2=0.34
r254 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.685 $Y=0.425
+ $X2=2.77 $Y2=0.34
r255 31 32 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.685 $Y=0.425
+ $X2=2.685 $Y2=1.12
r256 30 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.205
+ $X2=2.07 $Y2=1.205
r257 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.6 $Y=1.205
+ $X2=2.685 $Y2=1.12
r258 29 30 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.6 $Y=1.205
+ $X2=2.155 $Y2=1.205
r259 27 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.29
+ $X2=2.07 $Y2=1.205
r260 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=1.29
+ $X2=2.07 $Y2=1.96
r261 25 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.205
+ $X2=2.07 $Y2=1.205
r262 25 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.985 $Y=1.205
+ $X2=1.69 $Y2=1.205
r263 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=2.045
+ $X2=2.07 $Y2=1.96
r264 23 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.985 $Y=2.045
+ $X2=1.655 $Y2=2.045
r265 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=2.13
+ $X2=1.655 $Y2=2.045
r266 21 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.57 $Y=2.13
+ $X2=1.57 $Y2=2.3
r267 20 26 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=1.587 $Y=1.12
+ $X2=1.69 $Y2=1.205
r268 19 63 4.51862 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=0.955
+ $X2=1.587 $Y2=0.79
r269 19 20 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=0.955
+ $X2=1.587 $Y2=1.12
r270 15 61 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.53 $Y=2.425
+ $X2=1.53 $Y2=2.3
r271 15 17 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.53 $Y=2.425
+ $X2=1.53 $Y2=2.515
r272 4 66 600 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=2.32 $X2=6.505 $Y2=2.515
r273 3 17 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=2.32 $X2=1.57 $Y2=2.515
r274 2 56 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=6.74
+ $Y=0.625 $X2=6.95 $Y2=0.81
r275 1 63 91 $w=1.7e-07 $l=6.3e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.595 $X2=1.525 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%Q_N 1 2 9 15 19 20 23
r29 20 25 4.72801 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=15.545 $Y=1.665
+ $X2=15.545 $Y2=1.78
r30 20 23 5.0075 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=15.545 $Y=1.665
+ $X2=15.545 $Y2=1.55
r31 19 23 16.1832 $w=2.33e-07 $l=3.3e-07 $layer=LI1_cond $X=15.492 $Y=1.22
+ $X2=15.492 $Y2=1.55
r32 15 17 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.5 $Y=1.985
+ $X2=15.5 $Y2=2.815
r33 15 25 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=15.5 $Y=1.985
+ $X2=15.5 $Y2=1.78
r34 7 19 6.73378 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.445 $Y=1.055
+ $X2=15.445 $Y2=1.22
r35 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=15.445 $Y=1.055
+ $X2=15.445 $Y2=0.515
r36 2 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=15.405
+ $Y=1.84 $X2=15.54 $Y2=2.815
r37 2 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=15.405
+ $Y=1.84 $X2=15.54 $Y2=1.985
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.305
+ $Y=0.37 $X2=15.445 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%Q 1 2 9 13 14 20 26
r28 17 20 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=17.55 $Y=1.975
+ $X2=17.55 $Y2=1.985
r29 14 17 0.483283 $w=3.08e-07 $l=1.3e-08 $layer=LI1_cond $X=17.55 $Y=1.962
+ $X2=17.55 $Y2=1.975
r30 14 26 7.61225 $w=3.08e-07 $l=1.42e-07 $layer=LI1_cond $X=17.55 $Y=1.962
+ $X2=17.55 $Y2=1.82
r31 14 23 28.5508 $w=3.08e-07 $l=7.68e-07 $layer=LI1_cond $X=17.55 $Y=2.047
+ $X2=17.55 $Y2=2.815
r32 14 20 2.30489 $w=3.08e-07 $l=6.2e-08 $layer=LI1_cond $X=17.55 $Y=2.047
+ $X2=17.55 $Y2=1.985
r33 13 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=17.62 $Y=1.05
+ $X2=17.62 $Y2=1.82
r34 7 13 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=17.537 $Y=0.883
+ $X2=17.537 $Y2=1.05
r35 7 9 12.6597 $w=3.33e-07 $l=3.68e-07 $layer=LI1_cond $X=17.537 $Y=0.883
+ $X2=17.537 $Y2=0.515
r36 2 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=17.375
+ $Y=1.84 $X2=17.51 $Y2=2.815
r37 2 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=17.375
+ $Y=1.84 $X2=17.51 $Y2=1.985
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.395
+ $Y=0.37 $X2=17.535 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%VGND 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 51 55 59 63 67 69 72 73 75 76 78 79 80 89 96 101 119 123 132 135 138 148 152
r191 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=0 $X2=18
+ $Y2=0
r192 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r193 139 143 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.76 $Y2=0
r194 138 139 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r195 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r196 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r197 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r198 127 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=18 $Y2=0
r199 127 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=17.04 $Y2=0
r200 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r201 124 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.2 $Y=0
+ $X2=17.035 $Y2=0
r202 124 126 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=17.2 $Y=0
+ $X2=17.52 $Y2=0
r203 123 151 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=17.88 $Y=0
+ $X2=18.06 $Y2=0
r204 123 126 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=17.88 $Y=0
+ $X2=17.52 $Y2=0
r205 122 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.04 $Y2=0
r206 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r207 119 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.87 $Y=0
+ $X2=17.035 $Y2=0
r208 119 121 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=16.87 $Y=0
+ $X2=16.56 $Y2=0
r209 118 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.56 $Y2=0
r210 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r211 115 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.6 $Y2=0
r212 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r213 112 115 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=14.64 $Y2=0
r214 112 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r215 111 114 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=14.64 $Y2=0
r216 111 112 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r217 109 111 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=12.24 $Y2=0
r218 107 108 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r219 105 108 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6 $Y=0 $X2=8.88
+ $Y2=0
r220 105 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r221 104 107 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.88
+ $Y2=0
r222 104 105 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6
+ $Y2=0
r223 102 135 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.72 $Y=0
+ $X2=5.585 $Y2=0
r224 102 104 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.72 $Y=0 $X2=6
+ $Y2=0
r225 101 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.055 $Y=0
+ $X2=9.22 $Y2=0
r226 101 107 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.055 $Y=0
+ $X2=8.88 $Y2=0
r227 100 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.52 $Y2=0
r228 100 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r229 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r230 97 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=0
+ $X2=4.055 $Y2=0
r231 97 99 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.56
+ $Y2=0
r232 96 135 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.45 $Y=0
+ $X2=5.585 $Y2=0
r233 96 99 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.45 $Y=0 $X2=4.56
+ $Y2=0
r234 95 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r235 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r236 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r237 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r238 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r239 89 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.93 $Y=0
+ $X2=4.055 $Y2=0
r240 89 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.6
+ $Y2=0
r241 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r242 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r243 85 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r244 85 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r245 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r246 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r247 82 129 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0
+ $X2=0.235 $Y2=0
r248 82 84 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r249 80 139 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=9.36 $Y2=0
r250 80 108 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=8.88 $Y2=0
r251 78 117 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=15.78 $Y=0
+ $X2=15.6 $Y2=0
r252 78 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.78 $Y=0
+ $X2=15.945 $Y2=0
r253 77 121 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=16.11 $Y=0
+ $X2=16.56 $Y2=0
r254 77 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.11 $Y=0
+ $X2=15.945 $Y2=0
r255 75 114 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=14.825 $Y=0
+ $X2=14.64 $Y2=0
r256 75 76 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=14.825 $Y=0
+ $X2=14.967 $Y2=0
r257 74 117 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=15.11 $Y=0
+ $X2=15.6 $Y2=0
r258 74 76 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=15.11 $Y=0
+ $X2=14.967 $Y2=0
r259 72 87 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.16
+ $Y2=0
r260 72 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.305
+ $Y2=0
r261 71 91 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.64
+ $Y2=0
r262 71 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.305
+ $Y2=0
r263 67 151 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=18.005 $Y=0.085
+ $X2=18.06 $Y2=0
r264 67 69 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=18.005 $Y=0.085
+ $X2=18.005 $Y2=0.515
r265 63 65 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.035 $Y=0.515
+ $X2=17.035 $Y2=0.885
r266 61 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.035 $Y=0.085
+ $X2=17.035 $Y2=0
r267 61 63 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=17.035 $Y=0.085
+ $X2=17.035 $Y2=0.515
r268 57 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.945 $Y=0.085
+ $X2=15.945 $Y2=0
r269 57 59 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.945 $Y=0.085
+ $X2=15.945 $Y2=0.515
r270 53 76 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=14.967 $Y=0.085
+ $X2=14.967 $Y2=0
r271 53 55 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=14.967 $Y=0.085
+ $X2=14.967 $Y2=0.515
r272 52 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.385 $Y=0
+ $X2=9.22 $Y2=0
r273 51 145 10.6025 $w=3.73e-07 $l=3.45e-07 $layer=LI1_cond $X=11.867 $Y=0
+ $X2=11.867 $Y2=0.345
r274 51 109 5.38787 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=11.867 $Y=0
+ $X2=12.055 $Y2=0
r275 51 143 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r276 51 52 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=11.68 $Y=0
+ $X2=9.385 $Y2=0
r277 47 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0
r278 47 49 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=9.22 $Y=0.085
+ $X2=9.22 $Y2=0.77
r279 43 135 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=0.085
+ $X2=5.585 $Y2=0
r280 43 45 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.585 $Y=0.085
+ $X2=5.585 $Y2=0.505
r281 39 132 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0
r282 39 41 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0.325
r283 35 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0
r284 35 37 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0.76
r285 31 129 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.235 $Y2=0
r286 31 33 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.305 $Y2=0.765
r287 10 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.825
+ $Y=0.37 $X2=17.965 $Y2=0.515
r288 9 65 182 $w=1.7e-07 $l=5.21368e-07 $layer=licon1_NDIFF $count=1 $X=16.795
+ $Y=0.47 $X2=17.035 $Y2=0.885
r289 9 63 182 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_NDIFF $count=1 $X=16.795
+ $Y=0.47 $X2=17.035 $Y2=0.515
r290 8 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.735
+ $Y=0.37 $X2=15.875 $Y2=0.515
r291 7 55 91 $w=1.7e-07 $l=9.12414e-07 $layer=licon1_NDIFF $count=2 $X=14.275
+ $Y=0.9 $X2=15.015 $Y2=0.515
r292 6 145 182 $w=1.7e-07 $l=2.70555e-07 $layer=licon1_NDIFF $count=1 $X=11.625
+ $Y=0.41 $X2=11.865 $Y2=0.345
r293 5 49 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=9.01
+ $Y=0.625 $X2=9.22 $Y2=0.77
r294 4 45 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.36 $X2=5.545 $Y2=0.505
r295 3 41 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.49 $X2=4.095 $Y2=0.325
r296 2 37 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.205
+ $Y=0.595 $X2=2.345 $Y2=0.76
r297 1 33 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_1473_73# 1 2 7 10 11 19
c40 19 0 8.54043e-20 $X=8.665 $Y=0.77
r41 16 19 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=0.77
+ $X2=8.665 $Y2=0.77
r42 11 14 4.33861 $w=4.23e-07 $l=1.6e-07 $layer=LI1_cond $X=7.557 $Y=0.35
+ $X2=7.557 $Y2=0.51
r43 10 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=0.605
+ $X2=8.535 $Y2=0.77
r44 9 10 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.535 $Y=0.435
+ $X2=8.535 $Y2=0.605
r45 8 11 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=7.77 $Y=0.35
+ $X2=7.557 $Y2=0.35
r46 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.45 $Y=0.35
+ $X2=8.535 $Y2=0.435
r47 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.45 $Y=0.35 $X2=7.77
+ $Y2=0.35
r48 2 19 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=8.405
+ $Y=0.625 $X2=8.665 $Y2=0.77
r49 1 14 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.365 $X2=7.555 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_MS__SDFBBN_2%A_2452_74# 1 2 9 15 16
c24 16 0 6.88126e-20 $X=13.265 $Y=0.375
r25 15 16 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=13.43 $Y=0.375
+ $X2=13.265 $Y2=0.375
r26 9 12 4.80185 $w=4.18e-07 $l=1.75e-07 $layer=LI1_cond $X=12.445 $Y=0.34
+ $X2=12.445 $Y2=0.515
r27 8 9 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=12.655 $Y=0.34
+ $X2=12.445 $Y2=0.34
r28 8 16 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=12.655 $Y=0.34
+ $X2=13.265 $Y2=0.34
r29 2 15 182 $w=1.7e-07 $l=2.39165e-07 $layer=licon1_NDIFF $count=1 $X=13.21
+ $Y=0.37 $X2=13.43 $Y2=0.41
r30 1 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=12.26
+ $Y=0.37 $X2=12.445 $Y2=0.515
.ends


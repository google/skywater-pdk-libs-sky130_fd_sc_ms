# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a2bb2oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__a2bb2oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.285000 0.435000 0.670000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.570000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.320000 3.735000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.716800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.080000 0.390000 2.250000 0.980000 ;
        RECT 2.080000 0.980000 3.795000 1.150000 ;
        RECT 2.525000 1.150000 3.235000 1.410000 ;
        RECT 2.525000 1.410000 2.780000 2.735000 ;
        RECT 3.465000 0.770000 3.795000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.580000  1.940000 0.910000 3.245000 ;
      RECT 0.605000  0.085000 0.855000 1.170000 ;
      RECT 1.035000  0.490000 1.330000 1.110000 ;
      RECT 1.035000  1.110000 1.910000 1.280000 ;
      RECT 1.420000  1.950000 1.910000 2.980000 ;
      RECT 1.570000  0.085000 1.900000 0.940000 ;
      RECT 1.740000  1.280000 1.910000 1.320000 ;
      RECT 1.740000  1.320000 2.205000 1.650000 ;
      RECT 1.740000  1.650000 1.910000 1.950000 ;
      RECT 2.080000  1.820000 2.330000 2.905000 ;
      RECT 2.080000  2.905000 3.230000 3.075000 ;
      RECT 2.430000  0.085000 2.760000 0.810000 ;
      RECT 2.980000  1.820000 3.230000 1.950000 ;
      RECT 2.980000  1.950000 5.110000 2.120000 ;
      RECT 2.980000  2.120000 3.230000 2.905000 ;
      RECT 3.035000  0.350000 4.145000 0.600000 ;
      RECT 3.430000  2.290000 3.760000 3.245000 ;
      RECT 3.960000  2.120000 4.130000 2.980000 ;
      RECT 3.975000  0.600000 4.145000 1.010000 ;
      RECT 3.975000  1.010000 5.085000 1.180000 ;
      RECT 4.325000  0.085000 4.575000 0.840000 ;
      RECT 4.330000  2.290000 4.660000 3.245000 ;
      RECT 4.755000  0.350000 5.085000 1.010000 ;
      RECT 4.860000  1.820000 5.110000 1.950000 ;
      RECT 4.860000  2.120000 5.110000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_ms__a2bb2oi_2

* File: sky130_fd_sc_ms__or3b_4.spice
* Created: Fri Aug 28 18:08:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or3b_4.pex.spice"
.subckt sky130_fd_sc_ms__or3b_4  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_C_N_M1015_g N_A_27_392#_M1015_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.66075 AS=0.1824 PD=3.58 PS=1.85 NRD=183.264 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_A_27_392#_M1009_g N_A_412_392#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2072 PD=1.09 PS=2.04 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003 A=0.111 P=1.78 MULT=1
MM1006 N_A_412_392#_M1006_d N_B_M1006_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_A_412_392#_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.1036 PD=1.1 PS=1.02 NRD=12.156 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_412_392#_M1001_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.1332 PD=1.045 PS=1.1 NRD=4.044 NRS=0.804 M=1 R=4.93333
+ SA=75001.6 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1001_d N_A_412_392#_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.1221 PD=1.045 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1007_d N_A_412_392#_M1007_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75002.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_X_M1007_d N_A_412_392#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_C_N_M1005_g N_A_27_392#_M1005_s VPB PSHORT L=0.18 W=1
+ AD=0.165 AS=0.275 PD=1.33 PS=2.55 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1005_d N_A_M1000_g N_A_220_392#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=10.8153 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1010 N_A_220_392#_M1000_s N_B_M1010_g N_A_310_392#_M1010_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.165 PD=1.27 PS=1.33 NRD=0 NRS=10.8153 M=1 R=5.55556
+ SA=90001.1 SB=90004 A=0.18 P=2.36 MULT=1
MM1004 N_A_412_392#_M1004_d N_A_27_392#_M1004_g N_A_310_392#_M1010_s VPB PSHORT
+ L=0.18 W=1 AD=0.1475 AS=0.165 PD=1.295 PS=1.33 NRD=0.9653 NRS=0 M=1 R=5.55556
+ SA=90001.7 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1008 N_A_412_392#_M1004_d N_A_27_392#_M1008_g N_A_310_392#_M1008_s VPB PSHORT
+ L=0.18 W=1 AD=0.1475 AS=0.135 PD=1.295 PS=1.27 NRD=1.9503 NRS=0 M=1 R=5.55556
+ SA=90002.1 SB=90003 A=0.18 P=2.36 MULT=1
MM1013 N_A_220_392#_M1013_d N_B_M1013_g N_A_310_392#_M1008_s VPB PSHORT L=0.18
+ W=1 AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90002.6 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_A_220_392#_M1013_d VPB PSHORT L=0.18 W=1
+ AD=0.169811 AS=0.165 PD=1.36792 PS=1.33 NRD=6.8753 NRS=0.9653 M=1 R=5.55556
+ SA=90003.1 SB=90002 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1011_d N_A_412_392#_M1003_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.190189 AS=0.1512 PD=1.53208 PS=1.39 NRD=2.6201 NRS=0 M=1 R=6.22222
+ SA=90003.2 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_412_392#_M1014_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1014_d N_A_412_392#_M1016_g N_X_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1017_d N_A_412_392#_M1017_g N_X_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX19_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__or3b_4.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__fahcin_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__fahcin_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.350000 0.835000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.807000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.875000 1.180000 5.205000 1.585000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.588600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705000 1.155000 9.035000 1.485000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  1.934600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 0.440000 8.035000 0.985000 ;
        RECT 6.640000 0.985000 7.070000 1.310000 ;
        RECT 6.820000 2.335000 7.615000 2.665000 ;
        RECT 6.900000 1.310000 7.070000 2.335000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515000 0.440000 12.845000 0.840000 ;
        RECT 12.595000 0.840000 12.845000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.120000  0.350000  0.450000 1.010000 ;
      RECT  0.120000  1.010000  1.290000 1.180000 ;
      RECT  0.120000  1.180000  0.375000 2.980000 ;
      RECT  0.575000  1.950000  0.825000 3.245000 ;
      RECT  0.620000  0.085000  0.950000 0.840000 ;
      RECT  1.005000  1.180000  1.290000 1.300000 ;
      RECT  1.005000  1.300000  1.445000 1.630000 ;
      RECT  1.005000  1.630000  1.175000 2.905000 ;
      RECT  1.005000  2.905000  3.935000 3.075000 ;
      RECT  1.120000  0.255000  2.835000 0.425000 ;
      RECT  1.120000  0.425000  1.290000 1.010000 ;
      RECT  1.345000  1.820000  1.835000 2.565000 ;
      RECT  1.345000  2.565000  2.980000 2.735000 ;
      RECT  1.475000  0.615000  1.835000 1.020000 ;
      RECT  1.615000  1.020000  1.835000 1.820000 ;
      RECT  2.045000  1.890000  2.415000 2.070000 ;
      RECT  2.045000  2.070000  2.485000 2.395000 ;
      RECT  2.165000  0.615000  2.415000 1.890000 ;
      RECT  2.585000  0.425000  2.835000 0.750000 ;
      RECT  2.655000  2.045000  2.980000 2.565000 ;
      RECT  2.810000  0.920000  3.175000 1.090000 ;
      RECT  2.810000  1.090000  2.980000 2.045000 ;
      RECT  3.005000  0.255000  3.945000 0.425000 ;
      RECT  3.005000  0.425000  3.175000 0.920000 ;
      RECT  3.185000  1.875000  3.515000 1.880000 ;
      RECT  3.185000  1.880000  4.275000 2.050000 ;
      RECT  3.185000  2.050000  3.515000 2.735000 ;
      RECT  3.345000  0.595000  3.515000 1.875000 ;
      RECT  3.685000  1.380000  4.285000 1.550000 ;
      RECT  3.685000  1.550000  3.990000 1.710000 ;
      RECT  3.685000  2.250000  3.935000 2.905000 ;
      RECT  3.695000  0.425000  3.945000 1.125000 ;
      RECT  4.105000  2.050000  4.275000 2.905000 ;
      RECT  4.105000  2.905000  5.045000 3.075000 ;
      RECT  4.115000  0.255000  5.295000 0.425000 ;
      RECT  4.115000  0.425000  4.285000 1.380000 ;
      RECT  4.445000  1.875000  4.705000 2.735000 ;
      RECT  4.455000  0.670000  4.705000 1.875000 ;
      RECT  4.875000  2.390000  6.650000 2.560000 ;
      RECT  4.875000  2.560000  5.045000 2.905000 ;
      RECT  4.955000  1.820000  5.800000 1.990000 ;
      RECT  4.955000  1.990000  5.285000 2.220000 ;
      RECT  4.965000  0.425000  5.295000 0.840000 ;
      RECT  4.965000  0.840000  5.800000 1.010000 ;
      RECT  5.405000  2.730000  5.765000 3.245000 ;
      RECT  5.465000  0.085000  5.970000 0.635000 ;
      RECT  5.630000  1.010000  5.800000 1.255000 ;
      RECT  5.630000  1.255000  5.970000 1.585000 ;
      RECT  5.630000  1.585000  5.800000 1.820000 ;
      RECT  5.970000  1.820000  6.310000 2.220000 ;
      RECT  6.140000  0.385000  6.470000 1.065000 ;
      RECT  6.140000  1.065000  6.310000 1.820000 ;
      RECT  6.150000  2.560000  6.650000 2.905000 ;
      RECT  6.150000  2.905000  8.715000 3.075000 ;
      RECT  6.480000  1.510000  6.730000 1.840000 ;
      RECT  6.480000  1.840000  6.650000 2.390000 ;
      RECT  7.240000  1.170000  7.555000 2.150000 ;
      RECT  7.745000  1.155000  8.035000 1.485000 ;
      RECT  7.785000  1.485000  7.955000 2.905000 ;
      RECT  8.125000  1.820000  8.375000 2.735000 ;
      RECT  8.205000  0.385000  8.535000 1.065000 ;
      RECT  8.205000  1.065000  8.375000 1.820000 ;
      RECT  8.545000  1.655000  9.385000 1.825000 ;
      RECT  8.545000  1.825000  8.715000 2.905000 ;
      RECT  8.705000  0.085000  9.045000 0.985000 ;
      RECT  8.885000  1.995000  9.055000 3.245000 ;
      RECT  9.215000  0.255000 10.575000 0.570000 ;
      RECT  9.215000  0.570000  9.385000 1.655000 ;
      RECT  9.255000  1.995000  9.725000 2.905000 ;
      RECT  9.255000  2.905000 11.975000 3.075000 ;
      RECT  9.555000  0.740000  9.885000 1.340000 ;
      RECT  9.555000  1.340000  9.725000 1.995000 ;
      RECT  9.895000  1.900000 10.065000 2.400000 ;
      RECT  9.895000  2.400000 11.635000 2.570000 ;
      RECT  9.895000  2.570000 10.065000 2.735000 ;
      RECT 10.070000  0.740000 10.915000 1.260000 ;
      RECT 10.265000  1.260000 10.515000 2.230000 ;
      RECT 10.685000  1.430000 11.015000 2.150000 ;
      RECT 10.745000  0.320000 11.755000 0.490000 ;
      RECT 10.745000  0.490000 10.915000 0.740000 ;
      RECT 10.800000  2.740000 11.155000 2.905000 ;
      RECT 11.085000  0.660000 11.415000 1.220000 ;
      RECT 11.085000  1.220000 11.365000 1.250000 ;
      RECT 11.195000  1.250000 11.365000 1.850000 ;
      RECT 11.195000  1.850000 11.635000 2.400000 ;
      RECT 11.385000  2.570000 11.635000 2.735000 ;
      RECT 11.535000  1.350000 11.975000 1.680000 ;
      RECT 11.585000  0.490000 11.755000 1.010000 ;
      RECT 11.585000  1.010000 12.425000 1.180000 ;
      RECT 11.805000  1.680000 11.975000 2.905000 ;
      RECT 11.925000  0.085000 12.345000 0.810000 ;
      RECT 12.145000  1.180000 12.425000 1.680000 ;
      RECT 12.145000  1.850000 12.395000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.950000  2.245000 2.120000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  1.950000  4.645000 2.120000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.950000  7.525000 2.120000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
    LAYER met1 ;
      RECT  2.015000 1.920000  2.305000 1.965000 ;
      RECT  2.015000 1.965000 10.945000 2.105000 ;
      RECT  2.015000 2.105000  2.305000 2.150000 ;
      RECT  4.415000 1.920000  4.705000 1.965000 ;
      RECT  4.415000 2.105000  4.705000 2.150000 ;
      RECT  7.295000 1.920000  7.585000 1.965000 ;
      RECT  7.295000 2.105000  7.585000 2.150000 ;
      RECT 10.655000 1.920000 10.945000 1.965000 ;
      RECT 10.655000 2.105000 10.945000 2.150000 ;
  END
END sky130_fd_sc_ms__fahcin_1

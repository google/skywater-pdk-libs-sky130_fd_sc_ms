* File: sky130_fd_sc_ms__nand2_1.pxi.spice
* Created: Fri Aug 28 17:41:38 2020
* 
x_PM_SKY130_FD_SC_MS__NAND2_1%B N_B_M1001_g N_B_c_28_n N_B_M1003_g B N_B_c_30_n
+ PM_SKY130_FD_SC_MS__NAND2_1%B
x_PM_SKY130_FD_SC_MS__NAND2_1%A N_A_c_53_n N_A_M1000_g N_A_M1002_g A N_A_c_56_n
+ PM_SKY130_FD_SC_MS__NAND2_1%A
x_PM_SKY130_FD_SC_MS__NAND2_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_c_81_n
+ N_VPWR_c_82_n N_VPWR_c_83_n N_VPWR_c_84_n VPWR N_VPWR_c_85_n N_VPWR_c_80_n
+ PM_SKY130_FD_SC_MS__NAND2_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND2_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_103_n N_Y_c_104_n
+ Y Y Y Y Y Y N_Y_c_106_n PM_SKY130_FD_SC_MS__NAND2_1%Y
x_PM_SKY130_FD_SC_MS__NAND2_1%VGND N_VGND_M1003_s N_VGND_c_134_n N_VGND_c_135_n
+ VGND N_VGND_c_136_n N_VGND_c_137_n PM_SKY130_FD_SC_MS__NAND2_1%VGND
cc_1 VNB N_B_M1001_g 0.00933282f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_B_c_28_n 0.0207038f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_3 VNB B 0.00878284f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B_c_30_n 0.058145f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.385
cc_5 VNB N_A_c_53_n 0.0221784f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.55
cc_6 VNB N_A_M1002_g 0.00933282f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_7 VNB A 0.0096067f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_c_56_n 0.059425f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_9 VNB N_VPWR_c_80_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_Y_c_103_n 0.0070579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_104_n 0.0213168f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_12 VNB Y 0.00714178f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_Y_c_106_n 6.31494e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_134_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_135_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_16 VNB N_VGND_c_136_n 0.0306085f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_17 VNB N_VGND_c_137_n 0.119298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VPB N_B_M1001_g 0.0295103f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_19 VPB N_A_M1002_g 0.0295103f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_20 VPB N_VPWR_c_81_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_21 VPB N_VPWR_c_82_n 0.0552927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_83_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_23 VPB N_VPWR_c_84_n 0.0552927f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.385
cc_24 VPB N_VPWR_c_85_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_80_n 0.0473405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_26 VPB Y 0.00648934f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_27 N_B_c_28_n N_A_c_53_n 0.0329441f $X=0.51 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_28 N_B_M1001_g N_A_M1002_g 0.0184047f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_29 B N_A_c_56_n 2.30773e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_30 N_B_c_30_n N_A_c_56_n 0.0329441f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_31 N_B_M1001_g N_VPWR_c_82_n 0.0201908f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_32 B N_VPWR_c_82_n 0.0196739f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_33 N_B_c_30_n N_VPWR_c_82_n 0.00223706f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_34 N_B_M1001_g N_VPWR_c_84_n 6.38263e-19 $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_35 N_B_M1001_g N_VPWR_c_85_n 0.00460063f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_36 N_B_M1001_g N_VPWR_c_80_n 0.00908665f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_37 N_B_c_28_n N_Y_c_103_n 0.00129102f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_38 N_B_c_28_n N_Y_c_104_n 0.00138696f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_39 N_B_c_28_n Y 0.00535815f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_40 B Y 0.0285816f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 N_B_c_30_n Y 0.00535815f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_42 N_B_c_28_n N_Y_c_106_n 0.00382427f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_43 N_B_c_28_n N_VGND_c_135_n 0.0166171f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_44 B N_VGND_c_135_n 0.0241219f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_45 N_B_c_30_n N_VGND_c_135_n 0.00199226f $X=0.51 $Y=1.385 $X2=0 $Y2=0
cc_46 N_B_c_28_n N_VGND_c_136_n 0.00383152f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_47 N_B_c_28_n N_VGND_c_137_n 0.0075725f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_48 N_A_M1002_g N_VPWR_c_82_n 6.38263e-19 $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_VPWR_c_84_n 0.0201908f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_50 A N_VPWR_c_84_n 0.0196739f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A_c_56_n N_VPWR_c_84_n 0.00223706f $X=1.17 $Y=1.385 $X2=0 $Y2=0
cc_52 N_A_M1002_g N_VPWR_c_85_n 0.00460063f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_53 N_A_M1002_g N_VPWR_c_80_n 0.00908665f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_54 N_A_c_53_n N_Y_c_103_n 0.0126998f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_55 A N_Y_c_103_n 0.0207374f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_c_56_n N_Y_c_103_n 0.00167247f $X=1.17 $Y=1.385 $X2=0 $Y2=0
cc_57 N_A_c_53_n N_Y_c_104_n 0.00922372f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A_c_53_n Y 6.89533e-19 $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_59 N_A_M1002_g Y 0.00767761f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_60 A Y 0.0271114f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A_c_56_n Y 0.00769026f $X=1.17 $Y=1.385 $X2=0 $Y2=0
cc_62 N_A_c_53_n N_Y_c_106_n 0.00776809f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A_c_53_n N_VGND_c_135_n 0.00208984f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A_c_53_n N_VGND_c_136_n 0.00434272f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_65 N_A_c_53_n N_VGND_c_137_n 0.00451209f $X=0.9 $Y=1.22 $X2=0 $Y2=0
cc_66 N_VPWR_c_82_n Y 0.0450228f $X=0.27 $Y=1.985 $X2=0 $Y2=0
cc_67 N_VPWR_c_84_n Y 0.0450228f $X=1.17 $Y=1.985 $X2=0 $Y2=0
cc_68 N_VPWR_c_85_n Y 0.0101736f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_69 N_VPWR_c_80_n Y 0.0084208f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_70 N_Y_c_103_n N_VGND_c_135_n 0.0119089f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_71 N_Y_c_104_n N_VGND_c_135_n 0.0155235f $X=1.115 $Y=0.515 $X2=0 $Y2=0
cc_72 N_Y_c_104_n N_VGND_c_136_n 0.0142249f $X=1.115 $Y=0.515 $X2=0 $Y2=0
cc_73 N_Y_c_103_n N_VGND_c_137_n 0.00901755f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_74 N_Y_c_104_n N_VGND_c_137_n 0.011867f $X=1.115 $Y=0.515 $X2=0 $Y2=0
cc_75 N_Y_c_103_n A_117_74# 0.00390405f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_76 N_Y_c_106_n A_117_74# 0.00140851f $X=0.72 $Y=1.18 $X2=-0.19 $Y2=-0.245

* File: sky130_fd_sc_ms__o211a_4.pxi.spice
* Created: Wed Sep  2 12:20:26 2020
* 
x_PM_SKY130_FD_SC_MS__O211A_4%A_91_48# N_A_91_48#_M1015_s N_A_91_48#_M1010_s
+ N_A_91_48#_M1007_s N_A_91_48#_M1001_s N_A_91_48#_M1002_g N_A_91_48#_M1004_g
+ N_A_91_48#_M1013_g N_A_91_48#_M1006_g N_A_91_48#_M1016_g N_A_91_48#_M1008_g
+ N_A_91_48#_M1017_g N_A_91_48#_M1009_g N_A_91_48#_c_140_n N_A_91_48#_c_141_n
+ N_A_91_48#_c_151_n N_A_91_48#_c_209_p N_A_91_48#_c_152_n N_A_91_48#_c_142_n
+ N_A_91_48#_c_143_n N_A_91_48#_c_154_n N_A_91_48#_c_155_n N_A_91_48#_c_144_n
+ N_A_91_48#_c_156_n N_A_91_48#_c_157_n N_A_91_48#_c_145_n
+ PM_SKY130_FD_SC_MS__O211A_4%A_91_48#
x_PM_SKY130_FD_SC_MS__O211A_4%C1 N_C1_c_309_n N_C1_M1000_g N_C1_M1015_g
+ N_C1_c_310_n N_C1_M1007_g N_C1_M1020_g C1 N_C1_c_308_n
+ PM_SKY130_FD_SC_MS__O211A_4%C1
x_PM_SKY130_FD_SC_MS__O211A_4%B1 N_B1_c_357_n N_B1_c_358_n N_B1_c_359_n
+ N_B1_M1010_g N_B1_c_360_n N_B1_M1014_g N_B1_M1023_g N_B1_M1019_g N_B1_c_363_n
+ B1 N_B1_c_364_n PM_SKY130_FD_SC_MS__O211A_4%B1
x_PM_SKY130_FD_SC_MS__O211A_4%A2 N_A2_M1001_g N_A2_M1011_g N_A2_M1003_g
+ N_A2_M1021_g A2 A2 N_A2_c_440_n N_A2_c_441_n PM_SKY130_FD_SC_MS__O211A_4%A2
x_PM_SKY130_FD_SC_MS__O211A_4%A1 N_A1_c_486_n N_A1_M1005_g N_A1_M1012_g
+ N_A1_c_489_n N_A1_c_490_n N_A1_M1018_g N_A1_M1022_g A1 N_A1_c_493_n
+ PM_SKY130_FD_SC_MS__O211A_4%A1
x_PM_SKY130_FD_SC_MS__O211A_4%VPWR N_VPWR_M1004_s N_VPWR_M1006_s N_VPWR_M1009_s
+ N_VPWR_M1000_d N_VPWR_M1023_d N_VPWR_M1018_d N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n
+ N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n VPWR
+ N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n
+ N_VPWR_c_566_n N_VPWR_c_549_n PM_SKY130_FD_SC_MS__O211A_4%VPWR
x_PM_SKY130_FD_SC_MS__O211A_4%X N_X_M1002_s N_X_M1016_s N_X_M1004_d N_X_M1008_d
+ N_X_c_643_n N_X_c_644_n N_X_c_650_n N_X_c_651_n N_X_c_645_n N_X_c_652_n
+ N_X_c_646_n N_X_c_653_n N_X_c_647_n N_X_c_654_n N_X_c_648_n N_X_c_655_n X X
+ PM_SKY130_FD_SC_MS__O211A_4%X
x_PM_SKY130_FD_SC_MS__O211A_4%A_971_391# N_A_971_391#_M1005_s
+ N_A_971_391#_M1003_d N_A_971_391#_c_725_n N_A_971_391#_c_721_n
+ N_A_971_391#_c_722_n N_A_971_391#_c_723_n
+ PM_SKY130_FD_SC_MS__O211A_4%A_971_391#
x_PM_SKY130_FD_SC_MS__O211A_4%VGND N_VGND_M1002_d N_VGND_M1013_d N_VGND_M1017_d
+ N_VGND_M1012_d N_VGND_M1021_s N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n
+ N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n VGND N_VGND_c_753_n
+ N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n
+ N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ PM_SKY130_FD_SC_MS__O211A_4%VGND
x_PM_SKY130_FD_SC_MS__O211A_4%A_510_125# N_A_510_125#_M1014_d
+ N_A_510_125#_M1019_d N_A_510_125#_M1011_d N_A_510_125#_M1022_s
+ N_A_510_125#_c_835_n N_A_510_125#_c_836_n N_A_510_125#_c_837_n
+ N_A_510_125#_c_838_n N_A_510_125#_c_839_n N_A_510_125#_c_840_n
+ N_A_510_125#_c_841_n N_A_510_125#_c_842_n N_A_510_125#_c_843_n
+ N_A_510_125#_c_844_n PM_SKY130_FD_SC_MS__O211A_4%A_510_125#
x_PM_SKY130_FD_SC_MS__O211A_4%A_597_125# N_A_597_125#_M1014_s
+ N_A_597_125#_M1020_d N_A_597_125#_c_907_n N_A_597_125#_c_908_n
+ N_A_597_125#_c_909_n N_A_597_125#_c_910_n
+ PM_SKY130_FD_SC_MS__O211A_4%A_597_125#
cc_1 VNB N_A_91_48#_M1002_g 0.0225008f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_2 VNB N_A_91_48#_M1004_g 0.00168805f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_3 VNB N_A_91_48#_M1013_g 0.0212087f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_4 VNB N_A_91_48#_M1006_g 0.0016562f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_5 VNB N_A_91_48#_M1016_g 0.0217869f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.74
cc_6 VNB N_A_91_48#_M1008_g 0.0016556f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.4
cc_7 VNB N_A_91_48#_M1017_g 0.0216843f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.74
cc_8 VNB N_A_91_48#_M1009_g 0.00154244f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=2.4
cc_9 VNB N_A_91_48#_c_140_n 0.00579892f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.465
cc_10 VNB N_A_91_48#_c_141_n 4.52924e-19 $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.95
cc_11 VNB N_A_91_48#_c_142_n 0.00167683f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.195
cc_12 VNB N_A_91_48#_c_143_n 0.00329567f $X=-0.19 $Y=-0.245 $X2=4.035 $Y2=1.95
cc_13 VNB N_A_91_48#_c_144_n 0.00248665f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.105
cc_14 VNB N_A_91_48#_c_145_n 0.0916378f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=1.465
cc_15 VNB N_C1_M1015_g 0.0187808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_M1020_g 0.018993f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_17 VNB C1 9.25683e-19 $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_18 VNB N_C1_c_308_n 0.024686f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_19 VNB N_B1_c_357_n 0.0589691f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.955
cc_20 VNB N_B1_c_358_n 0.127671f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.955
cc_21 VNB N_B1_c_359_n 0.0123922f $X=-0.19 $Y=-0.245 $X2=5.305 $Y2=1.955
cc_22 VNB N_B1_c_360_n 0.0148688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_M1023_g 0.00923002f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_24 VNB N_B1_M1019_g 0.0280602f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_25 VNB N_B1_c_363_n 0.0146184f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.3
cc_26 VNB N_B1_c_364_n 0.0418929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_M1011_g 0.0192298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_M1021_g 0.0195968f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_29 VNB N_A2_c_440_n 0.00612267f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.63
cc_30 VNB N_A2_c_441_n 0.0262499f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_31 VNB N_A1_c_486_n 0.00620327f $X=-0.19 $Y=-0.245 $X2=3.415 $Y2=0.625
cc_32 VNB N_A1_M1005_g 0.0141775f $X=-0.19 $Y=-0.245 $X2=3.82 $Y2=1.955
cc_33 VNB N_A1_M1012_g 0.0266069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_c_489_n 0.102837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A1_c_490_n 0.00990222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A1_M1022_g 0.0458509f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_37 VNB A1 0.0115553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_493_n 0.0202529f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_39 VNB N_VPWR_c_549_n 0.283096f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=1.465
cc_40 VNB N_X_c_643_n 0.00150518f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_41 VNB N_X_c_644_n 0.00852127f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_42 VNB N_X_c_645_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_43 VNB N_X_c_646_n 0.00509139f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_44 VNB N_X_c_647_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.63
cc_45 VNB N_X_c_648_n 0.00184578f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=2.4
cc_46 VNB X 0.0268249f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.465
cc_47 VNB N_VGND_c_747_n 0.0117944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_748_n 0.0271311f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_49 VNB N_VGND_c_749_n 0.00495983f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_50 VNB N_VGND_c_750_n 0.0136768f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_51 VNB N_VGND_c_751_n 0.00381151f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.74
cc_52 VNB N_VGND_c_752_n 0.0081779f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.4
cc_53 VNB N_VGND_c_753_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.74
cc_54 VNB N_VGND_c_754_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=2.4
cc_55 VNB N_VGND_c_755_n 0.0602851f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.465
cc_56 VNB N_VGND_c_756_n 0.0157641f $X=-0.19 $Y=-0.245 $X2=2.285 $Y2=2.035
cc_57 VNB N_VGND_c_757_n 0.0191172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_758_n 0.351893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_759_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_760_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.105
cc_61 VNB N_VGND_c_761_n 0.00459433f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.195
cc_62 VNB N_VGND_c_762_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.955 $Y2=2.115
cc_63 VNB N_A_510_125#_c_835_n 0.0136664f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_64 VNB N_A_510_125#_c_836_n 0.0345039f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.63
cc_65 VNB N_A_510_125#_c_837_n 0.0029022f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_66 VNB N_A_510_125#_c_838_n 0.00395785f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_67 VNB N_A_510_125#_c_839_n 0.0042325f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_68 VNB N_A_510_125#_c_840_n 0.00458517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_510_125#_c_841_n 0.00252813f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_70 VNB N_A_510_125#_c_842_n 0.0152112f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.3
cc_71 VNB N_A_510_125#_c_843_n 0.0230853f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.63
cc_72 VNB N_A_510_125#_c_844_n 0.00182475f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=2.4
cc_73 VNB N_A_597_125#_c_907_n 0.00261948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_597_125#_c_908_n 0.00225846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_597_125#_c_909_n 0.0012438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_597_125#_c_910_n 0.00204411f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.3
cc_77 VPB N_A_91_48#_M1004_g 0.0240466f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_78 VPB N_A_91_48#_M1006_g 0.0232284f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_79 VPB N_A_91_48#_M1008_g 0.0232255f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=2.4
cc_80 VPB N_A_91_48#_M1009_g 0.0236404f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=2.4
cc_81 VPB N_A_91_48#_c_141_n 0.00314695f $X=-0.19 $Y=1.66 $X2=2.2 $Y2=1.95
cc_82 VPB N_A_91_48#_c_151_n 0.00229488f $X=-0.19 $Y=1.66 $X2=2.775 $Y2=2.035
cc_83 VPB N_A_91_48#_c_152_n 0.00542769f $X=-0.19 $Y=1.66 $X2=3.79 $Y2=2.035
cc_84 VPB N_A_91_48#_c_143_n 0.00227396f $X=-0.19 $Y=1.66 $X2=4.035 $Y2=1.95
cc_85 VPB N_A_91_48#_c_154_n 0.0106045f $X=-0.19 $Y=1.66 $X2=5.325 $Y2=2.035
cc_86 VPB N_A_91_48#_c_155_n 0.0082706f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=2.115
cc_87 VPB N_A_91_48#_c_156_n 0.00483655f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=2.115
cc_88 VPB N_A_91_48#_c_157_n 0.00236205f $X=-0.19 $Y=1.66 $X2=5.49 $Y2=2.115
cc_89 VPB N_C1_c_309_n 0.0169194f $X=-0.19 $Y=1.66 $X2=3.415 $Y2=0.625
cc_90 VPB N_C1_c_310_n 0.0169216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_C1_c_308_n 0.0383216f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_92 VPB N_B1_M1010_g 0.0253151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_B1_M1023_g 0.0290166f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_94 VPB B1 0.00163765f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_95 VPB N_B1_c_364_n 0.0189329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A2_M1001_g 0.0220393f $X=-0.19 $Y=1.66 $X2=3.82 $Y2=1.955
cc_97 VPB N_A2_M1003_g 0.0221158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A2_c_440_n 0.00407223f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.63
cc_99 VPB N_A2_c_441_n 0.0168855f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_100 VPB N_A1_M1005_g 0.0310594f $X=-0.19 $Y=1.66 $X2=3.82 $Y2=1.955
cc_101 VPB N_A1_M1018_g 0.0278614f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.3
cc_102 VPB A1 0.00733815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A1_c_493_n 0.0133096f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_104 VPB N_VPWR_c_550_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_105 VPB N_VPWR_c_551_n 0.0441655f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.3
cc_106 VPB N_VPWR_c_552_n 0.0083004f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.63
cc_107 VPB N_VPWR_c_553_n 0.0186948f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_108 VPB N_VPWR_c_554_n 0.015305f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=0.74
cc_109 VPB N_VPWR_c_555_n 0.0237863f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=1.3
cc_110 VPB N_VPWR_c_556_n 0.0155697f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.63
cc_111 VPB N_VPWR_c_557_n 0.0121872f $X=-0.19 $Y=1.66 $X2=2.115 $Y2=1.465
cc_112 VPB N_VPWR_c_558_n 0.0540252f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=1.465
cc_113 VPB N_VPWR_c_559_n 0.0244965f $X=-0.19 $Y=1.66 $X2=1.8 $Y2=1.465
cc_114 VPB N_VPWR_c_560_n 0.00632158f $X=-0.19 $Y=1.66 $X2=2.2 $Y2=1.63
cc_115 VPB N_VPWR_c_561_n 0.0186948f $X=-0.19 $Y=1.66 $X2=2.285 $Y2=2.035
cc_116 VPB N_VPWR_c_562_n 0.0209961f $X=-0.19 $Y=1.66 $X2=4.035 $Y2=1.28
cc_117 VPB N_VPWR_c_563_n 0.0389412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_564_n 0.00632158f $X=-0.19 $Y=1.66 $X2=5.49 $Y2=2.115
cc_119 VPB N_VPWR_c_565_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.78 $Y2=1.465
cc_120 VPB N_VPWR_c_566_n 0.00631788f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.465
cc_121 VPB N_VPWR_c_549_n 0.0916352f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=1.465
cc_122 VPB N_X_c_650_n 0.00160496f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_123 VPB N_X_c_651_n 0.00729281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_X_c_652_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_125 VPB N_X_c_653_n 0.00504941f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.3
cc_126 VPB N_X_c_654_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=1.3
cc_127 VPB N_X_c_655_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB X 0.00711055f $X=-0.19 $Y=1.66 $X2=2.115 $Y2=1.465
cc_129 VPB N_A_971_391#_c_721_n 0.00422885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_971_391#_c_722_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_971_391#_c_723_n 0.00379927f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_132 N_A_91_48#_c_152_n N_C1_c_309_n 0.0155473f $X=3.79 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_91_48#_c_155_n N_C1_c_309_n 0.0128865f $X=2.94 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_91_48#_c_156_n N_C1_c_309_n 8.15309e-19 $X=3.955 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_91_48#_c_144_n N_C1_M1015_g 0.00467806f $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_91_48#_c_152_n N_C1_c_310_n 0.0136394f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_137 N_A_91_48#_c_143_n N_C1_c_310_n 0.00150112f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_138 N_A_91_48#_c_155_n N_C1_c_310_n 8.78667e-19 $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_139 N_A_91_48#_c_156_n N_C1_c_310_n 0.013266f $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_140 N_A_91_48#_c_142_n N_C1_M1020_g 0.0100222f $X=3.95 $Y=1.195 $X2=0 $Y2=0
cc_141 N_A_91_48#_c_143_n N_C1_M1020_g 0.00848512f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_142 N_A_91_48#_c_144_n N_C1_M1020_g 0.00505149f $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_91_48#_c_152_n C1 0.0242535f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_144 N_A_91_48#_c_142_n C1 0.00423541f $X=3.95 $Y=1.195 $X2=0 $Y2=0
cc_145 N_A_91_48#_c_143_n C1 0.0247996f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_146 N_A_91_48#_c_144_n C1 0.0213982f $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A_91_48#_c_152_n N_C1_c_308_n 0.00705803f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_148 N_A_91_48#_c_144_n N_C1_c_308_n 7.38005e-19 $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A_91_48#_c_156_n N_C1_c_308_n 9.73339e-19 $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_150 N_A_91_48#_c_140_n N_B1_c_357_n 0.00639074f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_151 N_A_91_48#_c_145_n N_B1_c_357_n 0.0129206f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_152 N_A_91_48#_M1017_g N_B1_c_359_n 0.0209604f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_91_48#_M1009_g N_B1_M1010_g 0.0124997f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_91_48#_c_141_n N_B1_M1010_g 0.0032397f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_155 N_A_91_48#_c_151_n N_B1_M1010_g 0.0138664f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_156 N_A_91_48#_c_155_n N_B1_M1010_g 0.0151463f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_157 N_A_91_48#_c_143_n N_B1_M1023_g 0.0120142f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_158 N_A_91_48#_c_154_n N_B1_M1023_g 0.0179648f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_159 N_A_91_48#_c_156_n N_B1_M1023_g 0.0127326f $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_160 N_A_91_48#_c_142_n N_B1_M1019_g 0.0016974f $X=3.95 $Y=1.195 $X2=0 $Y2=0
cc_161 N_A_91_48#_c_143_n N_B1_M1019_g 0.00136361f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_162 N_A_91_48#_c_144_n N_B1_M1019_g 7.49792e-19 $X=3.555 $Y=1.105 $X2=0 $Y2=0
cc_163 N_A_91_48#_c_143_n N_B1_c_363_n 0.00452782f $X=4.035 $Y=1.95 $X2=0 $Y2=0
cc_164 N_A_91_48#_c_154_n N_B1_c_363_n 0.00229403f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_165 N_A_91_48#_c_140_n B1 0.013554f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_91_48#_c_141_n B1 0.00932184f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_91_48#_c_151_n B1 0.0202829f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_168 N_A_91_48#_c_155_n B1 0.00499989f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_169 N_A_91_48#_M1009_g N_B1_c_364_n 0.0129206f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A_91_48#_c_141_n N_B1_c_364_n 0.00113592f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_171 N_A_91_48#_c_151_n N_B1_c_364_n 0.00818805f $X=2.775 $Y=2.035 $X2=0 $Y2=0
cc_172 N_A_91_48#_c_155_n N_B1_c_364_n 0.0055656f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_173 N_A_91_48#_c_154_n N_A2_M1001_g 0.0141975f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_174 N_A_91_48#_c_157_n N_A2_M1003_g 0.0108929f $X=5.49 $Y=2.115 $X2=0 $Y2=0
cc_175 N_A_91_48#_c_154_n N_A2_c_440_n 0.0301772f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_176 N_A_91_48#_c_157_n N_A2_c_440_n 0.0276979f $X=5.49 $Y=2.115 $X2=0 $Y2=0
cc_177 N_A_91_48#_c_157_n N_A2_c_441_n 0.00330083f $X=5.49 $Y=2.115 $X2=0 $Y2=0
cc_178 N_A_91_48#_c_143_n N_A1_c_486_n 0.00270553f $X=4.035 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_91_48#_c_154_n N_A1_M1005_g 0.019481f $X=5.325 $Y=2.035 $X2=0 $Y2=0
cc_180 N_A_91_48#_c_156_n N_A1_M1005_g 7.03683e-19 $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_181 N_A_91_48#_c_141_n N_VPWR_M1009_s 0.00224929f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_182 N_A_91_48#_c_151_n N_VPWR_M1009_s 0.00958966f $X=2.775 $Y=2.035 $X2=0
+ $Y2=0
cc_183 N_A_91_48#_c_209_p N_VPWR_M1009_s 0.00271221f $X=2.285 $Y=2.035 $X2=0
+ $Y2=0
cc_184 N_A_91_48#_c_152_n N_VPWR_M1000_d 0.0031008f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_185 N_A_91_48#_c_154_n N_VPWR_M1023_d 0.00350187f $X=5.325 $Y=2.035 $X2=0
+ $Y2=0
cc_186 N_A_91_48#_M1004_g N_VPWR_c_551_n 0.00643907f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_91_48#_M1006_g N_VPWR_c_552_n 0.00275958f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_91_48#_M1008_g N_VPWR_c_552_n 0.00275958f $X=1.555 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_91_48#_M1008_g N_VPWR_c_553_n 0.005209f $X=1.555 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_91_48#_M1009_g N_VPWR_c_553_n 0.005209f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_91_48#_M1009_g N_VPWR_c_554_n 0.00410889f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_91_48#_c_151_n N_VPWR_c_554_n 0.0128995f $X=2.775 $Y=2.035 $X2=0
+ $Y2=0
cc_193 N_A_91_48#_c_209_p N_VPWR_c_554_n 0.0119464f $X=2.285 $Y=2.035 $X2=0
+ $Y2=0
cc_194 N_A_91_48#_c_155_n N_VPWR_c_554_n 0.0245367f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_195 N_A_91_48#_c_152_n N_VPWR_c_555_n 0.0220481f $X=3.79 $Y=2.035 $X2=0 $Y2=0
cc_196 N_A_91_48#_c_155_n N_VPWR_c_555_n 0.0204897f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_197 N_A_91_48#_c_156_n N_VPWR_c_555_n 0.0191531f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_198 N_A_91_48#_c_154_n N_VPWR_c_556_n 0.0236753f $X=5.325 $Y=2.035 $X2=0
+ $Y2=0
cc_199 N_A_91_48#_c_156_n N_VPWR_c_556_n 0.0176517f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_200 N_A_91_48#_c_155_n N_VPWR_c_559_n 0.008585f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_201 N_A_91_48#_M1004_g N_VPWR_c_561_n 0.005209f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_91_48#_M1006_g N_VPWR_c_561_n 0.005209f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_91_48#_c_156_n N_VPWR_c_562_n 0.008585f $X=3.955 $Y=2.115 $X2=0 $Y2=0
cc_204 N_A_91_48#_M1004_g N_VPWR_c_549_n 0.00985497f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_91_48#_M1006_g N_VPWR_c_549_n 0.00982526f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_91_48#_M1008_g N_VPWR_c_549_n 0.00982526f $X=1.555 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_91_48#_M1009_g N_VPWR_c_549_n 0.00986727f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_91_48#_c_155_n N_VPWR_c_549_n 0.0107951f $X=2.94 $Y=2.115 $X2=0 $Y2=0
cc_209 N_A_91_48#_c_156_n N_VPWR_c_549_n 0.0107951f $X=3.955 $Y=2.115 $X2=0
+ $Y2=0
cc_210 N_A_91_48#_M1002_g N_X_c_643_n 0.0143817f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_91_48#_M1004_g N_X_c_650_n 0.0166628f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_91_48#_c_145_n N_X_c_650_n 2.51395e-19 $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_213 N_A_91_48#_M1002_g N_X_c_645_n 0.0128625f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_91_48#_M1013_g N_X_c_645_n 3.97481e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_91_48#_M1004_g N_X_c_652_n 0.0184131f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A_91_48#_M1006_g N_X_c_652_n 0.0142049f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A_91_48#_M1008_g N_X_c_652_n 6.31736e-19 $X=1.555 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_91_48#_M1013_g N_X_c_646_n 0.0128832f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_91_48#_M1016_g N_X_c_646_n 0.0124641f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_91_48#_c_140_n N_X_c_646_n 0.0709823f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_221 N_A_91_48#_c_145_n N_X_c_646_n 0.00677187f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_222 N_A_91_48#_M1006_g N_X_c_653_n 0.0134861f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_91_48#_M1008_g N_X_c_653_n 0.0148403f $X=1.555 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A_91_48#_M1009_g N_X_c_653_n 0.00284761f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_91_48#_c_140_n N_X_c_653_n 0.0767299f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_226 N_A_91_48#_c_141_n N_X_c_653_n 0.00779205f $X=2.2 $Y=1.95 $X2=0 $Y2=0
cc_227 N_A_91_48#_c_145_n N_X_c_653_n 0.00702668f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_228 N_A_91_48#_M1013_g N_X_c_647_n 9.31498e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_91_48#_M1016_g N_X_c_647_n 0.00862472f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A_91_48#_M1017_g N_X_c_647_n 3.97481e-19 $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_91_48#_M1006_g N_X_c_654_n 6.31736e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_91_48#_M1008_g N_X_c_654_n 0.0142049f $X=1.555 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_91_48#_M1009_g N_X_c_654_n 0.0146729f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A_91_48#_M1002_g N_X_c_648_n 0.00132316f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_91_48#_c_140_n N_X_c_648_n 0.0181339f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_236 N_A_91_48#_c_145_n N_X_c_648_n 0.00248733f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_237 N_A_91_48#_M1004_g N_X_c_655_n 0.00135419f $X=0.555 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A_91_48#_M1006_g N_X_c_655_n 0.00135419f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_91_48#_c_140_n N_X_c_655_n 0.0275631f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_240 N_A_91_48#_c_145_n N_X_c_655_n 0.00221493f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_241 N_A_91_48#_M1002_g X 0.0109941f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_91_48#_c_140_n X 0.0194533f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_243 N_A_91_48#_c_145_n X 0.0118891f $X=1.89 $Y=1.465 $X2=0 $Y2=0
cc_244 N_A_91_48#_c_154_n N_A_971_391#_M1005_s 0.00165831f $X=5.325 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_245 N_A_91_48#_c_154_n N_A_971_391#_c_725_n 0.0170259f $X=5.325 $Y=2.035
+ $X2=0 $Y2=0
cc_246 N_A_91_48#_M1001_s N_A_971_391#_c_721_n 0.00218982f $X=5.305 $Y=1.955
+ $X2=0 $Y2=0
cc_247 N_A_91_48#_c_157_n N_A_971_391#_c_721_n 0.0177084f $X=5.49 $Y=2.115 $X2=0
+ $Y2=0
cc_248 N_A_91_48#_c_157_n N_A_971_391#_c_723_n 0.00642579f $X=5.49 $Y=2.115
+ $X2=0 $Y2=0
cc_249 N_A_91_48#_M1002_g N_VGND_c_748_n 0.00409307f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_91_48#_M1002_g N_VGND_c_749_n 5.04273e-19 $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_91_48#_M1013_g N_VGND_c_749_n 0.00935695f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_91_48#_M1016_g N_VGND_c_749_n 0.00397833f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_91_48#_M1016_g N_VGND_c_750_n 6.13182e-19 $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_91_48#_M1017_g N_VGND_c_750_n 0.013465f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_91_48#_c_140_n N_VGND_c_750_n 0.029036f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_256 N_A_91_48#_c_145_n N_VGND_c_750_n 0.00354118f $X=1.89 $Y=1.465 $X2=0
+ $Y2=0
cc_257 N_A_91_48#_M1002_g N_VGND_c_753_n 0.00434272f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_91_48#_M1013_g N_VGND_c_753_n 0.00383152f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_91_48#_M1016_g N_VGND_c_754_n 0.00434272f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_91_48#_M1017_g N_VGND_c_754_n 0.00383152f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_91_48#_M1002_g N_VGND_c_758_n 0.00824056f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_91_48#_M1013_g N_VGND_c_758_n 0.0075754f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_91_48#_M1016_g N_VGND_c_758_n 0.00820718f $X=1.46 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_91_48#_M1017_g N_VGND_c_758_n 0.0075754f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_91_48#_M1017_g N_A_510_125#_c_835_n 4.67658e-19 $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_91_48#_M1017_g N_A_510_125#_c_837_n 2.4306e-19 $X=1.89 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_91_48#_c_154_n N_A_510_125#_c_839_n 0.00670788f $X=5.325 $Y=2.035
+ $X2=0 $Y2=0
cc_268 N_A_91_48#_c_142_n N_A_510_125#_c_840_n 0.00537821f $X=3.95 $Y=1.195
+ $X2=0 $Y2=0
cc_269 N_A_91_48#_c_143_n N_A_510_125#_c_840_n 2.47868e-19 $X=4.035 $Y=1.95
+ $X2=0 $Y2=0
cc_270 N_A_91_48#_c_154_n N_A_510_125#_c_840_n 0.00812137f $X=5.325 $Y=2.035
+ $X2=0 $Y2=0
cc_271 N_A_91_48#_c_142_n N_A_597_125#_M1020_d 0.0041638f $X=3.95 $Y=1.195 $X2=0
+ $Y2=0
cc_272 N_A_91_48#_c_152_n N_A_597_125#_c_907_n 0.00298145f $X=3.79 $Y=2.035
+ $X2=0 $Y2=0
cc_273 N_A_91_48#_c_155_n N_A_597_125#_c_907_n 0.0021645f $X=2.94 $Y=2.115 $X2=0
+ $Y2=0
cc_274 N_A_91_48#_c_144_n N_A_597_125#_c_907_n 0.0128711f $X=3.555 $Y=1.105
+ $X2=0 $Y2=0
cc_275 N_A_91_48#_M1015_s N_A_597_125#_c_908_n 0.00169276f $X=3.415 $Y=0.625
+ $X2=0 $Y2=0
cc_276 N_A_91_48#_c_142_n N_A_597_125#_c_908_n 0.0048036f $X=3.95 $Y=1.195 $X2=0
+ $Y2=0
cc_277 N_A_91_48#_c_144_n N_A_597_125#_c_908_n 0.0161743f $X=3.555 $Y=1.105
+ $X2=0 $Y2=0
cc_278 N_A_91_48#_c_142_n N_A_597_125#_c_910_n 0.0182562f $X=3.95 $Y=1.195 $X2=0
+ $Y2=0
cc_279 N_C1_M1015_g N_B1_c_358_n 0.00737859f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_280 N_C1_M1020_g N_B1_c_358_n 0.00737859f $X=3.77 $Y=0.945 $X2=0 $Y2=0
cc_281 N_C1_c_308_n N_B1_M1010_g 0.0235877f $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_282 N_C1_M1015_g N_B1_c_360_n 0.00877012f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_283 N_C1_c_310_n N_B1_M1023_g 0.0159955f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_284 N_C1_c_308_n N_B1_M1023_g 0.0140334f $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_285 N_C1_M1020_g N_B1_M1019_g 0.0207562f $X=3.77 $Y=0.945 $X2=0 $Y2=0
cc_286 N_C1_M1020_g N_B1_c_363_n 0.0140334f $X=3.77 $Y=0.945 $X2=0 $Y2=0
cc_287 C1 N_B1_c_363_n 2.95263e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_288 N_C1_M1015_g B1 0.00140466f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_289 C1 B1 0.00858387f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_290 N_C1_c_308_n B1 3.40608e-19 $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_291 C1 N_B1_c_364_n 0.00105873f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_292 N_C1_c_308_n N_B1_c_364_n 0.0178595f $X=3.73 $Y=1.665 $X2=0 $Y2=0
cc_293 N_C1_c_309_n N_VPWR_c_555_n 0.00438901f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_294 N_C1_c_310_n N_VPWR_c_555_n 0.00646137f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_295 N_C1_c_309_n N_VPWR_c_559_n 0.00536648f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_296 N_C1_c_310_n N_VPWR_c_562_n 0.00536648f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_297 N_C1_c_309_n N_VPWR_c_549_n 0.0059403f $X=3.165 $Y=1.88 $X2=0 $Y2=0
cc_298 N_C1_c_310_n N_VPWR_c_549_n 0.0059403f $X=3.73 $Y=1.88 $X2=0 $Y2=0
cc_299 N_C1_M1015_g N_A_510_125#_c_836_n 0.00116683f $X=3.34 $Y=0.945 $X2=0
+ $Y2=0
cc_300 N_C1_M1020_g N_A_510_125#_c_836_n 0.00116683f $X=3.77 $Y=0.945 $X2=0
+ $Y2=0
cc_301 N_C1_M1015_g N_A_597_125#_c_907_n 2.23441e-19 $X=3.34 $Y=0.945 $X2=0
+ $Y2=0
cc_302 N_C1_c_308_n N_A_597_125#_c_907_n 0.00323873f $X=3.73 $Y=1.665 $X2=0
+ $Y2=0
cc_303 N_C1_M1015_g N_A_597_125#_c_908_n 0.0114956f $X=3.34 $Y=0.945 $X2=0 $Y2=0
cc_304 N_C1_M1020_g N_A_597_125#_c_908_n 0.00923977f $X=3.77 $Y=0.945 $X2=0
+ $Y2=0
cc_305 N_C1_M1020_g N_A_597_125#_c_910_n 4.44855e-19 $X=3.77 $Y=0.945 $X2=0
+ $Y2=0
cc_306 N_B1_c_363_n N_A1_c_486_n 0.00605855f $X=4.217 $Y=1.49 $X2=-0.19
+ $Y2=-0.245
cc_307 N_B1_M1023_g N_A1_M1005_g 0.029373f $X=4.18 $Y=2.375 $X2=0 $Y2=0
cc_308 N_B1_M1019_g N_A1_M1012_g 0.0132251f $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_309 N_B1_c_358_n N_A1_c_490_n 0.0132251f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_310 N_B1_M1010_g N_VPWR_c_554_n 0.0083306f $X=2.715 $Y=2.375 $X2=0 $Y2=0
cc_311 N_B1_M1023_g N_VPWR_c_556_n 0.00641497f $X=4.18 $Y=2.375 $X2=0 $Y2=0
cc_312 N_B1_M1010_g N_VPWR_c_559_n 0.00536648f $X=2.715 $Y=2.375 $X2=0 $Y2=0
cc_313 N_B1_M1023_g N_VPWR_c_562_n 0.00536648f $X=4.18 $Y=2.375 $X2=0 $Y2=0
cc_314 N_B1_M1010_g N_VPWR_c_549_n 0.0059403f $X=2.715 $Y=2.375 $X2=0 $Y2=0
cc_315 N_B1_M1023_g N_VPWR_c_549_n 0.0059403f $X=4.18 $Y=2.375 $X2=0 $Y2=0
cc_316 N_B1_M1010_g N_X_c_654_n 8.99627e-19 $X=2.715 $Y=2.375 $X2=0 $Y2=0
cc_317 N_B1_c_359_n N_VGND_c_750_n 0.0144891f $X=2.475 $Y=0.18 $X2=0 $Y2=0
cc_318 N_B1_c_358_n N_VGND_c_751_n 0.00107466f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_319 N_B1_M1019_g N_VGND_c_751_n 2.44756e-19 $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_320 N_B1_c_359_n N_VGND_c_755_n 0.045518f $X=2.475 $Y=0.18 $X2=0 $Y2=0
cc_321 N_B1_c_358_n N_VGND_c_758_n 0.047086f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_322 N_B1_c_359_n N_VGND_c_758_n 0.0114395f $X=2.475 $Y=0.18 $X2=0 $Y2=0
cc_323 N_B1_c_357_n N_A_510_125#_c_835_n 0.0110018f $X=2.4 $Y=1.34 $X2=0 $Y2=0
cc_324 N_B1_c_360_n N_A_510_125#_c_835_n 0.00295702f $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_325 B1 N_A_510_125#_c_835_n 0.0206962f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_326 N_B1_c_364_n N_A_510_125#_c_835_n 0.00530945f $X=2.715 $Y=1.552 $X2=0
+ $Y2=0
cc_327 N_B1_c_358_n N_A_510_125#_c_836_n 0.023808f $X=4.195 $Y=0.18 $X2=0 $Y2=0
cc_328 N_B1_c_360_n N_A_510_125#_c_836_n 0.00366331f $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_329 N_B1_M1019_g N_A_510_125#_c_836_n 0.0156653f $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_330 N_B1_c_357_n N_A_510_125#_c_837_n 0.00198754f $X=2.4 $Y=1.34 $X2=0 $Y2=0
cc_331 N_B1_c_358_n N_A_510_125#_c_837_n 0.00732085f $X=4.195 $Y=0.18 $X2=0
+ $Y2=0
cc_332 N_B1_M1019_g N_A_510_125#_c_838_n 0.0047697f $X=4.27 $Y=0.945 $X2=0 $Y2=0
cc_333 N_B1_M1019_g N_A_510_125#_c_840_n 2.13054e-19 $X=4.27 $Y=0.945 $X2=0
+ $Y2=0
cc_334 N_B1_c_360_n N_A_597_125#_c_907_n 4.5765e-19 $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_335 N_B1_c_360_n N_A_597_125#_c_909_n 2.90897e-19 $X=2.91 $Y=1.34 $X2=0 $Y2=0
cc_336 N_B1_M1019_g N_A_597_125#_c_910_n 0.00538803f $X=4.27 $Y=0.945 $X2=0
+ $Y2=0
cc_337 N_B1_c_363_n N_A_597_125#_c_910_n 0.00185774f $X=4.217 $Y=1.49 $X2=0
+ $Y2=0
cc_338 N_A2_c_441_n N_A1_c_486_n 0.0157564f $X=5.715 $Y=1.615 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A2_c_440_n N_A1_M1005_g 0.0102979f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_340 N_A2_c_441_n N_A1_M1005_g 0.0349674f $X=5.715 $Y=1.615 $X2=0 $Y2=0
cc_341 N_A2_M1011_g N_A1_M1012_g 0.0157564f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_342 N_A2_M1011_g N_A1_c_489_n 0.00902758f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_343 N_A2_M1021_g N_A1_c_489_n 0.00894529f $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_344 N_A2_M1003_g N_A1_M1018_g 0.0154921f $X=5.715 $Y=2.455 $X2=0 $Y2=0
cc_345 N_A2_M1021_g N_A1_M1022_g 0.0255078f $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_346 N_A2_c_440_n A1 0.0205984f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_347 N_A2_c_441_n A1 4.1393e-19 $X=5.715 $Y=1.615 $X2=0 $Y2=0
cc_348 N_A2_c_440_n N_A1_c_493_n 4.16072e-19 $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_349 N_A2_c_441_n N_A1_c_493_n 0.018249f $X=5.715 $Y=1.615 $X2=0 $Y2=0
cc_350 N_A2_M1001_g N_VPWR_c_563_n 0.0033082f $X=5.215 $Y=2.455 $X2=0 $Y2=0
cc_351 N_A2_M1003_g N_VPWR_c_563_n 0.00330849f $X=5.715 $Y=2.455 $X2=0 $Y2=0
cc_352 N_A2_M1001_g N_VPWR_c_549_n 0.00653145f $X=5.215 $Y=2.455 $X2=0 $Y2=0
cc_353 N_A2_M1003_g N_VPWR_c_549_n 0.00653145f $X=5.715 $Y=2.455 $X2=0 $Y2=0
cc_354 N_A2_M1001_g N_A_971_391#_c_725_n 0.00888608f $X=5.215 $Y=2.455 $X2=0
+ $Y2=0
cc_355 N_A2_M1003_g N_A_971_391#_c_725_n 8.58708e-19 $X=5.715 $Y=2.455 $X2=0
+ $Y2=0
cc_356 N_A2_M1001_g N_A_971_391#_c_721_n 0.0119072f $X=5.215 $Y=2.455 $X2=0
+ $Y2=0
cc_357 N_A2_M1003_g N_A_971_391#_c_721_n 0.014321f $X=5.715 $Y=2.455 $X2=0 $Y2=0
cc_358 N_A2_M1001_g N_A_971_391#_c_722_n 0.00196843f $X=5.215 $Y=2.455 $X2=0
+ $Y2=0
cc_359 N_A2_M1011_g N_VGND_c_751_n 0.00684563f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_360 N_A2_M1021_g N_VGND_c_751_n 4.05518e-19 $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_361 N_A2_M1011_g N_VGND_c_752_n 4.23833e-19 $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_362 N_A2_M1021_g N_VGND_c_752_n 0.00771226f $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_363 N_A2_M1011_g N_VGND_c_758_n 8.92987e-19 $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_364 N_A2_M1021_g N_VGND_c_758_n 7.97988e-19 $X=5.725 $Y=0.945 $X2=0 $Y2=0
cc_365 N_A2_M1011_g N_A_510_125#_c_839_n 0.0128053f $X=5.24 $Y=0.945 $X2=0 $Y2=0
cc_366 N_A2_c_440_n N_A_510_125#_c_839_n 0.0319578f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_367 N_A2_M1021_g N_A_510_125#_c_842_n 0.0125779f $X=5.725 $Y=0.945 $X2=0
+ $Y2=0
cc_368 N_A2_c_440_n N_A_510_125#_c_842_n 0.0174392f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_369 N_A2_c_441_n N_A_510_125#_c_842_n 8.04419e-19 $X=5.715 $Y=1.615 $X2=0
+ $Y2=0
cc_370 N_A2_M1021_g N_A_510_125#_c_843_n 8.30676e-19 $X=5.725 $Y=0.945 $X2=0
+ $Y2=0
cc_371 N_A2_c_440_n N_A_510_125#_c_844_n 0.0210724f $X=5.67 $Y=1.615 $X2=0 $Y2=0
cc_372 N_A2_c_441_n N_A_510_125#_c_844_n 0.00370253f $X=5.715 $Y=1.615 $X2=0
+ $Y2=0
cc_373 N_A1_M1005_g N_VPWR_c_556_n 0.00341369f $X=4.765 $Y=2.455 $X2=0 $Y2=0
cc_374 N_A1_M1018_g N_VPWR_c_558_n 0.00346677f $X=6.165 $Y=2.455 $X2=0 $Y2=0
cc_375 A1 N_VPWR_c_558_n 0.0276867f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_376 N_A1_c_493_n N_VPWR_c_558_n 0.0030998f $X=6.24 $Y=1.615 $X2=0 $Y2=0
cc_377 N_A1_M1005_g N_VPWR_c_563_n 0.00512529f $X=4.765 $Y=2.455 $X2=0 $Y2=0
cc_378 N_A1_M1018_g N_VPWR_c_563_n 0.00512529f $X=6.165 $Y=2.455 $X2=0 $Y2=0
cc_379 N_A1_M1005_g N_VPWR_c_549_n 0.00653145f $X=4.765 $Y=2.455 $X2=0 $Y2=0
cc_380 N_A1_M1018_g N_VPWR_c_549_n 0.00653145f $X=6.165 $Y=2.455 $X2=0 $Y2=0
cc_381 N_A1_M1005_g N_A_971_391#_c_725_n 0.00751518f $X=4.765 $Y=2.455 $X2=0
+ $Y2=0
cc_382 N_A1_M1018_g N_A_971_391#_c_721_n 0.00350328f $X=6.165 $Y=2.455 $X2=0
+ $Y2=0
cc_383 N_A1_M1005_g N_A_971_391#_c_722_n 0.00350107f $X=4.765 $Y=2.455 $X2=0
+ $Y2=0
cc_384 N_A1_M1018_g N_A_971_391#_c_723_n 0.0116237f $X=6.165 $Y=2.455 $X2=0
+ $Y2=0
cc_385 A1 N_A_971_391#_c_723_n 0.00231492f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_386 N_A1_M1012_g N_VGND_c_751_n 0.0139844f $X=4.78 $Y=0.945 $X2=0 $Y2=0
cc_387 N_A1_c_489_n N_VGND_c_751_n 0.0185436f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_388 N_A1_c_490_n N_VGND_c_751_n 0.00364942f $X=4.855 $Y=0.18 $X2=0 $Y2=0
cc_389 N_A1_c_489_n N_VGND_c_752_n 0.0232456f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_390 N_A1_M1022_g N_VGND_c_752_n 0.0151144f $X=6.225 $Y=0.945 $X2=0 $Y2=0
cc_391 N_A1_c_490_n N_VGND_c_755_n 0.00486043f $X=4.855 $Y=0.18 $X2=0 $Y2=0
cc_392 N_A1_c_489_n N_VGND_c_756_n 0.0184168f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_393 N_A1_c_489_n N_VGND_c_757_n 0.00730708f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_394 N_A1_c_489_n N_VGND_c_758_n 0.0323021f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_395 N_A1_c_490_n N_VGND_c_758_n 0.00859636f $X=4.855 $Y=0.18 $X2=0 $Y2=0
cc_396 N_A1_M1012_g N_A_510_125#_c_836_n 0.00157748f $X=4.78 $Y=0.945 $X2=0
+ $Y2=0
cc_397 N_A1_M1012_g N_A_510_125#_c_838_n 0.00421702f $X=4.78 $Y=0.945 $X2=0
+ $Y2=0
cc_398 N_A1_c_486_n N_A_510_125#_c_839_n 0.00107945f $X=4.765 $Y=1.43 $X2=0
+ $Y2=0
cc_399 N_A1_M1012_g N_A_510_125#_c_839_n 0.0167942f $X=4.78 $Y=0.945 $X2=0 $Y2=0
cc_400 N_A1_c_489_n N_A_510_125#_c_841_n 0.00490132f $X=6.15 $Y=0.18 $X2=0 $Y2=0
cc_401 N_A1_M1022_g N_A_510_125#_c_842_n 0.0124988f $X=6.225 $Y=0.945 $X2=0
+ $Y2=0
cc_402 A1 N_A_510_125#_c_842_n 0.0421713f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_403 N_A1_c_493_n N_A_510_125#_c_842_n 0.0044184f $X=6.24 $Y=1.615 $X2=0 $Y2=0
cc_404 N_A1_M1022_g N_A_510_125#_c_843_n 0.00759673f $X=6.225 $Y=0.945 $X2=0
+ $Y2=0
cc_405 N_VPWR_M1004_s N_X_c_650_n 5.5277e-19 $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_406 N_VPWR_c_551_n N_X_c_650_n 0.00427553f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_407 N_VPWR_M1004_s N_X_c_651_n 0.0035139f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_408 N_VPWR_c_551_n N_X_c_651_n 0.0207257f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_409 N_VPWR_c_551_n N_X_c_652_n 0.0323093f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_410 N_VPWR_c_552_n N_X_c_652_n 0.0323093f $X=1.28 $Y=2.305 $X2=0 $Y2=0
cc_411 N_VPWR_c_561_n N_X_c_652_n 0.0144623f $X=1.115 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_c_549_n N_X_c_652_n 0.0118344f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_413 N_VPWR_M1006_s N_X_c_653_n 0.00279273f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_414 N_VPWR_c_552_n N_X_c_653_n 0.0208278f $X=1.28 $Y=2.305 $X2=0 $Y2=0
cc_415 N_VPWR_c_552_n N_X_c_654_n 0.0323093f $X=1.28 $Y=2.305 $X2=0 $Y2=0
cc_416 N_VPWR_c_553_n N_X_c_654_n 0.0144623f $X=2.115 $Y=3.33 $X2=0 $Y2=0
cc_417 N_VPWR_c_554_n N_X_c_654_n 0.0266809f $X=2.28 $Y=2.405 $X2=0 $Y2=0
cc_418 N_VPWR_c_549_n N_X_c_654_n 0.0118344f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_419 N_VPWR_c_558_n N_A_971_391#_c_721_n 0.0121327f $X=6.44 $Y=2.115 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_563_n N_A_971_391#_c_721_n 0.0618604f $X=6.275 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_549_n N_A_971_391#_c_721_n 0.0343867f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_556_n N_A_971_391#_c_722_n 0.0121327f $X=4.49 $Y=2.41 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_563_n N_A_971_391#_c_722_n 0.0234458f $X=6.275 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_549_n N_A_971_391#_c_722_n 0.0125551f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_558_n N_A_971_391#_c_723_n 0.0344717f $X=6.44 $Y=2.115 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_558_n N_A_510_125#_c_842_n 3.21367e-19 $X=6.44 $Y=2.115 $X2=0
+ $Y2=0
cc_427 N_X_c_643_n N_VGND_M1002_d 4.46468e-19 $X=0.58 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_428 N_X_c_644_n N_VGND_M1002_d 0.00291902f $X=0.355 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_429 N_X_c_646_n N_VGND_M1013_d 0.00250873f $X=1.51 $Y=1.045 $X2=0 $Y2=0
cc_430 N_X_c_643_n N_VGND_c_748_n 0.00346194f $X=0.58 $Y=1.045 $X2=0 $Y2=0
cc_431 N_X_c_644_n N_VGND_c_748_n 0.0184602f $X=0.355 $Y=1.045 $X2=0 $Y2=0
cc_432 N_X_c_645_n N_VGND_c_748_n 0.0158413f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_433 N_X_c_645_n N_VGND_c_749_n 0.0164981f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_434 N_X_c_646_n N_VGND_c_749_n 0.0210288f $X=1.51 $Y=1.045 $X2=0 $Y2=0
cc_435 N_X_c_647_n N_VGND_c_749_n 0.0166127f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_436 N_X_c_646_n N_VGND_c_750_n 0.00697079f $X=1.51 $Y=1.045 $X2=0 $Y2=0
cc_437 N_X_c_647_n N_VGND_c_750_n 0.0225912f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_438 N_X_c_645_n N_VGND_c_753_n 0.0109942f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_439 N_X_c_647_n N_VGND_c_754_n 0.0109942f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_440 N_X_c_645_n N_VGND_c_758_n 0.00904371f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_441 N_X_c_647_n N_VGND_c_758_n 0.00904371f $X=1.675 $Y=0.515 $X2=0 $Y2=0
cc_442 N_A_971_391#_c_723_n N_A_510_125#_c_842_n 0.00707466f $X=5.94 $Y=2.115
+ $X2=0 $Y2=0
cc_443 N_VGND_c_750_n N_A_510_125#_c_835_n 0.0426691f $X=2.105 $Y=0.515 $X2=0
+ $Y2=0
cc_444 N_VGND_c_751_n N_A_510_125#_c_836_n 0.0137357f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_445 N_VGND_c_755_n N_A_510_125#_c_836_n 0.121756f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_758_n N_A_510_125#_c_836_n 0.0642692f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_750_n N_A_510_125#_c_837_n 0.011157f $X=2.105 $Y=0.515 $X2=0
+ $Y2=0
cc_448 N_VGND_c_755_n N_A_510_125#_c_837_n 0.0170431f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_758_n N_A_510_125#_c_837_n 0.00857552f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_751_n N_A_510_125#_c_838_n 0.0259901f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_451 N_VGND_M1012_d N_A_510_125#_c_839_n 0.00210887f $X=4.855 $Y=0.625 $X2=0
+ $Y2=0
cc_452 N_VGND_c_751_n N_A_510_125#_c_839_n 0.0179772f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_453 N_VGND_c_751_n N_A_510_125#_c_841_n 0.0132249f $X=5 $Y=0.77 $X2=0 $Y2=0
cc_454 N_VGND_c_752_n N_A_510_125#_c_841_n 0.0127348f $X=5.94 $Y=0.77 $X2=0
+ $Y2=0
cc_455 N_VGND_c_756_n N_A_510_125#_c_841_n 0.00533975f $X=5.775 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_c_758_n N_A_510_125#_c_841_n 0.00671154f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_M1021_s N_A_510_125#_c_842_n 0.00250873f $X=5.8 $Y=0.625 $X2=0
+ $Y2=0
cc_458 N_VGND_c_752_n N_A_510_125#_c_842_n 0.0209867f $X=5.94 $Y=0.77 $X2=0
+ $Y2=0
cc_459 N_VGND_c_752_n N_A_510_125#_c_843_n 0.0133605f $X=5.94 $Y=0.77 $X2=0
+ $Y2=0
cc_460 N_VGND_c_757_n N_A_510_125#_c_843_n 0.00701744f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_758_n N_A_510_125#_c_843_n 0.0100487f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_462 N_A_510_125#_c_836_n N_A_597_125#_c_908_n 0.0471472f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_463 N_A_510_125#_c_835_n N_A_597_125#_c_909_n 0.00186525f $X=2.695 $Y=0.76
+ $X2=0 $Y2=0
cc_464 N_A_510_125#_c_836_n N_A_597_125#_c_909_n 0.0134458f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_465 N_A_510_125#_c_836_n N_A_597_125#_c_910_n 0.0244253f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_466 N_A_510_125#_c_838_n N_A_597_125#_c_910_n 0.0134764f $X=4.485 $Y=0.77
+ $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_585_368# A2 a_177_48# VPB pshort w=1e+06u l=180000u
+  ad=3.3e+11p pd=2.66e+06u as=2.7e+11p ps=2.54e+06u
M1001 VGND a_177_48# X VNB nlowvt w=740000u l=150000u
+  ad=7.8915e+11p pd=6.84e+06u as=2.072e+11p ps=2.04e+06u
M1002 VPWR B1_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=1.4348e+12p pd=9.16e+06u as=2.352e+11p ps=2.24e+06u
M1003 VGND A2 a_487_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.07e+11p ps=4.06e+06u
M1004 X a_177_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VPWR a_177_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND B1_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5125e+11p ps=1.65e+06u
M1007 X a_177_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_487_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_585_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_177_48# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_487_74# a_27_74# a_177_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.035e+11p ps=2.03e+06u
.ends

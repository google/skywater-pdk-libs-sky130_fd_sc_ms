* File: sky130_fd_sc_ms__o311ai_2.pxi.spice
* Created: Fri Aug 28 18:01:42 2020
* 
x_PM_SKY130_FD_SC_MS__O311AI_2%A1 N_A1_M1003_g N_A1_M1005_g N_A1_M1014_g
+ N_A1_M1018_g A1 A1 N_A1_c_103_n PM_SKY130_FD_SC_MS__O311AI_2%A1
x_PM_SKY130_FD_SC_MS__O311AI_2%A2 N_A2_c_146_n N_A2_M1001_g N_A2_M1012_g
+ N_A2_M1013_g N_A2_M1002_g A2 A2 A2 N_A2_c_145_n
+ PM_SKY130_FD_SC_MS__O311AI_2%A2
x_PM_SKY130_FD_SC_MS__O311AI_2%A3 N_A3_M1009_g N_A3_M1016_g N_A3_c_202_n
+ N_A3_M1017_g N_A3_c_199_n N_A3_c_200_n N_A3_c_205_n N_A3_M1019_g A3 A3
+ PM_SKY130_FD_SC_MS__O311AI_2%A3
x_PM_SKY130_FD_SC_MS__O311AI_2%B1 N_B1_c_261_n N_B1_M1008_g N_B1_c_262_n
+ N_B1_c_263_n N_B1_c_264_n N_B1_M1015_g N_B1_M1000_g N_B1_c_265_n N_B1_M1006_g
+ N_B1_c_266_n B1 B1 N_B1_c_268_n PM_SKY130_FD_SC_MS__O311AI_2%B1
x_PM_SKY130_FD_SC_MS__O311AI_2%C1 N_C1_M1007_g N_C1_M1004_g N_C1_M1010_g
+ N_C1_M1011_g C1 C1 N_C1_c_336_n PM_SKY130_FD_SC_MS__O311AI_2%C1
x_PM_SKY130_FD_SC_MS__O311AI_2%A_28_368# N_A_28_368#_M1005_s N_A_28_368#_M1014_s
+ N_A_28_368#_M1002_s N_A_28_368#_c_382_n N_A_28_368#_c_383_n
+ N_A_28_368#_c_390_n N_A_28_368#_c_384_n N_A_28_368#_c_396_n
+ N_A_28_368#_c_400_n N_A_28_368#_c_385_n PM_SKY130_FD_SC_MS__O311AI_2%A_28_368#
x_PM_SKY130_FD_SC_MS__O311AI_2%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_M1007_d
+ N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n
+ VPWR N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_419_n N_VPWR_c_428_n
+ N_VPWR_c_429_n PM_SKY130_FD_SC_MS__O311AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O311AI_2%A_310_368# N_A_310_368#_M1001_d
+ N_A_310_368#_M1017_d N_A_310_368#_c_489_n N_A_310_368#_c_487_n
+ N_A_310_368#_c_488_n N_A_310_368#_c_507_p
+ PM_SKY130_FD_SC_MS__O311AI_2%A_310_368#
x_PM_SKY130_FD_SC_MS__O311AI_2%Y N_Y_M1004_s N_Y_M1011_s N_Y_M1017_s N_Y_M1019_s
+ N_Y_M1006_s N_Y_M1010_s N_Y_c_519_n N_Y_c_514_n N_Y_c_533_n N_Y_c_515_n
+ N_Y_c_510_n N_Y_c_553_n N_Y_c_516_n N_Y_c_517_n N_Y_c_511_n N_Y_c_518_n
+ N_Y_c_529_n N_Y_c_539_n Y Y Y Y PM_SKY130_FD_SC_MS__O311AI_2%Y
x_PM_SKY130_FD_SC_MS__O311AI_2%A_27_74# N_A_27_74#_M1003_d N_A_27_74#_M1018_d
+ N_A_27_74#_M1013_s N_A_27_74#_M1016_s N_A_27_74#_M1015_s N_A_27_74#_c_600_n
+ N_A_27_74#_c_601_n N_A_27_74#_c_602_n N_A_27_74#_c_603_n N_A_27_74#_c_604_n
+ N_A_27_74#_c_605_n N_A_27_74#_c_606_n N_A_27_74#_c_607_n N_A_27_74#_c_608_n
+ N_A_27_74#_c_609_n N_A_27_74#_c_610_n N_A_27_74#_c_611_n N_A_27_74#_c_612_n
+ PM_SKY130_FD_SC_MS__O311AI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O311AI_2%VGND N_VGND_M1003_s N_VGND_M1012_d N_VGND_M1009_d
+ N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n VGND N_VGND_c_684_n
+ N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n
+ N_VGND_c_690_n N_VGND_c_691_n PM_SKY130_FD_SC_MS__O311AI_2%VGND
x_PM_SKY130_FD_SC_MS__O311AI_2%A_670_74# N_A_670_74#_M1008_d N_A_670_74#_M1004_d
+ N_A_670_74#_c_763_n N_A_670_74#_c_748_n N_A_670_74#_c_749_n
+ N_A_670_74#_c_754_n PM_SKY130_FD_SC_MS__O311AI_2%A_670_74#
cc_1 VNB N_A1_M1003_g 0.0327337f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1018_g 0.0253298f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_3 VNB A1 0.0167148f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A1_c_103_n 0.0405875f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.515
cc_5 VNB N_A2_M1012_g 0.0240209f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_6 VNB N_A2_M1013_g 0.0237011f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_7 VNB A2 0.0105759f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_A2_c_145_n 0.0351858f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.515
cc_9 VNB N_A3_M1009_g 0.0246497f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A3_M1016_g 0.0238365f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_11 VNB N_A3_c_199_n 0.0138978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A3_c_200_n 0.0412373f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_13 VNB A3 0.00488881f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_14 VNB N_B1_c_261_n 0.0157815f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_15 VNB N_B1_c_262_n 0.0203202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_263_n 0.00814437f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.68
cc_17 VNB N_B1_c_264_n 0.0179631f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_18 VNB N_B1_c_265_n 0.027212f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_19 VNB N_B1_c_266_n 0.0143038f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB B1 0.006035f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_21 VNB N_B1_c_268_n 0.0170025f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_22 VNB N_C1_M1007_g 0.00141505f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_23 VNB N_C1_M1004_g 0.0239843f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_24 VNB N_C1_M1010_g 0.0017572f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_25 VNB N_C1_M1011_g 0.0291604f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_26 VNB C1 0.0152566f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_C1_c_336_n 0.0675406f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.515
cc_28 VNB N_VPWR_c_419_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_510_n 0.012331f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_30 VNB N_Y_c_511_n 0.0247743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB Y 0.0060107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.00619631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_600_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_A_27_74#_c_601_n 0.00612368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_602_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_36 VNB N_A_27_74#_c_603_n 0.00253842f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_37 VNB N_A_27_74#_c_604_n 0.00285384f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_38 VNB N_A_27_74#_c_605_n 0.00253214f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_39 VNB N_A_27_74#_c_606_n 0.00491768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_607_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_608_n 0.00725544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_609_n 0.00351892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_610_n 0.00234762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_74#_c_611_n 0.0028931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_74#_c_612_n 0.00155944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_681_n 0.00576795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_682_n 0.00276855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_683_n 0.00563529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_684_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_50 VNB N_VGND_c_685_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_686_n 0.016883f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_52 VNB N_VGND_c_687_n 0.0749446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_688_n 0.326435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_689_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_690_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_691_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_670_74#_c_748_n 0.0178206f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_58 VNB N_A_670_74#_c_749_n 0.00417668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_A1_M1005_g 0.0277014f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_60 VPB N_A1_M1014_g 0.0217773f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_61 VPB A1 0.010983f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_62 VPB N_A1_c_103_n 0.00522345f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.515
cc_63 VPB N_A2_c_146_n 0.0176103f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_64 VPB N_A2_M1002_g 0.0253379f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_65 VPB A2 0.00998577f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_66 VPB N_A2_c_145_n 0.0118258f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.515
cc_67 VPB N_A3_c_202_n 0.0225686f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.68
cc_68 VPB N_A3_c_199_n 0.00634024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A3_c_200_n 0.0273884f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.35
cc_70 VPB N_A3_c_205_n 0.0189996f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_71 VPB A3 0.00793647f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_72 VPB N_B1_M1000_g 0.0202409f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_73 VPB N_B1_c_265_n 0.00532161f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.35
cc_74 VPB N_B1_M1006_g 0.0202441f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_75 VPB B1 0.00514479f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_76 VPB N_C1_M1007_g 0.0212685f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_77 VPB N_C1_M1010_g 0.0288517f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_78 VPB C1 0.0107056f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_79 VPB N_A_28_368#_c_382_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_80 VPB N_A_28_368#_c_383_n 0.0352219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_28_368#_c_384_n 0.00275632f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_82 VPB N_A_28_368#_c_385_n 0.00730977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_420_n 0.00564953f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_84 VPB N_VPWR_c_421_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_85 VPB N_VPWR_c_422_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_423_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_87 VPB N_VPWR_c_424_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_88 VPB N_VPWR_c_425_n 0.0757789f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_426_n 0.0205835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_419_n 0.0808124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_428_n 0.0248432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_429_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_310_368#_c_487_n 0.0195444f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_94 VPB N_A_310_368#_c_488_n 0.00382902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_Y_c_514_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_96 VPB N_Y_c_515_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_Y_c_516_n 0.00723723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_Y_c_517_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_Y_c_518_n 0.00720753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 N_A1_M1018_g N_A2_M1012_g 0.0179972f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_101 A1 A2 0.0290771f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A1_c_103_n A2 0.00542073f $X=0.985 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A1_M1014_g N_A2_c_145_n 0.0151363f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_104 A1 N_A2_c_145_n 2.03322e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_105 N_A1_c_103_n N_A2_c_145_n 0.0179972f $X=0.985 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A1_M1005_g N_A_28_368#_c_382_n 8.84614e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_107 A1 N_A_28_368#_c_382_n 0.0259449f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A1_M1005_g N_A_28_368#_c_383_n 0.0122513f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A1_M1014_g N_A_28_368#_c_383_n 6.64069e-19 $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A1_M1005_g N_A_28_368#_c_390_n 0.0129934f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A1_M1014_g N_A_28_368#_c_390_n 0.0200914f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_112 A1 N_A_28_368#_c_390_n 0.0271227f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A1_c_103_n N_A_28_368#_c_390_n 5.45297e-19 $X=0.985 $Y=1.515 $X2=0
+ $Y2=0
cc_114 N_A1_M1005_g N_VPWR_c_420_n 0.00299709f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A1_M1014_g N_VPWR_c_420_n 0.0111632f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A1_M1014_g N_VPWR_c_425_n 0.00490827f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A1_M1005_g N_VPWR_c_419_n 0.00986126f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A1_M1014_g N_VPWR_c_419_n 0.00969246f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A1_M1005_g N_VPWR_c_428_n 0.005209f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A1_M1003_g N_A_27_74#_c_600_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A1_M1003_g N_A_27_74#_c_601_n 0.013995f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A1_M1018_g N_A_27_74#_c_601_n 0.0188629f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_123 A1 N_A_27_74#_c_601_n 0.0356901f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A1_c_103_n N_A_27_74#_c_601_n 0.00382368f $X=0.985 $Y=1.515 $X2=0 $Y2=0
cc_125 A1 N_A_27_74#_c_602_n 0.0216404f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A1_M1018_g N_A_27_74#_c_603_n 4.77375e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_M1003_g N_VGND_c_681_n 0.0133418f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A1_M1018_g N_VGND_c_681_n 0.00435015f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A1_M1018_g N_VGND_c_682_n 4.54333e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A1_M1003_g N_VGND_c_684_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A1_M1018_g N_VGND_c_685_n 0.00461464f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A1_M1003_g N_VGND_c_688_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A1_M1018_g N_VGND_c_688_n 0.00909082f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A2_M1013_g N_A3_M1009_g 0.0164357f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_135 A2 N_A3_c_202_n 2.03697e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_136 A2 N_A3_c_200_n 0.00413316f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_c_145_n N_A3_c_200_n 0.0205015f $X=1.915 $Y=1.56 $X2=0 $Y2=0
cc_138 N_A2_M1002_g A3 2.73266e-19 $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_139 A2 A3 0.0288737f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A2_c_145_n A3 2.54568e-19 $X=1.915 $Y=1.56 $X2=0 $Y2=0
cc_141 N_A2_c_146_n N_A_28_368#_c_384_n 0.0120121f $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_142 N_A2_M1002_g N_A_28_368#_c_384_n 8.9936e-19 $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A2_c_146_n N_A_28_368#_c_396_n 0.0133349f $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_144 N_A2_M1002_g N_A_28_368#_c_396_n 0.0146602f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_145 A2 N_A_28_368#_c_396_n 0.049118f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A2_c_145_n N_A_28_368#_c_396_n 8.68948e-19 $X=1.915 $Y=1.56 $X2=0 $Y2=0
cc_147 N_A2_c_146_n N_A_28_368#_c_400_n 8.84614e-19 $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_148 A2 N_A_28_368#_c_400_n 0.0235982f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 A2 N_A_28_368#_c_385_n 0.0133874f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A2_c_146_n N_VPWR_c_420_n 6.94422e-19 $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_151 N_A2_c_146_n N_VPWR_c_425_n 0.005209f $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_152 N_A2_M1002_g N_VPWR_c_425_n 0.00333896f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A2_c_146_n N_VPWR_c_419_n 0.00984513f $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_154 N_A2_M1002_g N_VPWR_c_419_n 0.00428489f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A2_M1002_g N_A_310_368#_c_489_n 0.0134366f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A2_M1002_g N_A_310_368#_c_487_n 0.0137576f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A2_c_146_n N_A_310_368#_c_488_n 0.00364522f $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_158 N_A2_M1002_g N_A_310_368#_c_488_n 0.0019608f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_159 A2 N_A_27_74#_c_601_n 0.0023919f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A2_M1012_g N_A_27_74#_c_603_n 0.00348659f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A2_M1012_g N_A_27_74#_c_604_n 0.014989f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A2_M1013_g N_A_27_74#_c_604_n 0.0132249f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_163 A2 N_A_27_74#_c_604_n 0.0511151f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A2_c_145_n N_A_27_74#_c_604_n 0.00401672f $X=1.915 $Y=1.56 $X2=0 $Y2=0
cc_165 N_A2_M1013_g N_A_27_74#_c_605_n 4.39117e-19 $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_166 A2 N_A_27_74#_c_610_n 0.0225421f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 A2 N_A_27_74#_c_611_n 0.0206318f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A2_c_145_n N_A_27_74#_c_611_n 6.80996e-19 $X=1.915 $Y=1.56 $X2=0 $Y2=0
cc_169 N_A2_M1012_g N_VGND_c_682_n 0.00983261f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_M1013_g N_VGND_c_682_n 0.0105836f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1012_g N_VGND_c_685_n 0.00413917f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_M1013_g N_VGND_c_686_n 0.00383152f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_VGND_c_688_n 0.00818158f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A2_M1013_g N_VGND_c_688_n 0.00757998f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A3_M1016_g N_B1_c_261_n 0.0198315f $X=2.845 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A3_c_199_n N_B1_c_263_n 0.0197387f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_177 A3 N_B1_c_263_n 3.30527e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A3_c_199_n N_B1_M1000_g 0.0180942f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_179 N_A3_c_199_n N_B1_c_265_n 0.00581932f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_180 N_A3_c_199_n B1 0.00529037f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_181 N_A3_c_200_n B1 9.24619e-19 $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_182 N_A3_c_205_n B1 0.00199223f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_183 A3 B1 0.029057f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_184 A3 N_B1_c_268_n 9.7564e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A3_c_202_n N_A_28_368#_c_385_n 0.00115119f $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_186 N_A3_c_200_n N_A_28_368#_c_385_n 0.00273636f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_187 N_A3_c_205_n N_VPWR_c_421_n 5.97691e-19 $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_188 N_A3_c_202_n N_VPWR_c_425_n 0.00333926f $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_189 N_A3_c_205_n N_VPWR_c_425_n 0.005209f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_190 N_A3_c_202_n N_VPWR_c_419_n 0.0042782f $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_191 N_A3_c_205_n N_VPWR_c_419_n 0.00983474f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_192 N_A3_c_202_n N_A_310_368#_c_487_n 0.0158247f $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_193 N_A3_c_205_n N_A_310_368#_c_487_n 0.0017347f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_194 N_A3_c_202_n N_Y_c_519_n 0.012931f $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_195 N_A3_c_199_n N_Y_c_519_n 0.001207f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_196 N_A3_c_205_n N_Y_c_519_n 0.0136492f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_197 A3 N_Y_c_519_n 0.0211864f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A3_c_202_n N_Y_c_514_n 6.61291e-19 $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_199 N_A3_c_205_n N_Y_c_514_n 0.011873f $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_200 N_A3_c_202_n N_Y_c_518_n 0.011119f $X=2.99 $Y=1.725 $X2=0 $Y2=0
cc_201 N_A3_c_200_n N_Y_c_518_n 0.0018814f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_202 N_A3_c_205_n N_Y_c_518_n 5.73047e-19 $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_203 A3 N_Y_c_518_n 0.0263952f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A3_c_205_n N_Y_c_529_n 8.71663e-19 $X=3.44 $Y=1.725 $X2=0 $Y2=0
cc_205 N_A3_M1009_g N_A_27_74#_c_605_n 4.73925e-19 $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1009_g N_A_27_74#_c_606_n 0.018337f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_M1016_g N_A_27_74#_c_606_n 0.0132506f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_c_200_n N_A_27_74#_c_606_n 0.00321928f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_209 A3 N_A_27_74#_c_606_n 0.034156f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A3_M1016_g N_A_27_74#_c_607_n 3.97481e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_c_199_n N_A_27_74#_c_608_n 0.00221944f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_212 A3 N_A_27_74#_c_608_n 7.38037e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A3_c_200_n N_A_27_74#_c_612_n 0.00106083f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_214 A3 N_A_27_74#_c_612_n 0.0224275f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_215 N_A3_M1009_g N_VGND_c_682_n 4.69274e-19 $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A3_M1009_g N_VGND_c_683_n 0.00227662f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A3_M1016_g N_VGND_c_683_n 0.0103163f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A3_M1009_g N_VGND_c_686_n 0.00461464f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A3_M1016_g N_VGND_c_687_n 0.00383152f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A3_M1009_g N_VGND_c_688_n 0.00907963f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A3_M1016_g N_VGND_c_688_n 0.00757637f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B1_M1006_g N_C1_M1007_g 0.0110944f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_223 N_B1_c_266_n N_C1_M1004_g 0.00126295f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_224 N_B1_c_265_n N_C1_c_336_n 0.0110944f $X=4.34 $Y=1.68 $X2=0 $Y2=0
cc_225 N_B1_c_266_n N_C1_c_336_n 0.00317238f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_226 B1 N_C1_c_336_n 5.56058e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B1_M1000_g N_VPWR_c_421_n 0.0129315f $X=3.89 $Y=2.4 $X2=0 $Y2=0
cc_228 N_B1_M1006_g N_VPWR_c_421_n 0.0127835f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B1_M1006_g N_VPWR_c_422_n 5.43099e-19 $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_230 N_B1_M1006_g N_VPWR_c_423_n 0.00460063f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_231 N_B1_M1000_g N_VPWR_c_425_n 0.00460063f $X=3.89 $Y=2.4 $X2=0 $Y2=0
cc_232 N_B1_M1000_g N_VPWR_c_419_n 0.00908665f $X=3.89 $Y=2.4 $X2=0 $Y2=0
cc_233 N_B1_M1006_g N_VPWR_c_419_n 0.00908665f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_234 N_B1_c_262_n N_Y_c_519_n 4.87111e-19 $X=3.77 $Y=1.26 $X2=0 $Y2=0
cc_235 N_B1_c_263_n N_Y_c_519_n 5.76785e-19 $X=3.35 $Y=1.26 $X2=0 $Y2=0
cc_236 B1 N_Y_c_519_n 0.00106056f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_237 N_B1_M1000_g N_Y_c_533_n 0.0142562f $X=3.89 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B1_c_265_n N_Y_c_533_n 4.94024e-19 $X=4.34 $Y=1.68 $X2=0 $Y2=0
cc_239 N_B1_M1006_g N_Y_c_533_n 0.0161344f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_240 B1 N_Y_c_533_n 0.0302485f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B1_M1006_g N_Y_c_515_n 3.62369e-19 $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_242 B1 N_Y_c_529_n 0.0189744f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_243 N_B1_M1006_g N_Y_c_539_n 0.00191786f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_244 N_B1_c_264_n Y 0.00117611f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_245 N_B1_c_264_n Y 3.14144e-19 $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_246 N_B1_M1000_g Y 8.8406e-19 $X=3.89 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B1_c_265_n Y 0.00520009f $X=4.34 $Y=1.68 $X2=0 $Y2=0
cc_248 N_B1_M1006_g Y 0.00622411f $X=4.34 $Y=2.4 $X2=0 $Y2=0
cc_249 N_B1_c_266_n Y 0.00415302f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_250 B1 Y 0.031504f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B1_c_268_n Y 6.27941e-19 $X=3.935 $Y=1.515 $X2=0 $Y2=0
cc_252 N_B1_c_261_n N_A_27_74#_c_607_n 0.00944442f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_253 N_B1_c_264_n N_A_27_74#_c_607_n 6.66923e-19 $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_254 N_B1_c_261_n N_A_27_74#_c_608_n 0.011964f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_255 N_B1_c_262_n N_A_27_74#_c_608_n 0.0063964f $X=3.77 $Y=1.26 $X2=0 $Y2=0
cc_256 N_B1_c_264_n N_A_27_74#_c_608_n 0.0129915f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_257 N_B1_c_265_n N_A_27_74#_c_608_n 0.00165823f $X=4.34 $Y=1.68 $X2=0 $Y2=0
cc_258 N_B1_c_266_n N_A_27_74#_c_608_n 0.0058838f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_259 B1 N_A_27_74#_c_608_n 0.0579009f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_260 N_B1_c_261_n N_A_27_74#_c_609_n 5.80141e-19 $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_261 N_B1_c_264_n N_A_27_74#_c_609_n 0.0077283f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_262 N_B1_c_261_n N_A_27_74#_c_612_n 0.0014099f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_263 N_B1_c_261_n N_VGND_c_683_n 5.57463e-19 $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_264 N_B1_c_261_n N_VGND_c_687_n 0.00434272f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_265 N_B1_c_264_n N_VGND_c_687_n 0.00278271f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_266 N_B1_c_261_n N_VGND_c_688_n 0.00822601f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_267 N_B1_c_264_n N_VGND_c_688_n 0.00359661f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_268 N_B1_c_264_n N_A_670_74#_c_748_n 0.0132715f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_269 N_B1_c_261_n N_A_670_74#_c_749_n 0.00220721f $X=3.275 $Y=1.185 $X2=0
+ $Y2=0
cc_270 N_C1_M1007_g N_VPWR_c_421_n 5.41206e-19 $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_271 N_C1_M1007_g N_VPWR_c_422_n 0.0124151f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_272 N_C1_M1010_g N_VPWR_c_422_n 0.002979f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_273 N_C1_M1007_g N_VPWR_c_423_n 0.00460063f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_274 N_C1_M1010_g N_VPWR_c_426_n 0.005209f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_275 N_C1_M1007_g N_VPWR_c_419_n 0.00908665f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_276 N_C1_M1010_g N_VPWR_c_419_n 0.00986059f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_277 N_C1_M1007_g N_Y_c_515_n 3.62369e-19 $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_278 N_C1_M1004_g N_Y_c_510_n 0.0160709f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_279 N_C1_M1011_g N_Y_c_510_n 0.0126386f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_280 C1 N_Y_c_510_n 0.0567145f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_281 N_C1_c_336_n N_Y_c_510_n 0.00951757f $X=5.43 $Y=1.465 $X2=0 $Y2=0
cc_282 N_C1_M1007_g N_Y_c_553_n 0.0165525f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_283 N_C1_M1010_g N_Y_c_553_n 0.012931f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_284 C1 N_Y_c_553_n 0.0265889f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_285 N_C1_c_336_n N_Y_c_553_n 4.37856e-19 $X=5.43 $Y=1.465 $X2=0 $Y2=0
cc_286 N_C1_M1010_g N_Y_c_516_n 8.84614e-19 $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_287 C1 N_Y_c_516_n 0.0266343f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_288 N_C1_c_336_n N_Y_c_516_n 0.00133528f $X=5.43 $Y=1.465 $X2=0 $Y2=0
cc_289 N_C1_M1007_g N_Y_c_517_n 6.74232e-19 $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_290 N_C1_M1010_g N_Y_c_517_n 0.0122988f $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_291 N_C1_M1011_g N_Y_c_511_n 0.00159289f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_292 N_C1_M1007_g N_Y_c_539_n 0.00191786f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_293 N_C1_M1007_g Y 0.00736012f $X=4.79 $Y=2.4 $X2=0 $Y2=0
cc_294 N_C1_M1004_g Y 0.0060753f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_295 N_C1_M1010_g Y 9.18997e-19 $X=5.24 $Y=2.4 $X2=0 $Y2=0
cc_296 C1 Y 0.0349366f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_297 N_C1_c_336_n Y 0.011288f $X=5.43 $Y=1.465 $X2=0 $Y2=0
cc_298 N_C1_M1004_g N_A_27_74#_c_608_n 4.45329e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_299 N_C1_M1004_g N_VGND_c_687_n 0.00278247f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_300 N_C1_M1011_g N_VGND_c_687_n 0.00430908f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_301 N_C1_M1004_g N_VGND_c_688_n 0.00358425f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_302 N_C1_M1011_g N_VGND_c_688_n 0.00820326f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_303 N_C1_M1004_g N_A_670_74#_c_748_n 0.0117594f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_304 N_C1_M1011_g N_A_670_74#_c_748_n 0.00685665f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_305 N_C1_M1004_g N_A_670_74#_c_754_n 0.0100975f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_306 N_C1_M1011_g N_A_670_74#_c_754_n 0.00461693f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_28_368#_c_390_n N_VPWR_M1005_d 0.00333697f $X=1.07 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_308 N_A_28_368#_c_383_n N_VPWR_c_420_n 0.0234083f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_309 N_A_28_368#_c_390_n N_VPWR_c_420_n 0.0149107f $X=1.07 $Y=2.035 $X2=0
+ $Y2=0
cc_310 N_A_28_368#_c_384_n N_VPWR_c_420_n 0.0256025f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_311 N_A_28_368#_c_384_n N_VPWR_c_425_n 0.014549f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_312 N_A_28_368#_c_383_n N_VPWR_c_419_n 0.0119743f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_313 N_A_28_368#_c_384_n N_VPWR_c_419_n 0.0119743f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_314 N_A_28_368#_c_383_n N_VPWR_c_428_n 0.014549f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_315 N_A_28_368#_c_396_n N_A_310_368#_M1001_d 0.00449621f $X=2.12 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_316 N_A_28_368#_c_396_n N_A_310_368#_c_489_n 0.020554f $X=2.12 $Y=2.035 $X2=0
+ $Y2=0
cc_317 N_A_28_368#_M1002_s N_A_310_368#_c_487_n 0.00266942f $X=2.07 $Y=1.84
+ $X2=0 $Y2=0
cc_318 N_A_28_368#_c_385_n N_A_310_368#_c_487_n 0.0184743f $X=2.205 $Y=2.115
+ $X2=0 $Y2=0
cc_319 N_A_28_368#_c_384_n N_A_310_368#_c_488_n 0.00340372f $X=1.235 $Y=2.815
+ $X2=0 $Y2=0
cc_320 N_A_28_368#_c_385_n N_Y_c_518_n 0.0534093f $X=2.205 $Y=2.115 $X2=0 $Y2=0
cc_321 N_VPWR_c_421_n N_A_310_368#_c_487_n 0.00286526f $X=4.115 $Y=2.455 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_425_n N_A_310_368#_c_487_n 0.0891169f $X=3.95 $Y=3.33 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_419_n N_A_310_368#_c_487_n 0.0505934f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_425_n N_A_310_368#_c_488_n 0.0235512f $X=3.95 $Y=3.33 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_419_n N_A_310_368#_c_488_n 0.0126924f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_421_n N_Y_c_514_n 0.0234083f $X=4.115 $Y=2.455 $X2=0 $Y2=0
cc_327 N_VPWR_c_425_n N_Y_c_514_n 0.0109793f $X=3.95 $Y=3.33 $X2=0 $Y2=0
cc_328 N_VPWR_c_419_n N_Y_c_514_n 0.00901959f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_329 N_VPWR_M1000_d N_Y_c_533_n 0.00314376f $X=3.98 $Y=1.84 $X2=0 $Y2=0
cc_330 N_VPWR_c_421_n N_Y_c_533_n 0.0170259f $X=4.115 $Y=2.455 $X2=0 $Y2=0
cc_331 N_VPWR_c_421_n N_Y_c_515_n 0.0233699f $X=4.115 $Y=2.455 $X2=0 $Y2=0
cc_332 N_VPWR_c_422_n N_Y_c_515_n 0.022423f $X=5.015 $Y=2.455 $X2=0 $Y2=0
cc_333 N_VPWR_c_423_n N_Y_c_515_n 0.00749631f $X=4.85 $Y=3.33 $X2=0 $Y2=0
cc_334 N_VPWR_c_419_n N_Y_c_515_n 0.0062048f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_M1007_d N_Y_c_553_n 0.00315967f $X=4.88 $Y=1.84 $X2=0 $Y2=0
cc_336 N_VPWR_c_422_n N_Y_c_553_n 0.0148589f $X=5.015 $Y=2.455 $X2=0 $Y2=0
cc_337 N_VPWR_c_422_n N_Y_c_517_n 0.0234083f $X=5.015 $Y=2.455 $X2=0 $Y2=0
cc_338 N_VPWR_c_426_n N_Y_c_517_n 0.014549f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_c_419_n N_Y_c_517_n 0.0119743f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_340 N_A_310_368#_c_487_n N_Y_M1017_s 0.00266942f $X=3.13 $Y=2.99 $X2=0 $Y2=0
cc_341 N_A_310_368#_M1017_d N_Y_c_519_n 0.00342674f $X=3.08 $Y=1.84 $X2=0 $Y2=0
cc_342 N_A_310_368#_c_507_p N_Y_c_519_n 0.0126919f $X=3.215 $Y=2.455 $X2=0 $Y2=0
cc_343 N_A_310_368#_c_487_n N_Y_c_514_n 0.00316698f $X=3.13 $Y=2.99 $X2=0 $Y2=0
cc_344 N_A_310_368#_c_487_n N_Y_c_518_n 0.0205035f $X=3.13 $Y=2.99 $X2=0 $Y2=0
cc_345 Y N_A_27_74#_c_608_n 0.011013f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_346 Y N_A_27_74#_c_608_n 0.00429194f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_347 Y N_A_27_74#_c_609_n 0.0338529f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_348 N_Y_c_511_n N_VGND_c_687_n 0.011066f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_349 N_Y_c_511_n N_VGND_c_688_n 0.00915947f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_350 N_Y_c_510_n N_A_670_74#_M1004_d 0.00176461f $X=5.395 $Y=1.045 $X2=0 $Y2=0
cc_351 N_Y_M1004_s N_A_670_74#_c_748_n 0.00273752f $X=4.475 $Y=0.37 $X2=0 $Y2=0
cc_352 N_Y_c_510_n N_A_670_74#_c_748_n 0.0032855f $X=5.395 $Y=1.045 $X2=0 $Y2=0
cc_353 N_Y_c_511_n N_A_670_74#_c_748_n 0.00374778f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_354 Y N_A_670_74#_c_748_n 0.0232003f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_355 N_Y_c_510_n N_A_670_74#_c_754_n 0.0168291f $X=5.395 $Y=1.045 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_601_n N_VGND_M1003_s 0.00240242f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_357 N_A_27_74#_c_604_n N_VGND_M1012_d 0.00187091f $X=2.045 $Y=1.095 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_606_n N_VGND_M1009_d 0.00208352f $X=2.975 $Y=1.095 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_600_n N_VGND_c_681_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_601_n N_VGND_c_681_n 0.0202152f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_603_n N_VGND_c_681_n 0.00121634f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_603_n N_VGND_c_682_n 0.0191439f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_604_n N_VGND_c_682_n 0.0172138f $X=2.045 $Y=1.095 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_605_n N_VGND_c_682_n 0.0182902f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_605_n N_VGND_c_683_n 0.00154841f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_606_n N_VGND_c_683_n 0.0177745f $X=2.975 $Y=1.095 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_607_n N_VGND_c_683_n 0.0182902f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_600_n N_VGND_c_684_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_603_n N_VGND_c_685_n 0.011066f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_605_n N_VGND_c_686_n 0.011066f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_607_n N_VGND_c_687_n 0.0109942f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_600_n N_VGND_c_688_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_373 N_A_27_74#_c_603_n N_VGND_c_688_n 0.00915947f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_605_n N_VGND_c_688_n 0.00915947f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_375 N_A_27_74#_c_607_n N_VGND_c_688_n 0.00904371f $X=3.06 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_608_n N_A_670_74#_M1008_d 0.00358162f $X=3.895 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_377 N_A_27_74#_c_608_n N_A_670_74#_c_763_n 0.0245925f $X=3.895 $Y=1.095 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_M1015_s N_A_670_74#_c_748_n 0.00273752f $X=3.92 $Y=0.37 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_c_608_n N_A_670_74#_c_748_n 0.00304353f $X=3.895 $Y=1.095
+ $X2=0 $Y2=0
cc_380 N_A_27_74#_c_609_n N_A_670_74#_c_748_n 0.0203278f $X=4.06 $Y=0.86 $X2=0
+ $Y2=0
cc_381 N_A_27_74#_c_607_n N_A_670_74#_c_749_n 0.00359554f $X=3.06 $Y=0.515 $X2=0
+ $Y2=0
cc_382 N_VGND_c_687_n N_A_670_74#_c_748_n 0.096935f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_688_n N_A_670_74#_c_748_n 0.0548766f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_683_n N_A_670_74#_c_749_n 0.00306547f $X=2.63 $Y=0.595 $X2=0
+ $Y2=0
cc_385 N_VGND_c_687_n N_A_670_74#_c_749_n 0.023391f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_688_n N_A_670_74#_c_749_n 0.0127797f $X=5.52 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o21bai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o21bai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.350000 2.580000 1.950000 ;
        RECT 2.250000 1.950000 3.715000 2.120000 ;
        RECT 3.485000 1.320000 4.055000 1.650000 ;
        RECT 3.485000 1.650000 3.715000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.820000 1.350000 3.235000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.460000 1.350000 0.835000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.812000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.180000 1.865000 2.290000 ;
        RECT 1.530000 2.290000 3.220000 2.460000 ;
        RECT 1.530000 2.460000 1.780000 2.980000 ;
        RECT 1.615000 0.615000 1.865000 1.180000 ;
        RECT 3.050000 2.460000 3.220000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 1.010000 ;
      RECT 0.115000  1.010000 1.360000 1.180000 ;
      RECT 0.115000  1.180000 0.285000 1.950000 ;
      RECT 0.115000  1.950000 0.640000 2.860000 ;
      RECT 0.545000  0.085000 0.875000 0.840000 ;
      RECT 1.005000  1.820000 1.335000 3.245000 ;
      RECT 1.030000  1.180000 1.360000 1.550000 ;
      RECT 1.105000  0.255000 2.365000 0.425000 ;
      RECT 1.105000  0.425000 1.435000 0.840000 ;
      RECT 1.980000  2.650000 2.350000 3.245000 ;
      RECT 2.035000  0.425000 2.365000 1.010000 ;
      RECT 2.035000  1.010000 4.185000 1.150000 ;
      RECT 2.035000  1.150000 3.245000 1.180000 ;
      RECT 2.520000  2.630000 2.850000 2.905000 ;
      RECT 2.520000  2.905000 3.755000 3.075000 ;
      RECT 2.535000  0.085000 2.865000 0.840000 ;
      RECT 3.075000  0.350000 3.245000 0.980000 ;
      RECT 3.075000  0.980000 4.185000 1.010000 ;
      RECT 3.420000  2.290000 3.755000 2.905000 ;
      RECT 3.425000  0.085000 3.755000 0.810000 ;
      RECT 3.935000  0.350000 4.185000 0.980000 ;
      RECT 3.955000  1.820000 4.205000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__o21bai_2

* NGSPICE file created from sky130_fd_sc_ms__o22ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_145_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=2.688e+11p ps=2.72e+06u
M1001 VPWR A1 a_343_368# VPB pshort w=1.12e+06u l=180000u
+  ad=7.616e+11p pd=5.84e+06u as=4.368e+11p ps=3.02e+06u
M1002 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=6.808e+11p ps=6.28e+06u
M1003 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.255e+11p ps=2.63e+06u
M1004 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_145_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_343_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


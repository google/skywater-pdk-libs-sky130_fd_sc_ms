* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR D1 a_239_368# VPB pshort w=1e+06u l=180000u
+  ad=1.9396e+12p pd=1.222e+07u as=7.1e+11p ps=5.42e+06u
M1001 VPWR a_239_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1002 a_239_368# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_54_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.217e+11p pd=4.37e+06u as=7.955e+11p ps=6.59e+06u
M1004 VGND a_239_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1005 a_461_74# C1 a_369_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=2.294e+11p ps=2.1e+06u
M1006 a_155_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND A1 a_54_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_239_368# D1 a_461_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 X a_239_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_239_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_239_368# A2 a_155_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_239_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_369_74# B1 a_54_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

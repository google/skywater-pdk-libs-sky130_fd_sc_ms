* File: sky130_fd_sc_ms__or4b_2.spice
* Created: Fri Aug 28 18:09:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4b_2.pex.spice"
.subckt sky130_fd_sc_ms__or4b_2  VNB VPB D_N A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_D_N_M1010_g N_A_27_368#_M1010_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.109083 AS=0.15675 PD=0.942248 PS=1.67 NRD=18.54 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.5 A=0.0825 P=1.4 MULT=1
MM1005 N_X_M1005_d N_A_190_48#_M1005_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.146767 PD=1.02 PS=1.26775 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.6 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1005_d N_A_190_48#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.164409 PD=1.02 PS=1.26551 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75001 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1004 N_A_190_48#_M1004_d N_A_M1004_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1408 AS=0.142191 PD=1.08 PS=1.09449 NRD=14.988 NRS=8.436 M=1 R=4.26667
+ SA=75001.7 SB=75002 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_A_190_48#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1584 AS=0.1408 PD=1.135 PS=1.08 NRD=17.808 NRS=14.988 M=1 R=4.26667
+ SA=75002.3 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_190_48#_M1002_d N_C_M1002_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.104 AS=0.1584 PD=0.965 PS=1.135 NRD=8.436 NRS=22.488 M=1 R=4.26667
+ SA=75002.9 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A_27_368#_M1011_g N_A_190_48#_M1002_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2272 AS=0.104 PD=1.99 PS=0.965 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_D_N_M1003_g N_A_27_368#_M1003_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1614 AS=0.2352 PD=1.26429 PS=2.24 NRD=32.1504 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003.2 A=0.1512 P=2.04 MULT=1
MM1009 N_X_M1009_d N_A_190_48#_M1009_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2152 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1009_d N_A_190_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.287925 PD=1.39 PS=1.72755 NRD=0 NRS=20.2122 M=1 R=6.22222
+ SA=90001 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1000 A_455_392# N_A_M1000_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.257075 PD=1.24 PS=1.54245 NRD=12.7853 NRS=23.6203 M=1 R=5.55556
+ SA=90001.7 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1007 A_539_392# N_B_M1007_g A_455_392# VPB PSHORT L=0.18 W=1 AD=0.165 AS=0.12
+ PD=1.33 PS=1.24 NRD=21.6503 NRS=12.7853 M=1 R=5.55556 SA=90002.1 SB=90001.4
+ A=0.18 P=2.36 MULT=1
MM1001 A_641_392# N_C_M1001_g A_539_392# VPB PSHORT L=0.18 W=1 AD=0.18 AS=0.165
+ PD=1.36 PS=1.33 NRD=24.6053 NRS=21.6503 M=1 R=5.55556 SA=90002.7 SB=90000.9
+ A=0.18 P=2.36 MULT=1
MM1006 N_A_190_48#_M1006_d N_A_27_368#_M1006_g A_641_392# VPB PSHORT L=0.18 W=1
+ AD=0.43 AS=0.18 PD=2.86 PS=1.36 NRD=28.5453 NRS=24.6053 M=1 R=5.55556
+ SA=90003.2 SB=90000.3 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_53 VNB 0 1.7764e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__or4b_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a41o_2.pxi.spice
* Created: Fri Aug 28 17:09:33 2020
* 
x_PM_SKY130_FD_SC_MS__A41O_2%A4 N_A4_M1002_g N_A4_c_82_n N_A4_M1005_g A4
+ N_A4_c_84_n PM_SKY130_FD_SC_MS__A41O_2%A4
x_PM_SKY130_FD_SC_MS__A41O_2%A3 N_A3_M1004_g N_A3_M1008_g A3 A3 A3 N_A3_c_110_n
+ N_A3_c_111_n PM_SKY130_FD_SC_MS__A41O_2%A3
x_PM_SKY130_FD_SC_MS__A41O_2%A2 N_A2_M1006_g N_A2_M1010_g A2 A2 A2 N_A2_c_146_n
+ N_A2_c_147_n PM_SKY130_FD_SC_MS__A41O_2%A2
x_PM_SKY130_FD_SC_MS__A41O_2%A1 N_A1_M1007_g N_A1_M1013_g A1 N_A1_c_182_n
+ PM_SKY130_FD_SC_MS__A41O_2%A1
x_PM_SKY130_FD_SC_MS__A41O_2%B1 N_B1_M1003_g N_B1_M1001_g B1 N_B1_c_221_n
+ N_B1_c_222_n PM_SKY130_FD_SC_MS__A41O_2%B1
x_PM_SKY130_FD_SC_MS__A41O_2%A_441_74# N_A_441_74#_M1007_d N_A_441_74#_M1001_d
+ N_A_441_74#_c_257_n N_A_441_74#_M1009_g N_A_441_74#_M1000_g
+ N_A_441_74#_c_259_n N_A_441_74#_M1012_g N_A_441_74#_M1011_g
+ N_A_441_74#_c_261_n N_A_441_74#_c_262_n N_A_441_74#_c_263_n
+ N_A_441_74#_c_264_n N_A_441_74#_c_265_n N_A_441_74#_c_266_n
+ N_A_441_74#_c_272_n N_A_441_74#_c_267_n N_A_441_74#_c_273_n
+ N_A_441_74#_c_268_n N_A_441_74#_c_269_n PM_SKY130_FD_SC_MS__A41O_2%A_441_74#
x_PM_SKY130_FD_SC_MS__A41O_2%A_27_392# N_A_27_392#_M1002_s N_A_27_392#_M1008_d
+ N_A_27_392#_M1013_d N_A_27_392#_c_341_n N_A_27_392#_c_342_n
+ N_A_27_392#_c_343_n N_A_27_392#_c_344_n N_A_27_392#_c_345_n
+ N_A_27_392#_c_346_n N_A_27_392#_c_347_n N_A_27_392#_c_348_n
+ PM_SKY130_FD_SC_MS__A41O_2%A_27_392#
x_PM_SKY130_FD_SC_MS__A41O_2%VPWR N_VPWR_M1002_d N_VPWR_M1010_d N_VPWR_M1000_d
+ N_VPWR_M1011_d N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n
+ N_VPWR_c_403_n N_VPWR_c_404_n VPWR N_VPWR_c_405_n N_VPWR_c_406_n
+ N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_398_n
+ PM_SKY130_FD_SC_MS__A41O_2%VPWR
x_PM_SKY130_FD_SC_MS__A41O_2%X N_X_M1009_d N_X_M1000_s N_X_c_458_n N_X_c_455_n
+ N_X_c_456_n N_X_c_468_n N_X_c_453_n X PM_SKY130_FD_SC_MS__A41O_2%X
x_PM_SKY130_FD_SC_MS__A41O_2%VGND N_VGND_M1005_s N_VGND_M1003_d N_VGND_M1012_s
+ N_VGND_c_489_n N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n
+ VGND N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n
+ PM_SKY130_FD_SC_MS__A41O_2%VGND
cc_1 VNB N_A4_M1002_g 0.00976783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_2 VNB N_A4_c_82_n 0.0207173f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.22
cc_3 VNB A4 0.0082382f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A4_c_84_n 0.0581619f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_5 VNB N_A3_M1008_g 0.00659705f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_6 VNB A3 0.00532111f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_A3_c_110_n 0.0306953f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_8 VNB N_A3_c_111_n 0.0181058f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_9 VNB N_A2_M1010_g 0.00678988f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_10 VNB A2 0.0038768f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A2_c_146_n 0.0391047f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.385
cc_12 VNB N_A2_c_147_n 0.0200799f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_13 VNB N_A1_M1007_g 0.0334159f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_14 VNB A1 0.00316184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_182_n 0.0205628f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_16 VNB N_B1_M1003_g 0.0325672f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_17 VNB N_B1_c_221_n 0.0185267f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_18 VNB N_B1_c_222_n 0.00357093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_441_74#_c_257_n 0.0187608f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_20 VNB N_A_441_74#_M1000_g 0.00691622f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_21 VNB N_A_441_74#_c_259_n 0.0197849f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_22 VNB N_A_441_74#_M1011_g 0.00871317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_441_74#_c_261_n 0.0165285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_441_74#_c_262_n 0.0397326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_441_74#_c_263_n 0.0565216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_441_74#_c_264_n 0.0033626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_441_74#_c_265_n 0.00990139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_441_74#_c_266_n 0.0065138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_441_74#_c_267_n 0.00557865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_441_74#_c_268_n 0.00197732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_441_74#_c_269_n 0.00285482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_398_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_453_n 0.00545204f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_34 VNB X 0.00329372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_489_n 0.0131437f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_36 VNB N_VGND_c_490_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_37 VNB N_VGND_c_491_n 0.00985577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_492_n 0.0655012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_493_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_40 VNB N_VGND_c_494_n 0.0217179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_495_n 0.0492105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_496_n 0.292499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A4_M1002_g 0.0383644f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_44 VPB N_A3_M1008_g 0.0294155f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_45 VPB N_A2_M1010_g 0.0321404f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_46 VPB N_A1_M1013_g 0.0259847f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_47 VPB A1 0.00137218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A1_c_182_n 0.0135374f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_49 VPB N_B1_M1001_g 0.025876f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_50 VPB N_B1_c_221_n 0.0131725f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_51 VPB N_B1_c_222_n 0.0024806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_441_74#_M1000_g 0.0248893f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_53 VPB N_A_441_74#_M1011_g 0.0273944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_441_74#_c_272_n 0.011878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_441_74#_c_273_n 0.0120258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_441_74#_c_268_n 0.00720913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_392#_c_341_n 0.0442448f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_58 VPB N_A_27_392#_c_342_n 0.0135978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_27_392#_c_343_n 0.00985309f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.295
cc_60 VPB N_A_27_392#_c_344_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_61 VPB N_A_27_392#_c_345_n 0.010042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_392#_c_346_n 0.00379931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_392#_c_347_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_392#_c_348_n 0.00560004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_399_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.385
cc_66 VPB N_VPWR_c_400_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_401_n 0.0109541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_402_n 0.0166496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_403_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_404_n 0.0695565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_405_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_406_n 0.0339528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_407_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_408_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_409_n 0.00978383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_410_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_398_n 0.0717866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_X_c_455_n 0.00415743f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_79 VPB N_X_c_456_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_X_c_453_n 0.00148895f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_81 N_A4_M1002_g N_A3_M1008_g 0.0174197f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_82 N_A4_c_82_n A3 0.00462195f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_83 A4 A3 0.0147682f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_84 A4 N_A3_c_110_n 9.67587e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A4_c_84_n N_A3_c_110_n 0.033243f $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_86 N_A4_c_82_n N_A3_c_111_n 0.033243f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_87 N_A4_M1002_g N_A_27_392#_c_341_n 0.0160655f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_88 N_A4_M1002_g N_A_27_392#_c_342_n 0.0177353f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_89 A4 N_A_27_392#_c_342_n 6.17992e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A4_c_84_n N_A_27_392#_c_342_n 4.15062e-19 $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_91 N_A4_M1002_g N_A_27_392#_c_343_n 0.0043353f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_92 A4 N_A_27_392#_c_343_n 0.0271109f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A4_c_84_n N_A_27_392#_c_343_n 0.00228736f $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_94 N_A4_M1002_g N_A_27_392#_c_348_n 5.60475e-19 $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_95 N_A4_M1002_g N_VPWR_c_399_n 0.00343717f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_96 N_A4_M1002_g N_VPWR_c_405_n 0.005209f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_97 N_A4_M1002_g N_VPWR_c_398_n 0.00986318f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_98 N_A4_c_82_n N_VGND_c_490_n 0.0159948f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_99 A4 N_VGND_c_490_n 0.0241219f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A4_c_84_n N_VGND_c_490_n 0.00199143f $X=0.53 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A4_c_82_n N_VGND_c_492_n 0.00383152f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A4_c_82_n N_VGND_c_496_n 0.0075725f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A3_M1008_g N_A2_M1010_g 0.0263684f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_104 A3 A2 0.0892488f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A3_c_110_n A2 2.90162e-19 $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A3_c_111_n A2 5.869e-19 $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A3_c_110_n N_A2_c_146_n 0.0174537f $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_108 A3 N_A2_c_147_n 0.00916629f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A3_c_111_n N_A2_c_147_n 0.0245047f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_110 N_A3_M1008_g N_A_27_392#_c_341_n 4.81978e-19 $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_111 N_A3_M1008_g N_A_27_392#_c_342_n 0.0139943f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_112 A3 N_A_27_392#_c_342_n 0.0209363f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_113 N_A3_c_110_n N_A_27_392#_c_342_n 8.27684e-19 $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_114 N_A3_M1008_g N_A_27_392#_c_344_n 0.0102485f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_115 N_A3_M1008_g N_A_27_392#_c_348_n 0.00840213f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_116 A3 N_A_27_392#_c_348_n 0.0181535f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A3_c_110_n N_A_27_392#_c_348_n 2.37442e-19 $X=1.01 $Y=1.385 $X2=0 $Y2=0
cc_118 N_A3_M1008_g N_VPWR_c_399_n 0.00203999f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_119 N_A3_M1008_g N_VPWR_c_400_n 0.005209f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_120 N_A3_M1008_g N_VPWR_c_398_n 0.00982687f $X=1.055 $Y=2.46 $X2=0 $Y2=0
cc_121 A3 N_VGND_c_490_n 0.0237984f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A3_c_111_n N_VGND_c_490_n 0.00251629f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_123 A3 N_VGND_c_492_n 0.0137277f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 N_A3_c_111_n N_VGND_c_492_n 0.00304348f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_125 A3 N_VGND_c_496_n 0.0155751f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_126 N_A3_c_111_n N_VGND_c_496_n 0.00371612f $X=1.01 $Y=1.22 $X2=0 $Y2=0
cc_127 A3 A_199_74# 0.0136602f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_128 A2 N_A1_M1007_g 0.00887723f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_129 N_A2_c_146_n N_A1_M1007_g 0.0127399f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_130 N_A2_c_147_n N_A1_M1007_g 0.0197473f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A2_M1010_g N_A1_M1013_g 0.0223977f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_132 N_A2_M1010_g A1 0.0012121f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_133 A2 A1 0.00633735f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 N_A2_c_146_n A1 3.61063e-19 $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A2_M1010_g N_A1_c_182_n 0.00678722f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_136 A2 N_A1_c_182_n 3.48291e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A2_c_146_n N_A1_c_182_n 0.006184f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_138 A2 N_A_441_74#_c_266_n 0.00778382f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A2_M1010_g N_A_27_392#_c_344_n 0.016064f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_140 N_A2_M1010_g N_A_27_392#_c_345_n 0.0168178f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_141 A2 N_A_27_392#_c_345_n 0.0133431f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_142 N_A2_c_146_n N_A_27_392#_c_345_n 0.00127627f $X=1.65 $Y=1.385 $X2=0 $Y2=0
cc_143 N_A2_M1010_g N_A_27_392#_c_348_n 0.0139552f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_144 N_A2_M1010_g N_VPWR_c_400_n 0.005209f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_145 N_A2_M1010_g N_VPWR_c_401_n 0.00799135f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_146 N_A2_M1010_g N_VPWR_c_398_n 0.00983908f $X=1.505 $Y=2.46 $X2=0 $Y2=0
cc_147 A2 N_VGND_c_492_n 0.0094108f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A2_c_147_n N_VGND_c_492_n 0.00378161f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_149 A2 N_VGND_c_496_n 0.0110426f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A2_c_147_n N_VGND_c_496_n 0.00629143f $X=1.615 $Y=1.22 $X2=0 $Y2=0
cc_151 A2 A_313_74# 0.0135149f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_152 N_A1_M1007_g N_B1_M1003_g 0.0231835f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1013_g N_B1_M1001_g 0.0159878f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_154 A1 N_B1_c_221_n 3.62235e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A1_c_182_n N_B1_c_221_n 0.0174106f $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_156 A1 N_B1_c_222_n 0.0264884f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A1_c_182_n N_B1_c_222_n 0.00201746f $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_158 N_A1_M1007_g N_A_441_74#_c_264_n 9.25648e-19 $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A1_M1007_g N_A_441_74#_c_266_n 0.00253341f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_160 A1 N_A_441_74#_c_266_n 0.0105084f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A1_c_182_n N_A_441_74#_c_266_n 9.72452e-19 $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_162 N_A1_M1013_g N_A_27_392#_c_345_n 0.0140979f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_163 A1 N_A_27_392#_c_345_n 0.0197217f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A1_c_182_n N_A_27_392#_c_345_n 8.30414e-19 $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_165 N_A1_M1013_g N_A_27_392#_c_346_n 0.00100081f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_166 A1 N_A_27_392#_c_346_n 0.00486484f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A1_c_182_n N_A_27_392#_c_346_n 2.29527e-19 $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_168 N_A1_M1013_g N_A_27_392#_c_347_n 0.016064f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_169 A1 N_A_27_392#_c_348_n 0.00163617f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_c_182_n N_A_27_392#_c_348_n 2.03256e-19 $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_171 N_A1_M1013_g N_VPWR_c_401_n 0.00953257f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_172 N_A1_M1013_g N_VPWR_c_406_n 0.005209f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_173 N_A1_M1013_g N_VPWR_c_398_n 0.00983908f $X=2.235 $Y=2.46 $X2=0 $Y2=0
cc_174 N_A1_M1007_g N_VGND_c_492_n 0.00461464f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_M1007_g N_VGND_c_496_n 0.00912075f $X=2.13 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B1_M1003_g N_A_441_74#_c_257_n 0.0260862f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B1_c_221_n N_A_441_74#_c_261_n 0.00525612f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_178 N_B1_M1003_g N_A_441_74#_c_264_n 0.00451422f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B1_M1003_g N_A_441_74#_c_265_n 0.0160524f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_c_221_n N_A_441_74#_c_265_n 0.0041539f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_181 N_B1_c_222_n N_A_441_74#_c_265_n 0.0269774f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_182 N_B1_c_222_n N_A_441_74#_c_266_n 0.00309615f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_183 N_B1_M1001_g N_A_441_74#_c_273_n 7.22795e-19 $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_184 N_B1_c_221_n N_A_441_74#_c_273_n 0.00300514f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_185 N_B1_c_222_n N_A_441_74#_c_273_n 0.010879f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_186 N_B1_M1001_g N_A_441_74#_c_268_n 0.00503397f $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_187 N_B1_c_221_n N_A_441_74#_c_268_n 0.00161215f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_188 N_B1_c_222_n N_A_441_74#_c_268_n 0.0175146f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_189 N_B1_M1003_g N_A_441_74#_c_269_n 0.00398645f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B1_c_221_n N_A_441_74#_c_269_n 3.86402e-19 $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_191 N_B1_c_222_n N_A_441_74#_c_269_n 0.00850124f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_192 N_B1_M1001_g N_A_27_392#_c_346_n 0.00254175f $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_193 N_B1_c_222_n N_A_27_392#_c_346_n 0.00858705f $X=2.76 $Y=1.615 $X2=0 $Y2=0
cc_194 N_B1_M1001_g N_A_27_392#_c_347_n 0.0105904f $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_195 N_B1_M1001_g N_VPWR_c_402_n 0.00380477f $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_196 N_B1_M1001_g N_VPWR_c_406_n 0.005209f $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_197 N_B1_M1001_g N_VPWR_c_398_n 0.00988607f $X=2.685 $Y=2.46 $X2=0 $Y2=0
cc_198 N_B1_M1003_g N_VGND_c_491_n 0.00693601f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_199 N_B1_M1003_g N_VGND_c_492_n 0.00461464f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B1_M1003_g N_VGND_c_496_n 0.00910461f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_441_74#_c_266_n N_A_27_392#_c_346_n 0.00610935f $X=2.56 $Y=1.195
+ $X2=0 $Y2=0
cc_202 N_A_441_74#_c_273_n N_A_27_392#_c_346_n 0.00755776f $X=2.96 $Y=2.115
+ $X2=0 $Y2=0
cc_203 N_A_441_74#_c_272_n N_A_27_392#_c_347_n 0.0330222f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_204 N_A_441_74#_M1000_g N_VPWR_c_402_n 0.00488246f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_205 N_A_441_74#_c_272_n N_VPWR_c_402_n 0.0478677f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_206 N_A_441_74#_M1011_g N_VPWR_c_404_n 0.00546761f $X=4.245 $Y=2.4 $X2=0
+ $Y2=0
cc_207 N_A_441_74#_c_272_n N_VPWR_c_406_n 0.0146357f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_208 N_A_441_74#_M1000_g N_VPWR_c_407_n 0.005209f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_441_74#_M1011_g N_VPWR_c_407_n 0.005209f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_441_74#_M1000_g N_VPWR_c_398_n 0.00986727f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_441_74#_M1011_g N_VPWR_c_398_n 0.00985497f $X=4.245 $Y=2.4 $X2=0
+ $Y2=0
cc_212 N_A_441_74#_c_272_n N_VPWR_c_398_n 0.0121141f $X=2.96 $Y=2.815 $X2=0
+ $Y2=0
cc_213 N_A_441_74#_c_259_n N_X_c_458_n 0.0122008f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A_441_74#_c_263_n N_X_c_458_n 0.00376241f $X=4.245 $Y=1.385 $X2=0 $Y2=0
cc_215 N_A_441_74#_c_267_n N_X_c_458_n 0.0088769f $X=3.68 $Y=1.385 $X2=0 $Y2=0
cc_216 N_A_441_74#_M1000_g N_X_c_455_n 0.00532455f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A_441_74#_M1011_g N_X_c_455_n 0.00215936f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_441_74#_c_263_n N_X_c_455_n 0.00159703f $X=4.245 $Y=1.385 $X2=0 $Y2=0
cc_219 N_A_441_74#_c_268_n N_X_c_455_n 0.00459591f $X=3.03 $Y=1.95 $X2=0 $Y2=0
cc_220 N_A_441_74#_M1000_g N_X_c_456_n 0.0189694f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A_441_74#_M1011_g N_X_c_456_n 0.0127634f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_441_74#_c_273_n N_X_c_456_n 0.00459591f $X=2.96 $Y=2.115 $X2=0 $Y2=0
cc_223 N_A_441_74#_c_257_n N_X_c_468_n 0.00195381f $X=3.25 $Y=1.22 $X2=0 $Y2=0
cc_224 N_A_441_74#_c_262_n N_X_c_468_n 0.00136132f $X=3.705 $Y=1.385 $X2=0 $Y2=0
cc_225 N_A_441_74#_c_267_n N_X_c_468_n 0.0272424f $X=3.68 $Y=1.385 $X2=0 $Y2=0
cc_226 N_A_441_74#_M1000_g N_X_c_453_n 0.00585219f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_441_74#_c_259_n N_X_c_453_n 0.00825937f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_228 N_A_441_74#_M1011_g N_X_c_453_n 0.0128774f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A_441_74#_c_263_n N_X_c_453_n 0.0272944f $X=4.245 $Y=1.385 $X2=0 $Y2=0
cc_230 N_A_441_74#_c_267_n N_X_c_453_n 0.0337299f $X=3.68 $Y=1.385 $X2=0 $Y2=0
cc_231 N_A_441_74#_c_257_n X 0.0044265f $X=3.25 $Y=1.22 $X2=0 $Y2=0
cc_232 N_A_441_74#_c_269_n N_VGND_M1003_d 0.00279178f $X=3.18 $Y=1.33 $X2=0
+ $Y2=0
cc_233 N_A_441_74#_c_257_n N_VGND_c_491_n 0.00683054f $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_234 N_A_441_74#_c_264_n N_VGND_c_491_n 0.00127913f $X=2.395 $Y=0.515 $X2=0
+ $Y2=0
cc_235 N_A_441_74#_c_265_n N_VGND_c_491_n 0.0246062f $X=3.095 $Y=1.195 $X2=0
+ $Y2=0
cc_236 N_A_441_74#_c_269_n N_VGND_c_491_n 0.0021188f $X=3.18 $Y=1.33 $X2=0 $Y2=0
cc_237 N_A_441_74#_c_264_n N_VGND_c_492_n 0.0146357f $X=2.395 $Y=0.515 $X2=0
+ $Y2=0
cc_238 N_A_441_74#_c_257_n N_VGND_c_494_n 0.00461464f $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_239 N_A_441_74#_c_259_n N_VGND_c_494_n 0.00460063f $X=3.81 $Y=1.22 $X2=0
+ $Y2=0
cc_240 N_A_441_74#_c_257_n N_VGND_c_495_n 4.95096e-19 $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_241 N_A_441_74#_c_259_n N_VGND_c_495_n 0.00590656f $X=3.81 $Y=1.22 $X2=0
+ $Y2=0
cc_242 N_A_441_74#_c_263_n N_VGND_c_495_n 0.00518943f $X=4.245 $Y=1.385 $X2=0
+ $Y2=0
cc_243 N_A_441_74#_c_257_n N_VGND_c_496_n 0.00910813f $X=3.25 $Y=1.22 $X2=0
+ $Y2=0
cc_244 N_A_441_74#_c_259_n N_VGND_c_496_n 0.00442948f $X=3.81 $Y=1.22 $X2=0
+ $Y2=0
cc_245 N_A_441_74#_c_264_n N_VGND_c_496_n 0.0121141f $X=2.395 $Y=0.515 $X2=0
+ $Y2=0
cc_246 N_A_27_392#_c_345_n N_VPWR_M1010_d 0.0063069f $X=2.295 $Y=2.035 $X2=0
+ $Y2=0
cc_247 N_A_27_392#_c_341_n N_VPWR_c_399_n 0.0353111f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_248 N_A_27_392#_c_342_n N_VPWR_c_399_n 0.0238907f $X=1.115 $Y=1.805 $X2=0
+ $Y2=0
cc_249 N_A_27_392#_c_348_n N_VPWR_c_399_n 0.0352735f $X=1.28 $Y=1.805 $X2=0
+ $Y2=0
cc_250 N_A_27_392#_c_344_n N_VPWR_c_400_n 0.0144623f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_27_392#_c_344_n N_VPWR_c_401_n 0.0267347f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_252 N_A_27_392#_c_345_n N_VPWR_c_401_n 0.0354723f $X=2.295 $Y=2.035 $X2=0
+ $Y2=0
cc_253 N_A_27_392#_c_347_n N_VPWR_c_401_n 0.0267347f $X=2.46 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_A_27_392#_c_341_n N_VPWR_c_405_n 0.014549f $X=0.28 $Y=2.105 $X2=0 $Y2=0
cc_255 N_A_27_392#_c_347_n N_VPWR_c_406_n 0.0144623f $X=2.46 $Y=2.815 $X2=0
+ $Y2=0
cc_256 N_A_27_392#_c_341_n N_VPWR_c_398_n 0.0119743f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_257 N_A_27_392#_c_344_n N_VPWR_c_398_n 0.0118344f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_258 N_A_27_392#_c_347_n N_VPWR_c_398_n 0.0118344f $X=2.46 $Y=2.815 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_404_n N_X_c_455_n 0.0450694f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_260 N_VPWR_c_402_n N_X_c_456_n 0.0274314f $X=3.52 $Y=2.38 $X2=0 $Y2=0
cc_261 N_VPWR_c_407_n N_X_c_456_n 0.0144623f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_c_398_n N_X_c_456_n 0.0118344f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_263 N_X_c_458_n N_VGND_M1012_s 0.0123021f $X=4.015 $Y=0.855 $X2=0 $Y2=0
cc_264 N_X_c_453_n N_VGND_M1012_s 0.00901369f $X=4.02 $Y=1.82 $X2=0 $Y2=0
cc_265 X N_VGND_c_491_n 0.0127255f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_266 X N_VGND_c_494_n 0.0144853f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_267 N_X_c_458_n N_VGND_c_495_n 0.0205938f $X=4.015 $Y=0.855 $X2=0 $Y2=0
cc_268 X N_VGND_c_495_n 0.0123663f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_269 N_X_c_458_n N_VGND_c_496_n 0.00626145f $X=4.015 $Y=0.855 $X2=0 $Y2=0
cc_270 X N_VGND_c_496_n 0.0120561f $X=3.515 $Y=0.47 $X2=0 $Y2=0

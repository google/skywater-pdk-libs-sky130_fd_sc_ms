* File: sky130_fd_sc_ms__dlclkp_4.spice
* Created: Fri Aug 28 17:26:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlclkp_4.pex.spice"
.subckt sky130_fd_sc_ms__dlclkp_4  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_A_84_48#_M1020_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.258437 AS=0.2109 PD=1.55507 PS=2.05 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1017 A_286_80# N_GATE_M1017_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.223513 PD=0.88 PS=1.34493 NRD=12.18 NRS=75.936 M=1 R=4.26667
+ SA=75001.1 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_84_48#_M1018_d N_A_334_54#_M1018_g A_286_80# VNB NLOWVT L=0.15 W=0.64
+ AD=0.156196 AS=0.0768 PD=1.35849 PS=0.88 NRD=18.744 NRS=12.18 M=1 R=4.26667
+ SA=75001.5 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1011 A_491_124# N_A_334_338#_M1011_g N_A_84_48#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.118875 AS=0.102504 PD=1.195 PS=0.891509 NRD=65.148 NRS=30 M=1
+ R=2.8 SA=75002.1 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_27_74#_M1001_g A_491_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.11894 AS=0.118875 PD=0.945 PS=1.195 NRD=65.196 NRS=65.148 M=1 R=2.8
+ SA=75000.8 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1025 N_A_334_338#_M1025_d N_A_334_54#_M1025_g N_VGND_M1001_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2675 AS=0.20956 PD=2.66 PS=1.665 NRD=49.692 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_CLK_M1019_g N_A_334_54#_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2333 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1005 A_1047_74# N_CLK_M1005_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1036 PD=0.98 PS=1.02 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1021 N_A_1047_368#_M1021_d N_A_27_74#_M1021_g A_1047_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_GCLK_M1006_d N_A_1047_368#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2977 PD=1.02 PS=2.9 NRD=0 NRS=56.316 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 N_GCLK_M1006_d N_A_1047_368#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1013 N_GCLK_M1013_d N_A_1047_368#_M1013_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_GCLK_M1013_d N_A_1047_368#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_84_48#_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.311698 AS=0.3136 PD=1.77509 PS=2.8 NRD=23.7385 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1023 A_286_392# N_GATE_M1023_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.278302 PD=1.24 PS=1.58491 NRD=12.7853 NRS=28.565 M=1 R=5.55556 SA=90000.9
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1000 N_A_84_48#_M1000_d N_A_334_338#_M1000_g A_286_392# VPB PSHORT L=0.18 W=1
+ AD=0.281056 AS=0.12 PD=2.26056 PS=1.24 NRD=31.5003 NRS=12.7853 M=1 R=5.55556
+ SA=90001.3 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1024 A_527_508# N_A_334_54#_M1024_g N_A_84_48#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.118044 PD=0.66 PS=0.949437 NRD=30.4759 NRS=77.3816 M=1
+ R=2.33333 SA=90002.1 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_27_74#_M1002_g A_527_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1169 AS=0.0504 PD=0.993333 PS=0.66 NRD=39.8531 NRS=30.4759 M=1 R=2.33333
+ SA=90002.6 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1015 N_A_334_338#_M1015_d N_A_334_54#_M1015_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2338 PD=2.24 PS=1.98667 NRD=0 NRS=52.3626 M=1 R=4.66667
+ SA=90001.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_334_54#_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1686 AS=0.2352 PD=1.27714 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003.7 A=0.1512 P=2.04 MULT=1
MM1008 N_A_1047_368#_M1008_d N_CLK_M1008_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1708 AS=0.2248 PD=1.425 PS=1.70286 NRD=5.2599 NRS=1.7533 M=1
+ R=6.22222 SA=90000.6 SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_27_74#_M1014_g N_A_1047_368#_M1008_d VPB PSHORT L=0.18
+ W=1.12 AD=0.518 AS=0.1708 PD=2.045 PS=1.425 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1004 N_GCLK_M1004_d N_A_1047_368#_M1004_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1596 AS=0.518 PD=1.405 PS=2.045 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.2 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1007 N_GCLK_M1004_d N_A_1047_368#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1596 AS=0.1708 PD=1.405 PS=1.425 NRD=1.7533 NRS=5.2599 M=1
+ R=6.22222 SA=90002.7 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1010 N_GCLK_M1010_d N_A_1047_368#_M1010_g N_VPWR_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1708 PD=1.39 PS=1.425 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.1 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1022 N_GCLK_M1010_d N_A_1047_368#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX26_noxref VNB VPB NWDIODE A=16.3897 P=22.3
*
.include "sky130_fd_sc_ms__dlclkp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__clkinv_2.pxi.spice
* Created: Fri Aug 28 17:19:55 2020
* 
x_PM_SKY130_FD_SC_MS__CLKINV_2%A N_A_M1002_g N_A_M1000_g N_A_M1001_g N_A_M1003_g
+ N_A_M1004_g A A A N_A_c_34_n PM_SKY130_FD_SC_MS__CLKINV_2%A
x_PM_SKY130_FD_SC_MS__CLKINV_2%Y N_Y_M1002_s N_Y_M1000_s N_Y_M1001_s N_Y_c_82_n
+ N_Y_c_83_n N_Y_c_91_n N_Y_c_84_n N_Y_c_79_n N_Y_c_85_n N_Y_c_80_n N_Y_c_104_n
+ Y PM_SKY130_FD_SC_MS__CLKINV_2%Y
x_PM_SKY130_FD_SC_MS__CLKINV_2%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_c_128_n
+ N_VPWR_c_129_n N_VPWR_c_130_n VPWR N_VPWR_c_131_n N_VPWR_c_132_n
+ N_VPWR_c_127_n PM_SKY130_FD_SC_MS__CLKINV_2%VPWR
x_PM_SKY130_FD_SC_MS__CLKINV_2%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_c_155_n
+ N_VGND_c_156_n N_VGND_c_157_n N_VGND_c_158_n VGND N_VGND_c_159_n
+ N_VGND_c_160_n PM_SKY130_FD_SC_MS__CLKINV_2%VGND
cc_1 VNB N_A_M1002_g 0.0644232f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.61
cc_2 VNB N_A_M1004_g 0.0581471f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.61
cc_3 VNB A 0.0183006f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_A_c_34_n 0.0674526f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_5 VNB N_Y_c_79_n 0.0153843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_Y_c_80_n 0.0174246f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_7 VNB Y 0.0240108f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.515
cc_8 VNB N_VPWR_c_127_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_9 VNB N_VGND_c_155_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_10 VNB N_VGND_c_156_n 0.0338694f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.68
cc_11 VNB N_VGND_c_157_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_12 VNB N_VGND_c_158_n 0.0321896f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.68
cc_13 VNB N_VGND_c_159_n 0.0287859f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.35
cc_14 VNB N_VGND_c_160_n 0.143782f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_15 VPB N_A_M1000_g 0.027583f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_16 VPB N_A_M1001_g 0.0204961f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_17 VPB N_A_M1003_g 0.0227485f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_18 VPB A 0.0137513f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_19 VPB N_A_c_34_n 0.00850978f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.515
cc_20 VPB N_Y_c_82_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_21 VPB N_Y_c_83_n 0.0352219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_22 VPB N_Y_c_84_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.61
cc_23 VPB N_Y_c_85_n 0.00714919f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_24 VPB Y 0.0129485f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.515
cc_25 VPB N_VPWR_c_128_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_26 VPB N_VPWR_c_129_n 0.0108116f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.68
cc_27 VPB N_VPWR_c_130_n 0.0370432f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_28 VPB N_VPWR_c_131_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.61
cc_29 VPB N_VPWR_c_132_n 0.0234893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_127_n 0.0559442f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.515
cc_31 N_A_M1000_g N_Y_c_82_n 8.84614e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_32 A N_Y_c_82_n 0.0259449f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_33 N_A_M1000_g N_Y_c_83_n 0.0121004f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_34 N_A_M1001_g N_Y_c_83_n 6.50516e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_35 N_A_M1000_g N_Y_c_91_n 0.012931f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_36 N_A_M1001_g N_Y_c_91_n 0.012931f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_37 A N_Y_c_91_n 0.0391869f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_38 N_A_c_34_n N_Y_c_91_n 4.90767e-19 $X=1.425 $Y=1.515 $X2=0 $Y2=0
cc_39 N_A_M1000_g N_Y_c_84_n 6.50516e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_40 N_A_M1001_g N_Y_c_84_n 0.0119382f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_41 N_A_M1003_g N_Y_c_84_n 0.0166062f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_42 N_A_M1004_g N_Y_c_79_n 0.0223231f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_43 N_A_M1003_g N_Y_c_85_n 0.0189057f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_44 N_A_M1002_g N_Y_c_80_n 0.0223806f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_45 N_A_M1004_g N_Y_c_80_n 0.0144176f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_46 A N_Y_c_80_n 0.0596487f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_c_34_n N_Y_c_80_n 0.0155943f $X=1.425 $Y=1.515 $X2=0 $Y2=0
cc_48 N_A_M1001_g N_Y_c_104_n 8.84614e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_49 N_A_M1003_g N_Y_c_104_n 0.00196977f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_50 A N_Y_c_104_n 0.0209325f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_51 N_A_c_34_n N_Y_c_104_n 5.54777e-19 $X=1.425 $Y=1.515 $X2=0 $Y2=0
cc_52 N_A_M1004_g Y 0.0263051f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_53 A Y 0.0265979f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A_M1000_g N_VPWR_c_128_n 0.0027763f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_55 N_A_M1001_g N_VPWR_c_128_n 0.0027763f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_56 N_A_M1003_g N_VPWR_c_130_n 0.00501904f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A_M1001_g N_VPWR_c_131_n 0.005209f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_58 N_A_M1003_g N_VPWR_c_131_n 0.005209f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_59 N_A_M1000_g N_VPWR_c_132_n 0.005209f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_VPWR_c_127_n 0.00986025f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_VPWR_c_127_n 0.00982266f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A_M1003_g N_VPWR_c_127_n 0.00986025f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A_M1002_g N_VGND_c_156_n 0.0187336f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_64 A N_VGND_c_156_n 0.013195f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_M1004_g N_VGND_c_158_n 0.0184421f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_66 N_A_M1002_g N_VGND_c_159_n 0.00462012f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_67 N_A_M1004_g N_VGND_c_159_n 0.00462012f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_VGND_c_160_n 0.00450456f $X=0.495 $Y=0.61 $X2=0 $Y2=0
cc_69 N_A_M1004_g N_VGND_c_160_n 0.00450456f $X=1.425 $Y=0.61 $X2=0 $Y2=0
cc_70 N_Y_c_91_n N_VPWR_M1000_d 0.00314376f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_71 N_Y_c_85_n N_VPWR_M1003_d 0.00365063f $X=1.565 $Y=2.035 $X2=0 $Y2=0
cc_72 Y N_VPWR_M1003_d 0.00184872f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_73 N_Y_c_83_n N_VPWR_c_128_n 0.0233699f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_74 N_Y_c_91_n N_VPWR_c_128_n 0.0126919f $X=1.02 $Y=2.035 $X2=0 $Y2=0
cc_75 N_Y_c_84_n N_VPWR_c_128_n 0.0233699f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_76 N_Y_c_84_n N_VPWR_c_130_n 0.0234083f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_77 N_Y_c_85_n N_VPWR_c_130_n 0.0213127f $X=1.565 $Y=2.035 $X2=0 $Y2=0
cc_78 N_Y_c_84_n N_VPWR_c_131_n 0.0144623f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_79 N_Y_c_83_n N_VPWR_c_132_n 0.014549f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_80 N_Y_c_83_n N_VPWR_c_127_n 0.0119743f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_81 N_Y_c_84_n N_VPWR_c_127_n 0.0118344f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_82 N_Y_c_80_n N_VGND_c_156_n 0.0132912f $X=1.305 $Y=0.845 $X2=0 $Y2=0
cc_83 N_Y_c_79_n N_VGND_c_158_n 0.0288308f $X=1.565 $Y=1.095 $X2=0 $Y2=0
cc_84 N_Y_c_80_n N_VGND_c_158_n 0.0132912f $X=1.305 $Y=0.845 $X2=0 $Y2=0
cc_85 N_Y_c_80_n N_VGND_c_159_n 0.0175309f $X=1.305 $Y=0.845 $X2=0 $Y2=0
cc_86 N_Y_c_80_n N_VGND_c_160_n 0.0228888f $X=1.305 $Y=0.845 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dlclkp_1.spice
* Created: Wed Sep  2 12:04:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlclkp_1.pex.spice"
.subckt sky130_fd_sc_ms__dlclkp_1  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_A_83_260#_M1017_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.235647 AS=0.2109 PD=1.51754 PS=2.05 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1018 A_267_80# N_GATE_M1018_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.203803 PD=0.88 PS=1.31246 NRD=12.18 NRS=48.744 M=1 R=4.26667
+ SA=75001 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_83_260#_M1019_d N_A_315_54#_M1019_g A_267_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.162536 AS=0.0768 PD=1.38868 PS=0.88 NRD=21.552 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1001 A_477_124# N_A_309_338#_M1001_g N_A_83_260#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.106664 PD=0.66 PS=0.911321 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75002 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_27_74#_M1016_g A_477_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.102746 AS=0.0504 PD=0.89069 PS=0.66 NRD=28.56 NRS=18.564 M=1 R=2.8
+ SA=75002.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_309_338#_M1004_d N_A_315_54#_M1004_g N_VGND_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.181029 PD=2.05 PS=1.56931 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_CLK_M1002_g N_A_315_54#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13883 AS=0.2183 PD=1.17971 PS=2.07 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1012 A_984_125# N_CLK_M1012_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.12007 PD=0.88 PS=1.02029 NRD=12.18 NRS=14.988 M=1 R=4.26667
+ SA=75000.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_990_393#_M1009_d N_A_27_74#_M1009_g A_984_125# VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_GCLK_M1013_d N_A_990_393#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_83_260#_M1006_g N_A_27_74#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.295849 AS=0.3136 PD=1.7434 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1000 A_261_392# N_GATE_M1000_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.264151 PD=1.24 PS=1.5566 NRD=12.7853 NRS=40.3653 M=1 R=5.55556 SA=90000.9
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1003 N_A_83_260#_M1003_d N_A_309_338#_M1003_g A_261_392# VPB PSHORT L=0.18 W=1
+ AD=0.258873 AS=0.12 PD=2.15493 PS=1.24 NRD=24.6053 NRS=12.7853 M=1 R=5.55556
+ SA=90001.3 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1007 A_487_508# N_A_315_54#_M1007_g N_A_83_260#_M1003_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.108727 PD=0.66 PS=0.90507 NRD=30.4759 NRS=58.6272 M=1
+ R=2.33333 SA=90002 SB=90001 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_74#_M1010_g A_487_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0936833 AS=0.0504 PD=0.89 PS=0.66 NRD=2.3443 NRS=30.4759 M=1 R=2.33333
+ SA=90002.4 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1014 N_A_309_338#_M1014_d N_A_315_54#_M1014_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.187367 PD=2.24 PS=1.78 NRD=0 NRS=19.9167 M=1 R=4.66667
+ SA=90001.1 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1008_d N_CLK_M1008_g N_A_315_54#_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1512 AS=0.2352 PD=1.2 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90002 A=0.1512 P=2.04 MULT=1
MM1015 N_A_990_393#_M1015_d N_CLK_M1015_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=1.1623 NRS=8.1952 M=1 R=4.66667
+ SA=90000.7 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1011 N_VPWR_M1011_d N_A_27_74#_M1011_g N_A_990_393#_M1015_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2718 AS=0.1176 PD=1.51286 PS=1.12 NRD=75.4313 NRS=0 M=1 R=4.66667
+ SA=90001.2 SB=90001 A=0.1512 P=2.04 MULT=1
MM1005 N_GCLK_M1005_d N_A_990_393#_M1005_g N_VPWR_M1011_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3624 PD=2.8 PS=2.01714 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.9104 P=18.17
c_123 VPB 0 1.78419e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dlclkp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a21o_1.spice
* Created: Fri Aug 28 16:59:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21o_1.pex.spice"
.subckt sky130_fd_sc_ms__a21o_1  VNB VPB B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_81_264#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.152558 AS=0.1961 PD=1.22261 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1003 N_A_81_264#_M1003_d N_B1_M1003_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.131942 PD=0.92 PS=1.05739 NRD=0 NRS=22.488 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 A_452_136# N_A1_M1004_g N_A_81_264#_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.104 AS=0.0896 PD=0.965 PS=0.92 NRD=20.148 NRS=0 M=1 R=4.26667 SA=75001.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_452_136# VNB NLOWVT L=0.15 W=0.64 AD=0.1696
+ AS=0.104 PD=1.81 PS=0.965 NRD=0 NRS=20.148 M=1 R=4.26667 SA=75001.6 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_81_264#_M1005_g N_X_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1006 N_A_367_392#_M1006_d N_B1_M1006_g N_A_81_264#_M1006_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_367_392#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=1.9503 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1002 N_A_367_392#_M1002_d N_A2_M1002_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.15 PD=2.52 PS=1.3 NRD=0 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_34 VNB 0 1.84796e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a21o_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sdfxbp_2.spice
* Created: Wed Sep  2 12:31:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfxbp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfxbp_2  VNB VPB SCE D SCD CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1038 N_VGND_M1038_d N_SCE_M1038_g N_A_36_74#_M1038_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1017 A_223_74# N_A_36_74#_M1017_g N_VGND_M1038_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_301_74#_M1018_d N_D_M1018_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.12495 AS=0.0504 PD=1.015 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1033 A_450_74# N_SCE_M1033_g N_A_301_74#_M1018_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.12495 PD=0.66 PS=1.015 NRD=18.564 NRS=45.708 M=1 R=2.8
+ SA=75001.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_SCD_M1031_g A_450_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_630_74#_M1005_d N_CLK_M1005_g N_VGND_M1031_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_828_74#_M1015_d N_A_630_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.2109 PD=2.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_1021_97#_M1024_d N_A_630_74#_M1024_g N_A_301_74#_M1024_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1155 PD=1.03 PS=1.39 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1035 A_1173_97# N_A_828_74#_M1035_g N_A_1021_97#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.082125 AS=0.1281 PD=0.885 PS=1.03 NRD=40.152 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1243_48#_M1020_g A_1173_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125004 AS=0.082125 PD=1.00454 PS=0.885 NRD=0 NRS=40.152 M=1 R=2.8
+ SA=75001.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_1243_48#_M1025_d N_A_1021_97#_M1025_g N_VGND_M1020_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.163696 PD=0.83 PS=1.31546 NRD=0 NRS=72 M=1
+ R=3.66667 SA=75001.5 SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1039 N_A_1511_74#_M1039_d N_A_828_74#_M1039_g N_A_1243_48#_M1025_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.163696 AS=0.077 PD=1.31546 PS=0.83 NRD=72 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1012 A_1663_74# N_A_630_74#_M1012_g N_A_1511_74#_M1039_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.125004 PD=0.66 PS=1.00454 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1711_48#_M1013_g A_1663_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.139976 AS=0.0504 PD=1.06448 PS=0.66 NRD=79.5 NRS=18.564 M=1 R=2.8
+ SA=75003.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1032 N_A_1711_48#_M1032_d N_A_1511_74#_M1032_g N_VGND_M1013_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.246624 PD=2.05 PS=1.87552 NRD=0 NRS=45.12 M=1
+ R=4.93333 SA=75002.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_1711_48#_M1000_g N_Q_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1029_d N_A_1711_48#_M1029_g N_Q_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_1711_48#_M1027_g N_A_2322_368#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.12007 AS=0.1824 PD=1.02029 PS=1.85 NRD=12.648 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1027_d N_A_2322_368#_M1002_g N_Q_N_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13883 AS=0.10915 PD=1.17971 PS=1.035 NRD=2.424 NRS=0.804 M=1
+ R=4.93333 SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1026_d N_A_2322_368#_M1026_g N_Q_N_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1962 AS=0.10915 PD=2.05 PS=1.035 NRD=0 NRS=1.62 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_SCE_M1004_g N_A_36_74#_M1004_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.2336 PD=0.91 PS=2.01 NRD=0 NRS=24.6053 M=1 R=3.55556 SA=90000.3
+ SB=90003 A=0.1152 P=1.64 MULT=1
MM1006 A_241_453# N_SCE_M1006_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.0864 PD=0.88 PS=0.91 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90002.5 A=0.1152 P=1.64 MULT=1
MM1016 N_A_301_74#_M1016_d N_D_M1016_g A_241_453# VPB PSHORT L=0.18 W=0.64
+ AD=0.104 AS=0.0768 PD=0.965 PS=0.88 NRD=15.3857 NRS=19.9955 M=1 R=3.55556
+ SA=90001.1 SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1021 A_426_453# N_A_36_74#_M1021_g N_A_301_74#_M1016_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0976 AS=0.104 PD=0.945 PS=0.965 NRD=30.0031 NRS=0 M=1 R=3.55556
+ SA=90001.6 SB=90001.6 A=0.1152 P=1.64 MULT=1
MM1037 N_VPWR_M1037_d N_SCD_M1037_g A_426_453# VPB PSHORT L=0.18 W=0.64
+ AD=0.179373 AS=0.0976 PD=1.24364 PS=0.945 NRD=40.0107 NRS=30.0031 M=1
+ R=3.55556 SA=90002.1 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1007 N_A_630_74#_M1007_d N_CLK_M1007_g N_VPWR_M1037_d VPB PSHORT L=0.18 W=1.12
+ AD=0.5488 AS=0.313902 PD=3.22 PS=2.17636 NRD=0 NRS=22.852 M=1 R=6.22222
+ SA=90001.7 SB=90000.4 A=0.2016 P=2.6 MULT=1
MM1028 N_A_828_74#_M1028_d N_A_630_74#_M1028_g N_VPWR_M1028_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1023 N_A_1021_97#_M1023_d N_A_828_74#_M1023_g N_A_301_74#_M1023_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.07455 AS=0.1176 PD=0.775 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90004.1 A=0.0756 P=1.2 MULT=1
MM1008 A_1220_499# N_A_630_74#_M1008_g N_A_1021_97#_M1023_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.07455 PD=0.66 PS=0.775 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90000.7 SB=90003.5 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_1243_48#_M1011_g A_1220_499# VPB PSHORT L=0.18 W=0.42
+ AD=0.120075 AS=0.0504 PD=1.00333 PS=0.66 NRD=108.291 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1019 N_A_1243_48#_M1019_d N_A_1021_97#_M1019_g N_VPWR_M1011_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2583 AS=0.24015 PD=1.455 PS=2.00667 NRD=2.3443 NRS=54.1356
+ M=1 R=4.66667 SA=90001 SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1001 N_A_1511_74#_M1001_d N_A_630_74#_M1001_g N_A_1243_48#_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1778 AS=0.2583 PD=1.59333 PS=1.455 NRD=0 NRS=76.2193 M=1
+ R=4.66667 SA=90001.8 SB=90001 A=0.1512 P=2.04 MULT=1
MM1022 A_1694_508# N_A_828_74#_M1022_g N_A_1511_74#_M1001_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0889 PD=0.66 PS=0.796667 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90002.9 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1003 N_VPWR_M1003_d N_A_1711_48#_M1003_g A_1694_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.112454 AS=0.0504 PD=0.922817 PS=0.66 NRD=53.9386 NRS=30.4759 M=1
+ R=2.33333 SA=90003.4 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1014 N_A_1711_48#_M1014_d N_A_1511_74#_M1014_g N_VPWR_M1003_d VPB PSHORT
+ L=0.18 W=1 AD=0.27 AS=0.267746 PD=2.54 PS=2.19718 NRD=0 NRS=32.4853 M=1
+ R=5.55556 SA=90001.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1009 N_Q_M1009_d N_A_1711_48#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_Q_M1009_d N_A_1711_48#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1030 N_VPWR_M1030_d N_A_1711_48#_M1030_g N_A_2322_368#_M1030_s VPB PSHORT
+ L=0.18 W=1 AD=0.178019 AS=0.27 PD=1.38208 PS=2.54 NRD=14.1052 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1034 N_Q_N_M1034_d N_A_2322_368#_M1034_g N_VPWR_M1030_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.199381 PD=1.39 PS=1.54792 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1036 N_Q_N_M1034_d N_A_2322_368#_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.7052 P=31.36
c_147 VNB 0 1.47924e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sdfxbp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o221a_2.pxi.spice
* Created: Fri Aug 28 17:56:43 2020
* 
x_PM_SKY130_FD_SC_MS__O221A_2%C1 N_C1_M1006_g N_C1_c_85_n N_C1_M1007_g C1
+ N_C1_c_87_n PM_SKY130_FD_SC_MS__O221A_2%C1
x_PM_SKY130_FD_SC_MS__O221A_2%B1 N_B1_M1009_g N_B1_c_116_n N_B1_M1011_g B1
+ N_B1_c_114_n N_B1_c_115_n PM_SKY130_FD_SC_MS__O221A_2%B1
x_PM_SKY130_FD_SC_MS__O221A_2%B2 N_B2_c_153_n N_B2_M1003_g N_B2_c_154_n
+ N_B2_M1002_g B2 B2 N_B2_c_156_n N_B2_c_157_n PM_SKY130_FD_SC_MS__O221A_2%B2
x_PM_SKY130_FD_SC_MS__O221A_2%A2 N_A2_M1001_g N_A2_M1010_g A2 N_A2_c_195_n
+ N_A2_c_196_n PM_SKY130_FD_SC_MS__O221A_2%A2
x_PM_SKY130_FD_SC_MS__O221A_2%A1 N_A1_M1005_g N_A1_M1004_g A1 N_A1_c_229_n
+ N_A1_c_230_n PM_SKY130_FD_SC_MS__O221A_2%A1
x_PM_SKY130_FD_SC_MS__O221A_2%A_27_368# N_A_27_368#_M1007_s N_A_27_368#_M1006_s
+ N_A_27_368#_M1002_d N_A_27_368#_M1000_g N_A_27_368#_M1012_g
+ N_A_27_368#_c_273_n N_A_27_368#_M1008_g N_A_27_368#_M1013_g
+ N_A_27_368#_c_276_n N_A_27_368#_c_285_n N_A_27_368#_c_277_n
+ N_A_27_368#_c_278_n N_A_27_368#_c_296_n N_A_27_368#_c_287_n
+ N_A_27_368#_c_317_n N_A_27_368#_c_279_n N_A_27_368#_c_289_n
+ N_A_27_368#_c_280_n N_A_27_368#_c_313_n N_A_27_368#_c_281_n
+ N_A_27_368#_c_282_n PM_SKY130_FD_SC_MS__O221A_2%A_27_368#
x_PM_SKY130_FD_SC_MS__O221A_2%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_M1013_s
+ N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_393_n VPWR
+ N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n
+ N_VPWR_c_389_n PM_SKY130_FD_SC_MS__O221A_2%VPWR
x_PM_SKY130_FD_SC_MS__O221A_2%X N_X_M1000_s N_X_M1012_d N_X_c_442_n N_X_c_443_n
+ N_X_c_439_n X X N_X_c_440_n X PM_SKY130_FD_SC_MS__O221A_2%X
x_PM_SKY130_FD_SC_MS__O221A_2%A_165_74# N_A_165_74#_M1007_d N_A_165_74#_M1003_d
+ N_A_165_74#_c_474_n N_A_165_74#_c_475_n N_A_165_74#_c_476_n
+ PM_SKY130_FD_SC_MS__O221A_2%A_165_74#
x_PM_SKY130_FD_SC_MS__O221A_2%A_264_74# N_A_264_74#_M1009_d N_A_264_74#_M1010_d
+ N_A_264_74#_c_500_n N_A_264_74#_c_501_n N_A_264_74#_c_502_n
+ PM_SKY130_FD_SC_MS__O221A_2%A_264_74#
x_PM_SKY130_FD_SC_MS__O221A_2%VGND N_VGND_M1010_s N_VGND_M1004_d N_VGND_M1008_d
+ N_VGND_c_535_n N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n
+ N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n VGND N_VGND_c_543_n
+ N_VGND_c_544_n PM_SKY130_FD_SC_MS__O221A_2%VGND
cc_1 VNB N_C1_M1006_g 0.0100079f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_2 VNB N_C1_c_85_n 0.0227378f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.22
cc_3 VNB C1 0.0159976f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_C1_c_87_n 0.0813779f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.385
cc_5 VNB N_B1_M1009_g 0.0263143f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_6 VNB N_B1_c_114_n 0.00333483f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_7 VNB N_B1_c_115_n 0.0397528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_c_153_n 0.0181556f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_9 VNB N_B2_c_154_n 0.0318298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB B2 0.00636131f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.385
cc_11 VNB N_B2_c_156_n 0.0122502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B2_c_157_n 0.00898421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1010_g 0.027284f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_14 VNB N_A2_c_195_n 0.0269948f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_15 VNB N_A2_c_196_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1004_g 0.0261039f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_17 VNB N_A1_c_229_n 0.0247509f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_18 VNB N_A1_c_230_n 0.00552033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_368#_M1000_g 0.0241917f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_20 VNB N_A_27_368#_M1012_g 5.20588e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_368#_c_273_n 0.00638712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_368#_M1008_g 0.0251809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_368#_M1013_g 0.0150953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_368#_c_276_n 0.0206797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_c_277_n 0.0204696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_368#_c_278_n 0.00460576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_368#_c_279_n 2.18704e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_368#_c_280_n 0.00797994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_368#_c_281_n 0.00257315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_368#_c_282_n 0.0272958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_389_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_439_n 0.00795141f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.385
cc_33 VNB N_X_c_440_n 0.00274256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.00577223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_165_74#_c_474_n 0.00342538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_165_74#_c_475_n 0.00716791f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_37 VNB N_A_165_74#_c_476_n 0.00704577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_264_74#_c_500_n 0.0300192f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.74
cc_39 VNB N_A_264_74#_c_501_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_40 VNB N_A_264_74#_c_502_n 0.00313103f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_41 VNB N_VGND_c_535_n 0.0106116f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_42 VNB N_VGND_c_536_n 0.017767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_537_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_538_n 0.0506881f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_45 VNB N_VGND_c_539_n 0.0648512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_540_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_541_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_542_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_543_n 0.0221763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_544_n 0.299576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_C1_M1006_g 0.0319821f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_52 VPB N_B1_c_116_n 0.0214444f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.22
cc_53 VPB N_B1_c_114_n 0.00384703f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_54 VPB N_B1_c_115_n 0.0183381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_B2_M1002_g 0.0210678f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_56 VPB B2 0.00471405f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.385
cc_57 VPB N_B2_c_157_n 0.00544883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A2_M1001_g 0.0233423f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_59 VPB N_A2_c_195_n 0.00566547f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_60 VPB N_A2_c_196_n 0.00203931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A1_M1005_g 0.023745f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_62 VPB N_A1_c_229_n 0.0056412f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_63 VPB N_A1_c_230_n 0.0033526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_368#_M1012_g 0.0245837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_368#_M1013_g 0.0274013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_368#_c_285_n 0.0313441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_368#_c_278_n 0.00441313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_368#_c_287_n 0.0034139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_368#_c_279_n 0.00289029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_368#_c_289_n 0.0159288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_390_n 0.025885f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_72 VPB N_VPWR_c_391_n 0.0143413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_392_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_74 VPB N_VPWR_c_393_n 0.0644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_394_n 0.0196898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_395_n 0.0577377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_396_n 0.0194151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_397_n 0.0174777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_398_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_389_n 0.108289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_X_c_442_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_X_c_443_n 0.00459114f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_83 VPB N_X_c_439_n 8.51836e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.385
cc_84 N_C1_c_85_n N_B1_M1009_g 0.024596f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_85 N_C1_c_87_n N_B1_c_114_n 8.785e-19 $X=0.75 $Y=1.385 $X2=0 $Y2=0
cc_86 N_C1_M1006_g N_B1_c_115_n 0.00332362f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_87 N_C1_c_87_n N_B1_c_115_n 0.0111125f $X=0.75 $Y=1.385 $X2=0 $Y2=0
cc_88 N_C1_M1006_g N_A_27_368#_c_285_n 0.0150376f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_89 N_C1_c_85_n N_A_27_368#_c_277_n 0.00869286f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C1_M1006_g N_A_27_368#_c_278_n 0.00886683f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_91 N_C1_c_85_n N_A_27_368#_c_278_n 0.00554011f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_92 C1 N_A_27_368#_c_278_n 0.0267371f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_C1_c_87_n N_A_27_368#_c_278_n 0.018301f $X=0.75 $Y=1.385 $X2=0 $Y2=0
cc_94 N_C1_c_87_n N_A_27_368#_c_296_n 0.00161321f $X=0.75 $Y=1.385 $X2=0 $Y2=0
cc_95 N_C1_M1006_g N_A_27_368#_c_289_n 0.0266395f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_96 C1 N_A_27_368#_c_289_n 0.0178783f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_97 N_C1_c_87_n N_A_27_368#_c_289_n 0.00303699f $X=0.75 $Y=1.385 $X2=0 $Y2=0
cc_98 N_C1_c_85_n N_A_27_368#_c_280_n 0.00306847f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_99 C1 N_A_27_368#_c_280_n 0.00555399f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_100 N_C1_c_87_n N_A_27_368#_c_280_n 0.00825166f $X=0.75 $Y=1.385 $X2=0 $Y2=0
cc_101 N_C1_M1006_g N_VPWR_c_390_n 0.00590965f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_102 N_C1_M1006_g N_VPWR_c_394_n 0.00567889f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_103 N_C1_M1006_g N_VPWR_c_389_n 0.00610055f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_104 N_C1_c_85_n N_A_165_74#_c_475_n 0.005506f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_105 N_C1_c_85_n N_A_264_74#_c_502_n 2.32508e-19 $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_106 N_C1_c_85_n N_VGND_c_539_n 0.00349296f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_107 N_C1_c_85_n N_VGND_c_544_n 0.00551056f $X=0.75 $Y=1.22 $X2=0 $Y2=0
cc_108 N_B1_M1009_g N_B2_c_153_n 0.027221f $X=1.245 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_109 N_B1_c_116_n N_B2_M1002_g 0.0374383f $X=1.585 $Y=1.725 $X2=0 $Y2=0
cc_110 N_B1_c_116_n B2 0.00302504f $X=1.585 $Y=1.725 $X2=0 $Y2=0
cc_111 N_B1_c_114_n B2 0.0354777f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B1_c_115_n B2 0.00955028f $X=1.245 $Y=1.537 $X2=0 $Y2=0
cc_113 N_B1_M1009_g N_B2_c_156_n 3.78334e-19 $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_c_114_n N_B2_c_156_n 2.50692e-19 $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_115 N_B1_c_115_n N_B2_c_156_n 0.00382197f $X=1.245 $Y=1.537 $X2=0 $Y2=0
cc_116 N_B1_c_115_n N_B2_c_157_n 0.0374383f $X=1.245 $Y=1.537 $X2=0 $Y2=0
cc_117 N_B1_M1009_g N_A_27_368#_c_277_n 0.00133362f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B1_c_114_n N_A_27_368#_c_278_n 0.0211588f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B1_c_115_n N_A_27_368#_c_278_n 0.00217035f $X=1.245 $Y=1.537 $X2=0
+ $Y2=0
cc_120 N_B1_c_116_n N_A_27_368#_c_296_n 0.0200624f $X=1.585 $Y=1.725 $X2=0 $Y2=0
cc_121 N_B1_c_114_n N_A_27_368#_c_296_n 0.0262472f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_122 N_B1_c_115_n N_A_27_368#_c_296_n 0.00430646f $X=1.245 $Y=1.537 $X2=0
+ $Y2=0
cc_123 N_B1_c_116_n N_A_27_368#_c_287_n 0.00243009f $X=1.585 $Y=1.725 $X2=0
+ $Y2=0
cc_124 N_B1_c_116_n N_VPWR_c_390_n 0.016942f $X=1.585 $Y=1.725 $X2=0 $Y2=0
cc_125 N_B1_c_116_n N_VPWR_c_395_n 0.00492916f $X=1.585 $Y=1.725 $X2=0 $Y2=0
cc_126 N_B1_c_116_n N_VPWR_c_389_n 0.00511769f $X=1.585 $Y=1.725 $X2=0 $Y2=0
cc_127 N_B1_M1009_g N_A_165_74#_c_474_n 0.0123547f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B1_M1009_g N_A_165_74#_c_475_n 4.59233e-19 $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B1_c_114_n N_A_165_74#_c_475_n 0.00341112f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_130 N_B1_c_115_n N_A_165_74#_c_475_n 3.67352e-19 $X=1.245 $Y=1.537 $X2=0
+ $Y2=0
cc_131 N_B1_M1009_g N_A_165_74#_c_476_n 0.00133243f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B1_c_115_n N_A_264_74#_c_500_n 2.28236e-19 $X=1.245 $Y=1.537 $X2=0
+ $Y2=0
cc_133 N_B1_M1009_g N_A_264_74#_c_502_n 0.00591218f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B1_c_114_n N_A_264_74#_c_502_n 0.00797323f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B1_c_115_n N_A_264_74#_c_502_n 0.00626205f $X=1.245 $Y=1.537 $X2=0
+ $Y2=0
cc_136 N_B1_M1009_g N_VGND_c_539_n 0.00291649f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B1_M1009_g N_VGND_c_544_n 0.00360544f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B2_M1002_g N_A2_M1001_g 0.0222225f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_139 N_B2_c_154_n N_A2_M1010_g 0.00639049f $X=2.08 $Y=1.335 $X2=0 $Y2=0
cc_140 B2 N_A2_c_195_n 0.00294479f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_141 N_B2_c_156_n N_A2_c_195_n 0.0174954f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_142 B2 N_A2_c_196_n 0.0308891f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_B2_c_156_n N_A2_c_196_n 3.95877e-19 $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_144 N_B2_M1002_g N_A_27_368#_c_296_n 0.0127019f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_145 B2 N_A_27_368#_c_296_n 0.0339127f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_B2_M1002_g N_A_27_368#_c_287_n 0.0143201f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_147 N_B2_M1002_g N_A_27_368#_c_313_n 8.84614e-19 $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_148 B2 N_A_27_368#_c_313_n 0.0157526f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B2_c_157_n N_A_27_368#_c_313_n 7.76119e-19 $X=2.08 $Y=1.68 $X2=0 $Y2=0
cc_150 N_B2_M1002_g N_VPWR_c_390_n 0.00212941f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_151 N_B2_M1002_g N_VPWR_c_395_n 0.00567889f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_152 N_B2_M1002_g N_VPWR_c_389_n 0.00610055f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_153 N_B2_c_153_n N_A_165_74#_c_474_n 0.00917015f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_154 N_B2_c_153_n N_A_165_74#_c_476_n 0.0096459f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_155 N_B2_c_153_n N_A_264_74#_c_500_n 0.0116015f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_156 N_B2_c_154_n N_A_264_74#_c_500_n 0.0123197f $X=2.08 $Y=1.335 $X2=0 $Y2=0
cc_157 B2 N_A_264_74#_c_500_n 0.0510553f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_158 B2 N_A_264_74#_c_502_n 0.00465791f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B2_c_153_n N_VGND_c_535_n 0.00383008f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_160 N_B2_c_153_n N_VGND_c_539_n 0.00292759f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_161 N_B2_c_153_n N_VGND_c_544_n 0.00363909f $X=1.75 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A2_M1001_g N_A1_M1005_g 0.0440971f $X=2.575 $Y=2.34 $X2=0 $Y2=0
cc_163 N_A2_c_196_n N_A1_M1005_g 3.45791e-19 $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A2_M1010_g N_A1_M1004_g 0.0195038f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A2_c_195_n N_A1_c_229_n 0.0174484f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_166 N_A2_c_196_n N_A1_c_229_n 3.82036e-19 $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A2_M1001_g N_A1_c_230_n 2.83567e-19 $X=2.575 $Y=2.34 $X2=0 $Y2=0
cc_168 N_A2_c_195_n N_A1_c_230_n 0.00203158f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A2_c_196_n N_A1_c_230_n 0.0320815f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A2_M1001_g N_A_27_368#_c_287_n 0.0203086f $X=2.575 $Y=2.34 $X2=0 $Y2=0
cc_171 N_A2_M1001_g N_A_27_368#_c_317_n 0.0182755f $X=2.575 $Y=2.34 $X2=0 $Y2=0
cc_172 N_A2_c_195_n N_A_27_368#_c_317_n 6.98124e-19 $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A2_c_196_n N_A_27_368#_c_317_n 0.0229716f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A2_M1001_g N_VPWR_c_395_n 0.0059286f $X=2.575 $Y=2.34 $X2=0 $Y2=0
cc_175 N_A2_M1001_g N_VPWR_c_389_n 0.00610055f $X=2.575 $Y=2.34 $X2=0 $Y2=0
cc_176 N_A2_M1010_g N_A_165_74#_c_476_n 0.00109581f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A2_M1010_g N_A_264_74#_c_500_n 0.0151035f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_c_195_n N_A_264_74#_c_500_n 0.001245f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A2_c_196_n N_A_264_74#_c_500_n 0.0247243f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A2_M1010_g N_A_264_74#_c_501_n 3.97481e-19 $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A2_M1010_g N_VGND_c_535_n 0.0124788f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A2_M1010_g N_VGND_c_541_n 0.00383152f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A2_M1010_g N_VGND_c_544_n 0.00757637f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A1_M1004_g N_A_27_368#_M1000_g 0.0233513f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_M1005_g N_A_27_368#_M1012_g 0.0156104f $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_186 N_A1_c_229_n N_A_27_368#_M1012_g 7.51971e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_187 N_A1_M1005_g N_A_27_368#_c_317_n 0.0186995f $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_188 N_A1_c_229_n N_A_27_368#_c_317_n 7.07929e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A1_c_230_n N_A_27_368#_c_317_n 0.0251787f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A1_M1005_g N_A_27_368#_c_279_n 0.00348845f $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_191 N_A1_c_229_n N_A_27_368#_c_279_n 2.18308e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_192 N_A1_c_230_n N_A_27_368#_c_279_n 0.009884f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A1_M1004_g N_A_27_368#_c_281_n 5.96621e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_c_229_n N_A_27_368#_c_281_n 0.00170854f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A1_c_230_n N_A_27_368#_c_281_n 0.0231673f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A1_M1004_g N_A_27_368#_c_282_n 9.38887e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_c_229_n N_A_27_368#_c_282_n 0.0188248f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A1_c_230_n N_A_27_368#_c_282_n 3.50433e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A1_M1005_g N_VPWR_c_391_n 0.0177557f $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_200 N_A1_M1005_g N_VPWR_c_395_n 0.0059286f $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_201 N_A1_M1005_g N_VPWR_c_389_n 0.00610055f $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_202 N_A1_M1005_g N_X_c_442_n 8.2737e-19 $X=3.145 $Y=2.34 $X2=0 $Y2=0
cc_203 N_A1_M1004_g N_A_264_74#_c_500_n 0.00351804f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_c_229_n N_A_264_74#_c_500_n 3.1281e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_205 N_A1_c_230_n N_A_264_74#_c_500_n 0.00993544f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A1_M1004_g N_A_264_74#_c_501_n 0.00775604f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A1_M1004_g N_VGND_c_535_n 5.14838e-19 $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1004_g N_VGND_c_536_n 0.00657843f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A1_c_229_n N_VGND_c_536_n 7.12986e-19 $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A1_c_230_n N_VGND_c_536_n 0.00660905f $X=3.22 $Y=1.515 $X2=0 $Y2=0
cc_211 N_A1_M1004_g N_VGND_c_541_n 0.00434272f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A1_M1004_g N_VGND_c_544_n 0.0082141f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_27_368#_c_296_n N_VPWR_M1006_d 0.0252601f $X=2.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_27_368#_c_289_n N_VPWR_M1006_d 0.00627503f $X=0.775 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_27_368#_c_317_n N_VPWR_M1005_d 0.0177764f $X=3.565 $Y=2.035 $X2=0
+ $Y2=0
cc_216 N_A_27_368#_c_279_n N_VPWR_M1005_d 0.00223621f $X=3.65 $Y=1.95 $X2=0
+ $Y2=0
cc_217 N_A_27_368#_c_285_n N_VPWR_c_390_n 0.0222698f $X=0.28 $Y=2.695 $X2=0
+ $Y2=0
cc_218 N_A_27_368#_c_287_n N_VPWR_c_390_n 0.0175472f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_219 N_A_27_368#_c_289_n N_VPWR_c_390_n 0.0664764f $X=0.775 $Y=1.97 $X2=0
+ $Y2=0
cc_220 N_A_27_368#_M1012_g N_VPWR_c_391_n 0.00521714f $X=3.845 $Y=2.4 $X2=0
+ $Y2=0
cc_221 N_A_27_368#_c_317_n N_VPWR_c_391_n 0.0245287f $X=3.565 $Y=2.035 $X2=0
+ $Y2=0
cc_222 N_A_27_368#_c_282_n N_VPWR_c_391_n 3.83802e-19 $X=3.765 $Y=1.395 $X2=0
+ $Y2=0
cc_223 N_A_27_368#_M1013_g N_VPWR_c_393_n 0.00647357f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_27_368#_c_285_n N_VPWR_c_394_n 0.00975961f $X=0.28 $Y=2.695 $X2=0
+ $Y2=0
cc_225 N_A_27_368#_c_287_n N_VPWR_c_395_n 0.00975961f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_226 N_A_27_368#_M1012_g N_VPWR_c_396_n 0.005209f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_27_368#_M1013_g N_VPWR_c_396_n 0.0048691f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A_27_368#_M1012_g N_VPWR_c_389_n 0.00986727f $X=3.845 $Y=2.4 $X2=0
+ $Y2=0
cc_229 N_A_27_368#_M1013_g N_VPWR_c_389_n 0.00875947f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_230 N_A_27_368#_c_285_n N_VPWR_c_389_n 0.0111753f $X=0.28 $Y=2.695 $X2=0
+ $Y2=0
cc_231 N_A_27_368#_c_287_n N_VPWR_c_389_n 0.0111753f $X=2.23 $Y=2.375 $X2=0
+ $Y2=0
cc_232 N_A_27_368#_c_296_n A_335_368# 0.0060399f $X=2.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_233 N_A_27_368#_c_317_n A_533_368# 0.0186283f $X=3.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_234 N_A_27_368#_M1012_g N_X_c_442_n 0.0143207f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_27_368#_M1013_g N_X_c_442_n 0.0149161f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A_27_368#_M1012_g N_X_c_443_n 0.00304813f $X=3.845 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_27_368#_c_273_n N_X_c_443_n 0.00277677f $X=4.095 $Y=1.395 $X2=0 $Y2=0
cc_238 N_A_27_368#_M1013_g N_X_c_443_n 0.00270934f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_27_368#_c_279_n N_X_c_443_n 0.00565814f $X=3.65 $Y=1.95 $X2=0 $Y2=0
cc_240 N_A_27_368#_c_281_n N_X_c_443_n 0.00151667f $X=3.76 $Y=1.485 $X2=0 $Y2=0
cc_241 N_A_27_368#_M1000_g N_X_c_439_n 8.79499e-19 $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_27_368#_M1008_g N_X_c_439_n 0.00708533f $X=4.17 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_27_368#_M1013_g N_X_c_439_n 0.0178909f $X=4.295 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_27_368#_c_276_n N_X_c_439_n 0.0110677f $X=4.24 $Y=1.395 $X2=0 $Y2=0
cc_245 N_A_27_368#_c_279_n N_X_c_439_n 0.00535845f $X=3.65 $Y=1.95 $X2=0 $Y2=0
cc_246 N_A_27_368#_c_281_n N_X_c_439_n 0.0243803f $X=3.76 $Y=1.485 $X2=0 $Y2=0
cc_247 N_A_27_368#_c_282_n N_X_c_439_n 0.00206575f $X=3.765 $Y=1.395 $X2=0 $Y2=0
cc_248 N_A_27_368#_M1000_g N_X_c_440_n 0.00675574f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_27_368#_M1008_g N_X_c_440_n 0.0177451f $X=4.17 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_27_368#_M1000_g X 0.00303662f $X=3.74 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_27_368#_M1008_g X 0.00692602f $X=4.17 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_27_368#_c_281_n X 0.0102861f $X=3.76 $Y=1.485 $X2=0 $Y2=0
cc_253 N_A_27_368#_c_282_n X 0.00430299f $X=3.765 $Y=1.395 $X2=0 $Y2=0
cc_254 N_A_27_368#_c_277_n N_A_165_74#_c_475_n 0.0593848f $X=0.535 $Y=0.515
+ $X2=0 $Y2=0
cc_255 N_A_27_368#_M1000_g N_A_264_74#_c_500_n 2.49809e-19 $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_27_368#_c_278_n N_A_264_74#_c_502_n 0.00142925f $X=0.69 $Y=1.82 $X2=0
+ $Y2=0
cc_257 N_A_27_368#_M1000_g N_VGND_c_536_n 0.00805013f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_258 N_A_27_368#_c_281_n N_VGND_c_536_n 0.00431466f $X=3.76 $Y=1.485 $X2=0
+ $Y2=0
cc_259 N_A_27_368#_c_282_n N_VGND_c_536_n 5.53507e-19 $X=3.765 $Y=1.395 $X2=0
+ $Y2=0
cc_260 N_A_27_368#_M1008_g N_VGND_c_538_n 0.00925276f $X=4.17 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_27_368#_c_277_n N_VGND_c_539_n 0.0176636f $X=0.535 $Y=0.515 $X2=0
+ $Y2=0
cc_262 N_A_27_368#_M1000_g N_VGND_c_543_n 0.00434272f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_263 N_A_27_368#_M1008_g N_VGND_c_543_n 0.00291513f $X=4.17 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_27_368#_M1000_g N_VGND_c_544_n 0.00821312f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_265 N_A_27_368#_M1008_g N_VGND_c_544_n 0.00363054f $X=4.17 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_27_368#_c_277_n N_VGND_c_544_n 0.0143978f $X=0.535 $Y=0.515 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_391_n N_X_c_442_n 0.027028f $X=3.57 $Y=2.455 $X2=0 $Y2=0
cc_268 N_VPWR_c_396_n N_X_c_442_n 0.0157112f $X=4.435 $Y=3.33 $X2=0 $Y2=0
cc_269 N_VPWR_c_389_n N_X_c_442_n 0.0127977f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_270 N_VPWR_c_393_n N_X_c_443_n 0.0455874f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_271 N_X_c_440_n N_VGND_c_536_n 0.0324855f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_272 N_X_c_440_n N_VGND_c_538_n 0.0317393f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_273 N_X_c_440_n N_VGND_c_543_n 0.0205856f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_274 N_X_c_440_n N_VGND_c_544_n 0.0166302f $X=3.955 $Y=0.515 $X2=0 $Y2=0
cc_275 N_A_165_74#_c_474_n N_A_264_74#_M1009_d 0.00321664f $X=1.8 $Y=0.435
+ $X2=-0.19 $Y2=-0.245
cc_276 N_A_165_74#_M1003_d N_A_264_74#_c_500_n 0.0030579f $X=1.825 $Y=0.37 $X2=0
+ $Y2=0
cc_277 N_A_165_74#_c_474_n N_A_264_74#_c_500_n 0.00356375f $X=1.8 $Y=0.435 $X2=0
+ $Y2=0
cc_278 N_A_165_74#_c_476_n N_A_264_74#_c_500_n 0.020435f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_279 N_A_165_74#_c_474_n N_A_264_74#_c_502_n 0.0127762f $X=1.8 $Y=0.435 $X2=0
+ $Y2=0
cc_280 N_A_165_74#_c_475_n N_A_264_74#_c_502_n 0.0124866f $X=1.03 $Y=0.515 $X2=0
+ $Y2=0
cc_281 N_A_165_74#_c_476_n N_VGND_c_535_n 0.0323609f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_282 N_A_165_74#_c_474_n N_VGND_c_539_n 0.0269436f $X=1.8 $Y=0.435 $X2=0 $Y2=0
cc_283 N_A_165_74#_c_475_n N_VGND_c_539_n 0.00758556f $X=1.03 $Y=0.515 $X2=0
+ $Y2=0
cc_284 N_A_165_74#_c_476_n N_VGND_c_539_n 0.0142041f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_285 N_A_165_74#_c_474_n N_VGND_c_544_n 0.0229064f $X=1.8 $Y=0.435 $X2=0 $Y2=0
cc_286 N_A_165_74#_c_475_n N_VGND_c_544_n 0.00627867f $X=1.03 $Y=0.515 $X2=0
+ $Y2=0
cc_287 N_A_165_74#_c_476_n N_VGND_c_544_n 0.011859f $X=1.965 $Y=0.435 $X2=0
+ $Y2=0
cc_288 N_A_264_74#_c_500_n N_VGND_M1010_s 0.0030579f $X=2.87 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_264_74#_c_500_n N_VGND_c_535_n 0.02102f $X=2.87 $Y=1.095 $X2=0 $Y2=0
cc_290 N_A_264_74#_c_501_n N_VGND_c_535_n 0.0179318f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_291 N_A_264_74#_c_500_n N_VGND_c_536_n 0.00584871f $X=2.87 $Y=1.095 $X2=0
+ $Y2=0
cc_292 N_A_264_74#_c_501_n N_VGND_c_536_n 0.0244878f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_293 N_A_264_74#_c_501_n N_VGND_c_541_n 0.0109942f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_294 N_A_264_74#_c_501_n N_VGND_c_544_n 0.00904371f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_27_74# a_398_74# a_612_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X1 a_1225_74# a_398_74# a_1324_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_1514_88# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_1223_347# a_225_74# a_1324_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_27_74# a_225_74# a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 a_1436_88# a_1484_62# a_1514_88# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 VGND a_1940_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_767_402# a_612_74# a_1035_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X8 a_612_74# a_225_74# a_719_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X9 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_1035_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_612_74# a_398_74# a_732_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 a_719_463# a_767_402# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X13 Q a_1940_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_1483_508# a_1484_62# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 a_1940_74# a_1324_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_1940_74# a_1324_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X17 VPWR a_1940_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_1324_392# a_225_74# a_1436_88# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X20 VPWR a_612_74# a_767_402# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X21 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_1324_392# a_398_74# a_1483_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X23 VPWR a_1324_392# a_1484_62# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X24 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X25 a_767_402# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X26 Q a_1940_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND a_612_74# a_1225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VPWR a_612_74# a_1223_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X30 VPWR a_1324_392# a_1940_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X31 VPWR a_1940_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 VGND a_1324_392# a_1484_62# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 VPWR SET_B a_1324_392# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X34 a_732_74# a_767_402# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 Q a_1940_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 VGND a_1940_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 Q a_1940_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

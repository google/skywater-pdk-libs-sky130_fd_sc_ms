* File: sky130_fd_sc_ms__einvn_2.pxi.spice
* Created: Fri Aug 28 17:33:10 2020
* 
x_PM_SKY130_FD_SC_MS__EINVN_2%TE_B N_TE_B_c_68_n N_TE_B_c_73_n N_TE_B_M1006_g
+ N_TE_B_M1009_g N_TE_B_c_75_n N_TE_B_c_76_n N_TE_B_c_77_n N_TE_B_M1002_g
+ N_TE_B_c_78_n N_TE_B_c_79_n N_TE_B_M1003_g N_TE_B_c_80_n TE_B TE_B
+ N_TE_B_c_70_n N_TE_B_c_71_n PM_SKY130_FD_SC_MS__EINVN_2%TE_B
x_PM_SKY130_FD_SC_MS__EINVN_2%A_117_74# N_A_117_74#_M1009_d N_A_117_74#_M1006_d
+ N_A_117_74#_c_131_n N_A_117_74#_M1000_g N_A_117_74#_c_133_n
+ N_A_117_74#_M1007_g N_A_117_74#_c_135_n N_A_117_74#_c_141_n
+ N_A_117_74#_c_136_n N_A_117_74#_c_137_n N_A_117_74#_c_138_n
+ N_A_117_74#_c_139_n N_A_117_74#_c_140_n PM_SKY130_FD_SC_MS__EINVN_2%A_117_74#
x_PM_SKY130_FD_SC_MS__EINVN_2%A N_A_c_190_n N_A_M1001_g N_A_M1004_g N_A_c_192_n
+ N_A_M1008_g N_A_M1005_g N_A_c_194_n A A N_A_c_196_n N_A_c_197_n
+ PM_SKY130_FD_SC_MS__EINVN_2%A
x_PM_SKY130_FD_SC_MS__EINVN_2%VPWR N_VPWR_M1006_s N_VPWR_M1002_d N_VPWR_c_242_n
+ N_VPWR_c_243_n N_VPWR_c_244_n VPWR N_VPWR_c_245_n N_VPWR_c_246_n
+ N_VPWR_c_241_n N_VPWR_c_248_n PM_SKY130_FD_SC_MS__EINVN_2%VPWR
x_PM_SKY130_FD_SC_MS__EINVN_2%A_227_368# N_A_227_368#_M1002_s
+ N_A_227_368#_M1003_s N_A_227_368#_M1005_s N_A_227_368#_c_279_n
+ N_A_227_368#_c_280_n N_A_227_368#_c_281_n N_A_227_368#_c_282_n
+ N_A_227_368#_c_292_n N_A_227_368#_c_283_n N_A_227_368#_c_284_n
+ N_A_227_368#_c_285_n PM_SKY130_FD_SC_MS__EINVN_2%A_227_368#
x_PM_SKY130_FD_SC_MS__EINVN_2%Z N_Z_M1001_s N_Z_M1004_d Z Z Z Z Z
+ PM_SKY130_FD_SC_MS__EINVN_2%Z
x_PM_SKY130_FD_SC_MS__EINVN_2%VGND N_VGND_M1009_s N_VGND_M1000_d N_VGND_c_355_n
+ N_VGND_c_356_n N_VGND_c_357_n VGND N_VGND_c_358_n N_VGND_c_359_n
+ N_VGND_c_360_n N_VGND_c_361_n PM_SKY130_FD_SC_MS__EINVN_2%VGND
x_PM_SKY130_FD_SC_MS__EINVN_2%A_231_74# N_A_231_74#_M1000_s N_A_231_74#_M1007_s
+ N_A_231_74#_M1008_d N_A_231_74#_c_392_n N_A_231_74#_c_393_n
+ N_A_231_74#_c_394_n N_A_231_74#_c_395_n N_A_231_74#_c_396_n
+ PM_SKY130_FD_SC_MS__EINVN_2%A_231_74#
cc_1 VNB N_TE_B_c_68_n 0.0305908f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.948
cc_2 VNB N_TE_B_M1009_g 0.0431726f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_3 VNB N_TE_B_c_70_n 0.0227507f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_4 VNB N_TE_B_c_71_n 0.0261838f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_5 VNB N_A_117_74#_c_131_n 0.0174569f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.12
cc_6 VNB N_A_117_74#_M1000_g 0.0270981f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=3.11
cc_7 VNB N_A_117_74#_c_133_n 0.0224188f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=3.035
cc_8 VNB N_A_117_74#_M1007_g 0.021718f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=3.11
cc_9 VNB N_A_117_74#_c_135_n 0.00513534f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_10 VNB N_A_117_74#_c_136_n 0.0111828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_117_74#_c_137_n 0.0121801f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.12
cc_12 VNB N_A_117_74#_c_138_n 7.13956e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.965
cc_13 VNB N_A_117_74#_c_139_n 0.0095065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_117_74#_c_140_n 0.0497031f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.965
cc_15 VNB N_A_c_190_n 0.0172813f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.302
cc_16 VNB N_A_M1004_g 0.0200758f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.64
cc_17 VNB N_A_c_192_n 0.020506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_M1005_g 0.00913677f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_19 VNB N_A_c_194_n 0.00694111f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=3.11
cc_20 VNB A 0.02299f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=3.035
cc_21 VNB N_A_c_196_n 0.0135987f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_c_197_n 0.0587014f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.285
cc_23 VNB N_VPWR_c_241_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_24 VNB Z 5.654e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.12
cc_25 VNB Z 0.00184709f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_26 VNB N_VGND_c_355_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.12
cc_27 VNB N_VGND_c_356_n 0.0310923f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.58
cc_28 VNB N_VGND_c_357_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=3.035
cc_29 VNB N_VGND_c_358_n 0.0329878f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=3.11
cc_30 VNB N_VGND_c_359_n 0.0398307f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_31 VNB N_VGND_c_360_n 0.21764f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.285
cc_32 VNB N_VGND_c_361_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_231_74#_c_392_n 0.00810194f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=3.11
cc_34 VNB N_A_231_74#_c_393_n 0.0085596f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_35 VNB N_A_231_74#_c_394_n 0.00413418f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_36 VNB N_A_231_74#_c_395_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=3.11
cc_37 VNB N_A_231_74#_c_396_n 0.015961f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_38 VPB N_TE_B_c_68_n 0.0262002f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.948
cc_39 VPB N_TE_B_c_73_n 0.0356711f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.28
cc_40 VPB N_TE_B_M1006_g 0.00919986f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.64
cc_41 VPB N_TE_B_c_75_n 0.06053f $X=-0.19 $Y=1.66 $X2=1.415 $Y2=3.11
cc_42 VPB N_TE_B_c_76_n 0.013638f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=3.11
cc_43 VPB N_TE_B_c_77_n 0.0170338f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=3.035
cc_44 VPB N_TE_B_c_78_n 0.0277408f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=3.11
cc_45 VPB N_TE_B_c_79_n 0.014211f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=3.035
cc_46 VPB N_TE_B_c_80_n 0.00887809f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=3.11
cc_47 VPB N_TE_B_c_71_n 0.0223278f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_48 VPB N_A_117_74#_c_141_n 0.0133719f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_49 VPB N_A_117_74#_c_138_n 0.0138267f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.965
cc_50 VPB N_A_M1004_g 0.0226013f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.64
cc_51 VPB N_A_M1005_g 0.0286915f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_52 VPB N_VPWR_c_242_n 0.0104926f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.12
cc_53 VPB N_VPWR_c_243_n 0.0392007f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.58
cc_54 VPB N_VPWR_c_244_n 0.00196645f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=3.035
cc_55 VPB N_VPWR_c_245_n 0.0332027f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=3.11
cc_56 VPB N_VPWR_c_246_n 0.0386225f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_57 VPB N_VPWR_c_241_n 0.0531475f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.285
cc_58 VPB N_VPWR_c_248_n 0.00345125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_227_368#_c_279_n 0.00455148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_227_368#_c_280_n 0.0106796f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=3.11
cc_61 VPB N_A_227_368#_c_281_n 0.00313047f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_62 VPB N_A_227_368#_c_282_n 0.00565977f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=3.11
cc_63 VPB N_A_227_368#_c_283_n 0.0117061f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_64 VPB N_A_227_368#_c_284_n 0.00181992f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=3.11
cc_65 VPB N_A_227_368#_c_285_n 0.0427455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB Z 0.00153131f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.58
cc_67 N_TE_B_c_77_n N_A_117_74#_c_131_n 0.0112153f $X=1.505 $Y=3.035 $X2=0 $Y2=0
cc_68 N_TE_B_c_79_n N_A_117_74#_c_133_n 0.00981278f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_69 N_TE_B_M1006_g N_A_117_74#_c_141_n 0.0110866f $X=0.5 $Y=2.64 $X2=0 $Y2=0
cc_70 N_TE_B_c_75_n N_A_117_74#_c_141_n 0.00520959f $X=1.415 $Y=3.11 $X2=0 $Y2=0
cc_71 N_TE_B_M1009_g N_A_117_74#_c_136_n 0.0157368f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_72 N_TE_B_c_71_n N_A_117_74#_c_136_n 0.0152878f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_73 N_TE_B_M1009_g N_A_117_74#_c_137_n 0.00786676f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_74 N_TE_B_c_68_n N_A_117_74#_c_138_n 0.0135983f $X=0.402 $Y=1.948 $X2=0 $Y2=0
cc_75 N_TE_B_c_73_n N_A_117_74#_c_138_n 0.00397887f $X=0.5 $Y=2.28 $X2=0 $Y2=0
cc_76 N_TE_B_c_77_n N_A_117_74#_c_138_n 0.00295653f $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_77 N_TE_B_c_71_n N_A_117_74#_c_138_n 0.0367453f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_78 N_TE_B_c_68_n N_A_117_74#_c_139_n 0.00223631f $X=0.402 $Y=1.948 $X2=0
+ $Y2=0
cc_79 N_TE_B_c_71_n N_A_117_74#_c_139_n 0.0271789f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_80 N_TE_B_c_68_n N_A_117_74#_c_140_n 0.0170189f $X=0.402 $Y=1.948 $X2=0 $Y2=0
cc_81 N_TE_B_c_71_n N_A_117_74#_c_140_n 3.17368e-19 $X=0.385 $Y=1.285 $X2=0
+ $Y2=0
cc_82 N_TE_B_c_79_n N_A_M1004_g 0.0146013f $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_83 N_TE_B_c_73_n N_VPWR_c_243_n 0.00108702f $X=0.5 $Y=2.28 $X2=0 $Y2=0
cc_84 N_TE_B_M1006_g N_VPWR_c_243_n 0.00945243f $X=0.5 $Y=2.64 $X2=0 $Y2=0
cc_85 N_TE_B_c_71_n N_VPWR_c_243_n 0.0212001f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_86 N_TE_B_c_77_n N_VPWR_c_244_n 0.0129118f $X=1.505 $Y=3.035 $X2=0 $Y2=0
cc_87 N_TE_B_c_78_n N_VPWR_c_244_n 0.0121909f $X=1.865 $Y=3.11 $X2=0 $Y2=0
cc_88 N_TE_B_c_79_n N_VPWR_c_244_n 0.00100539f $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_89 N_TE_B_c_80_n N_VPWR_c_244_n 0.00515868f $X=1.505 $Y=3.11 $X2=0 $Y2=0
cc_90 N_TE_B_c_76_n N_VPWR_c_245_n 0.032251f $X=0.59 $Y=3.11 $X2=0 $Y2=0
cc_91 N_TE_B_c_78_n N_VPWR_c_246_n 0.00790132f $X=1.865 $Y=3.11 $X2=0 $Y2=0
cc_92 N_TE_B_c_75_n N_VPWR_c_241_n 0.0276032f $X=1.415 $Y=3.11 $X2=0 $Y2=0
cc_93 N_TE_B_c_76_n N_VPWR_c_241_n 0.011317f $X=0.59 $Y=3.11 $X2=0 $Y2=0
cc_94 N_TE_B_c_78_n N_VPWR_c_241_n 0.0145046f $X=1.865 $Y=3.11 $X2=0 $Y2=0
cc_95 N_TE_B_c_80_n N_VPWR_c_241_n 0.0100223f $X=1.505 $Y=3.11 $X2=0 $Y2=0
cc_96 N_TE_B_M1006_g N_A_227_368#_c_280_n 0.00122589f $X=0.5 $Y=2.64 $X2=0 $Y2=0
cc_97 N_TE_B_c_75_n N_A_227_368#_c_280_n 0.00521258f $X=1.415 $Y=3.11 $X2=0
+ $Y2=0
cc_98 N_TE_B_c_77_n N_A_227_368#_c_280_n 0.00152914f $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_99 N_TE_B_c_77_n N_A_227_368#_c_281_n 0.0155988f $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_100 N_TE_B_c_79_n N_A_227_368#_c_281_n 0.0133819f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_101 N_TE_B_c_79_n N_A_227_368#_c_282_n 0.00122083f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_102 N_TE_B_c_77_n N_A_227_368#_c_292_n 7.19888e-19 $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_79_n N_A_227_368#_c_292_n 0.0126556f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_104 N_TE_B_c_78_n N_A_227_368#_c_284_n 0.00143645f $X=1.865 $Y=3.11 $X2=0
+ $Y2=0
cc_105 N_TE_B_c_79_n N_A_227_368#_c_284_n 0.00237275f $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_106 N_TE_B_c_79_n Z 5.21901e-19 $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_107 N_TE_B_c_79_n Z 2.7754e-19 $X=1.955 $Y=3.035 $X2=0 $Y2=0
cc_108 N_TE_B_M1009_g N_VGND_c_356_n 0.00589946f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_109 N_TE_B_c_70_n N_VGND_c_356_n 0.00115809f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_110 N_TE_B_c_71_n N_VGND_c_356_n 0.0145115f $X=0.385 $Y=1.285 $X2=0 $Y2=0
cc_111 N_TE_B_M1009_g N_VGND_c_358_n 0.00434272f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_112 N_TE_B_M1009_g N_VGND_c_360_n 0.00828991f $X=0.51 $Y=0.58 $X2=0 $Y2=0
cc_113 N_TE_B_M1009_g N_A_231_74#_c_392_n 9.23906e-19 $X=0.51 $Y=0.58 $X2=0
+ $Y2=0
cc_114 N_TE_B_c_77_n N_A_231_74#_c_393_n 4.36843e-19 $X=1.505 $Y=3.035 $X2=0
+ $Y2=0
cc_115 N_TE_B_c_79_n N_A_231_74#_c_393_n 9.30886e-19 $X=1.955 $Y=3.035 $X2=0
+ $Y2=0
cc_116 N_A_117_74#_M1007_g N_A_c_190_n 0.0104506f $X=1.945 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_117_74#_c_133_n N_A_M1004_g 0.00490479f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_118 N_A_117_74#_c_133_n N_A_c_194_n 0.0104506f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_119 N_A_117_74#_c_141_n N_VPWR_c_243_n 0.0237219f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_117_74#_c_141_n N_VPWR_c_245_n 0.0145399f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_117_74#_c_141_n N_VPWR_c_241_n 0.010749f $X=0.725 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_117_74#_c_131_n N_A_227_368#_c_279_n 0.00507112f $X=1.44 $Y=1.395
+ $X2=0 $Y2=0
cc_123 N_A_117_74#_c_138_n N_A_227_368#_c_279_n 0.0117903f $X=0.725 $Y=2.3 $X2=0
+ $Y2=0
cc_124 N_A_117_74#_c_139_n N_A_227_368#_c_279_n 0.003795f $X=0.995 $Y=1.485
+ $X2=0 $Y2=0
cc_125 N_A_117_74#_c_140_n N_A_227_368#_c_279_n 0.0010483f $X=0.995 $Y=1.395
+ $X2=0 $Y2=0
cc_126 N_A_117_74#_c_138_n N_A_227_368#_c_280_n 0.0659094f $X=0.725 $Y=2.3 $X2=0
+ $Y2=0
cc_127 N_A_117_74#_c_131_n N_A_227_368#_c_281_n 9.88525e-19 $X=1.44 $Y=1.395
+ $X2=0 $Y2=0
cc_128 N_A_117_74#_c_133_n N_A_227_368#_c_281_n 0.00679491f $X=1.87 $Y=1.395
+ $X2=0 $Y2=0
cc_129 N_A_117_74#_M1007_g Z 0.00127446f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_117_74#_c_137_n N_VGND_c_356_n 0.0179429f $X=0.725 $Y=0.58 $X2=0
+ $Y2=0
cc_131 N_A_117_74#_M1000_g N_VGND_c_357_n 0.012411f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_117_74#_M1007_g N_VGND_c_357_n 0.00950277f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_133 N_A_117_74#_M1000_g N_VGND_c_358_n 0.00383152f $X=1.515 $Y=0.74 $X2=0
+ $Y2=0
cc_134 N_A_117_74#_c_137_n N_VGND_c_358_n 0.0143708f $X=0.725 $Y=0.58 $X2=0
+ $Y2=0
cc_135 N_A_117_74#_M1007_g N_VGND_c_359_n 0.00383152f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_117_74#_M1000_g N_VGND_c_360_n 0.00762539f $X=1.515 $Y=0.74 $X2=0
+ $Y2=0
cc_137 N_A_117_74#_M1007_g N_VGND_c_360_n 0.00757637f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_117_74#_c_137_n N_VGND_c_360_n 0.011923f $X=0.725 $Y=0.58 $X2=0 $Y2=0
cc_139 N_A_117_74#_M1000_g N_A_231_74#_c_392_n 0.00159319f $X=1.515 $Y=0.74
+ $X2=0 $Y2=0
cc_140 N_A_117_74#_c_137_n N_A_231_74#_c_392_n 0.039239f $X=0.725 $Y=0.58 $X2=0
+ $Y2=0
cc_141 N_A_117_74#_c_131_n N_A_231_74#_c_393_n 0.00129671f $X=1.44 $Y=1.395
+ $X2=0 $Y2=0
cc_142 N_A_117_74#_M1000_g N_A_231_74#_c_393_n 0.0141996f $X=1.515 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_117_74#_c_133_n N_A_231_74#_c_393_n 0.00240153f $X=1.87 $Y=1.395
+ $X2=0 $Y2=0
cc_144 N_A_117_74#_M1007_g N_A_231_74#_c_393_n 0.0138232f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_117_74#_c_136_n N_A_231_74#_c_394_n 0.0111139f $X=0.805 $Y=1.32 $X2=0
+ $Y2=0
cc_146 N_A_117_74#_c_139_n N_A_231_74#_c_394_n 0.00210833f $X=0.995 $Y=1.485
+ $X2=0 $Y2=0
cc_147 N_A_117_74#_c_140_n N_A_231_74#_c_394_n 0.00660264f $X=0.995 $Y=1.395
+ $X2=0 $Y2=0
cc_148 N_A_M1004_g N_VPWR_c_246_n 0.00333926f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_M1005_g N_VPWR_c_246_n 0.00333926f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1004_g N_VPWR_c_241_n 0.00422798f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_M1005_g N_VPWR_c_241_n 0.00426429f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_M1004_g N_A_227_368#_c_283_n 0.0139961f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_M1005_g N_A_227_368#_c_283_n 0.0149887f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_M1005_g N_A_227_368#_c_285_n 0.00151667f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_155 A N_A_227_368#_c_285_n 0.0175067f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_156 N_A_c_197_n N_A_227_368#_c_285_n 0.00207994f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_157 N_A_c_190_n Z 0.00549559f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A_c_192_n Z 0.00558139f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_159 A Z 0.0443015f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_160 N_A_c_190_n Z 0.00212163f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_M1004_g Z 0.0188477f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_c_192_n Z 0.00179582f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A_M1005_g Z 0.0075403f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_c_194_n Z 0.00290588f $X=2.397 $Y=1.295 $X2=0 $Y2=0
cc_165 N_A_c_196_n Z 0.0115492f $X=2.735 $Y=1.385 $X2=0 $Y2=0
cc_166 N_A_c_197_n Z 0.00756257f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A_M1004_g Z 0.00206313f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A_M1005_g Z 0.0036649f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_c_197_n Z 4.34692e-19 $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_170 N_A_M1004_g Z 0.00874145f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_M1005_g Z 0.00919522f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_c_190_n N_VGND_c_357_n 6.35276e-19 $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_173 N_A_c_190_n N_VGND_c_359_n 0.00291649f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A_c_192_n N_VGND_c_359_n 0.00291649f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_c_190_n N_VGND_c_360_n 0.00359269f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_176 N_A_c_192_n N_VGND_c_360_n 0.00363003f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_177 A N_VGND_c_360_n 0.00283239f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_178 A N_A_231_74#_M1008_d 0.00476174f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_179 N_A_c_190_n N_A_231_74#_c_393_n 3.43633e-19 $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_180 N_A_c_190_n N_A_231_74#_c_396_n 0.0142515f $X=2.375 $Y=1.22 $X2=0 $Y2=0
cc_181 N_A_c_192_n N_A_231_74#_c_396_n 0.0145459f $X=2.81 $Y=1.22 $X2=0 $Y2=0
cc_182 A N_A_231_74#_c_396_n 0.017603f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_183 N_A_c_196_n N_A_231_74#_c_396_n 3.11327e-19 $X=2.735 $Y=1.385 $X2=0 $Y2=0
cc_184 N_A_c_197_n N_A_231_74#_c_396_n 8.44951e-19 $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_185 N_VPWR_c_244_n N_A_227_368#_c_280_n 0.0286421f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_245_n N_A_227_368#_c_280_n 0.0126187f $X=1.58 $Y=3.33 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_241_n N_A_227_368#_c_280_n 0.00931741f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_188 N_VPWR_M1002_d N_A_227_368#_c_281_n 0.00165831f $X=1.595 $Y=1.84 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_244_n N_A_227_368#_c_281_n 0.0137163f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_246_n N_A_227_368#_c_283_n 0.0621263f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_241_n N_A_227_368#_c_283_n 0.03443f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_192 N_VPWR_c_244_n N_A_227_368#_c_284_n 0.0101196f $X=1.73 $Y=2.325 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_246_n N_A_227_368#_c_284_n 0.0199669f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_241_n N_A_227_368#_c_284_n 0.0107485f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_A_227_368#_c_283_n N_Z_M1004_d 0.00165831f $X=2.965 $Y=2.99 $X2=0 $Y2=0
cc_196 N_A_227_368#_c_282_n Z 0.00725715f $X=2.155 $Y=1.99 $X2=0 $Y2=0
cc_197 N_A_227_368#_c_285_n Z 0.0350665f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_227_368#_c_283_n Z 0.0159318f $X=2.965 $Y=2.99 $X2=0 $Y2=0
cc_199 N_A_227_368#_c_279_n N_A_231_74#_c_393_n 4.64785e-19 $X=1.257 $Y=1.99
+ $X2=0 $Y2=0
cc_200 N_A_227_368#_c_281_n N_A_231_74#_c_393_n 0.0153714f $X=2.015 $Y=1.905
+ $X2=0 $Y2=0
cc_201 N_A_227_368#_c_282_n N_A_231_74#_c_393_n 0.00784312f $X=2.155 $Y=1.99
+ $X2=0 $Y2=0
cc_202 N_A_227_368#_c_279_n N_A_231_74#_c_394_n 0.0079427f $X=1.257 $Y=1.99
+ $X2=0 $Y2=0
cc_203 Z N_A_231_74#_c_393_n 0.00625076f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_204 Z N_A_231_74#_c_393_n 0.00142622f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_205 N_Z_M1001_s N_A_231_74#_c_396_n 0.00174803f $X=2.45 $Y=0.37 $X2=0 $Y2=0
cc_206 Z N_A_231_74#_c_396_n 0.0168802f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_207 N_VGND_c_357_n N_A_231_74#_c_392_n 0.0164982f $X=1.73 $Y=0.61 $X2=0 $Y2=0
cc_208 N_VGND_c_358_n N_A_231_74#_c_392_n 0.011066f $X=1.565 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_360_n N_A_231_74#_c_392_n 0.00915947f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_M1000_d N_A_231_74#_c_393_n 0.00184993f $X=1.59 $Y=0.37 $X2=0
+ $Y2=0
cc_211 N_VGND_c_357_n N_A_231_74#_c_393_n 0.0156953f $X=1.73 $Y=0.61 $X2=0 $Y2=0
cc_212 N_VGND_c_357_n N_A_231_74#_c_395_n 0.00985092f $X=1.73 $Y=0.61 $X2=0
+ $Y2=0
cc_213 N_VGND_c_359_n N_A_231_74#_c_395_n 0.00758556f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_214 N_VGND_c_360_n N_A_231_74#_c_395_n 0.00627867f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_359_n N_A_231_74#_c_396_n 0.038742f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_360_n N_A_231_74#_c_396_n 0.0327013f $X=3.12 $Y=0 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlxtp_1 D GATE VGND VNB VPB VPWR Q
M1000 Q a_386_326# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.60698e+12p ps=1.245e+07u
M1001 VGND a_119_88# a_239_85# VNB nlowvt w=740000u l=150000u
+  ad=1.47895e+12p pd=1.06e+07u as=4.458e+11p ps=4.22e+06u
M1002 a_422_392# a_386_326# VPWR VPB pshort w=420000u l=180000u
+  ad=3.0425e+11p pd=3.2e+06u as=0p ps=0u
M1003 a_685_59# a_562_123# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 a_592_149# a_562_123# a_514_149# VNB nlowvt w=420000u l=150000u
+  ad=2.753e+11p pd=2.41e+06u as=1.008e+11p ps=1.32e+06u
M1005 Q a_386_326# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_119_88# D VGND VNB nlowvt w=550000u l=150000u
+  ad=1.815e+11p pd=1.76e+06u as=0p ps=0u
M1007 VPWR a_119_88# a_229_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1008 a_119_88# D VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1009 VGND a_592_149# a_386_326# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1010 VPWR a_592_149# a_386_326# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.528e+11p ps=2.87e+06u
M1011 a_685_59# a_562_123# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 VPWR GATE a_562_123# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 a_592_149# a_562_123# a_229_392# VPB pshort w=1e+06u l=180000u
+  ad=3.115e+11p pd=2.71e+06u as=0p ps=0u
M1014 a_514_149# a_386_326# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_239_85# a_685_59# a_592_149# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND GATE a_562_123# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.22e+11p ps=2.08e+06u
M1017 a_422_392# a_685_59# a_592_149# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

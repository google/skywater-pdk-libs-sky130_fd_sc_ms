* File: sky130_fd_sc_ms__einvp_2.pxi.spice
* Created: Fri Aug 28 17:34:07 2020
* 
x_PM_SKY130_FD_SC_MS__EINVP_2%A N_A_M1003_g N_A_c_73_n N_A_M1001_g N_A_M1004_g
+ N_A_c_75_n N_A_M1009_g A N_A_c_77_n PM_SKY130_FD_SC_MS__EINVP_2%A
x_PM_SKY130_FD_SC_MS__EINVP_2%A_263_323# N_A_263_323#_M1000_s
+ N_A_263_323#_M1002_s N_A_263_323#_c_122_n N_A_263_323#_M1005_g
+ N_A_263_323#_c_115_n N_A_263_323#_c_116_n N_A_263_323#_c_125_n
+ N_A_263_323#_M1006_g N_A_263_323#_c_117_n N_A_263_323#_c_118_n
+ N_A_263_323#_c_119_n N_A_263_323#_c_120_n N_A_263_323#_c_121_n
+ PM_SKY130_FD_SC_MS__EINVP_2%A_263_323#
x_PM_SKY130_FD_SC_MS__EINVP_2%TE N_TE_c_174_n N_TE_M1007_g N_TE_c_175_n
+ N_TE_c_176_n N_TE_c_177_n N_TE_M1008_g N_TE_c_178_n N_TE_c_179_n N_TE_c_186_n
+ N_TE_M1002_g N_TE_M1000_g N_TE_c_181_n N_TE_c_182_n N_TE_c_188_n N_TE_c_183_n
+ TE N_TE_c_184_n N_TE_c_185_n PM_SKY130_FD_SC_MS__EINVP_2%TE
x_PM_SKY130_FD_SC_MS__EINVP_2%A_27_368# N_A_27_368#_M1003_s N_A_27_368#_M1004_s
+ N_A_27_368#_M1006_s N_A_27_368#_c_240_n N_A_27_368#_c_241_n
+ N_A_27_368#_c_242_n N_A_27_368#_c_243_n N_A_27_368#_c_238_n
+ N_A_27_368#_c_239_n N_A_27_368#_c_244_n PM_SKY130_FD_SC_MS__EINVP_2%A_27_368#
x_PM_SKY130_FD_SC_MS__EINVP_2%Z N_Z_M1001_s N_Z_M1003_d N_Z_c_286_n Z Z Z Z Z
+ PM_SKY130_FD_SC_MS__EINVP_2%Z
x_PM_SKY130_FD_SC_MS__EINVP_2%VPWR N_VPWR_M1005_d N_VPWR_M1002_d N_VPWR_c_310_n
+ N_VPWR_c_311_n N_VPWR_c_312_n VPWR N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_315_n N_VPWR_c_309_n PM_SKY130_FD_SC_MS__EINVP_2%VPWR
x_PM_SKY130_FD_SC_MS__EINVP_2%A_36_74# N_A_36_74#_M1001_d N_A_36_74#_M1009_d
+ N_A_36_74#_M1008_s N_A_36_74#_c_345_n N_A_36_74#_c_346_n N_A_36_74#_c_347_n
+ N_A_36_74#_c_348_n N_A_36_74#_c_349_n N_A_36_74#_c_350_n N_A_36_74#_c_351_n
+ PM_SKY130_FD_SC_MS__EINVP_2%A_36_74#
x_PM_SKY130_FD_SC_MS__EINVP_2%VGND N_VGND_M1007_d N_VGND_M1000_d N_VGND_c_393_n
+ N_VGND_c_394_n N_VGND_c_395_n VGND N_VGND_c_396_n N_VGND_c_397_n
+ N_VGND_c_398_n N_VGND_c_399_n PM_SKY130_FD_SC_MS__EINVP_2%VGND
cc_1 VNB N_A_M1003_g 0.00913677f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_c_73_n 0.0203982f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.22
cc_3 VNB N_A_M1004_g 0.00570466f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_4 VNB N_A_c_75_n 0.0159117f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.22
cc_5 VNB A 0.0113831f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A_c_77_n 0.0876648f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.385
cc_7 VNB N_A_263_323#_c_115_n 0.00485002f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_8 VNB N_A_263_323#_c_116_n 0.00403751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_263_323#_c_117_n 0.00324064f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_10 VNB N_A_263_323#_c_118_n 0.0160163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_263_323#_c_119_n 0.0164879f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_12 VNB N_A_263_323#_c_120_n 0.00526886f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_A_263_323#_c_121_n 0.00987396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_TE_c_174_n 0.0145546f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_15 VNB N_TE_c_175_n 0.0126935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_TE_c_176_n 0.00751923f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.22
cc_17 VNB N_TE_c_177_n 0.0161538f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_18 VNB N_TE_c_178_n 0.026203f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_19 VNB N_TE_c_179_n 0.0333291f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.22
cc_20 VNB N_TE_M1000_g 0.0120118f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_21 VNB N_TE_c_181_n 0.0251423f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_22 VNB N_TE_c_182_n 0.00535066f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.385
cc_23 VNB N_TE_c_183_n 0.0342067f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_24 VNB N_TE_c_184_n 0.0588596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_TE_c_185_n 0.00566583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_368#_c_238_n 0.00845447f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.385
cc_27 VNB N_A_27_368#_c_239_n 0.00299021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Z_c_286_n 6.47547e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_29 VNB Z 0.0033102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_309_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_36_74#_c_345_n 0.0222939f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.22
cc_32 VNB N_A_36_74#_c_346_n 0.00449328f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_33 VNB N_A_36_74#_c_347_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_A_36_74#_c_348_n 4.66303e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_35 VNB N_A_36_74#_c_349_n 0.00668482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_36_74#_c_350_n 0.00289968f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_37 VNB N_A_36_74#_c_351_n 0.00892448f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.385
cc_38 VNB N_VGND_c_393_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_39 VNB N_VGND_c_394_n 0.0109649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_395_n 0.0418368f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_41 VNB N_VGND_c_396_n 0.0374035f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_42 VNB N_VGND_c_397_n 0.0327804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_398_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_399_n 0.215736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_M1003_g 0.0287872f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_46 VPB N_A_M1004_g 0.0211045f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_47 VPB N_A_263_323#_c_122_n 0.0164048f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=0.74
cc_48 VPB N_A_263_323#_c_115_n 0.00490076f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_49 VPB N_A_263_323#_c_116_n 0.00403299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_263_323#_c_125_n 0.0206017f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.22
cc_51 VPB N_A_263_323#_c_117_n 0.00200584f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_52 VPB N_A_263_323#_c_118_n 0.0236283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_263_323#_c_119_n 0.0242097f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_54 VPB N_A_263_323#_c_121_n 0.0232301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_TE_c_186_n 0.0238811f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=0.74
cc_56 VPB N_TE_c_181_n 0.0347972f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_57 VPB N_TE_c_188_n 0.0335451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_27_368#_c_240_n 0.0419704f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.22
cc_59 VPB N_A_27_368#_c_241_n 0.00472187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_368#_c_242_n 0.00929469f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_61 VPB N_A_27_368#_c_243_n 0.00280583f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_62 VPB N_A_27_368#_c_244_n 0.00261492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB Z 0.00199987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_310_n 0.00714653f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_65 VPB N_VPWR_c_311_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=0.74
cc_66 VPB N_VPWR_c_312_n 0.0415571f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_67 VPB N_VPWR_c_313_n 0.0374994f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_68 VPB N_VPWR_c_314_n 0.0334651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_315_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_309_n 0.0706486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_A_263_323#_c_116_n 0.0167059f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A_c_75_n N_TE_c_174_n 0.00855951f $X=0.97 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_73 N_A_c_77_n N_TE_c_176_n 0.00855951f $X=0.97 $Y=1.385 $X2=0 $Y2=0
cc_74 N_A_M1003_g N_A_27_368#_c_240_n 0.00148512f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_75 A N_A_27_368#_c_240_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_c_77_n N_A_27_368#_c_240_n 0.00185549f $X=0.97 $Y=1.385 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_A_27_368#_c_241_n 0.0158369f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_A_27_368#_c_241_n 0.0129371f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_M1004_g N_A_27_368#_c_243_n 0.00157246f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_c_77_n N_A_27_368#_c_239_n 0.00404856f $X=0.97 $Y=1.385 $X2=0 $Y2=0
cc_81 N_A_c_73_n N_Z_c_286_n 0.00215527f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_82 N_A_c_75_n N_Z_c_286_n 0.00757448f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A_M1003_g Z 0.00877997f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_c_73_n Z 0.00131177f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_85 N_A_M1004_g Z 0.0208268f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_c_75_n Z 8.7164e-19 $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_87 A Z 0.0277568f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A_c_77_n Z 0.0264139f $X=0.97 $Y=1.385 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VPWR_c_313_n 0.00333926f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_M1004_g N_VPWR_c_313_n 0.00333926f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VPWR_c_309_n 0.00426429f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_M1004_g N_VPWR_c_309_n 0.00422798f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A_c_73_n N_A_36_74#_c_345_n 0.00929919f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A_c_75_n N_A_36_74#_c_345_n 6.05004e-19 $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_95 A N_A_36_74#_c_345_n 0.0228393f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A_c_77_n N_A_36_74#_c_345_n 0.00186408f $X=0.97 $Y=1.385 $X2=0 $Y2=0
cc_97 N_A_c_73_n N_A_36_74#_c_346_n 0.0100245f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_98 N_A_c_75_n N_A_36_74#_c_346_n 0.0120332f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_99 N_A_c_73_n N_A_36_74#_c_347_n 0.00282152f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_100 N_A_c_75_n N_A_36_74#_c_348_n 4.60747e-19 $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A_c_75_n N_A_36_74#_c_350_n 0.0015676f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A_c_73_n N_VGND_c_396_n 0.00278247f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_103 N_A_c_75_n N_VGND_c_396_n 0.00278271f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_104 N_A_c_73_n N_VGND_c_399_n 0.00357229f $X=0.54 $Y=1.22 $X2=0 $Y2=0
cc_105 N_A_c_75_n N_VGND_c_399_n 0.00353526f $X=0.97 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A_263_323#_c_115_n N_TE_c_175_n 0.0126826f $X=1.765 $Y=1.69 $X2=0 $Y2=0
cc_107 N_A_263_323#_c_116_n N_TE_c_176_n 0.0126826f $X=1.495 $Y=1.69 $X2=0 $Y2=0
cc_108 N_A_263_323#_c_118_n N_TE_c_178_n 0.00297448f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_109 N_A_263_323#_c_121_n N_TE_c_178_n 0.0126826f $X=2.415 $Y=1.72 $X2=0 $Y2=0
cc_110 N_A_263_323#_c_120_n N_TE_c_179_n 0.00297448f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_111 N_A_263_323#_c_118_n N_TE_M1000_g 0.00628076f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_112 N_A_263_323#_c_120_n N_TE_M1000_g 0.00915681f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_113 N_A_263_323#_c_118_n N_TE_c_181_n 0.0103964f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_114 N_A_263_323#_c_119_n N_TE_c_181_n 0.0190575f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_115 N_A_263_323#_c_117_n N_TE_c_182_n 0.0126826f $X=1.855 $Y=1.69 $X2=0 $Y2=0
cc_116 N_A_263_323#_c_118_n N_TE_c_188_n 0.0106318f $X=2.58 $Y=1.72 $X2=0 $Y2=0
cc_117 N_A_263_323#_c_120_n N_TE_c_184_n 0.00115908f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_118 N_A_263_323#_c_120_n N_TE_c_185_n 0.0247075f $X=2.635 $Y=0.95 $X2=0 $Y2=0
cc_119 N_A_263_323#_c_122_n N_A_27_368#_c_241_n 0.00101073f $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_120 N_A_263_323#_c_116_n N_A_27_368#_c_243_n 0.00274331f $X=1.495 $Y=1.69
+ $X2=0 $Y2=0
cc_121 N_A_263_323#_c_115_n N_A_27_368#_c_238_n 0.00743586f $X=1.765 $Y=1.69
+ $X2=0 $Y2=0
cc_122 N_A_263_323#_c_116_n N_A_27_368#_c_238_n 0.00931127f $X=1.495 $Y=1.69
+ $X2=0 $Y2=0
cc_123 N_A_263_323#_c_117_n N_A_27_368#_c_238_n 0.00842343f $X=1.855 $Y=1.69
+ $X2=0 $Y2=0
cc_124 N_A_263_323#_c_118_n N_A_27_368#_c_238_n 0.0109091f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_125 N_A_263_323#_c_119_n N_A_27_368#_c_238_n 0.00133801f $X=2.58 $Y=1.72
+ $X2=0 $Y2=0
cc_126 N_A_263_323#_c_121_n N_A_27_368#_c_238_n 0.00286087f $X=2.415 $Y=1.72
+ $X2=0 $Y2=0
cc_127 N_A_263_323#_c_122_n N_A_27_368#_c_244_n 5.70219e-19 $X=1.405 $Y=1.765
+ $X2=0 $Y2=0
cc_128 N_A_263_323#_c_125_n N_A_27_368#_c_244_n 0.0173866f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_129 N_A_263_323#_c_117_n N_A_27_368#_c_244_n 0.00331335f $X=1.855 $Y=1.69
+ $X2=0 $Y2=0
cc_130 N_A_263_323#_c_118_n N_A_27_368#_c_244_n 0.0796667f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_131 N_A_263_323#_c_119_n N_A_27_368#_c_244_n 9.96973e-19 $X=2.58 $Y=1.72
+ $X2=0 $Y2=0
cc_132 N_A_263_323#_c_121_n N_A_27_368#_c_244_n 0.00954193f $X=2.415 $Y=1.72
+ $X2=0 $Y2=0
cc_133 N_A_263_323#_c_116_n Z 3.52663e-19 $X=1.495 $Y=1.69 $X2=0 $Y2=0
cc_134 N_A_263_323#_c_122_n N_VPWR_c_310_n 0.0179164f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_263_323#_c_115_n N_VPWR_c_310_n 0.00207325f $X=1.765 $Y=1.69 $X2=0
+ $Y2=0
cc_136 N_A_263_323#_c_125_n N_VPWR_c_310_n 0.00334711f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_263_323#_c_118_n N_VPWR_c_312_n 0.0270962f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_138 N_A_263_323#_c_122_n N_VPWR_c_313_n 0.00460063f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_263_323#_c_125_n N_VPWR_c_314_n 0.005209f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_263_323#_c_118_n N_VPWR_c_314_n 0.0146357f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_141 N_A_263_323#_c_122_n N_VPWR_c_309_n 0.00908665f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_263_323#_c_125_n N_VPWR_c_309_n 0.00987399f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_263_323#_c_118_n N_VPWR_c_309_n 0.0121141f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_144 N_A_263_323#_c_116_n N_A_36_74#_c_349_n 6.55318e-19 $X=1.495 $Y=1.69
+ $X2=0 $Y2=0
cc_145 N_A_263_323#_c_118_n N_A_36_74#_c_349_n 0.0125516f $X=2.58 $Y=1.72 $X2=0
+ $Y2=0
cc_146 N_A_263_323#_c_121_n N_A_36_74#_c_349_n 4.74394e-19 $X=2.415 $Y=1.72
+ $X2=0 $Y2=0
cc_147 N_A_263_323#_c_120_n N_A_36_74#_c_351_n 0.0217181f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_148 N_A_263_323#_c_120_n N_VGND_c_399_n 0.0031213f $X=2.635 $Y=0.95 $X2=0
+ $Y2=0
cc_149 N_TE_c_176_n N_A_27_368#_c_238_n 0.00415283f $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_150 N_TE_c_178_n N_A_27_368#_c_238_n 0.00179693f $X=2.265 $Y=1.26 $X2=0 $Y2=0
cc_151 N_TE_c_174_n N_Z_c_286_n 2.18758e-19 $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_152 N_TE_c_176_n Z 2.10146e-19 $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_153 N_TE_c_186_n N_VPWR_c_312_n 0.0176457f $X=2.855 $Y=2.245 $X2=0 $Y2=0
cc_154 N_TE_c_188_n N_VPWR_c_312_n 0.0100919f $X=3.06 $Y=2.17 $X2=0 $Y2=0
cc_155 N_TE_c_186_n N_VPWR_c_314_n 0.00460063f $X=2.855 $Y=2.245 $X2=0 $Y2=0
cc_156 N_TE_c_186_n N_VPWR_c_309_n 0.00913687f $X=2.855 $Y=2.245 $X2=0 $Y2=0
cc_157 N_TE_c_174_n N_A_36_74#_c_346_n 9.48753e-19 $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_158 N_TE_c_174_n N_A_36_74#_c_348_n 9.29165e-19 $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_159 N_TE_c_174_n N_A_36_74#_c_349_n 0.00741157f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_160 N_TE_c_175_n N_A_36_74#_c_349_n 0.00615573f $X=1.755 $Y=1.26 $X2=0 $Y2=0
cc_161 N_TE_c_176_n N_A_36_74#_c_349_n 0.00364399f $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_162 N_TE_c_177_n N_A_36_74#_c_349_n 0.00753496f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_163 N_TE_c_178_n N_A_36_74#_c_349_n 0.0112425f $X=2.265 $Y=1.26 $X2=0 $Y2=0
cc_164 N_TE_c_179_n N_A_36_74#_c_349_n 4.36766e-19 $X=2.34 $Y=1.185 $X2=0 $Y2=0
cc_165 N_TE_c_182_n N_A_36_74#_c_349_n 0.00251882f $X=1.83 $Y=1.26 $X2=0 $Y2=0
cc_166 N_TE_c_177_n N_A_36_74#_c_351_n 0.00130964f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_167 N_TE_c_184_n N_A_36_74#_c_351_n 0.0106764f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_168 N_TE_c_185_n N_A_36_74#_c_351_n 0.0179335f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_169 N_TE_c_174_n N_VGND_c_393_n 0.0100283f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_170 N_TE_c_175_n N_VGND_c_393_n 7.11061e-19 $X=1.755 $Y=1.26 $X2=0 $Y2=0
cc_171 N_TE_c_177_n N_VGND_c_393_n 0.0134095f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_172 N_TE_c_183_n N_VGND_c_395_n 0.00727925f $X=3.06 $Y=1.27 $X2=0 $Y2=0
cc_173 N_TE_c_184_n N_VGND_c_395_n 0.0124285f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_174 N_TE_c_185_n N_VGND_c_395_n 0.0318479f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_175 N_TE_c_174_n N_VGND_c_396_n 0.00383152f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_176 N_TE_c_177_n N_VGND_c_397_n 0.00383152f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_177 N_TE_c_184_n N_VGND_c_397_n 0.0128697f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_178 N_TE_c_185_n N_VGND_c_397_n 0.0208821f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_179 N_TE_c_174_n N_VGND_c_399_n 0.00757637f $X=1.4 $Y=1.185 $X2=0 $Y2=0
cc_180 N_TE_c_177_n N_VGND_c_399_n 0.00762539f $X=1.83 $Y=1.185 $X2=0 $Y2=0
cc_181 N_TE_c_184_n N_VGND_c_399_n 0.011158f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_182 N_TE_c_185_n N_VGND_c_399_n 0.0123609f $X=2.645 $Y=0.425 $X2=0 $Y2=0
cc_183 N_A_27_368#_c_241_n N_Z_M1003_d 0.00165831f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_184 N_A_27_368#_c_240_n Z 0.00121195f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_27_368#_c_241_n Z 0.015684f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_186 N_A_27_368#_c_243_n Z 0.0464232f $X=1.18 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_27_368#_c_239_n Z 0.0139434f $X=1.265 $Y=1.565 $X2=0 $Y2=0
cc_188 N_A_27_368#_c_241_n N_VPWR_c_310_n 0.010126f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_189 N_A_27_368#_c_243_n N_VPWR_c_310_n 0.0348943f $X=1.18 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_27_368#_c_238_n N_VPWR_c_310_n 0.0198461f $X=1.915 $Y=1.565 $X2=0
+ $Y2=0
cc_191 N_A_27_368#_c_244_n N_VPWR_c_310_n 0.0379768f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_27_368#_c_241_n N_VPWR_c_313_n 0.0580334f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_193 N_A_27_368#_c_242_n N_VPWR_c_313_n 0.0179217f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_194 N_A_27_368#_c_244_n N_VPWR_c_314_n 0.0109793f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_27_368#_c_241_n N_VPWR_c_309_n 0.0323988f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_196 N_A_27_368#_c_242_n N_VPWR_c_309_n 0.00971942f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_197 N_A_27_368#_c_244_n N_VPWR_c_309_n 0.00901959f $X=2.08 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_27_368#_c_238_n N_A_36_74#_c_349_n 0.0681198f $X=1.915 $Y=1.565 $X2=0
+ $Y2=0
cc_199 N_A_27_368#_c_238_n N_A_36_74#_c_350_n 3.84494e-19 $X=1.915 $Y=1.565
+ $X2=0 $Y2=0
cc_200 N_A_27_368#_c_239_n N_A_36_74#_c_350_n 0.0154601f $X=1.265 $Y=1.565 $X2=0
+ $Y2=0
cc_201 N_Z_M1001_s N_A_36_74#_c_346_n 0.00189202f $X=0.615 $Y=0.37 $X2=0 $Y2=0
cc_202 N_Z_c_286_n N_A_36_74#_c_346_n 0.0124268f $X=0.755 $Y=0.82 $X2=0 $Y2=0
cc_203 N_Z_c_286_n N_A_36_74#_c_348_n 0.0187012f $X=0.755 $Y=0.82 $X2=0 $Y2=0
cc_204 N_Z_c_286_n N_A_36_74#_c_350_n 0.0135667f $X=0.755 $Y=0.82 $X2=0 $Y2=0
cc_205 N_A_36_74#_c_346_n N_VGND_c_393_n 0.0112234f $X=1.1 $Y=0.34 $X2=0 $Y2=0
cc_206 N_A_36_74#_c_349_n N_VGND_c_393_n 0.0216086f $X=1.95 $Y=1.225 $X2=0 $Y2=0
cc_207 N_A_36_74#_c_351_n N_VGND_c_393_n 0.0240263f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_A_36_74#_c_346_n N_VGND_c_396_n 0.050626f $X=1.1 $Y=0.34 $X2=0 $Y2=0
cc_209 N_A_36_74#_c_347_n N_VGND_c_396_n 0.0235688f $X=0.49 $Y=0.34 $X2=0 $Y2=0
cc_210 N_A_36_74#_c_351_n N_VGND_c_397_n 0.0115122f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0
cc_211 N_A_36_74#_c_346_n N_VGND_c_399_n 0.028285f $X=1.1 $Y=0.34 $X2=0 $Y2=0
cc_212 N_A_36_74#_c_347_n N_VGND_c_399_n 0.0127152f $X=0.49 $Y=0.34 $X2=0 $Y2=0
cc_213 N_A_36_74#_c_351_n N_VGND_c_399_n 0.0095288f $X=2.045 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__nand2b_1.spice
* Created: Fri Aug 28 17:42:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand2b_1.pex.spice"
.subckt sky130_fd_sc_ms__nand2b_1  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_N_M1003_g N_A_27_112#_M1003_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.191114 AS=0.15675 PD=1.16395 PS=1.67 NRD=1.08 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1001 A_269_74# N_B_M1001_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.257136 PD=0.98 PS=1.56605 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_112#_M1000_g A_269_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.3182 AS=0.0888 PD=2.34 PS=0.98 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75001.2 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A_N_M1002_g N_A_27_112#_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2262 AS=0.2352 PD=1.38 PS=2.24 NRD=19.9167 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12 AD=0.1792
+ AS=0.3016 PD=1.44 PS=1.84 NRD=0 NRS=21.9852 M=1 R=6.22222 SA=90000.7
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_27_112#_M1005_g N_Y_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3192 AS=0.1792 PD=2.81 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
c_25 VNB 0 1.74227e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__nand2b_1.pxi.spice"
*
.ends
*
*

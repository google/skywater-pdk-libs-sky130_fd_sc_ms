* File: sky130_fd_sc_ms__sdfrtn_1.pxi.spice
* Created: Wed Sep  2 12:30:26 2020
* 
x_PM_SKY130_FD_SC_MS__SDFRTN_1%SCE N_SCE_M1011_g N_SCE_M1037_g N_SCE_c_269_n
+ N_SCE_M1012_g N_SCE_M1006_g N_SCE_c_271_n N_SCE_c_272_n N_SCE_c_273_n
+ N_SCE_c_274_n SCE N_SCE_c_275_n N_SCE_c_276_n PM_SKY130_FD_SC_MS__SDFRTN_1%SCE
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_27_88# N_A_27_88#_M1037_s N_A_27_88#_M1011_s
+ N_A_27_88#_M1018_g N_A_27_88#_M1015_g N_A_27_88#_c_338_n N_A_27_88#_c_339_n
+ N_A_27_88#_c_348_n N_A_27_88#_c_349_n N_A_27_88#_c_350_n N_A_27_88#_c_340_n
+ N_A_27_88#_c_341_n N_A_27_88#_c_352_n N_A_27_88#_c_342_n N_A_27_88#_c_343_n
+ N_A_27_88#_c_344_n N_A_27_88#_c_345_n PM_SKY130_FD_SC_MS__SDFRTN_1%A_27_88#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%D N_D_M1034_g N_D_c_428_n N_D_c_429_n N_D_M1020_g
+ D D N_D_c_431_n N_D_c_432_n PM_SKY130_FD_SC_MS__SDFRTN_1%D
x_PM_SKY130_FD_SC_MS__SDFRTN_1%SCD N_SCD_c_468_n N_SCD_M1036_g N_SCD_c_469_n
+ N_SCD_M1032_g N_SCD_c_470_n SCD SCD N_SCD_c_467_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%SCD
x_PM_SKY130_FD_SC_MS__SDFRTN_1%CLK_N N_CLK_N_c_516_n N_CLK_N_M1000_g
+ N_CLK_N_c_513_n N_CLK_N_M1007_g N_CLK_N_c_514_n N_CLK_N_c_515_n CLK_N
+ PM_SKY130_FD_SC_MS__SDFRTN_1%CLK_N
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_1069_74# N_A_1069_74#_M1008_d
+ N_A_1069_74#_M1029_d N_A_1069_74#_M1021_g N_A_1069_74#_c_575_n
+ N_A_1069_74#_M1024_g N_A_1069_74#_M1031_g N_A_1069_74#_c_560_n
+ N_A_1069_74#_M1026_g N_A_1069_74#_c_562_n N_A_1069_74#_c_638_p
+ N_A_1069_74#_c_563_n N_A_1069_74#_c_564_n N_A_1069_74#_c_565_n
+ N_A_1069_74#_c_566_n N_A_1069_74#_c_567_n N_A_1069_74#_c_568_n
+ N_A_1069_74#_c_581_p N_A_1069_74#_c_598_p N_A_1069_74#_c_569_n
+ N_A_1069_74#_c_570_n N_A_1069_74#_c_571_n N_A_1069_74#_c_594_p
+ N_A_1069_74#_c_595_p N_A_1069_74#_c_572_n N_A_1069_74#_c_579_n
+ N_A_1069_74#_c_573_n N_A_1069_74#_c_614_p N_A_1069_74#_c_649_p
+ N_A_1069_74#_c_574_n PM_SKY130_FD_SC_MS__SDFRTN_1%A_1069_74#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_1417_294# N_A_1417_294#_M1035_d
+ N_A_1417_294#_M1038_d N_A_1417_294#_M1033_g N_A_1417_294#_M1016_g
+ N_A_1417_294#_c_743_n N_A_1417_294#_c_744_n N_A_1417_294#_c_745_n
+ N_A_1417_294#_c_751_n N_A_1417_294#_c_746_n N_A_1417_294#_c_747_n
+ N_A_1417_294#_c_748_n N_A_1417_294#_c_776_n N_A_1417_294#_c_787_p
+ N_A_1417_294#_c_749_n PM_SKY130_FD_SC_MS__SDFRTN_1%A_1417_294#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%RESET_B N_RESET_B_M1002_g N_RESET_B_M1023_g
+ N_RESET_B_c_840_n N_RESET_B_c_857_n N_RESET_B_c_858_n N_RESET_B_M1003_g
+ N_RESET_B_M1030_g N_RESET_B_M1009_g N_RESET_B_M1019_g N_RESET_B_c_843_n
+ N_RESET_B_c_861_n N_RESET_B_c_844_n N_RESET_B_c_845_n N_RESET_B_c_846_n
+ N_RESET_B_c_847_n N_RESET_B_c_848_n RESET_B N_RESET_B_c_849_n
+ N_RESET_B_c_850_n N_RESET_B_c_851_n N_RESET_B_c_852_n N_RESET_B_c_853_n
+ N_RESET_B_c_854_n PM_SKY130_FD_SC_MS__SDFRTN_1%RESET_B
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_1273_131# N_A_1273_131#_M1021_d
+ N_A_1273_131#_M1001_d N_A_1273_131#_M1030_d N_A_1273_131#_c_1060_n
+ N_A_1273_131#_M1035_g N_A_1273_131#_M1038_g N_A_1273_131#_c_1061_n
+ N_A_1273_131#_c_1062_n N_A_1273_131#_c_1067_n N_A_1273_131#_c_1068_n
+ N_A_1273_131#_c_1069_n N_A_1273_131#_c_1070_n N_A_1273_131#_c_1063_n
+ N_A_1273_131#_c_1110_n N_A_1273_131#_c_1064_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%A_1273_131#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_859_347# N_A_859_347#_M1007_s
+ N_A_859_347#_M1000_s N_A_859_347#_c_1165_n N_A_859_347#_M1008_g
+ N_A_859_347#_c_1183_n N_A_859_347#_M1029_g N_A_859_347#_c_1166_n
+ N_A_859_347#_c_1167_n N_A_859_347#_c_1168_n N_A_859_347#_c_1169_n
+ N_A_859_347#_c_1185_n N_A_859_347#_c_1186_n N_A_859_347#_c_1187_n
+ N_A_859_347#_M1001_g N_A_859_347#_M1028_g N_A_859_347#_c_1171_n
+ N_A_859_347#_M1039_g N_A_859_347#_M1005_g N_A_859_347#_c_1174_n
+ N_A_859_347#_c_1196_n N_A_859_347#_c_1199_n N_A_859_347#_c_1200_n
+ N_A_859_347#_c_1202_n N_A_859_347#_c_1189_n N_A_859_347#_c_1175_n
+ N_A_859_347#_c_1176_n N_A_859_347#_c_1177_n N_A_859_347#_c_1178_n
+ N_A_859_347#_c_1179_n N_A_859_347#_c_1180_n N_A_859_347#_c_1181_n
+ N_A_859_347#_c_1182_n PM_SKY130_FD_SC_MS__SDFRTN_1%A_859_347#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_2087_410# N_A_2087_410#_M1010_d
+ N_A_2087_410#_M1019_d N_A_2087_410#_M1013_g N_A_2087_410#_M1004_g
+ N_A_2087_410#_c_1372_n N_A_2087_410#_c_1373_n N_A_2087_410#_c_1368_n
+ N_A_2087_410#_c_1374_n N_A_2087_410#_c_1369_n N_A_2087_410#_c_1376_n
+ N_A_2087_410#_c_1377_n N_A_2087_410#_c_1378_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%A_2087_410#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_1827_144# N_A_1827_144#_M1039_d
+ N_A_1827_144#_M1031_d N_A_1827_144#_c_1458_n N_A_1827_144#_M1010_g
+ N_A_1827_144#_c_1459_n N_A_1827_144#_c_1460_n N_A_1827_144#_M1022_g
+ N_A_1827_144#_c_1470_n N_A_1827_144#_c_1461_n N_A_1827_144#_c_1471_n
+ N_A_1827_144#_M1025_g N_A_1827_144#_c_1462_n N_A_1827_144#_M1027_g
+ N_A_1827_144#_c_1463_n N_A_1827_144#_c_1472_n N_A_1827_144#_c_1464_n
+ N_A_1827_144#_c_1473_n N_A_1827_144#_c_1474_n N_A_1827_144#_c_1475_n
+ N_A_1827_144#_c_1465_n N_A_1827_144#_c_1476_n N_A_1827_144#_c_1466_n
+ N_A_1827_144#_c_1467_n N_A_1827_144#_c_1478_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%A_1827_144#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_2492_424# N_A_2492_424#_M1027_s
+ N_A_2492_424#_M1025_s N_A_2492_424#_M1014_g N_A_2492_424#_M1017_g
+ N_A_2492_424#_c_1604_n N_A_2492_424#_c_1605_n N_A_2492_424#_c_1606_n
+ N_A_2492_424#_c_1611_n N_A_2492_424#_c_1607_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%A_2492_424#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%VPWR N_VPWR_M1011_d N_VPWR_M1036_d N_VPWR_M1000_d
+ N_VPWR_M1033_d N_VPWR_M1038_s N_VPWR_M1013_d N_VPWR_M1022_d N_VPWR_M1025_d
+ N_VPWR_c_1648_n N_VPWR_c_1649_n N_VPWR_c_1650_n N_VPWR_c_1651_n
+ N_VPWR_c_1652_n N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n VPWR
+ N_VPWR_c_1656_n N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n
+ N_VPWR_c_1660_n N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n
+ N_VPWR_c_1647_n N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1667_n
+ N_VPWR_c_1668_n N_VPWR_c_1669_n N_VPWR_c_1670_n N_VPWR_c_1671_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%VPWR
x_PM_SKY130_FD_SC_MS__SDFRTN_1%A_287_464# N_A_287_464#_M1020_d
+ N_A_287_464#_M1021_s N_A_287_464#_M1034_d N_A_287_464#_M1002_d
+ N_A_287_464#_M1001_s N_A_287_464#_c_1801_n N_A_287_464#_c_1792_n
+ N_A_287_464#_c_1787_n N_A_287_464#_c_1788_n N_A_287_464#_c_1789_n
+ N_A_287_464#_c_1790_n N_A_287_464#_c_1794_n N_A_287_464#_c_1795_n
+ N_A_287_464#_c_1791_n N_A_287_464#_c_1797_n N_A_287_464#_c_1798_n
+ N_A_287_464#_c_1799_n N_A_287_464#_c_1807_n N_A_287_464#_c_1812_n
+ N_A_287_464#_c_1835_n N_A_287_464#_c_1800_n
+ PM_SKY130_FD_SC_MS__SDFRTN_1%A_287_464#
x_PM_SKY130_FD_SC_MS__SDFRTN_1%Q N_Q_M1017_d N_Q_M1014_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__SDFRTN_1%Q
x_PM_SKY130_FD_SC_MS__SDFRTN_1%VGND N_VGND_M1037_d N_VGND_M1023_d N_VGND_M1007_d
+ N_VGND_M1003_d N_VGND_M1004_d N_VGND_M1027_d N_VGND_c_1933_n N_VGND_c_1934_n
+ N_VGND_c_1935_n N_VGND_c_1936_n N_VGND_c_1937_n N_VGND_c_1938_n
+ N_VGND_c_1939_n N_VGND_c_1940_n VGND N_VGND_c_1941_n N_VGND_c_1942_n
+ N_VGND_c_1943_n N_VGND_c_1944_n N_VGND_c_1945_n N_VGND_c_1946_n
+ N_VGND_c_1947_n N_VGND_c_1948_n N_VGND_c_1949_n N_VGND_c_1950_n
+ N_VGND_c_1951_n N_VGND_c_1952_n PM_SKY130_FD_SC_MS__SDFRTN_1%VGND
x_PM_SKY130_FD_SC_MS__SDFRTN_1%noxref_24 N_noxref_24_M1018_s N_noxref_24_M1032_d
+ N_noxref_24_c_2058_n N_noxref_24_c_2059_n N_noxref_24_c_2060_n
+ N_noxref_24_c_2063_n PM_SKY130_FD_SC_MS__SDFRTN_1%noxref_24
cc_1 VNB N_SCE_M1037_g 0.05663f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_2 VNB N_SCE_c_269_n 0.00333779f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.93
cc_3 VNB N_SCE_M1006_g 0.0185275f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.615
cc_4 VNB N_SCE_c_271_n 0.00276011f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_5 VNB N_SCE_c_272_n 0.0317749f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_6 VNB N_SCE_c_273_n 0.0256442f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.267
cc_7 VNB N_SCE_c_274_n 0.00942789f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.267
cc_8 VNB N_SCE_c_275_n 0.0114065f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_9 VNB N_SCE_c_276_n 0.046047f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.12
cc_10 VNB N_A_27_88#_c_338_n 0.0276281f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.615
cc_11 VNB N_A_27_88#_c_339_n 0.0210999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_88#_c_340_n 0.0146482f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.575
cc_13 VNB N_A_27_88#_c_341_n 0.0108567f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_14 VNB N_A_27_88#_c_342_n 0.00647888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_88#_c_343_n 0.03765f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.12
cc_16 VNB N_A_27_88#_c_344_n 0.0215459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_88#_c_345_n 0.0189579f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_18 VNB N_D_M1020_g 0.0631098f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.632
cc_19 VNB N_SCD_M1032_g 0.0483128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB SCD 0.00419665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_SCD_c_467_n 0.0148775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_CLK_N_c_513_n 0.0209351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_CLK_N_c_514_n 0.04335f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_24 VNB N_CLK_N_c_515_n 0.0137811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_1069_74#_M1021_g 0.0246055f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.632
cc_26 VNB N_A_1069_74#_M1031_g 0.0262807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_1069_74#_c_560_n 0.0294946f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.495
cc_28 VNB N_A_1069_74#_M1026_g 0.0246368f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_29 VNB N_A_1069_74#_c_562_n 0.0104354f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.267
cc_30 VNB N_A_1069_74#_c_563_n 0.00979101f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_31 VNB N_A_1069_74#_c_564_n 0.00332707f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_32 VNB N_A_1069_74#_c_565_n 0.00553606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1069_74#_c_566_n 0.06504f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.182
cc_34 VNB N_A_1069_74#_c_567_n 0.0170828f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_35 VNB N_A_1069_74#_c_568_n 0.00338164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1069_74#_c_569_n 0.0021081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1069_74#_c_570_n 0.0117821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1069_74#_c_571_n 0.0027073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1069_74#_c_572_n 0.00739436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1069_74#_c_573_n 6.24913e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1069_74#_c_574_n 0.0381518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1417_294#_M1016_g 0.0313938f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_43 VNB N_A_1417_294#_c_743_n 0.00868114f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_44 VNB N_A_1417_294#_c_744_n 0.00206132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1417_294#_c_745_n 0.00140633f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.495
cc_46 VNB N_A_1417_294#_c_746_n 0.00443149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1417_294#_c_747_n 0.0234461f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.575
cc_48 VNB N_A_1417_294#_c_748_n 0.00166205f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.41
cc_49 VNB N_A_1417_294#_c_749_n 0.00331528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_M1023_g 0.0457804f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_51 VNB N_RESET_B_c_840_n 0.00905985f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.93
cc_52 VNB N_RESET_B_M1003_g 0.0341098f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.955
cc_53 VNB N_RESET_B_M1009_g 0.0335346f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.495
cc_54 VNB N_RESET_B_c_843_n 0.0059249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_RESET_B_c_844_n 0.020734f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.41
cc_56 VNB N_RESET_B_c_845_n 4.19263e-19 $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_57 VNB N_RESET_B_c_846_n 0.01806f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_58 VNB N_RESET_B_c_847_n 8.92608e-19 $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_59 VNB N_RESET_B_c_848_n 0.00211188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_RESET_B_c_849_n 0.0194896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_c_850_n 0.0016999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_RESET_B_c_851_n 0.0261837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_RESET_B_c_852_n 0.00155453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_c_853_n 0.0293012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_RESET_B_c_854_n 0.00982208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1273_131#_c_1060_n 0.0189491f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.93
cc_67 VNB N_A_1273_131#_c_1061_n 0.00174337f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_68 VNB N_A_1273_131#_c_1062_n 0.00674844f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.495
cc_69 VNB N_A_1273_131#_c_1063_n 0.00106086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1273_131#_c_1064_n 0.0361833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_859_347#_c_1165_n 0.0181083f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_72 VNB N_A_859_347#_c_1166_n 0.0502825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_859_347#_c_1167_n 0.0040226f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_74 VNB N_A_859_347#_c_1168_n 0.0684595f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_75 VNB N_A_859_347#_c_1169_n 0.0123819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_859_347#_M1028_g 0.0400594f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.182
cc_77 VNB N_A_859_347#_c_1171_n 0.149807f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.267
cc_78 VNB N_A_859_347#_M1039_g 0.0440711f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_79 VNB N_A_859_347#_M1005_g 0.00205879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_859_347#_c_1174_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_859_347#_c_1175_n 0.00234601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_859_347#_c_1176_n 0.00108736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_859_347#_c_1177_n 0.00490328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_859_347#_c_1178_n 0.0237915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_859_347#_c_1179_n 0.00247817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_859_347#_c_1180_n 0.0340098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_859_347#_c_1181_n 0.00888046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_859_347#_c_1182_n 0.0552357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2087_410#_M1004_g 0.0626814f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_90 VNB N_A_2087_410#_c_1368_n 0.00234211f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.495
cc_91 VNB N_A_2087_410#_c_1369_n 0.0133151f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.267
cc_92 VNB N_A_1827_144#_c_1458_n 0.0218114f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.65
cc_93 VNB N_A_1827_144#_c_1459_n 0.0200739f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.08
cc_94 VNB N_A_1827_144#_c_1460_n 0.00490842f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_95 VNB N_A_1827_144#_c_1461_n 0.0770594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1827_144#_c_1462_n 0.0208776f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_97 VNB N_A_1827_144#_c_1463_n 0.0175897f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.267
cc_98 VNB N_A_1827_144#_c_1464_n 0.00837077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1827_144#_c_1465_n 0.0322706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1827_144#_c_1466_n 0.00113131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1827_144#_c_1467_n 0.0199884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2492_424#_M1017_g 0.0336704f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_103 VNB N_A_2492_424#_c_1604_n 0.0509652f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.955
cc_104 VNB N_A_2492_424#_c_1605_n 0.016189f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=0.615
cc_105 VNB N_A_2492_424#_c_1606_n 0.0173592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2492_424#_c_1607_n 0.00257436f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.182
cc_107 VNB N_VPWR_c_1647_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_287_464#_c_1787_n 0.00241686f $X=-0.19 $Y=-0.245 $X2=0.7
+ $Y2=1.575
cc_109 VNB N_A_287_464#_c_1788_n 0.0317474f $X=-0.19 $Y=-0.245 $X2=2.045
+ $Y2=1.182
cc_110 VNB N_A_287_464#_c_1789_n 0.00549408f $X=-0.19 $Y=-0.245 $X2=1.875
+ $Y2=1.267
cc_111 VNB N_A_287_464#_c_1790_n 0.00997902f $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=1.21
cc_112 VNB N_A_287_464#_c_1791_n 0.0193201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB Q 0.0545639f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_114 VNB N_VGND_c_1933_n 0.0212574f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=1.495
cc_115 VNB N_VGND_c_1934_n 0.011956f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.575
cc_116 VNB N_VGND_c_1935_n 0.00961271f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_117 VNB N_VGND_c_1936_n 0.0122202f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.12
cc_118 VNB N_VGND_c_1937_n 0.00450109f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.12
cc_119 VNB N_VGND_c_1938_n 0.015381f $X=-0.19 $Y=-0.245 $X2=2.385 $Y2=1.182
cc_120 VNB N_VGND_c_1939_n 0.0652707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1940_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1941_n 0.0194805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1942_n 0.0246035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1943_n 0.0681991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1944_n 0.0662658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1945_n 0.0500113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1946_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1947_n 0.749405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1948_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1949_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1950_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1951_n 0.00865198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1952_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_noxref_24_c_2058_n 0.00347762f $X=-0.19 $Y=-0.245 $X2=0.642
+ $Y2=1.632
cc_135 VNB N_noxref_24_c_2059_n 0.0148302f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.08
cc_136 VNB N_noxref_24_c_2060_n 0.00461646f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_137 VPB N_SCE_M1011_g 0.0243208f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_138 VPB N_SCE_c_269_n 0.059182f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.93
cc_139 VPB N_SCE_M1012_g 0.0243754f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_140 VPB N_SCE_c_271_n 9.10905e-19 $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_141 VPB N_A_27_88#_M1015_g 0.0441455f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_142 VPB N_A_27_88#_c_339_n 0.0318758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_27_88#_c_348_n 0.0214727f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.495
cc_144 VPB N_A_27_88#_c_349_n 0.0182131f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_145 VPB N_A_27_88#_c_350_n 0.00325153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_27_88#_c_340_n 0.021371f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.575
cc_147 VPB N_A_27_88#_c_352_n 0.00716038f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_148 VPB N_D_M1034_g 0.0332759f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_149 VPB N_D_c_428_n 0.0146877f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.41
cc_150 VPB N_D_c_429_n 0.00881863f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_151 VPB N_D_M1020_g 0.00943149f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.632
cc_152 VPB N_D_c_431_n 0.0336862f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.615
cc_153 VPB N_D_c_432_n 0.0162449f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.615
cc_154 VPB N_SCD_c_468_n 0.0182698f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.17
cc_155 VPB N_SCD_c_469_n 0.0136324f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.41
cc_156 VPB N_SCD_c_470_n 0.0282331f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_157 VPB SCD 0.00642005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_SCD_c_467_n 0.0178291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_CLK_N_c_516_n 0.0200428f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.17
cc_160 VPB N_CLK_N_c_514_n 0.0235312f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_161 VPB N_CLK_N_c_515_n 0.00356384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_1069_74#_c_575_n 0.00641676f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_163 VPB N_A_1069_74#_M1024_g 0.021145f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.955
cc_164 VPB N_A_1069_74#_M1031_g 0.0295007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_1069_74#_c_562_n 0.0116039f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.267
cc_166 VPB N_A_1069_74#_c_579_n 7.04287e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_1069_74#_c_573_n 3.9332e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1417_294#_M1033_g 0.0346898f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.632
cc_169 VPB N_A_1417_294#_c_751_n 0.006734f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.267
cc_170 VPB N_A_1417_294#_c_746_n 0.00161036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_1417_294#_c_747_n 0.00547497f $X=-0.19 $Y=1.66 $X2=0.642
+ $Y2=1.575
cc_172 VPB N_A_1417_294#_c_749_n 0.00241226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_RESET_B_M1002_g 0.0151206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_RESET_B_c_840_n 0.0665332f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.93
cc_175 VPB N_RESET_B_c_857_n 0.331367f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.08
cc_176 VPB N_RESET_B_c_858_n 0.0139277f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_177 VPB N_RESET_B_M1030_g 0.0565314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_c_843_n 0.0349147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_RESET_B_c_861_n 0.0330294f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.575
cc_180 VPB N_RESET_B_c_844_n 0.00651387f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.41
cc_181 VPB N_RESET_B_c_845_n 4.37909e-19 $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_182 VPB N_RESET_B_c_846_n 0.00114121f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_183 VPB N_RESET_B_c_847_n 2.20425e-19 $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_184 VPB N_RESET_B_c_848_n 0.00221319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_RESET_B_c_850_n 0.00266259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_RESET_B_c_851_n 0.00642675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_RESET_B_c_852_n 3.06104e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_RESET_B_c_854_n 6.46864e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1273_131#_M1038_g 0.028796f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.955
cc_190 VPB N_A_1273_131#_c_1062_n 0.00262806f $X=-0.19 $Y=1.66 $X2=1.875
+ $Y2=1.495
cc_191 VPB N_A_1273_131#_c_1067_n 0.0189858f $X=-0.19 $Y=1.66 $X2=0.865
+ $Y2=1.495
cc_192 VPB N_A_1273_131#_c_1068_n 0.0065836f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.495
cc_193 VPB N_A_1273_131#_c_1069_n 0.0132333f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_194 VPB N_A_1273_131#_c_1070_n 0.00908245f $X=-0.19 $Y=1.66 $X2=2.045
+ $Y2=1.182
cc_195 VPB N_A_1273_131#_c_1063_n 0.00318229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1273_131#_c_1064_n 0.0124662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_859_347#_c_1183_n 0.0187075f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.93
cc_198 VPB N_A_859_347#_c_1167_n 0.0162001f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.615
cc_199 VPB N_A_859_347#_c_1185_n 0.0393737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_859_347#_c_1186_n 0.00952378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_859_347#_c_1187_n 0.0188508f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.495
cc_202 VPB N_A_859_347#_M1005_g 0.0597226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_859_347#_c_1189_n 0.00237373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_859_347#_c_1175_n 2.06527e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_859_347#_c_1177_n 0.00274696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_859_347#_c_1178_n 0.0106103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_859_347#_c_1182_n 0.0190283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_2087_410#_M1013_g 0.02279f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.632
cc_209 VPB N_A_2087_410#_M1004_g 0.0217533f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_210 VPB N_A_2087_410#_c_1372_n 0.010007f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.955
cc_211 VPB N_A_2087_410#_c_1373_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_2087_410#_c_1374_n 0.0106612f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.575
cc_213 VPB N_A_2087_410#_c_1369_n 0.00834784f $X=-0.19 $Y=1.66 $X2=2.045
+ $Y2=1.267
cc_214 VPB N_A_2087_410#_c_1376_n 0.00347726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_2087_410#_c_1377_n 0.0337684f $X=-0.19 $Y=1.66 $X2=0.642
+ $Y2=1.575
cc_216 VPB N_A_2087_410#_c_1378_n 0.00251499f $X=-0.19 $Y=1.66 $X2=2.385
+ $Y2=1.12
cc_217 VPB N_A_1827_144#_c_1460_n 0.0140687f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_218 VPB N_A_1827_144#_M1022_g 0.0446384f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=0.615
cc_219 VPB N_A_1827_144#_c_1470_n 0.0736424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1827_144#_c_1471_n 0.0205307f $X=-0.19 $Y=1.66 $X2=0.865
+ $Y2=1.495
cc_221 VPB N_A_1827_144#_c_1472_n 0.00569915f $X=-0.19 $Y=1.66 $X2=2.075
+ $Y2=1.21
cc_222 VPB N_A_1827_144#_c_1473_n 0.00400866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1827_144#_c_1474_n 0.0134162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1827_144#_c_1475_n 0.00336725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1827_144#_c_1476_n 0.01246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1827_144#_c_1466_n 0.0041497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1827_144#_c_1478_n 0.0081065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_2492_424#_M1014_g 0.0289694f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.632
cc_229 VPB N_A_2492_424#_c_1604_n 0.0194078f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.955
cc_230 VPB N_A_2492_424#_c_1605_n 0.00119105f $X=-0.19 $Y=1.66 $X2=2.615
+ $Y2=0.615
cc_231 VPB N_A_2492_424#_c_1611_n 0.0161255f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.495
cc_232 VPB N_A_2492_424#_c_1607_n 3.52822e-19 $X=-0.19 $Y=1.66 $X2=2.045
+ $Y2=1.182
cc_233 VPB N_VPWR_c_1648_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.875 $Y2=1.267
cc_234 VPB N_VPWR_c_1649_n 0.020001f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.575
cc_235 VPB N_VPWR_c_1650_n 0.012958f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=1.12
cc_236 VPB N_VPWR_c_1651_n 0.0145779f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.182
cc_237 VPB N_VPWR_c_1652_n 0.0126407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1653_n 0.0159801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1654_n 0.0187266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1655_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1656_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1657_n 0.0518169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1658_n 0.0465394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1659_n 0.0622721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1660_n 0.0212211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1661_n 0.0546438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1662_n 0.0215226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1663_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1647_n 0.120235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1665_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1666_n 0.013941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1667_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1668_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1669_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1670_n 0.0200143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1671_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_287_464#_c_1792_n 0.033187f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.495
cc_258 VPB N_A_287_464#_c_1790_n 0.0126396f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.21
cc_259 VPB N_A_287_464#_c_1794_n 0.00785257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_287_464#_c_1795_n 0.00462229f $X=-0.19 $Y=1.66 $X2=0.642 $Y2=1.41
cc_261 VPB N_A_287_464#_c_1791_n 0.00154534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_287_464#_c_1797_n 0.00387559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_287_464#_c_1798_n 0.00134275f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.182
cc_264 VPB N_A_287_464#_c_1799_n 0.00709212f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_287_464#_c_1800_n 0.00155579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB Q 0.0535067f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_267 N_SCE_M1037_g N_A_27_88#_c_338_n 0.0173492f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_268 N_SCE_M1037_g N_A_27_88#_c_339_n 0.0255944f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_269 N_SCE_c_269_n N_A_27_88#_c_339_n 0.00871119f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_270 N_SCE_c_271_n N_A_27_88#_c_339_n 0.0525665f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_271 N_SCE_M1011_g N_A_27_88#_c_348_n 4.69176e-19 $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_272 N_SCE_M1011_g N_A_27_88#_c_349_n 0.0183618f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_273 N_SCE_c_269_n N_A_27_88#_c_349_n 5.99745e-19 $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_274 N_SCE_M1012_g N_A_27_88#_c_349_n 0.0204478f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_275 N_SCE_c_271_n N_A_27_88#_c_349_n 0.0220875f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_276 N_SCE_c_275_n N_A_27_88#_c_350_n 0.0282051f $X=2.385 $Y=1.12 $X2=0 $Y2=0
cc_277 N_SCE_c_276_n N_A_27_88#_c_350_n 3.15902e-19 $X=2.615 $Y=1.12 $X2=0 $Y2=0
cc_278 N_SCE_c_274_n N_A_27_88#_c_340_n 6.75701e-19 $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_279 N_SCE_c_275_n N_A_27_88#_c_340_n 0.00373152f $X=2.385 $Y=1.12 $X2=0 $Y2=0
cc_280 N_SCE_c_276_n N_A_27_88#_c_340_n 0.0150192f $X=2.615 $Y=1.12 $X2=0 $Y2=0
cc_281 N_SCE_M1037_g N_A_27_88#_c_341_n 0.00558381f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_282 N_SCE_c_274_n N_A_27_88#_c_342_n 0.016963f $X=2.045 $Y=1.267 $X2=0 $Y2=0
cc_283 N_SCE_M1037_g N_A_27_88#_c_343_n 0.00404033f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_284 N_SCE_c_273_n N_A_27_88#_c_343_n 0.00396344f $X=1.875 $Y=1.267 $X2=0
+ $Y2=0
cc_285 N_SCE_c_274_n N_A_27_88#_c_343_n 4.95772e-19 $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_286 N_SCE_M1037_g N_A_27_88#_c_344_n 0.0161451f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_287 N_SCE_c_271_n N_A_27_88#_c_344_n 0.0264209f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_288 N_SCE_c_272_n N_A_27_88#_c_344_n 0.00206933f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_289 N_SCE_c_273_n N_A_27_88#_c_344_n 0.0568522f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_290 N_SCE_M1012_g N_D_M1034_g 0.0358851f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_291 N_SCE_c_269_n N_D_c_429_n 0.0358851f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_292 N_SCE_c_273_n N_D_c_429_n 0.00120253f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_293 N_SCE_M1006_g N_D_M1020_g 0.0146952f $X=2.615 $Y=0.615 $X2=0 $Y2=0
cc_294 N_SCE_c_273_n N_D_M1020_g 0.00734487f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_295 N_SCE_c_274_n N_D_M1020_g 0.027662f $X=2.045 $Y=1.267 $X2=0 $Y2=0
cc_296 N_SCE_c_276_n N_D_M1020_g 0.0181201f $X=2.615 $Y=1.12 $X2=0 $Y2=0
cc_297 N_SCE_c_269_n N_D_c_431_n 3.94848e-19 $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_298 N_SCE_c_273_n N_D_c_431_n 0.00395715f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_299 N_SCE_c_269_n N_D_c_432_n 0.00643854f $X=0.642 $Y=1.93 $X2=0 $Y2=0
cc_300 N_SCE_c_271_n N_D_c_432_n 0.0207563f $X=0.7 $Y=1.575 $X2=0 $Y2=0
cc_301 N_SCE_c_273_n N_D_c_432_n 0.0621482f $X=1.875 $Y=1.267 $X2=0 $Y2=0
cc_302 N_SCE_M1006_g N_SCD_M1032_g 0.0518638f $X=2.615 $Y=0.615 $X2=0 $Y2=0
cc_303 N_SCE_c_275_n N_SCD_M1032_g 0.0046975f $X=2.385 $Y=1.12 $X2=0 $Y2=0
cc_304 N_SCE_M1011_g N_VPWR_c_1648_n 0.0116339f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_305 N_SCE_M1012_g N_VPWR_c_1648_n 0.0107737f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_306 N_SCE_M1011_g N_VPWR_c_1656_n 0.00460063f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_307 N_SCE_M1012_g N_VPWR_c_1657_n 0.00460063f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_308 N_SCE_M1011_g N_VPWR_c_1647_n 0.00912296f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_309 N_SCE_M1012_g N_VPWR_c_1647_n 0.00908061f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_310 N_SCE_M1006_g N_A_287_464#_c_1801_n 0.0148189f $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_311 N_SCE_c_274_n N_A_287_464#_c_1801_n 0.0386304f $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_312 N_SCE_c_276_n N_A_287_464#_c_1801_n 0.00694878f $X=2.615 $Y=1.12 $X2=0
+ $Y2=0
cc_313 N_SCE_M1006_g N_A_287_464#_c_1787_n 0.00344346f $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_314 N_SCE_c_275_n N_A_287_464#_c_1789_n 0.020046f $X=2.385 $Y=1.12 $X2=0
+ $Y2=0
cc_315 N_SCE_c_276_n N_A_287_464#_c_1789_n 0.00204275f $X=2.615 $Y=1.12 $X2=0
+ $Y2=0
cc_316 N_SCE_M1012_g N_A_287_464#_c_1807_n 8.90742e-19 $X=0.955 $Y=2.64 $X2=0
+ $Y2=0
cc_317 N_SCE_M1037_g N_VGND_c_1933_n 0.0137116f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_318 N_SCE_M1006_g N_VGND_c_1939_n 9.15902e-19 $X=2.615 $Y=0.615 $X2=0 $Y2=0
cc_319 N_SCE_M1037_g N_VGND_c_1941_n 0.00504315f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_320 N_SCE_M1037_g N_VGND_c_1947_n 0.00523671f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_321 N_SCE_M1006_g N_noxref_24_c_2059_n 0.0105907f $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_322 N_SCE_c_274_n N_noxref_24_c_2059_n 0.00237332f $X=2.045 $Y=1.267 $X2=0
+ $Y2=0
cc_323 N_SCE_M1006_g N_noxref_24_c_2063_n 9.6581e-19 $X=2.615 $Y=0.615 $X2=0
+ $Y2=0
cc_324 N_A_27_88#_c_349_n N_D_M1034_g 0.0176962f $X=2.215 $Y=2.375 $X2=0 $Y2=0
cc_325 N_A_27_88#_c_349_n N_D_c_428_n 0.00373424f $X=2.215 $Y=2.375 $X2=0 $Y2=0
cc_326 N_A_27_88#_c_343_n N_D_c_429_n 0.00329011f $X=1.455 $Y=1.1 $X2=0 $Y2=0
cc_327 N_A_27_88#_c_350_n N_D_M1020_g 0.00125677f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_328 N_A_27_88#_c_340_n N_D_M1020_g 0.0173599f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_329 N_A_27_88#_c_342_n N_D_M1020_g 0.00101912f $X=1.455 $Y=1.1 $X2=0 $Y2=0
cc_330 N_A_27_88#_c_345_n N_D_M1020_g 0.0606403f $X=1.455 $Y=0.935 $X2=0 $Y2=0
cc_331 N_A_27_88#_M1015_g N_D_c_431_n 0.0173599f $X=2.28 $Y=2.64 $X2=0 $Y2=0
cc_332 N_A_27_88#_c_350_n N_D_c_431_n 3.97221e-19 $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_333 N_A_27_88#_c_349_n N_D_c_432_n 0.0697007f $X=2.215 $Y=2.375 $X2=0 $Y2=0
cc_334 N_A_27_88#_c_350_n N_D_c_432_n 0.0208146f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_335 N_A_27_88#_c_340_n N_D_c_432_n 0.00108531f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_336 N_A_27_88#_c_349_n N_SCD_c_468_n 0.00141562f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_337 N_A_27_88#_M1015_g N_SCD_c_469_n 0.00468854f $X=2.28 $Y=2.64 $X2=0 $Y2=0
cc_338 N_A_27_88#_c_350_n N_SCD_c_469_n 0.0015238f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_339 N_A_27_88#_M1015_g N_SCD_c_470_n 0.0629564f $X=2.28 $Y=2.64 $X2=0 $Y2=0
cc_340 N_A_27_88#_c_350_n N_SCD_c_470_n 0.00430208f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_341 N_A_27_88#_M1015_g SCD 2.48643e-19 $X=2.28 $Y=2.64 $X2=0 $Y2=0
cc_342 N_A_27_88#_c_350_n SCD 0.0326702f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_343 N_A_27_88#_c_340_n SCD 0.00133605f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_344 N_A_27_88#_c_350_n N_SCD_c_467_n 0.00113065f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_345 N_A_27_88#_c_340_n N_SCD_c_467_n 0.0160213f $X=2.38 $Y=1.72 $X2=0 $Y2=0
cc_346 N_A_27_88#_c_349_n N_VPWR_M1011_d 0.00165831f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_347 N_A_27_88#_c_348_n N_VPWR_c_1648_n 0.0122069f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_348 N_A_27_88#_c_349_n N_VPWR_c_1648_n 0.0170259f $X=2.215 $Y=2.375 $X2=0
+ $Y2=0
cc_349 N_A_27_88#_c_348_n N_VPWR_c_1656_n 0.011066f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_350 N_A_27_88#_M1015_g N_VPWR_c_1657_n 0.00422272f $X=2.28 $Y=2.64 $X2=0
+ $Y2=0
cc_351 N_A_27_88#_M1015_g N_VPWR_c_1647_n 0.00638283f $X=2.28 $Y=2.64 $X2=0
+ $Y2=0
cc_352 N_A_27_88#_c_348_n N_VPWR_c_1647_n 0.00915947f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_353 N_A_27_88#_c_349_n A_209_464# 0.00366293f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_354 N_A_27_88#_c_349_n N_A_287_464#_M1034_d 0.00986957f $X=2.215 $Y=2.375
+ $X2=0 $Y2=0
cc_355 N_A_27_88#_c_345_n N_A_287_464#_c_1801_n 4.55233e-19 $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_356 N_A_27_88#_M1015_g N_A_287_464#_c_1792_n 0.00771663f $X=2.28 $Y=2.64
+ $X2=0 $Y2=0
cc_357 N_A_27_88#_c_349_n N_A_287_464#_c_1807_n 0.0527651f $X=2.215 $Y=2.375
+ $X2=0 $Y2=0
cc_358 N_A_27_88#_M1015_g N_A_287_464#_c_1812_n 0.00419974f $X=2.28 $Y=2.64
+ $X2=0 $Y2=0
cc_359 N_A_27_88#_c_349_n N_A_287_464#_c_1812_n 0.0199552f $X=2.215 $Y=2.375
+ $X2=0 $Y2=0
cc_360 N_A_27_88#_c_349_n A_474_464# 0.00106497f $X=2.215 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_361 N_A_27_88#_c_338_n N_VGND_c_1933_n 0.0188413f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_362 N_A_27_88#_c_344_n N_VGND_c_1933_n 0.0279144f $X=1.29 $Y=1.087 $X2=0
+ $Y2=0
cc_363 N_A_27_88#_c_345_n N_VGND_c_1933_n 0.00400291f $X=1.455 $Y=0.935 $X2=0
+ $Y2=0
cc_364 N_A_27_88#_c_345_n N_VGND_c_1939_n 9.34861e-19 $X=1.455 $Y=0.935 $X2=0
+ $Y2=0
cc_365 N_A_27_88#_c_338_n N_VGND_c_1941_n 0.0113438f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_366 N_A_27_88#_c_338_n N_VGND_c_1947_n 0.011567f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_367 N_A_27_88#_c_342_n N_noxref_24_c_2058_n 0.0138157f $X=1.455 $Y=1.1 $X2=0
+ $Y2=0
cc_368 N_A_27_88#_c_343_n N_noxref_24_c_2058_n 0.00399118f $X=1.455 $Y=1.1 $X2=0
+ $Y2=0
cc_369 N_A_27_88#_c_344_n N_noxref_24_c_2058_n 0.00699077f $X=1.29 $Y=1.087
+ $X2=0 $Y2=0
cc_370 N_A_27_88#_c_345_n N_noxref_24_c_2058_n 0.0059422f $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_371 N_A_27_88#_c_342_n N_noxref_24_c_2059_n 0.00360351f $X=1.455 $Y=1.1 $X2=0
+ $Y2=0
cc_372 N_A_27_88#_c_345_n N_noxref_24_c_2059_n 0.00794258f $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_373 N_A_27_88#_c_345_n N_noxref_24_c_2060_n 0.00331383f $X=1.455 $Y=0.935
+ $X2=0 $Y2=0
cc_374 N_D_M1034_g N_VPWR_c_1648_n 0.00155004f $X=1.345 $Y=2.64 $X2=0 $Y2=0
cc_375 N_D_M1034_g N_VPWR_c_1657_n 0.00520332f $X=1.345 $Y=2.64 $X2=0 $Y2=0
cc_376 N_D_M1034_g N_VPWR_c_1647_n 0.00984812f $X=1.345 $Y=2.64 $X2=0 $Y2=0
cc_377 N_D_M1020_g N_A_287_464#_c_1801_n 0.00653506f $X=1.905 $Y=0.615 $X2=0
+ $Y2=0
cc_378 N_D_M1034_g N_A_287_464#_c_1807_n 0.00660409f $X=1.345 $Y=2.64 $X2=0
+ $Y2=0
cc_379 N_D_M1020_g N_VGND_c_1939_n 9.15902e-19 $X=1.905 $Y=0.615 $X2=0 $Y2=0
cc_380 N_D_M1020_g N_noxref_24_c_2058_n 0.00131656f $X=1.905 $Y=0.615 $X2=0
+ $Y2=0
cc_381 N_D_M1020_g N_noxref_24_c_2059_n 0.0127325f $X=1.905 $Y=0.615 $X2=0 $Y2=0
cc_382 N_SCD_c_468_n N_RESET_B_M1002_g 0.0223391f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_383 N_SCD_M1032_g N_RESET_B_M1023_g 0.0388967f $X=3.005 $Y=0.615 $X2=0 $Y2=0
cc_384 N_SCD_c_469_n N_RESET_B_c_840_n 0.00563201f $X=2.875 $Y=2.095 $X2=0 $Y2=0
cc_385 N_SCD_c_470_n N_RESET_B_c_840_n 0.00865744f $X=2.875 $Y=2.17 $X2=0 $Y2=0
cc_386 SCD N_RESET_B_c_840_n 0.00370213f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_387 SCD N_RESET_B_c_845_n 0.00160474f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_388 SCD N_RESET_B_c_849_n 0.00478487f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_389 N_SCD_c_467_n N_RESET_B_c_849_n 0.0173672f $X=2.965 $Y=1.69 $X2=0 $Y2=0
cc_390 N_SCD_M1032_g N_RESET_B_c_850_n 9.76155e-19 $X=3.005 $Y=0.615 $X2=0 $Y2=0
cc_391 SCD N_RESET_B_c_850_n 0.0388123f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_392 N_SCD_c_467_n N_RESET_B_c_850_n 3.23745e-19 $X=2.965 $Y=1.69 $X2=0 $Y2=0
cc_393 N_SCD_c_468_n N_VPWR_c_1657_n 0.0037725f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_394 N_SCD_c_468_n N_VPWR_c_1647_n 0.00466028f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_395 N_SCD_c_468_n N_VPWR_c_1666_n 0.00349255f $X=2.67 $Y=2.245 $X2=0 $Y2=0
cc_396 N_SCD_c_468_n N_A_287_464#_c_1792_n 0.0178602f $X=2.67 $Y=2.245 $X2=0
+ $Y2=0
cc_397 N_SCD_c_470_n N_A_287_464#_c_1792_n 0.00391719f $X=2.875 $Y=2.17 $X2=0
+ $Y2=0
cc_398 SCD N_A_287_464#_c_1792_n 0.0148645f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_399 N_SCD_M1032_g N_A_287_464#_c_1787_n 0.00339631f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_400 N_SCD_M1032_g N_A_287_464#_c_1788_n 0.014248f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_401 SCD N_A_287_464#_c_1788_n 0.0164273f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_402 N_SCD_c_467_n N_A_287_464#_c_1788_n 5.59028e-19 $X=2.965 $Y=1.69 $X2=0
+ $Y2=0
cc_403 SCD N_A_287_464#_c_1789_n 0.00463754f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_404 N_SCD_c_467_n N_A_287_464#_c_1789_n 6.23418e-19 $X=2.965 $Y=1.69 $X2=0
+ $Y2=0
cc_405 SCD N_A_287_464#_c_1790_n 0.00365391f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_406 N_SCD_c_468_n N_A_287_464#_c_1812_n 7.62723e-19 $X=2.67 $Y=2.245 $X2=0
+ $Y2=0
cc_407 N_SCD_M1032_g N_VGND_c_1939_n 9.34905e-19 $X=3.005 $Y=0.615 $X2=0 $Y2=0
cc_408 N_SCD_M1032_g N_noxref_24_c_2059_n 0.0107848f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_409 N_SCD_M1032_g N_noxref_24_c_2063_n 0.0049663f $X=3.005 $Y=0.615 $X2=0
+ $Y2=0
cc_410 N_CLK_N_c_514_n N_RESET_B_M1023_g 0.00177089f $X=4.62 $Y=1.435 $X2=0
+ $Y2=0
cc_411 N_CLK_N_c_516_n N_RESET_B_c_857_n 0.0121828f $X=4.71 $Y=1.66 $X2=0 $Y2=0
cc_412 N_CLK_N_c_516_n N_RESET_B_c_844_n 0.00390613f $X=4.71 $Y=1.66 $X2=0 $Y2=0
cc_413 N_CLK_N_c_514_n N_RESET_B_c_844_n 0.0135682f $X=4.62 $Y=1.435 $X2=0 $Y2=0
cc_414 N_CLK_N_c_515_n N_RESET_B_c_844_n 0.00314445f $X=4.71 $Y=1.435 $X2=0
+ $Y2=0
cc_415 CLK_N N_RESET_B_c_844_n 0.0110696f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_416 N_CLK_N_c_514_n N_RESET_B_c_849_n 0.00816712f $X=4.62 $Y=1.435 $X2=0
+ $Y2=0
cc_417 N_CLK_N_c_513_n N_A_859_347#_c_1165_n 0.0196943f $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_418 N_CLK_N_c_516_n N_A_859_347#_c_1183_n 0.0327358f $X=4.71 $Y=1.66 $X2=0
+ $Y2=0
cc_419 N_CLK_N_c_516_n N_A_859_347#_c_1196_n 0.0110526f $X=4.71 $Y=1.66 $X2=0
+ $Y2=0
cc_420 N_CLK_N_c_514_n N_A_859_347#_c_1196_n 0.00572759f $X=4.62 $Y=1.435 $X2=0
+ $Y2=0
cc_421 CLK_N N_A_859_347#_c_1196_n 0.0107345f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_422 N_CLK_N_c_513_n N_A_859_347#_c_1199_n 0.00558688f $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_423 N_CLK_N_c_513_n N_A_859_347#_c_1200_n 0.0120157f $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_424 CLK_N N_A_859_347#_c_1200_n 8.89317e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_425 N_CLK_N_c_513_n N_A_859_347#_c_1202_n 2.94796e-19 $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_426 N_CLK_N_c_514_n N_A_859_347#_c_1202_n 0.00775189f $X=4.62 $Y=1.435 $X2=0
+ $Y2=0
cc_427 CLK_N N_A_859_347#_c_1202_n 0.0210647f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_428 N_CLK_N_c_516_n N_A_859_347#_c_1189_n 0.00461919f $X=4.71 $Y=1.66 $X2=0
+ $Y2=0
cc_429 N_CLK_N_c_515_n N_A_859_347#_c_1175_n 0.00461919f $X=4.71 $Y=1.435 $X2=0
+ $Y2=0
cc_430 N_CLK_N_c_513_n N_A_859_347#_c_1176_n 0.00461919f $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_431 CLK_N N_A_859_347#_c_1176_n 0.0196445f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_432 N_CLK_N_c_515_n N_A_859_347#_c_1182_n 0.0238821f $X=4.71 $Y=1.435 $X2=0
+ $Y2=0
cc_433 CLK_N N_A_859_347#_c_1182_n 3.02818e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_434 N_CLK_N_c_516_n N_VPWR_c_1649_n 0.00495808f $X=4.71 $Y=1.66 $X2=0 $Y2=0
cc_435 N_CLK_N_c_516_n N_VPWR_c_1647_n 0.00112709f $X=4.71 $Y=1.66 $X2=0 $Y2=0
cc_436 N_CLK_N_c_513_n N_A_287_464#_c_1788_n 0.00360967f $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_437 N_CLK_N_c_516_n N_A_287_464#_c_1790_n 0.00488914f $X=4.71 $Y=1.66 $X2=0
+ $Y2=0
cc_438 N_CLK_N_c_513_n N_A_287_464#_c_1790_n 5.39083e-19 $X=4.725 $Y=1.21 $X2=0
+ $Y2=0
cc_439 N_CLK_N_c_514_n N_A_287_464#_c_1790_n 0.00690074f $X=4.62 $Y=1.435 $X2=0
+ $Y2=0
cc_440 CLK_N N_A_287_464#_c_1790_n 0.0229056f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_441 N_CLK_N_c_514_n N_A_287_464#_c_1794_n 0.00379856f $X=4.62 $Y=1.435 $X2=0
+ $Y2=0
cc_442 CLK_N N_A_287_464#_c_1794_n 4.23593e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_443 N_CLK_N_c_516_n N_A_287_464#_c_1795_n 0.0174245f $X=4.71 $Y=1.66 $X2=0
+ $Y2=0
cc_444 N_CLK_N_c_516_n N_A_287_464#_c_1835_n 0.00886305f $X=4.71 $Y=1.66 $X2=0
+ $Y2=0
cc_445 N_CLK_N_c_513_n N_VGND_c_1934_n 0.00314573f $X=4.725 $Y=1.21 $X2=0 $Y2=0
cc_446 N_CLK_N_c_513_n N_VGND_c_1935_n 0.00534919f $X=4.725 $Y=1.21 $X2=0 $Y2=0
cc_447 N_CLK_N_c_513_n N_VGND_c_1942_n 0.00451627f $X=4.725 $Y=1.21 $X2=0 $Y2=0
cc_448 N_CLK_N_c_513_n N_VGND_c_1947_n 0.00454582f $X=4.725 $Y=1.21 $X2=0 $Y2=0
cc_449 N_A_1069_74#_c_581_p N_A_1417_294#_M1035_d 0.00239218f $X=8.39 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_450 N_A_1069_74#_c_569_n N_A_1417_294#_M1035_d 6.37056e-19 $X=8.475 $Y=0.79
+ $X2=-0.19 $Y2=-0.245
cc_451 N_A_1069_74#_c_575_n N_A_1417_294#_M1033_g 0.0456844f $X=6.815 $Y=2.055
+ $X2=0 $Y2=0
cc_452 N_A_1069_74#_c_562_n N_A_1417_294#_M1033_g 0.00769677f $X=6.815 $Y=1.965
+ $X2=0 $Y2=0
cc_453 N_A_1069_74#_c_566_n N_A_1417_294#_M1016_g 0.00312043f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_454 N_A_1069_74#_c_568_n N_A_1417_294#_M1016_g 0.00336294f $X=7.175 $Y=0.79
+ $X2=0 $Y2=0
cc_455 N_A_1069_74#_c_581_p N_A_1417_294#_M1016_g 0.00839835f $X=8.39 $Y=0.875
+ $X2=0 $Y2=0
cc_456 N_A_1069_74#_c_581_p N_A_1417_294#_c_743_n 0.0681288f $X=8.39 $Y=0.875
+ $X2=0 $Y2=0
cc_457 N_A_1069_74#_c_570_n N_A_1417_294#_c_743_n 0.00503881f $X=9.07 $Y=0.445
+ $X2=0 $Y2=0
cc_458 N_A_1069_74#_c_581_p N_A_1417_294#_c_744_n 0.0116449f $X=8.39 $Y=0.875
+ $X2=0 $Y2=0
cc_459 N_A_1069_74#_c_581_p N_A_1417_294#_c_745_n 0.0138309f $X=8.39 $Y=0.875
+ $X2=0 $Y2=0
cc_460 N_A_1069_74#_c_569_n N_A_1417_294#_c_745_n 0.00655386f $X=8.475 $Y=0.79
+ $X2=0 $Y2=0
cc_461 N_A_1069_74#_c_570_n N_A_1417_294#_c_745_n 0.013545f $X=9.07 $Y=0.445
+ $X2=0 $Y2=0
cc_462 N_A_1069_74#_c_594_p N_A_1417_294#_c_745_n 0.0231598f $X=9.155 $Y=1.03
+ $X2=0 $Y2=0
cc_463 N_A_1069_74#_c_595_p N_A_1417_294#_c_745_n 0.00782335f $X=9.24 $Y=1.115
+ $X2=0 $Y2=0
cc_464 N_A_1069_74#_M1031_g N_A_1417_294#_c_751_n 5.12299e-19 $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_465 N_A_1069_74#_c_566_n N_A_1417_294#_c_746_n 0.00175583f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_466 N_A_1069_74#_c_598_p N_A_1417_294#_c_746_n 0.00434364f $X=7.26 $Y=0.875
+ $X2=0 $Y2=0
cc_467 N_A_1069_74#_c_566_n N_A_1417_294#_c_747_n 0.021484f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_468 N_A_1069_74#_c_598_p N_A_1417_294#_c_747_n 7.88542e-19 $X=7.26 $Y=0.875
+ $X2=0 $Y2=0
cc_469 N_A_1069_74#_c_566_n N_A_1417_294#_c_748_n 4.18248e-19 $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_470 N_A_1069_74#_c_595_p N_A_1417_294#_c_776_n 0.00611823f $X=9.24 $Y=1.115
+ $X2=0 $Y2=0
cc_471 N_A_1069_74#_M1031_g N_A_1417_294#_c_749_n 0.00357144f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_472 N_A_1069_74#_M1024_g N_RESET_B_c_857_n 0.0102711f $X=6.815 $Y=2.495 $X2=0
+ $Y2=0
cc_473 N_A_1069_74#_c_581_p N_RESET_B_M1003_g 0.0102621f $X=8.39 $Y=0.875 $X2=0
+ $Y2=0
cc_474 N_A_1069_74#_c_569_n N_RESET_B_M1003_g 7.6286e-19 $X=8.475 $Y=0.79 $X2=0
+ $Y2=0
cc_475 N_A_1069_74#_M1029_d N_RESET_B_c_844_n 5.99887e-19 $X=5.385 $Y=1.735
+ $X2=0 $Y2=0
cc_476 N_A_1069_74#_c_575_n N_RESET_B_c_844_n 8.06642e-19 $X=6.815 $Y=2.055
+ $X2=0 $Y2=0
cc_477 N_A_1069_74#_c_562_n N_RESET_B_c_844_n 9.24483e-19 $X=6.815 $Y=1.965
+ $X2=0 $Y2=0
cc_478 N_A_1069_74#_c_565_n N_RESET_B_c_844_n 0.0148121f $X=6.415 $Y=1.43 $X2=0
+ $Y2=0
cc_479 N_A_1069_74#_c_566_n N_RESET_B_c_844_n 0.0067912f $X=6.415 $Y=1.43 $X2=0
+ $Y2=0
cc_480 N_A_1069_74#_c_579_n N_RESET_B_c_844_n 0.00536125f $X=5.525 $Y=1.915
+ $X2=0 $Y2=0
cc_481 N_A_1069_74#_c_573_n N_RESET_B_c_844_n 0.025807f $X=5.547 $Y=1.745 $X2=0
+ $Y2=0
cc_482 N_A_1069_74#_c_614_p N_RESET_B_c_844_n 5.77133e-19 $X=5.587 $Y=1.09 $X2=0
+ $Y2=0
cc_483 N_A_1069_74#_M1031_g N_RESET_B_c_846_n 0.0112916f $X=9.62 $Y=2.46 $X2=0
+ $Y2=0
cc_484 N_A_1069_74#_c_595_p N_RESET_B_c_846_n 8.63692e-19 $X=9.24 $Y=1.115 $X2=0
+ $Y2=0
cc_485 N_A_1069_74#_c_572_n N_RESET_B_c_846_n 0.00134553f $X=9.66 $Y=1.115 $X2=0
+ $Y2=0
cc_486 N_A_1069_74#_c_565_n N_A_1273_131#_M1021_d 0.00383506f $X=6.415 $Y=1.43
+ $X2=-0.19 $Y2=-0.245
cc_487 N_A_1069_74#_c_581_p N_A_1273_131#_c_1060_n 0.0104263f $X=8.39 $Y=0.875
+ $X2=0 $Y2=0
cc_488 N_A_1069_74#_c_569_n N_A_1273_131#_c_1060_n 0.00662009f $X=8.475 $Y=0.79
+ $X2=0 $Y2=0
cc_489 N_A_1069_74#_M1021_g N_A_1273_131#_c_1061_n 0.00193761f $X=6.29 $Y=0.865
+ $X2=0 $Y2=0
cc_490 N_A_1069_74#_c_565_n N_A_1273_131#_c_1061_n 0.0755826f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_491 N_A_1069_74#_c_567_n N_A_1273_131#_c_1061_n 0.0196961f $X=7.09 $Y=0.36
+ $X2=0 $Y2=0
cc_492 N_A_1069_74#_c_568_n N_A_1273_131#_c_1061_n 0.00628856f $X=7.175 $Y=0.79
+ $X2=0 $Y2=0
cc_493 N_A_1069_74#_c_562_n N_A_1273_131#_c_1062_n 0.0127359f $X=6.815 $Y=1.965
+ $X2=0 $Y2=0
cc_494 N_A_1069_74#_c_566_n N_A_1273_131#_c_1062_n 0.0144475f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_495 N_A_1069_74#_c_575_n N_A_1273_131#_c_1067_n 0.00210344f $X=6.815 $Y=2.055
+ $X2=0 $Y2=0
cc_496 N_A_1069_74#_M1024_g N_A_1273_131#_c_1067_n 0.00440834f $X=6.815 $Y=2.495
+ $X2=0 $Y2=0
cc_497 N_A_1069_74#_c_575_n N_A_1273_131#_c_1068_n 0.00228851f $X=6.815 $Y=2.055
+ $X2=0 $Y2=0
cc_498 N_A_1069_74#_M1024_g N_A_1273_131#_c_1068_n 0.0174754f $X=6.815 $Y=2.495
+ $X2=0 $Y2=0
cc_499 N_A_1069_74#_c_565_n N_A_1273_131#_c_1068_n 0.00150496f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_500 N_A_1069_74#_c_566_n N_A_1273_131#_c_1068_n 0.00347443f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_501 N_A_1069_74#_c_564_n N_A_859_347#_c_1165_n 0.00173447f $X=5.735 $Y=0.36
+ $X2=0 $Y2=0
cc_502 N_A_1069_74#_c_573_n N_A_859_347#_c_1165_n 8.38974e-19 $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_503 N_A_1069_74#_c_579_n N_A_859_347#_c_1183_n 0.00356981f $X=5.525 $Y=1.915
+ $X2=0 $Y2=0
cc_504 N_A_1069_74#_c_573_n N_A_859_347#_c_1183_n 6.09784e-19 $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_505 N_A_1069_74#_M1021_g N_A_859_347#_c_1166_n 0.0138755f $X=6.29 $Y=0.865
+ $X2=0 $Y2=0
cc_506 N_A_1069_74#_c_638_p N_A_859_347#_c_1166_n 0.0117407f $X=5.525 $Y=0.56
+ $X2=0 $Y2=0
cc_507 N_A_1069_74#_c_563_n N_A_859_347#_c_1166_n 0.0130864f $X=6.33 $Y=0.36
+ $X2=0 $Y2=0
cc_508 N_A_1069_74#_c_564_n N_A_859_347#_c_1166_n 0.00276418f $X=5.735 $Y=0.36
+ $X2=0 $Y2=0
cc_509 N_A_1069_74#_c_565_n N_A_859_347#_c_1166_n 7.73946e-19 $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_510 N_A_1069_74#_c_573_n N_A_859_347#_c_1166_n 0.00249267f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_511 N_A_1069_74#_c_614_p N_A_859_347#_c_1166_n 0.00318247f $X=5.587 $Y=1.09
+ $X2=0 $Y2=0
cc_512 N_A_1069_74#_c_579_n N_A_859_347#_c_1167_n 0.00665735f $X=5.525 $Y=1.915
+ $X2=0 $Y2=0
cc_513 N_A_1069_74#_c_573_n N_A_859_347#_c_1167_n 0.00145048f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_514 N_A_1069_74#_M1021_g N_A_859_347#_c_1168_n 0.00902735f $X=6.29 $Y=0.865
+ $X2=0 $Y2=0
cc_515 N_A_1069_74#_c_563_n N_A_859_347#_c_1168_n 0.00670492f $X=6.33 $Y=0.36
+ $X2=0 $Y2=0
cc_516 N_A_1069_74#_c_567_n N_A_859_347#_c_1168_n 0.0072068f $X=7.09 $Y=0.36
+ $X2=0 $Y2=0
cc_517 N_A_1069_74#_c_649_p N_A_859_347#_c_1168_n 0.0036181f $X=6.415 $Y=0.36
+ $X2=0 $Y2=0
cc_518 N_A_1069_74#_M1024_g N_A_859_347#_c_1185_n 0.0188017f $X=6.815 $Y=2.495
+ $X2=0 $Y2=0
cc_519 N_A_1069_74#_c_565_n N_A_859_347#_c_1185_n 0.00160792f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_520 N_A_1069_74#_c_566_n N_A_859_347#_c_1185_n 0.00597277f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_521 N_A_1069_74#_M1021_g N_A_859_347#_M1028_g 0.0094641f $X=6.29 $Y=0.865
+ $X2=0 $Y2=0
cc_522 N_A_1069_74#_c_565_n N_A_859_347#_M1028_g 0.00210048f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_523 N_A_1069_74#_c_567_n N_A_859_347#_M1028_g 0.0191653f $X=7.09 $Y=0.36
+ $X2=0 $Y2=0
cc_524 N_A_1069_74#_c_568_n N_A_859_347#_M1028_g 0.00256248f $X=7.175 $Y=0.79
+ $X2=0 $Y2=0
cc_525 N_A_1069_74#_c_567_n N_A_859_347#_c_1171_n 0.00443325f $X=7.09 $Y=0.36
+ $X2=0 $Y2=0
cc_526 N_A_1069_74#_c_581_p N_A_859_347#_c_1171_n 0.00821493f $X=8.39 $Y=0.875
+ $X2=0 $Y2=0
cc_527 N_A_1069_74#_c_570_n N_A_859_347#_c_1171_n 0.00736464f $X=9.07 $Y=0.445
+ $X2=0 $Y2=0
cc_528 N_A_1069_74#_c_571_n N_A_859_347#_c_1171_n 0.00348338f $X=8.56 $Y=0.445
+ $X2=0 $Y2=0
cc_529 N_A_1069_74#_M1031_g N_A_859_347#_M1039_g 0.00578589f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_530 N_A_1069_74#_c_569_n N_A_859_347#_M1039_g 0.00193414f $X=8.475 $Y=0.79
+ $X2=0 $Y2=0
cc_531 N_A_1069_74#_c_570_n N_A_859_347#_M1039_g 0.0147282f $X=9.07 $Y=0.445
+ $X2=0 $Y2=0
cc_532 N_A_1069_74#_c_594_p N_A_859_347#_M1039_g 0.0152559f $X=9.155 $Y=1.03
+ $X2=0 $Y2=0
cc_533 N_A_1069_74#_c_595_p N_A_859_347#_M1039_g 0.00557926f $X=9.24 $Y=1.115
+ $X2=0 $Y2=0
cc_534 N_A_1069_74#_c_574_n N_A_859_347#_M1039_g 0.0118451f $X=9.66 $Y=1.005
+ $X2=0 $Y2=0
cc_535 N_A_1069_74#_c_638_p N_A_859_347#_c_1200_n 0.0163074f $X=5.525 $Y=0.56
+ $X2=0 $Y2=0
cc_536 N_A_1069_74#_c_573_n N_A_859_347#_c_1189_n 0.00686016f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_537 N_A_1069_74#_c_573_n N_A_859_347#_c_1175_n 0.0263792f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_538 N_A_1069_74#_c_573_n N_A_859_347#_c_1176_n 0.00877966f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_539 N_A_1069_74#_c_614_p N_A_859_347#_c_1176_n 0.00611922f $X=5.587 $Y=1.09
+ $X2=0 $Y2=0
cc_540 N_A_1069_74#_M1031_g N_A_859_347#_c_1177_n 0.00391639f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_541 N_A_1069_74#_c_595_p N_A_859_347#_c_1177_n 0.0115051f $X=9.24 $Y=1.115
+ $X2=0 $Y2=0
cc_542 N_A_1069_74#_c_572_n N_A_859_347#_c_1177_n 0.00828947f $X=9.66 $Y=1.115
+ $X2=0 $Y2=0
cc_543 N_A_1069_74#_M1031_g N_A_859_347#_c_1178_n 0.0211354f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_544 N_A_1069_74#_c_595_p N_A_859_347#_c_1178_n 5.03607e-19 $X=9.24 $Y=1.115
+ $X2=0 $Y2=0
cc_545 N_A_1069_74#_c_572_n N_A_859_347#_c_1178_n 4.33652e-19 $X=9.66 $Y=1.115
+ $X2=0 $Y2=0
cc_546 N_A_1069_74#_M1031_g N_A_859_347#_c_1179_n 4.66885e-19 $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_547 N_A_1069_74#_c_560_n N_A_859_347#_c_1179_n 0.00120212f $X=10.215 $Y=1.005
+ $X2=0 $Y2=0
cc_548 N_A_1069_74#_M1031_g N_A_859_347#_c_1180_n 0.041812f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_549 N_A_1069_74#_c_560_n N_A_859_347#_c_1180_n 0.0209009f $X=10.215 $Y=1.005
+ $X2=0 $Y2=0
cc_550 N_A_1069_74#_M1031_g N_A_859_347#_c_1181_n 0.0116557f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_551 N_A_1069_74#_c_560_n N_A_859_347#_c_1181_n 0.00433131f $X=10.215 $Y=1.005
+ $X2=0 $Y2=0
cc_552 N_A_1069_74#_c_572_n N_A_859_347#_c_1181_n 0.0321071f $X=9.66 $Y=1.115
+ $X2=0 $Y2=0
cc_553 N_A_1069_74#_c_574_n N_A_859_347#_c_1181_n 0.00374181f $X=9.66 $Y=1.005
+ $X2=0 $Y2=0
cc_554 N_A_1069_74#_c_566_n N_A_859_347#_c_1182_n 0.0138755f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_555 N_A_1069_74#_c_573_n N_A_859_347#_c_1182_n 0.0281923f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_556 N_A_1069_74#_c_614_p N_A_859_347#_c_1182_n 0.0010507f $X=5.587 $Y=1.09
+ $X2=0 $Y2=0
cc_557 N_A_1069_74#_M1026_g N_A_2087_410#_M1004_g 0.0421839f $X=10.29 $Y=0.58
+ $X2=0 $Y2=0
cc_558 N_A_1069_74#_c_570_n N_A_1827_144#_M1039_d 0.00791052f $X=9.07 $Y=0.445
+ $X2=-0.19 $Y2=-0.245
cc_559 N_A_1069_74#_c_594_p N_A_1827_144#_M1039_d 0.00742046f $X=9.155 $Y=1.03
+ $X2=-0.19 $Y2=-0.245
cc_560 N_A_1069_74#_c_595_p N_A_1827_144#_M1039_d 4.16738e-19 $X=9.24 $Y=1.115
+ $X2=-0.19 $Y2=-0.245
cc_561 N_A_1069_74#_c_572_n N_A_1827_144#_M1039_d 0.00680879f $X=9.66 $Y=1.115
+ $X2=-0.19 $Y2=-0.245
cc_562 N_A_1069_74#_c_560_n N_A_1827_144#_c_1464_n 0.0063315f $X=10.215 $Y=1.005
+ $X2=0 $Y2=0
cc_563 N_A_1069_74#_M1026_g N_A_1827_144#_c_1464_n 0.0175228f $X=10.29 $Y=0.58
+ $X2=0 $Y2=0
cc_564 N_A_1069_74#_c_594_p N_A_1827_144#_c_1464_n 0.0266854f $X=9.155 $Y=1.03
+ $X2=0 $Y2=0
cc_565 N_A_1069_74#_c_572_n N_A_1827_144#_c_1464_n 0.0319013f $X=9.66 $Y=1.115
+ $X2=0 $Y2=0
cc_566 N_A_1069_74#_c_574_n N_A_1827_144#_c_1464_n 0.0196311f $X=9.66 $Y=1.005
+ $X2=0 $Y2=0
cc_567 N_A_1069_74#_M1031_g N_A_1827_144#_c_1473_n 0.00248113f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_568 N_A_1069_74#_M1031_g N_A_1827_144#_c_1475_n 0.00388519f $X=9.62 $Y=2.46
+ $X2=0 $Y2=0
cc_569 N_A_1069_74#_M1024_g N_VPWR_c_1650_n 0.00156346f $X=6.815 $Y=2.495 $X2=0
+ $Y2=0
cc_570 N_A_1069_74#_M1031_g N_VPWR_c_1661_n 0.00553757f $X=9.62 $Y=2.46 $X2=0
+ $Y2=0
cc_571 N_A_1069_74#_M1024_g N_VPWR_c_1647_n 0.00113998f $X=6.815 $Y=2.495 $X2=0
+ $Y2=0
cc_572 N_A_1069_74#_M1031_g N_VPWR_c_1647_n 0.0109558f $X=9.62 $Y=2.46 $X2=0
+ $Y2=0
cc_573 N_A_1069_74#_M1029_d N_A_287_464#_c_1795_n 0.00576874f $X=5.385 $Y=1.735
+ $X2=0 $Y2=0
cc_574 N_A_1069_74#_c_579_n N_A_287_464#_c_1795_n 0.0247182f $X=5.525 $Y=1.915
+ $X2=0 $Y2=0
cc_575 N_A_1069_74#_M1021_g N_A_287_464#_c_1791_n 0.00499753f $X=6.29 $Y=0.865
+ $X2=0 $Y2=0
cc_576 N_A_1069_74#_c_562_n N_A_287_464#_c_1791_n 8.49879e-19 $X=6.815 $Y=1.965
+ $X2=0 $Y2=0
cc_577 N_A_1069_74#_c_638_p N_A_287_464#_c_1791_n 0.0340491f $X=5.525 $Y=0.56
+ $X2=0 $Y2=0
cc_578 N_A_1069_74#_c_563_n N_A_287_464#_c_1791_n 0.0200637f $X=6.33 $Y=0.36
+ $X2=0 $Y2=0
cc_579 N_A_1069_74#_c_565_n N_A_287_464#_c_1791_n 0.0592862f $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_580 N_A_1069_74#_c_562_n N_A_287_464#_c_1797_n 6.25019e-19 $X=6.815 $Y=1.965
+ $X2=0 $Y2=0
cc_581 N_A_1069_74#_c_566_n N_A_287_464#_c_1797_n 5.02733e-19 $X=6.415 $Y=1.43
+ $X2=0 $Y2=0
cc_582 N_A_1069_74#_c_614_p N_A_287_464#_c_1797_n 0.0340491f $X=5.587 $Y=1.09
+ $X2=0 $Y2=0
cc_583 N_A_1069_74#_c_575_n N_A_287_464#_c_1798_n 6.25019e-19 $X=6.815 $Y=2.055
+ $X2=0 $Y2=0
cc_584 N_A_1069_74#_c_573_n N_A_287_464#_c_1798_n 0.0340491f $X=5.547 $Y=1.745
+ $X2=0 $Y2=0
cc_585 N_A_1069_74#_c_581_p N_VGND_M1003_d 0.00871171f $X=8.39 $Y=0.875 $X2=0
+ $Y2=0
cc_586 N_A_1069_74#_c_564_n N_VGND_c_1935_n 0.0102123f $X=5.735 $Y=0.36 $X2=0
+ $Y2=0
cc_587 N_A_1069_74#_c_567_n N_VGND_c_1936_n 0.00743709f $X=7.09 $Y=0.36 $X2=0
+ $Y2=0
cc_588 N_A_1069_74#_c_568_n N_VGND_c_1936_n 0.00483194f $X=7.175 $Y=0.79 $X2=0
+ $Y2=0
cc_589 N_A_1069_74#_c_581_p N_VGND_c_1936_n 0.0260918f $X=8.39 $Y=0.875 $X2=0
+ $Y2=0
cc_590 N_A_1069_74#_c_569_n N_VGND_c_1936_n 0.00698435f $X=8.475 $Y=0.79 $X2=0
+ $Y2=0
cc_591 N_A_1069_74#_c_571_n N_VGND_c_1936_n 0.0150385f $X=8.56 $Y=0.445 $X2=0
+ $Y2=0
cc_592 N_A_1069_74#_M1026_g N_VGND_c_1937_n 0.00160614f $X=10.29 $Y=0.58 $X2=0
+ $Y2=0
cc_593 N_A_1069_74#_c_563_n N_VGND_c_1943_n 0.0384101f $X=6.33 $Y=0.36 $X2=0
+ $Y2=0
cc_594 N_A_1069_74#_c_564_n N_VGND_c_1943_n 0.0211124f $X=5.735 $Y=0.36 $X2=0
+ $Y2=0
cc_595 N_A_1069_74#_c_567_n N_VGND_c_1943_n 0.0496716f $X=7.09 $Y=0.36 $X2=0
+ $Y2=0
cc_596 N_A_1069_74#_c_649_p N_VGND_c_1943_n 0.0115893f $X=6.415 $Y=0.36 $X2=0
+ $Y2=0
cc_597 N_A_1069_74#_M1026_g N_VGND_c_1944_n 0.00315309f $X=10.29 $Y=0.58 $X2=0
+ $Y2=0
cc_598 N_A_1069_74#_c_570_n N_VGND_c_1944_n 0.0266206f $X=9.07 $Y=0.445 $X2=0
+ $Y2=0
cc_599 N_A_1069_74#_c_571_n N_VGND_c_1944_n 0.00722011f $X=8.56 $Y=0.445 $X2=0
+ $Y2=0
cc_600 N_A_1069_74#_M1026_g N_VGND_c_1947_n 0.00393098f $X=10.29 $Y=0.58 $X2=0
+ $Y2=0
cc_601 N_A_1069_74#_c_563_n N_VGND_c_1947_n 0.0199841f $X=6.33 $Y=0.36 $X2=0
+ $Y2=0
cc_602 N_A_1069_74#_c_564_n N_VGND_c_1947_n 0.0114232f $X=5.735 $Y=0.36 $X2=0
+ $Y2=0
cc_603 N_A_1069_74#_c_567_n N_VGND_c_1947_n 0.025617f $X=7.09 $Y=0.36 $X2=0
+ $Y2=0
cc_604 N_A_1069_74#_c_581_p N_VGND_c_1947_n 0.0255776f $X=8.39 $Y=0.875 $X2=0
+ $Y2=0
cc_605 N_A_1069_74#_c_570_n N_VGND_c_1947_n 0.0216892f $X=9.07 $Y=0.445 $X2=0
+ $Y2=0
cc_606 N_A_1069_74#_c_571_n N_VGND_c_1947_n 0.00553204f $X=8.56 $Y=0.445 $X2=0
+ $Y2=0
cc_607 N_A_1069_74#_c_649_p N_VGND_c_1947_n 0.00583135f $X=6.415 $Y=0.36 $X2=0
+ $Y2=0
cc_608 N_A_1069_74#_c_598_p A_1409_131# 0.00171413f $X=7.26 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_609 N_A_1069_74#_c_581_p A_1483_131# 0.00179164f $X=8.39 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_610 N_A_1417_294#_M1033_g N_RESET_B_c_857_n 0.0107325f $X=7.235 $Y=2.495
+ $X2=0 $Y2=0
cc_611 N_A_1417_294#_M1016_g N_RESET_B_M1003_g 0.0422504f $X=7.34 $Y=0.865 $X2=0
+ $Y2=0
cc_612 N_A_1417_294#_c_743_n N_RESET_B_M1003_g 0.0112845f $X=8.73 $Y=1.215 $X2=0
+ $Y2=0
cc_613 N_A_1417_294#_c_748_n N_RESET_B_M1003_g 0.00117015f $X=7.245 $Y=1.47
+ $X2=0 $Y2=0
cc_614 N_A_1417_294#_M1033_g N_RESET_B_M1030_g 0.0283629f $X=7.235 $Y=2.495
+ $X2=0 $Y2=0
cc_615 N_A_1417_294#_c_743_n N_RESET_B_c_844_n 0.00704635f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_616 N_A_1417_294#_c_746_n N_RESET_B_c_844_n 0.028548f $X=7.25 $Y=1.635 $X2=0
+ $Y2=0
cc_617 N_A_1417_294#_c_747_n N_RESET_B_c_844_n 6.94548e-19 $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_618 N_A_1417_294#_c_743_n N_RESET_B_c_846_n 0.0146017f $X=8.73 $Y=1.215 $X2=0
+ $Y2=0
cc_619 N_A_1417_294#_c_787_p N_RESET_B_c_846_n 0.0143525f $X=8.96 $Y=2.135 $X2=0
+ $Y2=0
cc_620 N_A_1417_294#_c_749_n N_RESET_B_c_846_n 0.0234363f $X=9.112 $Y=1.97 $X2=0
+ $Y2=0
cc_621 N_A_1417_294#_c_743_n N_RESET_B_c_847_n 0.00253594f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_622 N_A_1417_294#_c_746_n N_RESET_B_c_847_n 4.91583e-19 $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_623 N_A_1417_294#_c_743_n N_RESET_B_c_851_n 0.00549913f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_624 N_A_1417_294#_c_746_n N_RESET_B_c_851_n 0.00117015f $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_625 N_A_1417_294#_c_747_n N_RESET_B_c_851_n 0.0422504f $X=7.25 $Y=1.635 $X2=0
+ $Y2=0
cc_626 N_A_1417_294#_c_743_n N_RESET_B_c_852_n 0.0260743f $X=8.73 $Y=1.215 $X2=0
+ $Y2=0
cc_627 N_A_1417_294#_c_746_n N_RESET_B_c_852_n 0.0165906f $X=7.25 $Y=1.635 $X2=0
+ $Y2=0
cc_628 N_A_1417_294#_c_747_n N_RESET_B_c_852_n 0.00108705f $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_629 N_A_1417_294#_c_743_n N_A_1273_131#_c_1060_n 0.012315f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_630 N_A_1417_294#_c_745_n N_A_1273_131#_c_1060_n 0.0040669f $X=8.815 $Y=0.865
+ $X2=0 $Y2=0
cc_631 N_A_1417_294#_c_749_n N_A_1273_131#_c_1060_n 0.00333382f $X=9.112 $Y=1.97
+ $X2=0 $Y2=0
cc_632 N_A_1417_294#_c_751_n N_A_1273_131#_M1038_g 4.93842e-19 $X=8.96 $Y=2.815
+ $X2=0 $Y2=0
cc_633 N_A_1417_294#_c_787_p N_A_1273_131#_M1038_g 0.00529099f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_634 N_A_1417_294#_c_749_n N_A_1273_131#_M1038_g 0.00512316f $X=9.112 $Y=1.97
+ $X2=0 $Y2=0
cc_635 N_A_1417_294#_M1033_g N_A_1273_131#_c_1062_n 0.00103339f $X=7.235
+ $Y=2.495 $X2=0 $Y2=0
cc_636 N_A_1417_294#_M1016_g N_A_1273_131#_c_1062_n 0.00102076f $X=7.34 $Y=0.865
+ $X2=0 $Y2=0
cc_637 N_A_1417_294#_c_744_n N_A_1273_131#_c_1062_n 0.00815829f $X=7.415
+ $Y=1.215 $X2=0 $Y2=0
cc_638 N_A_1417_294#_c_746_n N_A_1273_131#_c_1062_n 0.0188831f $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_639 N_A_1417_294#_c_747_n N_A_1273_131#_c_1062_n 4.85805e-19 $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_640 N_A_1417_294#_c_748_n N_A_1273_131#_c_1062_n 0.00708115f $X=7.245 $Y=1.47
+ $X2=0 $Y2=0
cc_641 N_A_1417_294#_M1033_g N_A_1273_131#_c_1067_n 0.0180737f $X=7.235 $Y=2.495
+ $X2=0 $Y2=0
cc_642 N_A_1417_294#_c_743_n N_A_1273_131#_c_1067_n 0.00261875f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_643 N_A_1417_294#_c_746_n N_A_1273_131#_c_1067_n 0.0241092f $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_644 N_A_1417_294#_c_747_n N_A_1273_131#_c_1067_n 0.0010619f $X=7.25 $Y=1.635
+ $X2=0 $Y2=0
cc_645 N_A_1417_294#_M1033_g N_A_1273_131#_c_1068_n 0.00213524f $X=7.235
+ $Y=2.495 $X2=0 $Y2=0
cc_646 N_A_1417_294#_c_743_n N_A_1273_131#_c_1069_n 0.00205576f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_647 N_A_1417_294#_c_787_p N_A_1273_131#_c_1069_n 0.0121827f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_648 N_A_1417_294#_M1033_g N_A_1273_131#_c_1070_n 7.18596e-19 $X=7.235
+ $Y=2.495 $X2=0 $Y2=0
cc_649 N_A_1417_294#_c_743_n N_A_1273_131#_c_1063_n 0.0156786f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_650 N_A_1417_294#_c_749_n N_A_1273_131#_c_1063_n 0.0259649f $X=9.112 $Y=1.97
+ $X2=0 $Y2=0
cc_651 N_A_1417_294#_M1016_g N_A_1273_131#_c_1110_n 5.793e-19 $X=7.34 $Y=0.865
+ $X2=0 $Y2=0
cc_652 N_A_1417_294#_c_743_n N_A_1273_131#_c_1064_n 0.00989482f $X=8.73 $Y=1.215
+ $X2=0 $Y2=0
cc_653 N_A_1417_294#_c_749_n N_A_1273_131#_c_1064_n 0.00872479f $X=9.112 $Y=1.97
+ $X2=0 $Y2=0
cc_654 N_A_1417_294#_M1016_g N_A_859_347#_M1028_g 0.0392913f $X=7.34 $Y=0.865
+ $X2=0 $Y2=0
cc_655 N_A_1417_294#_c_744_n N_A_859_347#_M1028_g 6.51628e-19 $X=7.415 $Y=1.215
+ $X2=0 $Y2=0
cc_656 N_A_1417_294#_M1016_g N_A_859_347#_c_1171_n 0.00999433f $X=7.34 $Y=0.865
+ $X2=0 $Y2=0
cc_657 N_A_1417_294#_c_745_n N_A_859_347#_M1039_g 0.00125916f $X=8.815 $Y=0.865
+ $X2=0 $Y2=0
cc_658 N_A_1417_294#_c_749_n N_A_859_347#_M1039_g 0.00423916f $X=9.112 $Y=1.97
+ $X2=0 $Y2=0
cc_659 N_A_1417_294#_c_787_p N_A_859_347#_c_1177_n 0.0216168f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_660 N_A_1417_294#_c_749_n N_A_859_347#_c_1177_n 0.0309855f $X=9.112 $Y=1.97
+ $X2=0 $Y2=0
cc_661 N_A_1417_294#_c_787_p N_A_859_347#_c_1178_n 0.00612587f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_662 N_A_1417_294#_c_787_p N_A_859_347#_c_1181_n 0.00272068f $X=8.96 $Y=2.135
+ $X2=0 $Y2=0
cc_663 N_A_1417_294#_c_751_n N_A_1827_144#_c_1473_n 0.00131652f $X=8.96 $Y=2.815
+ $X2=0 $Y2=0
cc_664 N_A_1417_294#_M1033_g N_VPWR_c_1650_n 0.0101187f $X=7.235 $Y=2.495 $X2=0
+ $Y2=0
cc_665 N_A_1417_294#_c_751_n N_VPWR_c_1651_n 0.0260255f $X=8.96 $Y=2.815 $X2=0
+ $Y2=0
cc_666 N_A_1417_294#_c_751_n N_VPWR_c_1661_n 0.0311454f $X=8.96 $Y=2.815 $X2=0
+ $Y2=0
cc_667 N_A_1417_294#_M1033_g N_VPWR_c_1647_n 9.56319e-19 $X=7.235 $Y=2.495 $X2=0
+ $Y2=0
cc_668 N_A_1417_294#_c_751_n N_VPWR_c_1647_n 0.0257795f $X=8.96 $Y=2.815 $X2=0
+ $Y2=0
cc_669 N_A_1417_294#_c_743_n N_VGND_M1003_d 0.00610254f $X=8.73 $Y=1.215 $X2=0
+ $Y2=0
cc_670 N_A_1417_294#_M1016_g N_VGND_c_1947_n 9.39239e-19 $X=7.34 $Y=0.865 $X2=0
+ $Y2=0
cc_671 N_RESET_B_M1003_g N_A_1273_131#_c_1060_n 0.0214343f $X=7.7 $Y=0.865 $X2=0
+ $Y2=0
cc_672 N_RESET_B_c_844_n N_A_1273_131#_c_1062_n 0.0256788f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_673 N_RESET_B_M1030_g N_A_1273_131#_c_1067_n 0.0157308f $X=7.715 $Y=2.495
+ $X2=0 $Y2=0
cc_674 N_RESET_B_c_844_n N_A_1273_131#_c_1067_n 0.019501f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_RESET_B_c_852_n N_A_1273_131#_c_1067_n 0.00867656f $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_676 N_RESET_B_c_857_n N_A_1273_131#_c_1068_n 0.00513681f $X=7.625 $Y=3.15
+ $X2=0 $Y2=0
cc_677 N_RESET_B_c_844_n N_A_1273_131#_c_1068_n 0.00779596f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_RESET_B_M1030_g N_A_1273_131#_c_1069_n 0.00574918f $X=7.715 $Y=2.495
+ $X2=0 $Y2=0
cc_679 N_RESET_B_c_846_n N_A_1273_131#_c_1069_n 0.00484579f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_680 N_RESET_B_c_847_n N_A_1273_131#_c_1069_n 0.00310167f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_681 N_RESET_B_c_851_n N_A_1273_131#_c_1069_n 0.00489209f $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_682 N_RESET_B_c_852_n N_A_1273_131#_c_1069_n 0.0189906f $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_683 N_RESET_B_M1030_g N_A_1273_131#_c_1070_n 0.010638f $X=7.715 $Y=2.495
+ $X2=0 $Y2=0
cc_684 N_RESET_B_M1030_g N_A_1273_131#_c_1063_n 0.00477807f $X=7.715 $Y=2.495
+ $X2=0 $Y2=0
cc_685 N_RESET_B_c_846_n N_A_1273_131#_c_1063_n 0.0177544f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_686 N_RESET_B_c_847_n N_A_1273_131#_c_1063_n 0.00260992f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_687 N_RESET_B_c_851_n N_A_1273_131#_c_1063_n 4.82162e-19 $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_852_n N_A_1273_131#_c_1063_n 0.0209987f $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_844_n N_A_1273_131#_c_1110_n 0.00226953f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_846_n N_A_1273_131#_c_1064_n 0.00927046f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_691 N_RESET_B_c_847_n N_A_1273_131#_c_1064_n 0.00141062f $X=8.065 $Y=1.665
+ $X2=0 $Y2=0
cc_692 N_RESET_B_c_851_n N_A_1273_131#_c_1064_n 0.0220033f $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_852_n N_A_1273_131#_c_1064_n 0.00168155f $X=7.82 $Y=1.635
+ $X2=0 $Y2=0
cc_694 N_RESET_B_c_844_n N_A_859_347#_M1000_s 0.00243377f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_695 N_RESET_B_c_857_n N_A_859_347#_c_1183_n 0.0121828f $X=7.625 $Y=3.15 $X2=0
+ $Y2=0
cc_696 N_RESET_B_c_844_n N_A_859_347#_c_1183_n 0.00356343f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_844_n N_A_859_347#_c_1167_n 0.00278504f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_698 N_RESET_B_c_844_n N_A_859_347#_c_1185_n 0.00357158f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_699 N_RESET_B_c_857_n N_A_859_347#_c_1187_n 0.01074f $X=7.625 $Y=3.15 $X2=0
+ $Y2=0
cc_700 N_RESET_B_c_844_n N_A_859_347#_M1028_g 0.00367162f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_701 N_RESET_B_M1003_g N_A_859_347#_c_1171_n 0.00999433f $X=7.7 $Y=0.865 $X2=0
+ $Y2=0
cc_702 N_RESET_B_c_846_n N_A_859_347#_M1005_g 0.00138783f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_703 N_RESET_B_c_844_n N_A_859_347#_c_1196_n 0.0228322f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_704 N_RESET_B_c_844_n N_A_859_347#_c_1200_n 0.00742686f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_705 N_RESET_B_c_844_n N_A_859_347#_c_1189_n 0.0279904f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_844_n N_A_859_347#_c_1175_n 0.00384355f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_707 N_RESET_B_c_846_n N_A_859_347#_c_1177_n 0.0174731f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_708 N_RESET_B_c_846_n N_A_859_347#_c_1178_n 0.00494343f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_709 N_RESET_B_c_854_n N_A_859_347#_c_1179_n 0.0069234f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_710 N_RESET_B_c_846_n N_A_859_347#_c_1180_n 0.0048097f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_846_n N_A_859_347#_c_1181_n 0.0333185f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_844_n N_A_859_347#_c_1182_n 0.0143009f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_713 N_RESET_B_c_861_n N_A_2087_410#_M1013_g 0.0116941f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_714 N_RESET_B_M1009_g N_A_2087_410#_M1004_g 0.0291977f $X=11.25 $Y=0.58 $X2=0
+ $Y2=0
cc_715 N_RESET_B_c_843_n N_A_2087_410#_M1004_g 0.0115721f $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_716 N_RESET_B_c_846_n N_A_2087_410#_M1004_g 0.00407764f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_848_n N_A_2087_410#_M1004_g 6.26309e-19 $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_853_n N_A_2087_410#_M1004_g 0.0175496f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_854_n N_A_2087_410#_M1004_g 0.00284048f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_861_n N_A_2087_410#_c_1372_n 0.0153227f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_721 N_RESET_B_c_846_n N_A_2087_410#_c_1372_n 0.00166773f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_861_n N_A_2087_410#_c_1373_n 0.013977f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_723 N_RESET_B_M1009_g N_A_2087_410#_c_1368_n 7.40512e-19 $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_724 N_RESET_B_c_843_n N_A_2087_410#_c_1376_n 8.51156e-19 $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_725 N_RESET_B_c_846_n N_A_2087_410#_c_1376_n 0.00135183f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_726 N_RESET_B_c_861_n N_A_2087_410#_c_1377_n 0.0115721f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_727 N_RESET_B_c_861_n N_A_2087_410#_c_1378_n 0.00254182f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_728 N_RESET_B_M1009_g N_A_1827_144#_c_1458_n 0.0238259f $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_843_n N_A_1827_144#_c_1459_n 0.0238259f $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_730 N_RESET_B_c_854_n N_A_1827_144#_c_1459_n 0.00218879f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_843_n N_A_1827_144#_c_1460_n 0.0243914f $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_732 N_RESET_B_c_854_n N_A_1827_144#_c_1460_n 4.39803e-19 $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_861_n N_A_1827_144#_M1022_g 0.0193886f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_848_n N_A_1827_144#_c_1463_n 3.16322e-19 $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_846_n N_A_1827_144#_c_1464_n 0.00193276f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_846_n N_A_1827_144#_c_1474_n 0.0335295f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_846_n N_A_1827_144#_c_1475_n 0.0208335f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_738 N_RESET_B_M1009_g N_A_1827_144#_c_1465_n 0.0143997f $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_846_n N_A_1827_144#_c_1465_n 0.0102645f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_848_n N_A_1827_144#_c_1465_n 0.00174298f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_853_n N_A_1827_144#_c_1465_n 0.00126891f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_854_n N_A_1827_144#_c_1465_n 0.0296916f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_843_n N_A_1827_144#_c_1476_n 0.0105998f $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_861_n N_A_1827_144#_c_1476_n 0.00225328f $X=11.292 $Y=2.435
+ $X2=0 $Y2=0
cc_745 N_RESET_B_c_846_n N_A_1827_144#_c_1476_n 0.00297115f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_848_n N_A_1827_144#_c_1476_n 0.00466048f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_853_n N_A_1827_144#_c_1476_n 8.68178e-19 $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_854_n N_A_1827_144#_c_1476_n 0.0158387f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_749 N_RESET_B_M1009_g N_A_1827_144#_c_1466_n 0.00109112f $X=11.25 $Y=0.58
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_843_n N_A_1827_144#_c_1466_n 0.00231391f $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_848_n N_A_1827_144#_c_1466_n 0.00755838f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_853_n N_A_1827_144#_c_1466_n 3.9684e-19 $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_854_n N_A_1827_144#_c_1466_n 0.0432263f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_853_n N_A_1827_144#_c_1467_n 0.0238259f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_755 N_RESET_B_c_843_n N_A_1827_144#_c_1478_n 0.00258184f $X=11.292 $Y=2.285
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_846_n N_A_1827_144#_c_1478_n 0.00615148f $X=11.135 $Y=1.665
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_848_n N_A_1827_144#_c_1478_n 0.00137624f $X=11.28 $Y=1.665
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_854_n N_A_1827_144#_c_1478_n 0.00644897f $X=11.16 $Y=1.375
+ $X2=0 $Y2=0
cc_759 N_RESET_B_c_844_n N_VPWR_M1000_d 0.00118222f $X=7.775 $Y=1.665 $X2=0
+ $Y2=0
cc_760 N_RESET_B_c_857_n N_VPWR_c_1649_n 0.0257138f $X=7.625 $Y=3.15 $X2=0 $Y2=0
cc_761 N_RESET_B_c_857_n N_VPWR_c_1650_n 0.0205158f $X=7.625 $Y=3.15 $X2=0 $Y2=0
cc_762 N_RESET_B_M1030_g N_VPWR_c_1650_n 0.0143104f $X=7.715 $Y=2.495 $X2=0
+ $Y2=0
cc_763 N_RESET_B_M1030_g N_VPWR_c_1651_n 0.013377f $X=7.715 $Y=2.495 $X2=0 $Y2=0
cc_764 N_RESET_B_c_846_n N_VPWR_c_1651_n 0.00498743f $X=11.135 $Y=1.665 $X2=0
+ $Y2=0
cc_765 N_RESET_B_c_861_n N_VPWR_c_1654_n 0.005209f $X=11.292 $Y=2.435 $X2=0
+ $Y2=0
cc_766 N_RESET_B_c_858_n N_VPWR_c_1658_n 0.0450827f $X=3.38 $Y=3.15 $X2=0 $Y2=0
cc_767 N_RESET_B_c_857_n N_VPWR_c_1659_n 0.0673855f $X=7.625 $Y=3.15 $X2=0 $Y2=0
cc_768 N_RESET_B_c_857_n N_VPWR_c_1660_n 0.00990254f $X=7.625 $Y=3.15 $X2=0
+ $Y2=0
cc_769 N_RESET_B_c_857_n N_VPWR_c_1647_n 0.147563f $X=7.625 $Y=3.15 $X2=0 $Y2=0
cc_770 N_RESET_B_c_858_n N_VPWR_c_1647_n 0.00706166f $X=3.38 $Y=3.15 $X2=0 $Y2=0
cc_771 N_RESET_B_c_861_n N_VPWR_c_1647_n 0.00984155f $X=11.292 $Y=2.435 $X2=0
+ $Y2=0
cc_772 N_RESET_B_M1002_g N_VPWR_c_1666_n 0.00848413f $X=3.29 $Y=2.64 $X2=0 $Y2=0
cc_773 N_RESET_B_c_861_n N_VPWR_c_1670_n 0.00529834f $X=11.292 $Y=2.435 $X2=0
+ $Y2=0
cc_774 N_RESET_B_M1002_g N_A_287_464#_c_1792_n 0.0191546f $X=3.29 $Y=2.64 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_840_n N_A_287_464#_c_1792_n 0.0106472f $X=3.552 $Y=1.843
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_857_n N_A_287_464#_c_1792_n 0.0118132f $X=7.625 $Y=3.15 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_844_n N_A_287_464#_c_1792_n 0.00529241f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_778 N_RESET_B_c_845_n N_A_287_464#_c_1792_n 0.00184111f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_850_n N_A_287_464#_c_1792_n 0.0169788f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_780 N_RESET_B_M1023_g N_A_287_464#_c_1788_n 0.0203401f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_844_n N_A_287_464#_c_1788_n 0.00588465f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_782 N_RESET_B_c_845_n N_A_287_464#_c_1788_n 0.00176911f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_849_n N_A_287_464#_c_1788_n 0.00561437f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_784 N_RESET_B_c_850_n N_A_287_464#_c_1788_n 0.0251017f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_785 N_RESET_B_M1023_g N_A_287_464#_c_1790_n 0.00331613f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_840_n N_A_287_464#_c_1790_n 0.00331199f $X=3.552 $Y=1.843
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_844_n N_A_287_464#_c_1790_n 0.0267649f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_845_n N_A_287_464#_c_1790_n 0.00260304f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_849_n N_A_287_464#_c_1790_n 0.0035604f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_850_n N_A_287_464#_c_1790_n 0.048278f $X=3.57 $Y=1.52 $X2=0
+ $Y2=0
cc_791 N_RESET_B_c_857_n N_A_287_464#_c_1794_n 0.00759611f $X=7.625 $Y=3.15
+ $X2=0 $Y2=0
cc_792 N_RESET_B_c_844_n N_A_287_464#_c_1794_n 0.00963991f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_857_n N_A_287_464#_c_1795_n 0.0133905f $X=7.625 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_RESET_B_c_844_n N_A_287_464#_c_1795_n 0.0113075f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_844_n N_A_287_464#_c_1791_n 0.0275289f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_844_n N_A_287_464#_c_1797_n 0.00416538f $X=7.775 $Y=1.665
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_857_n N_A_287_464#_c_1799_n 0.00508475f $X=7.625 $Y=3.15
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_857_n N_A_287_464#_c_1800_n 0.00130391f $X=7.625 $Y=3.15
+ $X2=0 $Y2=0
cc_799 N_RESET_B_M1023_g N_VGND_c_1934_n 0.0109311f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_800 N_RESET_B_M1003_g N_VGND_c_1936_n 0.00378302f $X=7.7 $Y=0.865 $X2=0 $Y2=0
cc_801 N_RESET_B_M1009_g N_VGND_c_1937_n 0.0154281f $X=11.25 $Y=0.58 $X2=0 $Y2=0
cc_802 N_RESET_B_M1023_g N_VGND_c_1939_n 0.00490893f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_803 N_RESET_B_M1009_g N_VGND_c_1945_n 0.00383152f $X=11.25 $Y=0.58 $X2=0
+ $Y2=0
cc_804 N_RESET_B_M1023_g N_VGND_c_1947_n 0.00463377f $X=3.445 $Y=0.615 $X2=0
+ $Y2=0
cc_805 N_RESET_B_M1003_g N_VGND_c_1947_n 9.39239e-19 $X=7.7 $Y=0.865 $X2=0 $Y2=0
cc_806 N_RESET_B_M1009_g N_VGND_c_1947_n 0.0075725f $X=11.25 $Y=0.58 $X2=0 $Y2=0
cc_807 N_RESET_B_M1023_g N_noxref_24_c_2059_n 0.00396489f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_808 N_RESET_B_M1023_g N_noxref_24_c_2063_n 0.00479113f $X=3.445 $Y=0.615
+ $X2=0 $Y2=0
cc_809 N_A_1273_131#_c_1068_n N_A_859_347#_c_1185_n 0.00206229f $X=6.85 $Y=2.08
+ $X2=0 $Y2=0
cc_810 N_A_1273_131#_c_1068_n N_A_859_347#_c_1187_n 0.00681999f $X=6.85 $Y=2.08
+ $X2=0 $Y2=0
cc_811 N_A_1273_131#_c_1061_n N_A_859_347#_M1028_g 0.00483456f $X=6.795 $Y=0.95
+ $X2=0 $Y2=0
cc_812 N_A_1273_131#_c_1062_n N_A_859_347#_M1028_g 0.00247346f $X=6.76 $Y=1.97
+ $X2=0 $Y2=0
cc_813 N_A_1273_131#_c_1110_n N_A_859_347#_M1028_g 0.00253902f $X=6.795 $Y=1.075
+ $X2=0 $Y2=0
cc_814 N_A_1273_131#_c_1060_n N_A_859_347#_c_1171_n 0.00550586f $X=8.35 $Y=1.47
+ $X2=0 $Y2=0
cc_815 N_A_1273_131#_c_1060_n N_A_859_347#_M1039_g 0.00812321f $X=8.35 $Y=1.47
+ $X2=0 $Y2=0
cc_816 N_A_1273_131#_c_1064_n N_A_859_347#_c_1177_n 3.47459e-19 $X=8.685
+ $Y=1.635 $X2=0 $Y2=0
cc_817 N_A_1273_131#_c_1064_n N_A_859_347#_c_1178_n 0.021333f $X=8.685 $Y=1.635
+ $X2=0 $Y2=0
cc_818 N_A_1273_131#_c_1069_n N_VPWR_M1038_s 0.00470227f $X=7.955 $Y=2.19 $X2=0
+ $Y2=0
cc_819 N_A_1273_131#_c_1067_n N_VPWR_c_1650_n 0.0180884f $X=7.785 $Y=2.08 $X2=0
+ $Y2=0
cc_820 N_A_1273_131#_c_1068_n N_VPWR_c_1650_n 0.0119109f $X=6.85 $Y=2.08 $X2=0
+ $Y2=0
cc_821 N_A_1273_131#_c_1070_n N_VPWR_c_1650_n 0.0201628f $X=7.94 $Y=2.525 $X2=0
+ $Y2=0
cc_822 N_A_1273_131#_M1038_g N_VPWR_c_1651_n 0.0171974f $X=8.685 $Y=2.46 $X2=0
+ $Y2=0
cc_823 N_A_1273_131#_c_1069_n N_VPWR_c_1651_n 0.0171063f $X=7.955 $Y=2.19 $X2=0
+ $Y2=0
cc_824 N_A_1273_131#_c_1070_n N_VPWR_c_1651_n 0.0329654f $X=7.94 $Y=2.525 $X2=0
+ $Y2=0
cc_825 N_A_1273_131#_c_1064_n N_VPWR_c_1651_n 0.00305782f $X=8.685 $Y=1.635
+ $X2=0 $Y2=0
cc_826 N_A_1273_131#_c_1068_n N_VPWR_c_1659_n 0.00712102f $X=6.85 $Y=2.08 $X2=0
+ $Y2=0
cc_827 N_A_1273_131#_c_1070_n N_VPWR_c_1660_n 0.00613361f $X=7.94 $Y=2.525 $X2=0
+ $Y2=0
cc_828 N_A_1273_131#_M1038_g N_VPWR_c_1661_n 0.00460063f $X=8.685 $Y=2.46 $X2=0
+ $Y2=0
cc_829 N_A_1273_131#_M1038_g N_VPWR_c_1647_n 0.00913687f $X=8.685 $Y=2.46 $X2=0
+ $Y2=0
cc_830 N_A_1273_131#_c_1068_n N_VPWR_c_1647_n 0.0112138f $X=6.85 $Y=2.08 $X2=0
+ $Y2=0
cc_831 N_A_1273_131#_c_1070_n N_VPWR_c_1647_n 0.0102216f $X=7.94 $Y=2.525 $X2=0
+ $Y2=0
cc_832 N_A_1273_131#_c_1062_n N_A_287_464#_c_1791_n 0.00522841f $X=6.76 $Y=1.97
+ $X2=0 $Y2=0
cc_833 N_A_1273_131#_c_1062_n N_A_287_464#_c_1797_n 0.00538011f $X=6.76 $Y=1.97
+ $X2=0 $Y2=0
cc_834 N_A_1273_131#_c_1068_n N_A_287_464#_c_1797_n 0.00911583f $X=6.85 $Y=2.08
+ $X2=0 $Y2=0
cc_835 N_A_1273_131#_c_1068_n N_A_287_464#_c_1800_n 0.00846126f $X=6.85 $Y=2.08
+ $X2=0 $Y2=0
cc_836 N_A_1273_131#_c_1060_n N_VGND_c_1936_n 3.02776e-19 $X=8.35 $Y=1.47 $X2=0
+ $Y2=0
cc_837 N_A_1273_131#_c_1060_n N_VGND_c_1947_n 7.46714e-19 $X=8.35 $Y=1.47 $X2=0
+ $Y2=0
cc_838 N_A_859_347#_M1005_g N_A_2087_410#_M1013_g 0.0390717f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_839 N_A_859_347#_M1005_g N_A_2087_410#_M1004_g 0.0128858f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_840 N_A_859_347#_c_1179_n N_A_2087_410#_M1004_g 9.75712e-19 $X=10.23 $Y=1.455
+ $X2=0 $Y2=0
cc_841 N_A_859_347#_c_1180_n N_A_2087_410#_M1004_g 0.019448f $X=10.23 $Y=1.455
+ $X2=0 $Y2=0
cc_842 N_A_859_347#_M1005_g N_A_2087_410#_c_1376_n 0.00173995f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_843 N_A_859_347#_M1005_g N_A_2087_410#_c_1377_n 0.0198316f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_844 N_A_859_347#_M1039_g N_A_1827_144#_c_1464_n 0.00202292f $X=9.06 $Y=1.04
+ $X2=0 $Y2=0
cc_845 N_A_859_347#_c_1179_n N_A_1827_144#_c_1464_n 0.0136692f $X=10.23 $Y=1.455
+ $X2=0 $Y2=0
cc_846 N_A_859_347#_c_1180_n N_A_1827_144#_c_1464_n 0.0010837f $X=10.23 $Y=1.455
+ $X2=0 $Y2=0
cc_847 N_A_859_347#_c_1181_n N_A_1827_144#_c_1464_n 0.00873933f $X=10.065
+ $Y=1.415 $X2=0 $Y2=0
cc_848 N_A_859_347#_M1005_g N_A_1827_144#_c_1473_n 0.0278361f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_849 N_A_859_347#_M1005_g N_A_1827_144#_c_1474_n 0.0132833f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_850 N_A_859_347#_c_1179_n N_A_1827_144#_c_1474_n 0.0203927f $X=10.23 $Y=1.455
+ $X2=0 $Y2=0
cc_851 N_A_859_347#_c_1180_n N_A_1827_144#_c_1474_n 0.00326631f $X=10.23
+ $Y=1.455 $X2=0 $Y2=0
cc_852 N_A_859_347#_M1005_g N_A_1827_144#_c_1475_n 0.00247333f $X=10.135 $Y=2.75
+ $X2=0 $Y2=0
cc_853 N_A_859_347#_c_1177_n N_A_1827_144#_c_1475_n 0.00400591f $X=9.21 $Y=1.455
+ $X2=0 $Y2=0
cc_854 N_A_859_347#_c_1181_n N_A_1827_144#_c_1475_n 0.0218019f $X=10.065
+ $Y=1.415 $X2=0 $Y2=0
cc_855 N_A_859_347#_c_1196_n N_VPWR_M1000_d 0.00570078f $X=4.94 $Y=1.915 $X2=0
+ $Y2=0
cc_856 N_A_859_347#_c_1189_n N_VPWR_M1000_d 0.00100198f $X=5.065 $Y=1.82 $X2=0
+ $Y2=0
cc_857 N_A_859_347#_c_1183_n N_VPWR_c_1649_n 0.00499467f $X=5.295 $Y=1.66 $X2=0
+ $Y2=0
cc_858 N_A_859_347#_M1005_g N_VPWR_c_1661_n 0.0053223f $X=10.135 $Y=2.75 $X2=0
+ $Y2=0
cc_859 N_A_859_347#_c_1183_n N_VPWR_c_1647_n 0.00112709f $X=5.295 $Y=1.66 $X2=0
+ $Y2=0
cc_860 N_A_859_347#_c_1187_n N_VPWR_c_1647_n 0.00113998f $X=6.355 $Y=2.21 $X2=0
+ $Y2=0
cc_861 N_A_859_347#_M1005_g N_VPWR_c_1647_n 0.0102046f $X=10.135 $Y=2.75 $X2=0
+ $Y2=0
cc_862 N_A_859_347#_M1005_g N_VPWR_c_1670_n 0.00146736f $X=10.135 $Y=2.75 $X2=0
+ $Y2=0
cc_863 N_A_859_347#_c_1202_n N_A_287_464#_c_1788_n 0.00347682f $X=4.66 $Y=0.91
+ $X2=0 $Y2=0
cc_864 N_A_859_347#_c_1196_n N_A_287_464#_c_1790_n 0.012299f $X=4.94 $Y=1.915
+ $X2=0 $Y2=0
cc_865 N_A_859_347#_M1000_s N_A_287_464#_c_1794_n 5.00038e-19 $X=4.295 $Y=1.735
+ $X2=0 $Y2=0
cc_866 N_A_859_347#_M1000_s N_A_287_464#_c_1795_n 0.00130197f $X=4.295 $Y=1.735
+ $X2=0 $Y2=0
cc_867 N_A_859_347#_c_1183_n N_A_287_464#_c_1795_n 0.0188514f $X=5.295 $Y=1.66
+ $X2=0 $Y2=0
cc_868 N_A_859_347#_c_1185_n N_A_287_464#_c_1795_n 0.00128226f $X=6.265 $Y=2.135
+ $X2=0 $Y2=0
cc_869 N_A_859_347#_c_1186_n N_A_287_464#_c_1795_n 0.00661191f $X=5.875 $Y=2.135
+ $X2=0 $Y2=0
cc_870 N_A_859_347#_c_1196_n N_A_287_464#_c_1795_n 0.0164054f $X=4.94 $Y=1.915
+ $X2=0 $Y2=0
cc_871 N_A_859_347#_c_1175_n N_A_287_464#_c_1795_n 0.00111175f $X=5.215 $Y=1.41
+ $X2=0 $Y2=0
cc_872 N_A_859_347#_c_1182_n N_A_287_464#_c_1795_n 9.60145e-19 $X=5.8 $Y=1.435
+ $X2=0 $Y2=0
cc_873 N_A_859_347#_c_1166_n N_A_287_464#_c_1791_n 0.00866852f $X=5.8 $Y=1.21
+ $X2=0 $Y2=0
cc_874 N_A_859_347#_c_1182_n N_A_287_464#_c_1797_n 0.00866852f $X=5.8 $Y=1.435
+ $X2=0 $Y2=0
cc_875 N_A_859_347#_c_1183_n N_A_287_464#_c_1798_n 4.13018e-19 $X=5.295 $Y=1.66
+ $X2=0 $Y2=0
cc_876 N_A_859_347#_c_1185_n N_A_287_464#_c_1798_n 0.0149169f $X=6.265 $Y=2.135
+ $X2=0 $Y2=0
cc_877 N_A_859_347#_c_1183_n N_A_287_464#_c_1799_n 0.007817f $X=5.295 $Y=1.66
+ $X2=0 $Y2=0
cc_878 N_A_859_347#_M1000_s N_A_287_464#_c_1835_n 0.0115183f $X=4.295 $Y=1.735
+ $X2=0 $Y2=0
cc_879 N_A_859_347#_c_1196_n N_A_287_464#_c_1835_n 0.0364689f $X=4.94 $Y=1.915
+ $X2=0 $Y2=0
cc_880 N_A_859_347#_c_1185_n N_A_287_464#_c_1800_n 0.00838881f $X=6.265 $Y=2.135
+ $X2=0 $Y2=0
cc_881 N_A_859_347#_c_1187_n N_A_287_464#_c_1800_n 0.00308399f $X=6.355 $Y=2.21
+ $X2=0 $Y2=0
cc_882 N_A_859_347#_c_1200_n N_VGND_M1007_d 0.00507268f $X=4.94 $Y=0.91 $X2=0
+ $Y2=0
cc_883 N_A_859_347#_c_1176_n N_VGND_M1007_d 0.00125792f $X=5.12 $Y=1.22 $X2=0
+ $Y2=0
cc_884 N_A_859_347#_c_1199_n N_VGND_c_1934_n 0.0185922f $X=4.49 $Y=0.56 $X2=0
+ $Y2=0
cc_885 N_A_859_347#_c_1165_n N_VGND_c_1935_n 0.00169675f $X=5.27 $Y=1.21 $X2=0
+ $Y2=0
cc_886 N_A_859_347#_c_1169_n N_VGND_c_1935_n 0.00215328f $X=5.875 $Y=0.18 $X2=0
+ $Y2=0
cc_887 N_A_859_347#_c_1200_n N_VGND_c_1935_n 0.0239919f $X=4.94 $Y=0.91 $X2=0
+ $Y2=0
cc_888 N_A_859_347#_c_1182_n N_VGND_c_1935_n 3.5807e-19 $X=5.8 $Y=1.435 $X2=0
+ $Y2=0
cc_889 N_A_859_347#_c_1171_n N_VGND_c_1936_n 0.0251635f $X=8.985 $Y=0.18 $X2=0
+ $Y2=0
cc_890 N_A_859_347#_c_1199_n N_VGND_c_1942_n 0.0111284f $X=4.49 $Y=0.56 $X2=0
+ $Y2=0
cc_891 N_A_859_347#_c_1165_n N_VGND_c_1943_n 0.00461464f $X=5.27 $Y=1.21 $X2=0
+ $Y2=0
cc_892 N_A_859_347#_c_1169_n N_VGND_c_1943_n 0.0551781f $X=5.875 $Y=0.18 $X2=0
+ $Y2=0
cc_893 N_A_859_347#_c_1171_n N_VGND_c_1944_n 0.0228934f $X=8.985 $Y=0.18 $X2=0
+ $Y2=0
cc_894 N_A_859_347#_c_1165_n N_VGND_c_1947_n 0.0068352f $X=5.27 $Y=1.21 $X2=0
+ $Y2=0
cc_895 N_A_859_347#_c_1168_n N_VGND_c_1947_n 0.0239744f $X=6.895 $Y=0.18 $X2=0
+ $Y2=0
cc_896 N_A_859_347#_c_1169_n N_VGND_c_1947_n 0.00600144f $X=5.875 $Y=0.18 $X2=0
+ $Y2=0
cc_897 N_A_859_347#_c_1171_n N_VGND_c_1947_n 0.0479544f $X=8.985 $Y=0.18 $X2=0
+ $Y2=0
cc_898 N_A_859_347#_c_1174_n N_VGND_c_1947_n 0.00370846f $X=6.97 $Y=0.18 $X2=0
+ $Y2=0
cc_899 N_A_859_347#_c_1199_n N_VGND_c_1947_n 0.0118586f $X=4.49 $Y=0.56 $X2=0
+ $Y2=0
cc_900 N_A_859_347#_c_1200_n N_VGND_c_1947_n 0.010218f $X=4.94 $Y=0.91 $X2=0
+ $Y2=0
cc_901 N_A_2087_410#_c_1368_n N_A_1827_144#_c_1458_n 0.0105238f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_902 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1458_n 0.00492805f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_903 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1459_n 0.00675601f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_904 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1460_n 0.00165643f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_905 N_A_2087_410#_c_1373_n N_A_1827_144#_M1022_g 0.0133292f $X=11.545 $Y=2.75
+ $X2=0 $Y2=0
cc_906 N_A_2087_410#_c_1374_n N_A_1827_144#_M1022_g 0.0143046f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_907 N_A_2087_410#_c_1369_n N_A_1827_144#_M1022_g 0.00618531f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_908 N_A_2087_410#_c_1378_n N_A_1827_144#_M1022_g 0.00282772f $X=11.545
+ $Y=2.375 $X2=0 $Y2=0
cc_909 N_A_2087_410#_c_1374_n N_A_1827_144#_c_1470_n 0.00361662f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_910 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1470_n 0.0143738f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_911 N_A_2087_410#_c_1368_n N_A_1827_144#_c_1461_n 0.00530055f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_912 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1461_n 0.0145814f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_913 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1471_n 5.1349e-19 $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_914 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1462_n 7.30697e-19 $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_915 N_A_2087_410#_M1004_g N_A_1827_144#_c_1464_n 0.00519097f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_916 N_A_2087_410#_M1013_g N_A_1827_144#_c_1473_n 0.00188712f $X=10.545
+ $Y=2.75 $X2=0 $Y2=0
cc_917 N_A_2087_410#_M1004_g N_A_1827_144#_c_1473_n 7.38644e-19 $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_918 N_A_2087_410#_c_1376_n N_A_1827_144#_c_1473_n 0.0164475f $X=10.6 $Y=2.215
+ $X2=0 $Y2=0
cc_919 N_A_2087_410#_c_1377_n N_A_1827_144#_c_1473_n 9.05214e-19 $X=10.6
+ $Y=2.215 $X2=0 $Y2=0
cc_920 N_A_2087_410#_M1004_g N_A_1827_144#_c_1474_n 0.0120601f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_921 N_A_2087_410#_c_1372_n N_A_1827_144#_c_1474_n 0.00538841f $X=11.38
+ $Y=2.375 $X2=0 $Y2=0
cc_922 N_A_2087_410#_c_1376_n N_A_1827_144#_c_1474_n 0.017528f $X=10.6 $Y=2.215
+ $X2=0 $Y2=0
cc_923 N_A_2087_410#_c_1377_n N_A_1827_144#_c_1474_n 0.00124679f $X=10.6
+ $Y=2.215 $X2=0 $Y2=0
cc_924 N_A_2087_410#_M1004_g N_A_1827_144#_c_1465_n 0.0156553f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_925 N_A_2087_410#_c_1368_n N_A_1827_144#_c_1465_n 0.0151071f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_926 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1465_n 0.0135536f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_927 N_A_2087_410#_c_1372_n N_A_1827_144#_c_1476_n 0.024548f $X=11.38 $Y=2.375
+ $X2=0 $Y2=0
cc_928 N_A_2087_410#_c_1374_n N_A_1827_144#_c_1476_n 0.0143017f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_929 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1476_n 0.0135702f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_930 N_A_2087_410#_c_1378_n N_A_1827_144#_c_1476_n 0.0286194f $X=11.545
+ $Y=2.375 $X2=0 $Y2=0
cc_931 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1466_n 0.0689819f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_932 N_A_2087_410#_c_1368_n N_A_1827_144#_c_1467_n 0.0010568f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_933 N_A_2087_410#_c_1369_n N_A_1827_144#_c_1467_n 6.697e-19 $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_934 N_A_2087_410#_M1004_g N_A_1827_144#_c_1478_n 0.00514664f $X=10.69 $Y=0.58
+ $X2=0 $Y2=0
cc_935 N_A_2087_410#_c_1372_n N_A_1827_144#_c_1478_n 0.0132541f $X=11.38
+ $Y=2.375 $X2=0 $Y2=0
cc_936 N_A_2087_410#_c_1376_n N_A_1827_144#_c_1478_n 0.00515102f $X=10.6
+ $Y=2.215 $X2=0 $Y2=0
cc_937 N_A_2087_410#_c_1369_n N_A_2492_424#_c_1604_n 0.00119502f $X=12.15
+ $Y=2.29 $X2=0 $Y2=0
cc_938 N_A_2087_410#_c_1368_n N_A_2492_424#_c_1606_n 0.0191493f $X=12.065
+ $Y=0.575 $X2=0 $Y2=0
cc_939 N_A_2087_410#_c_1369_n N_A_2492_424#_c_1606_n 0.108701f $X=12.15 $Y=2.29
+ $X2=0 $Y2=0
cc_940 N_A_2087_410#_c_1374_n N_A_2492_424#_c_1611_n 0.013247f $X=12.065
+ $Y=2.375 $X2=0 $Y2=0
cc_941 N_A_2087_410#_c_1373_n N_VPWR_c_1652_n 0.0139233f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_942 N_A_2087_410#_c_1374_n N_VPWR_c_1652_n 0.026786f $X=12.065 $Y=2.375 $X2=0
+ $Y2=0
cc_943 N_A_2087_410#_c_1373_n N_VPWR_c_1654_n 0.0144776f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_944 N_A_2087_410#_M1013_g N_VPWR_c_1661_n 0.00461464f $X=10.545 $Y=2.75 $X2=0
+ $Y2=0
cc_945 N_A_2087_410#_M1013_g N_VPWR_c_1647_n 0.00908269f $X=10.545 $Y=2.75 $X2=0
+ $Y2=0
cc_946 N_A_2087_410#_c_1373_n N_VPWR_c_1647_n 0.0118404f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_947 N_A_2087_410#_M1013_g N_VPWR_c_1670_n 0.0176304f $X=10.545 $Y=2.75 $X2=0
+ $Y2=0
cc_948 N_A_2087_410#_c_1372_n N_VPWR_c_1670_n 0.0381798f $X=11.38 $Y=2.375 $X2=0
+ $Y2=0
cc_949 N_A_2087_410#_c_1373_n N_VPWR_c_1670_n 0.0132486f $X=11.545 $Y=2.75 $X2=0
+ $Y2=0
cc_950 N_A_2087_410#_c_1376_n N_VPWR_c_1670_n 0.00412564f $X=10.6 $Y=2.215 $X2=0
+ $Y2=0
cc_951 N_A_2087_410#_c_1377_n N_VPWR_c_1670_n 4.89906e-19 $X=10.6 $Y=2.215 $X2=0
+ $Y2=0
cc_952 N_A_2087_410#_M1004_g N_VGND_c_1937_n 0.0155907f $X=10.69 $Y=0.58 $X2=0
+ $Y2=0
cc_953 N_A_2087_410#_c_1368_n N_VGND_c_1937_n 0.00776169f $X=12.065 $Y=0.575
+ $X2=0 $Y2=0
cc_954 N_A_2087_410#_M1004_g N_VGND_c_1944_n 0.00352388f $X=10.69 $Y=0.58 $X2=0
+ $Y2=0
cc_955 N_A_2087_410#_c_1368_n N_VGND_c_1945_n 0.015221f $X=12.065 $Y=0.575 $X2=0
+ $Y2=0
cc_956 N_A_2087_410#_M1004_g N_VGND_c_1947_n 0.0069736f $X=10.69 $Y=0.58 $X2=0
+ $Y2=0
cc_957 N_A_2087_410#_c_1368_n N_VGND_c_1947_n 0.0182599f $X=12.065 $Y=0.575
+ $X2=0 $Y2=0
cc_958 N_A_1827_144#_c_1470_n N_A_2492_424#_M1014_g 0.0149035f $X=12.74 $Y=1.97
+ $X2=0 $Y2=0
cc_959 N_A_1827_144#_c_1462_n N_A_2492_424#_M1017_g 0.0139661f $X=12.845
+ $Y=0.995 $X2=0 $Y2=0
cc_960 N_A_1827_144#_c_1459_n N_A_2492_424#_c_1604_n 0.00295561f $X=11.73
+ $Y=1.405 $X2=0 $Y2=0
cc_961 N_A_1827_144#_c_1460_n N_A_2492_424#_c_1604_n 0.00131811f $X=11.755
+ $Y=1.895 $X2=0 $Y2=0
cc_962 N_A_1827_144#_c_1470_n N_A_2492_424#_c_1604_n 0.0301073f $X=12.74 $Y=1.97
+ $X2=0 $Y2=0
cc_963 N_A_1827_144#_c_1461_n N_A_2492_424#_c_1604_n 0.030045f $X=12.77 $Y=1.07
+ $X2=0 $Y2=0
cc_964 N_A_1827_144#_c_1461_n N_A_2492_424#_c_1606_n 0.0201885f $X=12.77 $Y=1.07
+ $X2=0 $Y2=0
cc_965 N_A_1827_144#_c_1462_n N_A_2492_424#_c_1606_n 0.012287f $X=12.845
+ $Y=0.995 $X2=0 $Y2=0
cc_966 N_A_1827_144#_M1022_g N_A_2492_424#_c_1611_n 0.00543931f $X=11.77 $Y=2.75
+ $X2=0 $Y2=0
cc_967 N_A_1827_144#_c_1470_n N_A_2492_424#_c_1611_n 0.0173743f $X=12.74 $Y=1.97
+ $X2=0 $Y2=0
cc_968 N_A_1827_144#_c_1471_n N_A_2492_424#_c_1611_n 0.0180942f $X=12.83
+ $Y=2.045 $X2=0 $Y2=0
cc_969 N_A_1827_144#_M1022_g N_VPWR_c_1652_n 0.00394849f $X=11.77 $Y=2.75 $X2=0
+ $Y2=0
cc_970 N_A_1827_144#_c_1470_n N_VPWR_c_1652_n 6.69985e-19 $X=12.74 $Y=1.97 $X2=0
+ $Y2=0
cc_971 N_A_1827_144#_c_1471_n N_VPWR_c_1652_n 0.00345749f $X=12.83 $Y=2.045
+ $X2=0 $Y2=0
cc_972 N_A_1827_144#_c_1470_n N_VPWR_c_1653_n 0.0107666f $X=12.74 $Y=1.97 $X2=0
+ $Y2=0
cc_973 N_A_1827_144#_M1022_g N_VPWR_c_1654_n 0.005209f $X=11.77 $Y=2.75 $X2=0
+ $Y2=0
cc_974 N_A_1827_144#_c_1473_n N_VPWR_c_1661_n 0.0145789f $X=9.845 $Y=2.135 $X2=0
+ $Y2=0
cc_975 N_A_1827_144#_c_1471_n N_VPWR_c_1662_n 0.00492575f $X=12.83 $Y=2.045
+ $X2=0 $Y2=0
cc_976 N_A_1827_144#_M1022_g N_VPWR_c_1647_n 0.00986837f $X=11.77 $Y=2.75 $X2=0
+ $Y2=0
cc_977 N_A_1827_144#_c_1471_n N_VPWR_c_1647_n 0.00897008f $X=12.83 $Y=2.045
+ $X2=0 $Y2=0
cc_978 N_A_1827_144#_c_1473_n N_VPWR_c_1647_n 0.0120225f $X=9.845 $Y=2.135 $X2=0
+ $Y2=0
cc_979 N_A_1827_144#_c_1473_n N_VPWR_c_1670_n 0.0100615f $X=9.845 $Y=2.135 $X2=0
+ $Y2=0
cc_980 N_A_1827_144#_c_1461_n Q 2.35526e-19 $X=12.77 $Y=1.07 $X2=0 $Y2=0
cc_981 N_A_1827_144#_c_1458_n N_VGND_c_1937_n 0.0017037f $X=11.64 $Y=0.9 $X2=0
+ $Y2=0
cc_982 N_A_1827_144#_c_1464_n N_VGND_c_1937_n 0.00833692f $X=10.305 $Y=0.695
+ $X2=0 $Y2=0
cc_983 N_A_1827_144#_c_1465_n N_VGND_c_1937_n 0.0305939f $X=11.565 $Y=0.955
+ $X2=0 $Y2=0
cc_984 N_A_1827_144#_c_1462_n N_VGND_c_1938_n 0.00901588f $X=12.845 $Y=0.995
+ $X2=0 $Y2=0
cc_985 N_A_1827_144#_c_1464_n N_VGND_c_1944_n 0.0235417f $X=10.305 $Y=0.695
+ $X2=0 $Y2=0
cc_986 N_A_1827_144#_c_1458_n N_VGND_c_1945_n 0.00435333f $X=11.64 $Y=0.9 $X2=0
+ $Y2=0
cc_987 N_A_1827_144#_c_1462_n N_VGND_c_1945_n 0.00434272f $X=12.845 $Y=0.995
+ $X2=0 $Y2=0
cc_988 N_A_1827_144#_c_1458_n N_VGND_c_1947_n 0.00824743f $X=11.64 $Y=0.9 $X2=0
+ $Y2=0
cc_989 N_A_1827_144#_c_1462_n N_VGND_c_1947_n 0.00826607f $X=12.845 $Y=0.995
+ $X2=0 $Y2=0
cc_990 N_A_1827_144#_c_1464_n N_VGND_c_1947_n 0.0330971f $X=10.305 $Y=0.695
+ $X2=0 $Y2=0
cc_991 N_A_1827_144#_c_1464_n A_2073_74# 0.00353391f $X=10.305 $Y=0.695
+ $X2=-0.19 $Y2=-0.245
cc_992 N_A_2492_424#_c_1611_n N_VPWR_c_1652_n 0.0237276f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_993 N_A_2492_424#_M1014_g N_VPWR_c_1653_n 0.00432096f $X=13.41 $Y=2.4 $X2=0
+ $Y2=0
cc_994 N_A_2492_424#_c_1604_n N_VPWR_c_1653_n 0.0151403f $X=13.32 $Y=1.52 $X2=0
+ $Y2=0
cc_995 N_A_2492_424#_c_1611_n N_VPWR_c_1653_n 0.0550307f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_996 N_A_2492_424#_c_1611_n N_VPWR_c_1662_n 0.0155898f $X=12.605 $Y=2.265
+ $X2=0 $Y2=0
cc_997 N_A_2492_424#_M1014_g N_VPWR_c_1663_n 0.00526565f $X=13.41 $Y=2.4 $X2=0
+ $Y2=0
cc_998 N_A_2492_424#_M1014_g N_VPWR_c_1647_n 0.010048f $X=13.41 $Y=2.4 $X2=0
+ $Y2=0
cc_999 N_A_2492_424#_c_1611_n N_VPWR_c_1647_n 0.012777f $X=12.605 $Y=2.265 $X2=0
+ $Y2=0
cc_1000 N_A_2492_424#_M1014_g Q 0.0234271f $X=13.41 $Y=2.4 $X2=0 $Y2=0
cc_1001 N_A_2492_424#_M1017_g Q 0.0241875f $X=13.425 $Y=0.74 $X2=0 $Y2=0
cc_1002 N_A_2492_424#_c_1605_n Q 0.0172016f $X=13.41 $Y=1.52 $X2=0 $Y2=0
cc_1003 N_A_2492_424#_c_1607_n Q 0.00799574f $X=12.645 $Y=1.52 $X2=0 $Y2=0
cc_1004 N_A_2492_424#_M1017_g N_VGND_c_1938_n 0.0060503f $X=13.425 $Y=0.74 $X2=0
+ $Y2=0
cc_1005 N_A_2492_424#_c_1604_n N_VGND_c_1938_n 0.0137394f $X=13.32 $Y=1.52 $X2=0
+ $Y2=0
cc_1006 N_A_2492_424#_c_1606_n N_VGND_c_1938_n 0.0373449f $X=12.63 $Y=0.645
+ $X2=0 $Y2=0
cc_1007 N_A_2492_424#_c_1606_n N_VGND_c_1945_n 0.0156794f $X=12.63 $Y=0.645
+ $X2=0 $Y2=0
cc_1008 N_A_2492_424#_M1017_g N_VGND_c_1946_n 0.00434272f $X=13.425 $Y=0.74
+ $X2=0 $Y2=0
cc_1009 N_A_2492_424#_M1017_g N_VGND_c_1947_n 0.00825042f $X=13.425 $Y=0.74
+ $X2=0 $Y2=0
cc_1010 N_A_2492_424#_c_1606_n N_VGND_c_1947_n 0.0129217f $X=12.63 $Y=0.645
+ $X2=0 $Y2=0
cc_1011 N_VPWR_M1036_d N_A_287_464#_c_1792_n 0.00929472f $X=2.76 $Y=2.32 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1657_n N_A_287_464#_c_1792_n 0.0102758f $X=2.815 $Y=3.33 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1658_n N_A_287_464#_c_1792_n 0.0220533f $X=4.84 $Y=3.33 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1647_n N_A_287_464#_c_1792_n 0.0414045f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1666_n N_A_287_464#_c_1792_n 0.0246631f $X=2.98 $Y=3.055 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1658_n N_A_287_464#_c_1794_n 0.00688698f $X=4.84 $Y=3.33 $X2=0
+ $Y2=0
cc_1017 N_VPWR_c_1647_n N_A_287_464#_c_1794_n 0.0104321f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1018 N_VPWR_M1000_d N_A_287_464#_c_1795_n 0.00629868f $X=4.8 $Y=1.735 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1649_n N_A_287_464#_c_1795_n 0.0239372f $X=5.005 $Y=2.635 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1659_n N_A_287_464#_c_1799_n 0.00504459f $X=7.295 $Y=3.33 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1647_n N_A_287_464#_c_1799_n 0.00713738f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1648_n N_A_287_464#_c_1807_n 0.01064f $X=0.73 $Y=2.805 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1657_n N_A_287_464#_c_1807_n 0.0289591f $X=2.815 $Y=3.33 $X2=0
+ $Y2=0
cc_1024 N_VPWR_c_1647_n N_A_287_464#_c_1807_n 0.02868f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1025 N_VPWR_c_1653_n Q 0.0451069f $X=13.14 $Y=1.985 $X2=0 $Y2=0
cc_1026 N_VPWR_c_1663_n Q 0.0145639f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1027 N_VPWR_c_1647_n Q 0.0119984f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1028 N_A_287_464#_c_1792_n A_474_464# 0.00248235f $X=3.43 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_1029 N_A_287_464#_c_1788_n N_VGND_c_1934_n 0.027068f $X=3.905 $Y=1.072 $X2=0
+ $Y2=0
cc_1030 N_A_287_464#_c_1801_n N_noxref_24_c_2058_n 0.00596172f $X=2.72 $Y=0.68
+ $X2=0 $Y2=0
cc_1031 N_A_287_464#_M1020_d N_noxref_24_c_2059_n 0.00467414f $X=1.98 $Y=0.405
+ $X2=0 $Y2=0
cc_1032 N_A_287_464#_c_1801_n N_noxref_24_c_2059_n 0.0511317f $X=2.72 $Y=0.68
+ $X2=0 $Y2=0
cc_1033 N_A_287_464#_c_1788_n N_noxref_24_c_2059_n 0.0041995f $X=3.905 $Y=1.072
+ $X2=0 $Y2=0
cc_1034 N_A_287_464#_c_1788_n N_noxref_24_c_2063_n 0.0209527f $X=3.905 $Y=1.072
+ $X2=0 $Y2=0
cc_1035 N_A_287_464#_c_1801_n noxref_26 0.00135313f $X=2.72 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_1036 Q N_VGND_c_1938_n 0.0308485f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1037 Q N_VGND_c_1946_n 0.0145639f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1038 Q N_VGND_c_1947_n 0.0119984f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1039 N_VGND_c_1933_n N_noxref_24_c_2058_n 0.0236042f $X=0.78 $Y=0.65 $X2=0
+ $Y2=0
cc_1040 N_VGND_c_1934_n N_noxref_24_c_2059_n 0.0102804f $X=3.82 $Y=0.615 $X2=0
+ $Y2=0
cc_1041 N_VGND_c_1939_n N_noxref_24_c_2059_n 0.12396f $X=3.655 $Y=0 $X2=0 $Y2=0
cc_1042 N_VGND_c_1947_n N_noxref_24_c_2059_n 0.0715772f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1043 N_VGND_c_1933_n N_noxref_24_c_2060_n 0.0125438f $X=0.78 $Y=0.65 $X2=0
+ $Y2=0
cc_1044 N_VGND_c_1939_n N_noxref_24_c_2060_n 0.0231539f $X=3.655 $Y=0 $X2=0
+ $Y2=0
cc_1045 N_VGND_c_1947_n N_noxref_24_c_2060_n 0.0127354f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1046 N_VGND_c_1934_n N_noxref_24_c_2063_n 0.0195812f $X=3.82 $Y=0.615 $X2=0
+ $Y2=0
cc_1047 N_noxref_24_c_2059_n noxref_25 0.00366293f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1048 N_noxref_24_c_2059_n noxref_26 0.0013394f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245

* File: sky130_fd_sc_ms__o32a_2.pex.spice
* Created: Wed Sep  2 12:26:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O32A_2%A_83_264# 1 2 9 13 17 21 24 25 26 29 31 35 36
+ 39 41 44 46
c113 46 0 1.0069e-19 $X=4.02 $Y=0.88
c114 21 0 1.28418e-20 $X=1.1 $Y=0.74
r115 48 49 60.5154 $w=2.27e-07 $l=2.85e-07 $layer=POLY_cond $X=0.67 $Y=1.47
+ $X2=0.955 $Y2=1.47
r116 39 51 12.7401 $w=2.27e-07 $l=6e-08 $layer=POLY_cond $X=1.04 $Y=1.47 $X2=1.1
+ $Y2=1.47
r117 39 49 18.0485 $w=2.27e-07 $l=8.5e-08 $layer=POLY_cond $X=1.04 $Y=1.47
+ $X2=0.955 $Y2=1.47
r118 38 41 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.04 $Y=1.485
+ $X2=1.15 $Y2=1.485
r119 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.485 $X2=1.04 $Y2=1.485
r120 35 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=1.045
+ $X2=4.1 $Y2=0.88
r121 35 36 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.1 $Y=1.045
+ $X2=4.1 $Y2=1.95
r122 32 44 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=3.11 $Y=2.035
+ $X2=2.892 $Y2=2.035
r123 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=2.035
+ $X2=4.1 $Y2=1.95
r124 31 32 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.015 $Y=2.035
+ $X2=3.11 $Y2=2.035
r125 27 44 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.892 $Y=2.12
+ $X2=2.892 $Y2=2.035
r126 27 29 15.7633 $w=4.33e-07 $l=5.95e-07 $layer=LI1_cond $X=2.892 $Y=2.12
+ $X2=2.892 $Y2=2.715
r127 25 44 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.675 $Y=2.035
+ $X2=2.892 $Y2=2.035
r128 25 26 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.675 $Y=2.035
+ $X2=1.235 $Y2=2.035
r129 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=1.95
+ $X2=1.235 $Y2=2.035
r130 23 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=1.65
+ $X2=1.15 $Y2=1.485
r131 23 24 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.15 $Y=1.65 $X2=1.15
+ $Y2=1.95
r132 19 51 12.4931 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.1 $Y=1.32 $X2=1.1
+ $Y2=1.47
r133 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.1 $Y=1.32 $X2=1.1
+ $Y2=0.74
r134 15 49 8.29035 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=0.955 $Y=1.65
+ $X2=0.955 $Y2=1.47
r135 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.955 $Y=1.65
+ $X2=0.955 $Y2=2.4
r136 11 48 12.4931 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.67 $Y=1.32
+ $X2=0.67 $Y2=1.47
r137 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.67 $Y=1.32
+ $X2=0.67 $Y2=0.74
r138 7 48 35.0352 $w=2.27e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.47
+ $X2=0.67 $Y2=1.47
r139 7 9 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=0.505 $Y=1.47 $X2=0.505
+ $Y2=2.4
r140 2 44 400 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.84 $X2=2.9 $Y2=2.035
r141 2 29 400 $w=1.7e-07 $l=9.676e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.84 $X2=2.9 $Y2=2.715
r142 1 46 91 $w=1.7e-07 $l=9.97935e-07 $layer=licon1_NDIFF $count=2 $X=3.245
+ $Y=0.37 $X2=4.02 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%A1 3 6 8 11 12 14
c39 14 0 1.17819e-19 $X=1.58 $Y=1.725
r40 11 14 48.5591 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.725
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.35
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.515 $X2=1.58 $Y2=1.515
r43 8 12 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=1.605 $Y=1.665
+ $X2=1.605 $Y2=1.515
r44 6 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.67 $Y=0.74 $X2=1.67
+ $Y2=1.35
r45 3 14 164.683 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=1.655 $Y=2.34
+ $X2=1.655 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%A2 3 7 9 12 13
c37 3 0 1.02106e-19 $X=2.075 $Y=2.34
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.515
+ $X2=2.15 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.515
+ $X2=2.15 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.515 $X2=2.15 $Y2=1.515
r41 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.15 $Y=1.665
+ $X2=2.15 $Y2=1.515
r42 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.1 $Y=0.74 $X2=2.1
+ $Y2=1.35
r43 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.075 $Y=2.34
+ $X2=2.075 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%A3 3 7 9 12 13
c37 13 0 1.02106e-19 $X=2.69 $Y=1.515
c38 7 0 1.0069e-19 $X=2.67 $Y=0.74
c39 3 0 1.01332e-19 $X=2.615 $Y=2.34
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.515
+ $X2=2.69 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.515
+ $X2=2.69 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.515 $X2=2.69 $Y2=1.515
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.69 $Y=1.665
+ $X2=2.69 $Y2=1.515
r44 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.67 $Y=0.74 $X2=2.67
+ $Y2=1.35
r45 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.615 $Y=2.34
+ $X2=2.615 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%B2 3 7 9 12
c36 9 0 1.01332e-19 $X=3.6 $Y=1.665
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.515
+ $X2=3.26 $Y2=1.68
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.515
+ $X2=3.26 $Y2=1.35
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.515 $X2=3.26 $Y2=1.515
r40 9 13 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.26
+ $Y2=1.565
r41 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.185 $Y=2.34
+ $X2=3.185 $Y2=1.68
r42 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.17 $Y=0.74 $X2=3.17
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%B1 3 5 6 7 9 11 12 13 14 15 16 23
r36 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=1.385 $X2=4.52 $Y2=1.385
r37 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.405
+ $X2=4.52 $Y2=2.775
r38 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.035
+ $X2=4.52 $Y2=2.405
r39 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=1.665
+ $X2=4.52 $Y2=2.035
r40 13 24 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.52 $Y=1.665
+ $X2=4.52 $Y2=1.385
r41 12 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.52 $Y=1.295 $X2=4.52
+ $Y2=1.385
r42 10 23 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.31 $Y=1.385
+ $X2=4.52 $Y2=1.385
r43 10 11 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.31 $Y=1.385
+ $X2=4.235 $Y2=1.385
r44 7 11 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.22
+ $X2=4.235 $Y2=1.385
r45 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.235 $Y=1.22 $X2=4.235
+ $Y2=0.74
r46 5 11 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.16 $Y=1.475
+ $X2=4.235 $Y2=1.385
r47 5 6 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.16 $Y=1.475
+ $X2=3.845 $Y2=1.475
r48 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.755 $Y=1.55
+ $X2=3.845 $Y2=1.475
r49 1 3 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=3.755 $Y=1.55
+ $X2=3.755 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%VPWR 1 2 3 10 12 18 22 25 26 27 29 42 43 49
r50 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r53 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r54 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r57 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 34 49 11.757 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=1.6 $Y=3.33 $X2=1.332
+ $Y2=3.33
r59 34 36 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=3.33 $X2=1.68
+ $Y2=3.33
r60 33 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 30 46 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r64 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 29 49 11.757 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.332 $Y2=3.33
r66 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 27 40 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r68 27 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 25 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.6 $Y2=3.33
r70 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.98 $Y2=3.33
r71 24 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=3.98 $Y2=3.33
r73 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=3.33
r74 20 22 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=2.375
r75 16 49 2.24534 $w=5.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.332 $Y=3.245
+ $X2=1.332 $Y2=3.33
r76 16 18 19.2267 $w=5.33e-07 $l=8.6e-07 $layer=LI1_cond $X=1.332 $Y=3.245
+ $X2=1.332 $Y2=2.385
r77 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r78 10 46 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r79 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r80 3 22 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.845
+ $Y=1.84 $X2=3.98 $Y2=2.375
r81 2 18 300 $w=1.7e-07 $l=7.10018e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.425 $Y2=2.385
r82 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r83 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%X 1 2 9 11 17 18 19 26 35
c39 17 0 1.17819e-19 $X=0.635 $Y=1.95
r40 24 26 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.715 $Y=2 $X2=0.715
+ $Y2=2.035
r41 18 19 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=2.405
+ $X2=0.715 $Y2=2.775
r42 17 24 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.715 $Y=1.975
+ $X2=0.715 $Y2=2
r43 17 35 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.715 $Y=1.975
+ $X2=0.715 $Y2=1.82
r44 17 18 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.715 $Y=2.06
+ $X2=0.715 $Y2=2.405
r45 17 26 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.715 $Y=2.06
+ $X2=0.715 $Y2=2.035
r46 9 13 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.885 $Y=1.045
+ $X2=0.62 $Y2=1.045
r47 9 11 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.885 $Y=0.96
+ $X2=0.885 $Y2=0.515
r48 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.62 $Y=1.13 $X2=0.62
+ $Y2=1.045
r49 7 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.62 $Y=1.13 $X2=0.62
+ $Y2=1.82
r50 2 17 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r51 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r52 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.745
+ $Y=0.37 $X2=0.885 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%VGND 1 2 3 10 13 16 20 24 26 28 29 31 32 33
+ 46 47
c60 16 0 1.28418e-20 $X=0.28 $Y=0.945
r61 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 44 47 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r64 43 46 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r65 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r67 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r68 38 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r69 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r70 35 50 5.62837 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.27
+ $Y2=0
r71 35 37 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=1.2
+ $Y2=0
r72 33 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r73 33 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r74 31 40 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.16
+ $Y2=0
r75 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.385
+ $Y2=0
r76 30 43 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.64
+ $Y2=0
r77 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.385
+ $Y2=0
r78 28 37 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.2
+ $Y2=0
r79 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.385
+ $Y2=0
r80 27 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=2.16
+ $Y2=0
r81 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.385
+ $Y2=0
r82 22 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0
r83 22 24 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0.675
r84 18 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=0.085
+ $X2=1.385 $Y2=0
r85 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.385 $Y=0.085
+ $X2=1.385 $Y2=0.515
r86 16 26 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=0.945
+ $X2=0.24 $Y2=0.79
r87 11 26 7.68649 $w=4.23e-07 $l=2.12e-07 $layer=LI1_cond $X=0.327 $Y=0.578
+ $X2=0.327 $Y2=0.79
r88 11 13 1.70833 $w=4.23e-07 $l=6.3e-08 $layer=LI1_cond $X=0.327 $Y=0.578
+ $X2=0.327 $Y2=0.515
r89 10 50 2.9601 $w=4.25e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.327 $Y=0.085
+ $X2=0.27 $Y2=0
r90 10 13 11.66 $w=4.23e-07 $l=4.3e-07 $layer=LI1_cond $X=0.327 $Y=0.085
+ $X2=0.327 $Y2=0.515
r91 3 24 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=2.175
+ $Y=0.37 $X2=2.385 $Y2=0.675
r92 2 20 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.175
+ $Y=0.37 $X2=1.385 $Y2=0.515
r93 1 16 182 $w=1.7e-07 $l=6.43428e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.945
r94 1 13 182 $w=1.7e-07 $l=3.85746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.455 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_2%A_349_74# 1 2 3 12 14 15 16 17 18 25
r46 19 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0.435
+ $X2=2.885 $Y2=0.435
r47 18 25 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.355 $Y=0.435
+ $X2=4.485 $Y2=0.435
r48 18 19 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=4.355 $Y=0.435
+ $X2=3.05 $Y2=0.435
r49 16 23 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0.52
+ $X2=2.885 $Y2=0.435
r50 16 17 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.885 $Y=0.52
+ $X2=2.885 $Y2=1.01
r51 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.72 $Y=1.095
+ $X2=2.885 $Y2=1.01
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.72 $Y=1.095
+ $X2=2.05 $Y2=1.095
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.885 $Y=1.01
+ $X2=2.05 $Y2=1.095
r54 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.885 $Y=1.01
+ $X2=1.885 $Y2=0.515
r55 3 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.37 $X2=4.45 $Y2=0.495
r56 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.37 $X2=2.885 $Y2=0.515
r57 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.745
+ $Y=0.37 $X2=1.885 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__o22ai_4.pxi.spice
* Created: Wed Sep  2 12:24:02 2020
* 
x_PM_SKY130_FD_SC_MS__O22AI_4%A1 N_A1_M1000_g N_A1_M1001_g N_A1_M1002_g
+ N_A1_M1015_g N_A1_M1027_g N_A1_M1003_g N_A1_M1012_g N_A1_M1030_g N_A1_c_132_n
+ N_A1_c_140_n N_A1_c_133_n N_A1_c_134_n A1 A1 N_A1_c_135_n N_A1_c_143_n
+ N_A1_c_144_n PM_SKY130_FD_SC_MS__O22AI_4%A1
x_PM_SKY130_FD_SC_MS__O22AI_4%A2 N_A2_M1004_g N_A2_c_255_n N_A2_M1008_g
+ N_A2_c_256_n N_A2_M1013_g N_A2_M1005_g N_A2_M1006_g N_A2_c_259_n N_A2_M1023_g
+ N_A2_c_260_n N_A2_M1009_g N_A2_c_262_n N_A2_M1031_g A2 A2 A2
+ PM_SKY130_FD_SC_MS__O22AI_4%A2
x_PM_SKY130_FD_SC_MS__O22AI_4%B1 N_B1_M1011_g N_B1_M1007_g N_B1_M1010_g
+ N_B1_M1019_g N_B1_M1018_g N_B1_M1025_g N_B1_M1026_g N_B1_M1029_g N_B1_c_352_n
+ N_B1_c_353_n N_B1_c_354_n N_B1_c_355_n B1 N_B1_c_356_n N_B1_c_357_n
+ N_B1_c_358_n PM_SKY130_FD_SC_MS__O22AI_4%B1
x_PM_SKY130_FD_SC_MS__O22AI_4%B2 N_B2_M1016_g N_B2_M1014_g N_B2_M1021_g
+ N_B2_M1017_g N_B2_M1024_g N_B2_M1020_g N_B2_M1022_g N_B2_M1028_g B2 B2
+ N_B2_c_480_n N_B2_c_475_n N_B2_c_482_n N_B2_c_502_n
+ PM_SKY130_FD_SC_MS__O22AI_4%B2
x_PM_SKY130_FD_SC_MS__O22AI_4%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1012_s
+ N_VPWR_M1010_s N_VPWR_M1026_s N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n
+ N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n VPWR
+ N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n
+ N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_557_n PM_SKY130_FD_SC_MS__O22AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O22AI_4%A_120_368# N_A_120_368#_M1001_d
+ N_A_120_368#_M1003_d N_A_120_368#_M1005_s N_A_120_368#_M1009_s
+ N_A_120_368#_c_654_n N_A_120_368#_c_663_n N_A_120_368#_c_667_n
+ N_A_120_368#_c_670_n N_A_120_368#_c_655_n N_A_120_368#_c_656_n
+ N_A_120_368#_c_657_n PM_SKY130_FD_SC_MS__O22AI_4%A_120_368#
x_PM_SKY130_FD_SC_MS__O22AI_4%Y N_Y_M1011_s N_Y_M1025_s N_Y_M1021_s N_Y_M1028_s
+ N_Y_M1004_d N_Y_M1006_d N_Y_M1014_s N_Y_M1020_s N_Y_c_713_n N_Y_c_719_n
+ N_Y_c_734_n N_Y_c_720_n N_Y_c_767_n N_Y_c_709_n N_Y_c_705_n N_Y_c_706_n
+ N_Y_c_722_n N_Y_c_750_n N_Y_c_752_n N_Y_c_781_n N_Y_c_756_n N_Y_c_788_n
+ N_Y_c_757_n Y Y N_Y_c_707_n Y N_Y_c_708_n PM_SKY130_FD_SC_MS__O22AI_4%Y
x_PM_SKY130_FD_SC_MS__O22AI_4%A_880_368# N_A_880_368#_M1007_d
+ N_A_880_368#_M1018_d N_A_880_368#_M1017_d N_A_880_368#_M1022_d
+ N_A_880_368#_c_852_n N_A_880_368#_c_885_n N_A_880_368#_c_846_n
+ N_A_880_368#_c_847_n N_A_880_368#_c_888_n N_A_880_368#_c_848_n
+ N_A_880_368#_c_856_n N_A_880_368#_c_849_n N_A_880_368#_c_850_n
+ PM_SKY130_FD_SC_MS__O22AI_4%A_880_368#
x_PM_SKY130_FD_SC_MS__O22AI_4%A_27_74# N_A_27_74#_M1000_d N_A_27_74#_M1015_d
+ N_A_27_74#_M1008_d N_A_27_74#_M1023_d N_A_27_74#_M1030_d N_A_27_74#_M1019_d
+ N_A_27_74#_M1016_d N_A_27_74#_M1024_d N_A_27_74#_M1029_d N_A_27_74#_c_895_n
+ N_A_27_74#_c_896_n N_A_27_74#_c_897_n N_A_27_74#_c_898_n N_A_27_74#_c_919_n
+ N_A_27_74#_c_899_n N_A_27_74#_c_935_n N_A_27_74#_c_900_n N_A_27_74#_c_901_n
+ N_A_27_74#_c_902_n N_A_27_74#_c_925_n N_A_27_74#_c_903_n N_A_27_74#_c_904_n
+ N_A_27_74#_c_944_n N_A_27_74#_c_947_n N_A_27_74#_c_905_n N_A_27_74#_c_906_n
+ N_A_27_74#_c_907_n N_A_27_74#_c_908_n N_A_27_74#_c_909_n
+ PM_SKY130_FD_SC_MS__O22AI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O22AI_4%VGND N_VGND_M1000_s N_VGND_M1027_s N_VGND_M1013_s
+ N_VGND_M1031_s N_VGND_c_1021_n N_VGND_c_1022_n N_VGND_c_1023_n N_VGND_c_1024_n
+ VGND N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n N_VGND_c_1028_n
+ N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n N_VGND_c_1032_n
+ N_VGND_c_1033_n N_VGND_c_1034_n PM_SKY130_FD_SC_MS__O22AI_4%VGND
cc_1 VNB N_A1_M1000_g 0.0318055f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1001_g 7.57144e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_3 VNB N_A1_M1002_g 4.95692e-19 $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_4 VNB N_A1_M1015_g 0.0221345f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_5 VNB N_A1_M1027_g 0.023347f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_6 VNB N_A1_M1003_g 5.13588e-19 $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.4
cc_7 VNB N_A1_M1030_g 0.0256089f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_8 VNB N_A1_c_132_n 5.80078e-19 $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.485
cc_9 VNB N_A1_c_133_n 0.00755711f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_10 VNB N_A1_c_134_n 0.0233046f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_11 VNB N_A1_c_135_n 0.0788835f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.485
cc_12 VNB N_A2_M1004_g 0.00108117f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_13 VNB N_A2_c_255_n 0.0171512f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.65
cc_14 VNB N_A2_c_256_n 0.0173859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1005_g 0.00602065f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.32
cc_16 VNB N_A2_M1006_g 0.00579868f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.32
cc_17 VNB N_A2_c_259_n 0.0172061f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_18 VNB N_A2_c_260_n 0.0937118f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.4
cc_19 VNB N_A2_M1009_g 0.00585302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_262_n 0.0187428f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.4
cc_21 VNB A2 0.00911391f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_22 VNB N_B1_M1011_g 0.0213686f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_23 VNB N_B1_M1007_g 0.00156875f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_24 VNB N_B1_M1010_g 0.00154279f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_25 VNB N_B1_M1019_g 0.0209615f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_26 VNB N_B1_M1018_g 0.00160611f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_27 VNB N_B1_M1025_g 0.0206172f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.4
cc_28 VNB N_B1_M1026_g 0.00689395f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.4
cc_29 VNB N_B1_c_352_n 0.00305806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_c_353_n 0.0164724f $X=-0.19 $Y=-0.245 $X2=3.64 $Y2=1.805
cc_31 VNB N_B1_c_354_n 0.00320503f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.485
cc_32 VNB N_B1_c_355_n 0.0345219f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.805
cc_33 VNB N_B1_c_356_n 0.0596685f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.485
cc_34 VNB N_B1_c_357_n 0.0197466f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.485
cc_35 VNB N_B1_c_358_n 0.00417394f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.485
cc_36 VNB N_B2_M1016_g 0.0212007f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_37 VNB N_B2_M1021_g 0.0225267f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_38 VNB N_B2_M1024_g 0.0235253f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_39 VNB N_B2_M1028_g 0.02313f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_40 VNB N_B2_c_475_n 0.0729709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_557_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_705_n 0.00775967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_706_n 0.0327392f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_44 VNB N_Y_c_707_n 0.00340136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_708_n 0.00141707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_895_n 0.0265694f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_47 VNB N_A_27_74#_c_896_n 0.00324652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_897_n 0.0138252f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.485
cc_49 VNB N_A_27_74#_c_898_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.485
cc_50 VNB N_A_27_74#_c_899_n 0.00206561f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.485
cc_51 VNB N_A_27_74#_c_900_n 0.00253097f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_52 VNB N_A_27_74#_c_901_n 0.0104547f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_53 VNB N_A_27_74#_c_902_n 0.00211111f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.95
cc_54 VNB N_A_27_74#_c_903_n 0.00757463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_74#_c_904_n 0.00184947f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.485
cc_56 VNB N_A_27_74#_c_905_n 9.8643e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_74#_c_906_n 0.00281291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_74#_c_907_n 0.00219607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_74#_c_908_n 0.0155228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_74#_c_909_n 0.00288497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1021_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_62 VNB N_VGND_c_1022_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_63 VNB N_VGND_c_1023_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.4
cc_64 VNB N_VGND_c_1024_n 0.00851143f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.4
cc_65 VNB N_VGND_c_1025_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_66 VNB N_VGND_c_1026_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.485
cc_67 VNB N_VGND_c_1027_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=3.235 $Y2=1.805
cc_68 VNB N_VGND_c_1028_n 0.016883f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.805
cc_69 VNB N_VGND_c_1029_n 0.10275f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.485
cc_70 VNB N_VGND_c_1030_n 0.42396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1031_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.485
cc_72 VNB N_VGND_c_1032_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.485
cc_73 VNB N_VGND_c_1033_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_74 VNB N_VGND_c_1034_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.935
cc_75 VPB N_A1_M1001_g 0.028089f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_76 VPB N_A1_M1002_g 0.0223304f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_77 VPB N_A1_M1003_g 0.0228376f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.4
cc_78 VPB N_A1_M1012_g 0.0223804f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=2.4
cc_79 VPB N_A1_c_140_n 0.0082105f $X=-0.19 $Y=1.66 $X2=3.64 $Y2=1.805
cc_80 VPB N_A1_c_133_n 0.0028448f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_81 VPB N_A1_c_134_n 0.00545774f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_82 VPB N_A1_c_143_n 0.0119906f $X=-0.19 $Y=1.66 $X2=2.525 $Y2=1.935
cc_83 VPB N_A1_c_144_n 0.00422601f $X=-0.19 $Y=1.66 $X2=3.235 $Y2=1.935
cc_84 VPB N_A2_M1004_g 0.0222509f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_85 VPB N_A2_M1005_g 0.0219539f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.32
cc_86 VPB N_A2_M1006_g 0.0213135f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.32
cc_87 VPB N_A2_M1009_g 0.0215907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_B1_M1007_g 0.0239727f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_89 VPB N_B1_M1010_g 0.0224355f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_90 VPB N_B1_M1018_g 0.0228857f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_91 VPB N_B1_M1026_g 0.0247992f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=2.4
cc_92 VPB N_B2_M1014_g 0.0213323f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_93 VPB N_B2_M1017_g 0.0204338f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_94 VPB N_B2_M1020_g 0.0197603f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.4
cc_95 VPB N_B2_M1022_g 0.0209391f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=2.4
cc_96 VPB N_B2_c_480_n 0.00245085f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.95
cc_97 VPB N_B2_c_475_n 0.0128823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_B2_c_482_n 0.00267097f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.485
cc_99 VPB N_VPWR_c_558_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_559_n 0.0580564f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_101 VPB N_VPWR_c_560_n 0.0057767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_561_n 0.00969292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_562_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_563_n 0.0136226f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.485
cc_105 VPB N_VPWR_c_564_n 0.0384762f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.485
cc_106 VPB N_VPWR_c_565_n 0.0182909f $X=-0.19 $Y=1.66 $X2=3.64 $Y2=1.805
cc_107 VPB N_VPWR_c_566_n 0.0631261f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=1.485
cc_108 VPB N_VPWR_c_567_n 0.0196495f $X=-0.19 $Y=1.66 $X2=3.035 $Y2=1.95
cc_109 VPB N_VPWR_c_568_n 0.0588138f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.485
cc_110 VPB N_VPWR_c_569_n 0.0061274f $X=-0.19 $Y=1.66 $X2=2.525 $Y2=1.935
cc_111 VPB N_VPWR_c_570_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_571_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_557_n 0.080431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_120_368#_c_654_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_115 VPB N_A_120_368#_c_655_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.65
cc_116 VPB N_A_120_368#_c_656_n 0.00957532f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=1.68
cc_117 VPB N_A_120_368#_c_657_n 0.00224125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_Y_c_709_n 0.0105186f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=1.485
cc_119 VPB N_Y_c_706_n 0.0132219f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_120 VPB N_A_880_368#_c_846_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_121 VPB N_A_880_368#_c_847_n 0.00296278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_880_368#_c_848_n 0.0045905f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=1.68
cc_123 VPB N_A_880_368#_c_849_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_880_368#_c_850_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.485
cc_125 N_A1_M1003_g N_A2_M1004_g 0.0200355f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A1_c_143_n N_A2_M1004_g 0.0183186f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_127 N_A1_M1027_g N_A2_c_255_n 0.0293754f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A1_c_143_n N_A2_M1005_g 0.01331f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_129 N_A1_c_144_n N_A2_M1006_g 0.0216811f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_130 N_A1_c_132_n N_A2_c_260_n 0.00218607f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_131 N_A1_c_133_n N_A2_c_260_n 0.00178991f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A1_c_134_n N_A2_c_260_n 0.0179433f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A1_c_135_n N_A2_c_260_n 0.0303199f $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_134 N_A1_c_143_n N_A2_c_260_n 0.00329647f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_135 N_A1_c_144_n N_A2_c_260_n 0.0041296f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_136 N_A1_M1012_g N_A2_M1009_g 0.0497057f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A1_c_140_n N_A2_M1009_g 0.0154909f $X=3.64 $Y=1.805 $X2=0 $Y2=0
cc_138 N_A1_c_133_n N_A2_M1009_g 7.63802e-19 $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_c_144_n N_A2_M1009_g 0.0106637f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_140 N_A1_M1030_g N_A2_c_262_n 0.0274388f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A1_M1027_g A2 7.61463e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A1_M1030_g A2 5.59403e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_c_132_n A2 0.0101061f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_144 N_A1_c_133_n A2 0.00788709f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_135_n A2 9.98877e-19 $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_146 N_A1_c_143_n A2 0.10443f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_147 N_A1_M1030_g N_B1_M1011_g 0.0199157f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A1_M1012_g N_B1_M1007_g 0.0289604f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A1_c_133_n N_B1_M1007_g 9.75149e-19 $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A1_M1030_g N_B1_c_352_n 2.59363e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A1_c_133_n N_B1_c_352_n 0.0134326f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A1_c_134_n N_B1_c_352_n 3.18267e-19 $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A1_c_133_n N_B1_c_356_n 0.00158937f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A1_c_134_n N_B1_c_356_n 0.0174817f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A1_M1001_g N_VPWR_c_559_n 0.00517389f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A1_M1001_g N_VPWR_c_560_n 5.10111e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A1_M1002_g N_VPWR_c_560_n 0.0111688f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A1_M1003_g N_VPWR_c_560_n 0.00334682f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A1_M1012_g N_VPWR_c_561_n 0.00345715f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A1_M1001_g N_VPWR_c_565_n 0.005209f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A1_M1002_g N_VPWR_c_565_n 0.00460063f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A1_M1003_g N_VPWR_c_566_n 0.00519767f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A1_M1012_g N_VPWR_c_566_n 0.00519794f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A1_M1001_g N_VPWR_c_557_n 0.00986025f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A1_M1002_g N_VPWR_c_557_n 0.00908554f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A1_M1003_g N_VPWR_c_557_n 0.00978524f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A1_M1012_g N_VPWR_c_557_n 0.0053431f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A1_c_143_n N_A_120_368#_M1003_d 0.00165831f $X=2.525 $Y=1.935 $X2=0
+ $Y2=0
cc_169 N_A1_c_144_n N_A_120_368#_M1005_s 0.001842f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_170 N_A1_c_140_n N_A_120_368#_M1009_s 0.00260026f $X=3.64 $Y=1.805 $X2=0
+ $Y2=0
cc_171 N_A1_M1001_g N_A_120_368#_c_654_n 0.0100782f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A1_M1002_g N_A_120_368#_c_654_n 2.69566e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_M1002_g N_A_120_368#_c_663_n 0.0146641f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A1_M1003_g N_A_120_368#_c_663_n 0.0132928f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A1_c_132_n N_A_120_368#_c_663_n 0.0258312f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_176 N_A1_c_135_n N_A_120_368#_c_663_n 0.00275393f $X=1.46 $Y=1.485 $X2=0
+ $Y2=0
cc_177 N_A1_M1003_g N_A_120_368#_c_667_n 8.8334e-19 $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A1_c_132_n N_A_120_368#_c_667_n 0.00242235f $X=1.38 $Y=1.485 $X2=0
+ $Y2=0
cc_179 N_A1_c_143_n N_A_120_368#_c_667_n 0.0149351f $X=2.525 $Y=1.935 $X2=0
+ $Y2=0
cc_180 N_A1_M1002_g N_A_120_368#_c_670_n 2.72638e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A1_M1003_g N_A_120_368#_c_670_n 0.00874072f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A1_M1003_g N_A_120_368#_c_655_n 0.00412402f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A1_M1012_g N_A_120_368#_c_656_n 0.00453342f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A1_M1001_g N_A_120_368#_c_657_n 0.00606807f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_M1002_g N_A_120_368#_c_657_n 0.00786471f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1003_g N_A_120_368#_c_657_n 0.00107422f $X=1.46 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_c_132_n N_A_120_368#_c_657_n 0.0293931f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_188 N_A1_c_135_n N_A_120_368#_c_657_n 0.00209661f $X=1.46 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A1_c_143_n N_Y_M1004_d 0.00218982f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_190 N_A1_c_144_n N_Y_M1006_d 0.00171048f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_191 N_A1_M1012_g N_Y_c_713_n 0.0150142f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A1_c_140_n N_Y_c_713_n 0.0109838f $X=3.64 $Y=1.805 $X2=0 $Y2=0
cc_193 N_A1_c_133_n N_Y_c_713_n 0.00822158f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A1_c_134_n N_Y_c_713_n 4.10665e-19 $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A1_c_143_n N_Y_c_713_n 0.00480209f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_196 N_A1_c_144_n N_Y_c_713_n 0.0385074f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_197 N_A1_M1012_g N_Y_c_719_n 0.00683809f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A1_M1012_g N_Y_c_720_n 0.00423453f $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A1_c_133_n N_Y_c_720_n 0.00349615f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A1_c_143_n N_Y_c_722_n 0.0182791f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_201 N_A1_M1012_g N_A_880_368#_c_849_n 7.61075e-19 $X=3.76 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A1_M1000_g N_A_27_74#_c_895_n 0.00980115f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A1_M1015_g N_A_27_74#_c_895_n 9.32548e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_M1000_g N_A_27_74#_c_896_n 0.0143535f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_M1015_g N_A_27_74#_c_896_n 0.01285f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A1_c_132_n N_A_27_74#_c_896_n 0.0432965f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_207 N_A1_c_135_n N_A_27_74#_c_896_n 0.00412669f $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A1_M1000_g N_A_27_74#_c_897_n 0.00247377f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A1_M1015_g N_A_27_74#_c_898_n 3.97481e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A1_M1027_g N_A_27_74#_c_898_n 0.00739853f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A1_M1027_g N_A_27_74#_c_919_n 0.0104473f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A1_c_132_n N_A_27_74#_c_919_n 0.0069724f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_213 N_A1_M1030_g N_A_27_74#_c_901_n 0.0131779f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_c_133_n N_A_27_74#_c_901_n 0.0146621f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A1_c_134_n N_A_27_74#_c_901_n 9.81106e-19 $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A1_M1030_g N_A_27_74#_c_902_n 0.00485335f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_M1030_g N_A_27_74#_c_925_n 0.00504463f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1027_g N_A_27_74#_c_904_n 0.00421845f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_c_132_n N_A_27_74#_c_904_n 0.0208089f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_220 N_A1_c_135_n N_A_27_74#_c_904_n 0.00232957f $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_221 N_A1_M1000_g N_VGND_c_1021_n 0.00555396f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1015_g N_VGND_c_1021_n 0.0098353f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1027_g N_VGND_c_1021_n 5.08869e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1027_g N_VGND_c_1022_n 0.00335277f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_M1030_g N_VGND_c_1024_n 0.00309798f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1000_g N_VGND_c_1025_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1015_g N_VGND_c_1026_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1027_g N_VGND_c_1026_n 0.00434272f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1030_g N_VGND_c_1029_n 0.00430908f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1000_g N_VGND_c_1030_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1015_g N_VGND_c_1030_n 0.0075754f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_M1027_g N_VGND_c_1030_n 0.00445549f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1030_g N_VGND_c_1030_n 0.00445992f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A2_M1004_g N_VPWR_c_566_n 0.00349951f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A2_M1005_g N_VPWR_c_566_n 0.00349978f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A2_M1006_g N_VPWR_c_566_n 0.00349978f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A2_M1009_g N_VPWR_c_566_n 0.00349978f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A2_M1004_g N_VPWR_c_557_n 0.00430096f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A2_M1005_g N_VPWR_c_557_n 0.0042906f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A2_M1006_g N_VPWR_c_557_n 0.00429518f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A2_M1009_g N_VPWR_c_557_n 0.00429629f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A2_M1004_g N_A_120_368#_c_667_n 0.00234398f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A2_M1004_g N_A_120_368#_c_670_n 0.00854839f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A2_M1005_g N_A_120_368#_c_670_n 8.63044e-19 $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A2_M1004_g N_A_120_368#_c_655_n 0.00138684f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A2_M1004_g N_A_120_368#_c_656_n 0.0172679f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A2_M1005_g N_A_120_368#_c_656_n 0.0140965f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A2_M1006_g N_A_120_368#_c_656_n 0.0135512f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A2_M1009_g N_A_120_368#_c_656_n 0.013547f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A2_M1005_g N_Y_c_713_n 0.0102852f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A2_M1006_g N_Y_c_713_n 0.00966931f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A2_M1009_g N_Y_c_713_n 0.0111323f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A2_M1005_g N_Y_c_722_n 0.00651862f $X=2.41 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A2_M1006_g N_Y_c_722_n 9.51697e-19 $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A2_c_255_n N_A_27_74#_c_898_n 7.18081e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_256 N_A2_c_255_n N_A_27_74#_c_919_n 0.0110188f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_257 A2 N_A_27_74#_c_919_n 0.0105847f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_258 N_A2_c_255_n N_A_27_74#_c_899_n 2.29136e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_259 N_A2_c_256_n N_A_27_74#_c_899_n 0.00703259f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_260 N_A2_c_259_n N_A_27_74#_c_899_n 7.13338e-19 $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_261 N_A2_c_256_n N_A_27_74#_c_935_n 0.00892313f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_262 N_A2_c_259_n N_A_27_74#_c_935_n 0.0100105f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_263 N_A2_c_260_n N_A_27_74#_c_935_n 0.00106692f $X=3.31 $Y=1.55 $X2=0 $Y2=0
cc_264 A2 N_A_27_74#_c_935_n 0.0454799f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_265 N_A2_c_259_n N_A_27_74#_c_900_n 2.49954e-19 $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_266 N_A2_c_262_n N_A_27_74#_c_900_n 2.68395e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_267 N_A2_c_262_n N_A_27_74#_c_901_n 0.0154305f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_268 N_A2_c_262_n N_A_27_74#_c_925_n 3.72705e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_269 N_A2_c_255_n N_A_27_74#_c_904_n 7.4692e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_270 N_A2_c_256_n N_A_27_74#_c_944_n 7.17169e-19 $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_271 N_A2_c_260_n N_A_27_74#_c_944_n 7.06072e-19 $X=3.31 $Y=1.55 $X2=0 $Y2=0
cc_272 A2 N_A_27_74#_c_944_n 0.0189543f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_273 N_A2_c_260_n N_A_27_74#_c_947_n 9.84341e-19 $X=3.31 $Y=1.55 $X2=0 $Y2=0
cc_274 A2 N_A_27_74#_c_947_n 0.0198393f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_275 N_A2_c_255_n N_VGND_c_1022_n 0.00771106f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_276 N_A2_c_256_n N_VGND_c_1022_n 4.39845e-19 $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A2_c_256_n N_VGND_c_1023_n 0.00335277f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A2_c_259_n N_VGND_c_1023_n 0.00775702f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_279 N_A2_c_262_n N_VGND_c_1023_n 4.2363e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_280 N_A2_c_262_n N_VGND_c_1024_n 0.00199261f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_281 N_A2_c_255_n N_VGND_c_1027_n 0.00383152f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_282 N_A2_c_256_n N_VGND_c_1027_n 0.00434272f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_283 N_A2_c_259_n N_VGND_c_1028_n 0.00383152f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A2_c_262_n N_VGND_c_1028_n 0.00461464f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_285 N_A2_c_255_n N_VGND_c_1030_n 0.00383967f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_286 N_A2_c_256_n N_VGND_c_1030_n 0.00445496f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_287 N_A2_c_259_n N_VGND_c_1030_n 0.00384354f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_288 N_A2_c_262_n N_VGND_c_1030_n 0.00463822f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_289 N_B1_M1025_g N_B2_M1016_g 0.0236783f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_290 N_B1_c_352_n N_B2_M1016_g 3.11251e-19 $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_291 N_B1_c_353_n N_B2_M1016_g 0.00788083f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_292 N_B1_c_358_n N_B2_M1016_g 0.00599736f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_293 N_B1_M1018_g N_B2_M1014_g 0.0266382f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_294 N_B1_c_353_n N_B2_M1021_g 0.0108858f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_295 N_B1_c_358_n N_B2_M1021_g 5.5004e-19 $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_296 N_B1_c_353_n N_B2_M1024_g 0.0112791f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_297 N_B1_c_353_n N_B2_M1028_g 0.0108342f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_298 N_B1_c_354_n N_B2_M1028_g 0.00185513f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_299 N_B1_c_355_n N_B2_M1028_g 0.0187736f $X=7.565 $Y=1.385 $X2=0 $Y2=0
cc_300 N_B1_c_357_n N_B2_M1028_g 0.0270173f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_301 N_B1_M1026_g N_B2_c_480_n 0.0013974f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_302 N_B1_c_354_n N_B2_c_480_n 0.0070832f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_303 N_B1_c_355_n N_B2_c_480_n 4.33934e-19 $X=7.565 $Y=1.385 $X2=0 $Y2=0
cc_304 N_B1_M1026_g N_B2_c_475_n 0.0361449f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_305 N_B1_c_353_n N_B2_c_475_n 0.0118333f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_306 N_B1_c_356_n N_B2_c_475_n 0.0236783f $X=5.225 $Y=1.465 $X2=0 $Y2=0
cc_307 N_B1_c_358_n N_B2_c_475_n 0.0106509f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_308 N_B1_c_353_n N_B2_c_502_n 0.0991186f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_309 N_B1_c_356_n N_B2_c_502_n 2.02701e-19 $X=5.225 $Y=1.465 $X2=0 $Y2=0
cc_310 N_B1_c_358_n N_B2_c_502_n 0.0154812f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_311 N_B1_M1007_g N_VPWR_c_561_n 0.00343717f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_312 N_B1_M1010_g N_VPWR_c_562_n 0.00315072f $X=4.76 $Y=2.4 $X2=0 $Y2=0
cc_313 N_B1_M1018_g N_VPWR_c_562_n 0.0089376f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_314 N_B1_M1026_g N_VPWR_c_564_n 0.00341401f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_315 N_B1_M1007_g N_VPWR_c_567_n 0.005209f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_316 N_B1_M1010_g N_VPWR_c_567_n 0.005209f $X=4.76 $Y=2.4 $X2=0 $Y2=0
cc_317 N_B1_M1018_g N_VPWR_c_568_n 0.00460063f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_318 N_B1_M1026_g N_VPWR_c_568_n 0.00517089f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_319 N_B1_M1007_g N_VPWR_c_557_n 0.00982576f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_320 N_B1_M1010_g N_VPWR_c_557_n 0.00982266f $X=4.76 $Y=2.4 $X2=0 $Y2=0
cc_321 N_B1_M1018_g N_VPWR_c_557_n 0.00909121f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_322 N_B1_M1026_g N_VPWR_c_557_n 0.00981313f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_323 N_B1_c_358_n N_Y_M1025_s 0.00148168f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_324 N_B1_c_353_n N_Y_M1021_s 0.00251484f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_325 N_B1_c_353_n N_Y_M1028_s 0.00199526f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_326 N_B1_c_354_n N_Y_M1028_s 6.17026e-19 $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_327 N_B1_M1007_g N_Y_c_713_n 0.00172597f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_328 N_B1_M1007_g N_Y_c_719_n 0.00532913f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_329 N_B1_M1007_g N_Y_c_734_n 0.0185532f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_330 N_B1_M1010_g N_Y_c_734_n 0.0119824f $X=4.76 $Y=2.4 $X2=0 $Y2=0
cc_331 N_B1_M1018_g N_Y_c_734_n 0.0122696f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_332 N_B1_c_352_n N_Y_c_734_n 0.0582548f $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_333 N_B1_c_353_n N_Y_c_734_n 0.00341175f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_334 N_B1_c_356_n N_Y_c_734_n 0.003941f $X=5.225 $Y=1.465 $X2=0 $Y2=0
cc_335 N_B1_c_358_n N_Y_c_734_n 0.0134413f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_336 N_B1_M1026_g N_Y_c_709_n 0.0196428f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_337 N_B1_c_354_n N_Y_c_709_n 0.0102433f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_338 N_B1_c_355_n N_Y_c_709_n 5.10201e-19 $X=7.565 $Y=1.385 $X2=0 $Y2=0
cc_339 N_B1_c_355_n N_Y_c_705_n 2.54483e-19 $X=7.565 $Y=1.385 $X2=0 $Y2=0
cc_340 N_B1_c_357_n N_Y_c_705_n 0.00967079f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_341 N_B1_M1026_g N_Y_c_706_n 0.0127994f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_342 N_B1_c_354_n N_Y_c_706_n 0.0350504f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_343 N_B1_c_355_n N_Y_c_706_n 0.00739878f $X=7.565 $Y=1.385 $X2=0 $Y2=0
cc_344 N_B1_c_357_n N_Y_c_706_n 0.00614976f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_345 N_B1_M1018_g N_Y_c_750_n 7.20807e-19 $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_346 N_B1_c_353_n N_Y_c_750_n 9.91556e-19 $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_347 N_B1_M1025_g N_Y_c_752_n 0.00725011f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_348 N_B1_c_352_n N_Y_c_752_n 0.00885985f $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_349 N_B1_c_353_n N_Y_c_752_n 0.09861f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_350 N_B1_c_358_n N_Y_c_752_n 0.0133434f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_351 N_B1_M1026_g N_Y_c_756_n 7.15369e-19 $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_352 N_B1_c_354_n N_Y_c_757_n 0.0163546f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_353 N_B1_c_355_n N_Y_c_757_n 4.69669e-19 $X=7.565 $Y=1.385 $X2=0 $Y2=0
cc_354 N_B1_c_357_n N_Y_c_757_n 0.00788319f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_355 N_B1_M1011_g N_Y_c_707_n 0.00203855f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_356 N_B1_M1019_g N_Y_c_707_n 0.0143968f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_357 N_B1_c_352_n N_Y_c_707_n 0.0593442f $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_358 N_B1_c_356_n N_Y_c_707_n 0.00656527f $X=5.225 $Y=1.465 $X2=0 $Y2=0
cc_359 N_B1_M1025_g N_Y_c_708_n 0.008409f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_360 N_B1_c_358_n N_Y_c_708_n 0.00235206f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_361 N_B1_M1010_g N_A_880_368#_c_852_n 0.012931f $X=4.76 $Y=2.4 $X2=0 $Y2=0
cc_362 N_B1_M1018_g N_A_880_368#_c_852_n 0.0142562f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_363 N_B1_M1018_g N_A_880_368#_c_847_n 0.00108516f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_364 N_B1_M1026_g N_A_880_368#_c_848_n 0.00361288f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_365 N_B1_M1026_g N_A_880_368#_c_856_n 0.00761611f $X=7.56 $Y=2.4 $X2=0 $Y2=0
cc_366 N_B1_M1007_g N_A_880_368#_c_849_n 0.0125891f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_367 N_B1_M1010_g N_A_880_368#_c_849_n 0.0109163f $X=4.76 $Y=2.4 $X2=0 $Y2=0
cc_368 N_B1_M1018_g N_A_880_368#_c_849_n 6.73157e-19 $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_369 N_B1_c_353_n N_A_27_74#_M1016_d 0.00176891f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_370 N_B1_c_353_n N_A_27_74#_M1024_d 0.00251484f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_371 N_B1_c_354_n N_A_27_74#_M1029_d 3.49062e-19 $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_372 N_B1_M1011_g N_A_27_74#_c_901_n 0.00376676f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_373 N_B1_M1011_g N_A_27_74#_c_902_n 0.00188298f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_374 N_B1_M1011_g N_A_27_74#_c_925_n 0.00469212f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_375 N_B1_M1019_g N_A_27_74#_c_925_n 7.81702e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_376 N_B1_M1011_g N_A_27_74#_c_903_n 0.0156461f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_377 N_B1_M1019_g N_A_27_74#_c_903_n 0.0132936f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_378 N_B1_M1025_g N_A_27_74#_c_903_n 0.0125475f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_379 N_B1_c_357_n N_A_27_74#_c_907_n 3.47155e-19 $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_380 N_B1_c_357_n N_A_27_74#_c_909_n 0.0118166f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_381 N_B1_M1011_g N_VGND_c_1029_n 0.00278257f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_382 N_B1_M1019_g N_VGND_c_1029_n 0.00278271f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_383 N_B1_M1025_g N_VGND_c_1029_n 0.00278271f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_384 N_B1_c_357_n N_VGND_c_1029_n 0.00278271f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_385 N_B1_M1011_g N_VGND_c_1030_n 0.00354187f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_386 N_B1_M1019_g N_VGND_c_1030_n 0.00354097f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_387 N_B1_M1025_g N_VGND_c_1030_n 0.00353625f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_388 N_B1_c_357_n N_VGND_c_1030_n 0.00358041f $X=7.565 $Y=1.22 $X2=0 $Y2=0
cc_389 N_B2_M1014_g N_VPWR_c_568_n 0.00333926f $X=5.71 $Y=2.4 $X2=0 $Y2=0
cc_390 N_B2_M1017_g N_VPWR_c_568_n 0.00333926f $X=6.16 $Y=2.4 $X2=0 $Y2=0
cc_391 N_B2_M1020_g N_VPWR_c_568_n 0.00333926f $X=6.61 $Y=2.4 $X2=0 $Y2=0
cc_392 N_B2_M1022_g N_VPWR_c_568_n 0.00333926f $X=7.07 $Y=2.4 $X2=0 $Y2=0
cc_393 N_B2_M1014_g N_VPWR_c_557_n 0.00423254f $X=5.71 $Y=2.4 $X2=0 $Y2=0
cc_394 N_B2_M1017_g N_VPWR_c_557_n 0.00422687f $X=6.16 $Y=2.4 $X2=0 $Y2=0
cc_395 N_B2_M1020_g N_VPWR_c_557_n 0.00422789f $X=6.61 $Y=2.4 $X2=0 $Y2=0
cc_396 N_B2_M1022_g N_VPWR_c_557_n 0.00423267f $X=7.07 $Y=2.4 $X2=0 $Y2=0
cc_397 N_B2_M1014_g N_Y_c_734_n 0.014983f $X=5.71 $Y=2.4 $X2=0 $Y2=0
cc_398 N_B2_M1017_g N_Y_c_767_n 0.0135066f $X=6.16 $Y=2.4 $X2=0 $Y2=0
cc_399 N_B2_M1020_g N_Y_c_767_n 0.012931f $X=6.61 $Y=2.4 $X2=0 $Y2=0
cc_400 N_B2_c_475_n N_Y_c_767_n 8.76993e-19 $X=7.085 $Y=1.515 $X2=0 $Y2=0
cc_401 N_B2_c_482_n N_Y_c_767_n 0.020799f $X=6.715 $Y=1.605 $X2=0 $Y2=0
cc_402 N_B2_c_502_n N_Y_c_767_n 0.0115474f $X=6.365 $Y=1.605 $X2=0 $Y2=0
cc_403 N_B2_M1022_g N_Y_c_709_n 0.0140141f $X=7.07 $Y=2.4 $X2=0 $Y2=0
cc_404 N_B2_c_480_n N_Y_c_709_n 0.0110877f $X=6.99 $Y=1.515 $X2=0 $Y2=0
cc_405 N_B2_M1014_g N_Y_c_750_n 0.0136375f $X=5.71 $Y=2.4 $X2=0 $Y2=0
cc_406 N_B2_M1017_g N_Y_c_750_n 0.013792f $X=6.16 $Y=2.4 $X2=0 $Y2=0
cc_407 N_B2_M1020_g N_Y_c_750_n 0.00104477f $X=6.61 $Y=2.4 $X2=0 $Y2=0
cc_408 N_B2_c_475_n N_Y_c_750_n 0.00233326f $X=7.085 $Y=1.515 $X2=0 $Y2=0
cc_409 N_B2_c_502_n N_Y_c_750_n 0.0188814f $X=6.365 $Y=1.605 $X2=0 $Y2=0
cc_410 N_B2_M1016_g N_Y_c_752_n 0.00841587f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_411 N_B2_M1021_g N_Y_c_752_n 0.0118672f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_412 N_B2_M1024_g N_Y_c_781_n 0.00427826f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_413 N_B2_M1028_g N_Y_c_781_n 2.63525e-19 $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_414 N_B2_M1017_g N_Y_c_756_n 5.73047e-19 $X=6.16 $Y=2.4 $X2=0 $Y2=0
cc_415 N_B2_M1020_g N_Y_c_756_n 0.0105882f $X=6.61 $Y=2.4 $X2=0 $Y2=0
cc_416 N_B2_M1022_g N_Y_c_756_n 0.00951555f $X=7.07 $Y=2.4 $X2=0 $Y2=0
cc_417 N_B2_c_475_n N_Y_c_756_n 6.16419e-19 $X=7.085 $Y=1.515 $X2=0 $Y2=0
cc_418 N_B2_c_482_n N_Y_c_756_n 0.0231433f $X=6.715 $Y=1.605 $X2=0 $Y2=0
cc_419 N_B2_M1024_g N_Y_c_788_n 0.00757292f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_420 N_B2_M1028_g N_Y_c_788_n 0.0121078f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_421 N_B2_M1016_g N_Y_c_708_n 5.9325e-19 $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_422 N_B2_M1014_g N_A_880_368#_c_846_n 0.0139924f $X=5.71 $Y=2.4 $X2=0 $Y2=0
cc_423 N_B2_M1017_g N_A_880_368#_c_846_n 0.0140221f $X=6.16 $Y=2.4 $X2=0 $Y2=0
cc_424 N_B2_M1020_g N_A_880_368#_c_848_n 0.0140846f $X=6.61 $Y=2.4 $X2=0 $Y2=0
cc_425 N_B2_M1022_g N_A_880_368#_c_848_n 0.0143433f $X=7.07 $Y=2.4 $X2=0 $Y2=0
cc_426 N_B2_M1016_g N_A_27_74#_c_903_n 0.0124925f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_427 N_B2_M1021_g N_A_27_74#_c_905_n 0.00528709f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_428 N_B2_M1024_g N_A_27_74#_c_905_n 3.43302e-19 $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B2_M1021_g N_A_27_74#_c_906_n 0.00644043f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_430 N_B2_M1024_g N_A_27_74#_c_906_n 0.0110646f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_431 N_B2_M1028_g N_A_27_74#_c_907_n 0.00557328f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_432 N_B2_M1028_g N_A_27_74#_c_909_n 0.00642625f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_433 N_B2_M1016_g N_VGND_c_1029_n 0.00278271f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_434 N_B2_M1021_g N_VGND_c_1029_n 0.00278271f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B2_M1024_g N_VGND_c_1029_n 0.00278271f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_436 N_B2_M1028_g N_VGND_c_1029_n 0.00278271f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_437 N_B2_M1016_g N_VGND_c_1030_n 0.00353526f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_438 N_B2_M1021_g N_VGND_c_1030_n 0.00354087f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_439 N_B2_M1024_g N_VGND_c_1030_n 0.00354745f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_440 N_B2_M1028_g N_VGND_c_1030_n 0.00354798f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_441 N_VPWR_c_560_n N_A_120_368#_c_654_n 0.022534f $X=1.185 $Y=2.485 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_565_n N_A_120_368#_c_654_n 0.0123179f $X=1.02 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_557_n N_A_120_368#_c_654_n 0.0101276f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_444 N_VPWR_M1002_s N_A_120_368#_c_663_n 0.00514066f $X=1.05 $Y=1.84 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_560_n N_A_120_368#_c_663_n 0.0189268f $X=1.185 $Y=2.485 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_560_n N_A_120_368#_c_655_n 0.0142735f $X=1.185 $Y=2.485 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_566_n N_A_120_368#_c_655_n 0.0145268f $X=3.87 $Y=3.33 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_557_n N_A_120_368#_c_655_n 0.0118929f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_561_n N_A_120_368#_c_656_n 0.0141475f $X=4.035 $Y=2.78 $X2=0
+ $Y2=0
cc_450 N_VPWR_c_566_n N_A_120_368#_c_656_n 0.0759519f $X=3.87 $Y=3.33 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_557_n N_A_120_368#_c_656_n 0.0631713f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_559_n N_A_120_368#_c_657_n 0.0389224f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_453 N_VPWR_M1012_s N_Y_c_713_n 0.00680331f $X=3.85 $Y=1.84 $X2=0 $Y2=0
cc_454 N_VPWR_c_561_n N_Y_c_713_n 0.0206672f $X=4.035 $Y=2.78 $X2=0 $Y2=0
cc_455 N_VPWR_c_557_n N_Y_c_713_n 0.00753174f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_456 N_VPWR_M1012_s N_Y_c_719_n 0.00758861f $X=3.85 $Y=1.84 $X2=0 $Y2=0
cc_457 N_VPWR_M1012_s N_Y_c_734_n 7.04873e-19 $X=3.85 $Y=1.84 $X2=0 $Y2=0
cc_458 N_VPWR_M1010_s N_Y_c_734_n 0.00329779f $X=4.85 $Y=1.84 $X2=0 $Y2=0
cc_459 N_VPWR_c_561_n N_Y_c_734_n 3.76314e-19 $X=4.035 $Y=2.78 $X2=0 $Y2=0
cc_460 N_VPWR_M1012_s N_Y_c_720_n 0.0101301f $X=3.85 $Y=1.84 $X2=0 $Y2=0
cc_461 N_VPWR_M1026_s N_Y_c_709_n 0.0110863f $X=7.65 $Y=1.84 $X2=0 $Y2=0
cc_462 N_VPWR_c_564_n N_Y_c_709_n 0.0246138f $X=7.835 $Y=2.455 $X2=0 $Y2=0
cc_463 N_VPWR_M1026_s N_Y_c_706_n 0.00181945f $X=7.65 $Y=1.84 $X2=0 $Y2=0
cc_464 N_VPWR_M1010_s N_A_880_368#_c_852_n 0.00322928f $X=4.85 $Y=1.84 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_562_n N_A_880_368#_c_852_n 0.014901f $X=4.985 $Y=2.755 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_568_n N_A_880_368#_c_846_n 0.0459191f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_557_n N_A_880_368#_c_846_n 0.0258001f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_562_n N_A_880_368#_c_847_n 0.0114567f $X=4.985 $Y=2.755 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_568_n N_A_880_368#_c_847_n 0.0179217f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_557_n N_A_880_368#_c_847_n 0.00971942f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_564_n N_A_880_368#_c_848_n 0.0119238f $X=7.835 $Y=2.455 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_568_n N_A_880_368#_c_848_n 0.0675378f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_557_n N_A_880_368#_c_848_n 0.0373646f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_561_n N_A_880_368#_c_849_n 0.0127976f $X=4.035 $Y=2.78 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_562_n N_A_880_368#_c_849_n 0.0155014f $X=4.985 $Y=2.755 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_567_n N_A_880_368#_c_849_n 0.0144623f $X=4.9 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_557_n N_A_880_368#_c_849_n 0.0118344f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_568_n N_A_880_368#_c_850_n 0.0121867f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_557_n N_A_880_368#_c_850_n 0.00660921f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_559_n N_A_27_74#_c_897_n 0.00886035f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_A_120_368#_c_656_n N_Y_M1004_d 0.00223287f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_482 N_A_120_368#_c_656_n N_Y_M1006_d 0.00169505f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_483 N_A_120_368#_M1005_s N_Y_c_713_n 0.00330209f $X=2.5 $Y=1.84 $X2=0 $Y2=0
cc_484 N_A_120_368#_M1009_s N_Y_c_713_n 0.00424f $X=3.4 $Y=1.84 $X2=0 $Y2=0
cc_485 N_A_120_368#_c_656_n N_Y_c_713_n 0.0721777f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_486 N_A_120_368#_c_656_n N_Y_c_722_n 0.018646f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_487 N_Y_c_734_n N_A_880_368#_M1007_d 0.00329375f $X=5.77 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_488 N_Y_c_734_n N_A_880_368#_M1018_d 0.00463012f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_489 N_Y_c_767_n N_A_880_368#_M1017_d 0.00327043f $X=6.67 $Y=2.035 $X2=0 $Y2=0
cc_490 N_Y_c_709_n N_A_880_368#_M1022_d 0.00926247f $X=7.9 $Y=2.035 $X2=0 $Y2=0
cc_491 N_Y_c_734_n N_A_880_368#_c_852_n 0.0336305f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_492 N_Y_c_734_n N_A_880_368#_c_885_n 0.0167599f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_493 N_Y_M1014_s N_A_880_368#_c_846_n 0.00165831f $X=5.8 $Y=1.84 $X2=0 $Y2=0
cc_494 N_Y_c_750_n N_A_880_368#_c_846_n 0.0159318f $X=5.935 $Y=2.015 $X2=0 $Y2=0
cc_495 N_Y_c_767_n N_A_880_368#_c_888_n 0.0126919f $X=6.67 $Y=2.035 $X2=0 $Y2=0
cc_496 N_Y_M1020_s N_A_880_368#_c_848_n 0.00176461f $X=6.7 $Y=1.84 $X2=0 $Y2=0
cc_497 N_Y_c_756_n N_A_880_368#_c_848_n 0.0159805f $X=6.835 $Y=2.115 $X2=0 $Y2=0
cc_498 N_Y_c_709_n N_A_880_368#_c_856_n 0.0181132f $X=7.9 $Y=2.035 $X2=0 $Y2=0
cc_499 N_Y_c_713_n N_A_880_368#_c_849_n 0.0116309f $X=3.98 $Y=2.405 $X2=0 $Y2=0
cc_500 N_Y_c_719_n N_A_880_368#_c_849_n 0.00833534f $X=4.065 $Y=2.32 $X2=0 $Y2=0
cc_501 N_Y_c_734_n N_A_880_368#_c_849_n 0.0171782f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_502 N_Y_c_707_n N_A_27_74#_M1019_d 5.0211e-19 $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_503 N_Y_c_708_n N_A_27_74#_M1019_d 0.00136745f $X=5.155 $Y=0.94 $X2=0 $Y2=0
cc_504 N_Y_c_752_n N_A_27_74#_M1016_d 0.00335829f $X=6.205 $Y=0.757 $X2=0 $Y2=0
cc_505 N_Y_c_788_n N_A_27_74#_M1024_d 0.00473528f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_506 N_Y_c_705_n N_A_27_74#_M1029_d 0.0115696f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_507 N_Y_c_706_n N_A_27_74#_M1029_d 0.00349433f $X=7.985 $Y=1.95 $X2=0 $Y2=0
cc_508 N_Y_c_707_n N_A_27_74#_c_901_n 0.01255f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_509 N_Y_M1011_s N_A_27_74#_c_903_n 0.00245681f $X=4.37 $Y=0.37 $X2=0 $Y2=0
cc_510 N_Y_M1025_s N_A_27_74#_c_903_n 0.00180456f $X=5.3 $Y=0.37 $X2=0 $Y2=0
cc_511 N_Y_c_707_n N_A_27_74#_c_903_n 0.0444771f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_512 N_Y_c_708_n N_A_27_74#_c_905_n 0.0444771f $X=5.155 $Y=0.94 $X2=0 $Y2=0
cc_513 N_Y_M1021_s N_A_27_74#_c_906_n 0.00251484f $X=6.16 $Y=0.37 $X2=0 $Y2=0
cc_514 N_Y_c_752_n N_A_27_74#_c_906_n 0.00265349f $X=6.205 $Y=0.757 $X2=0 $Y2=0
cc_515 N_Y_c_781_n N_A_27_74#_c_906_n 0.0185397f $X=6.535 $Y=0.757 $X2=0 $Y2=0
cc_516 N_Y_c_788_n N_A_27_74#_c_906_n 0.00247659f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_517 N_Y_c_788_n N_A_27_74#_c_907_n 0.0191051f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_518 N_Y_c_705_n N_A_27_74#_c_908_n 0.0254247f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_519 N_Y_M1028_s N_A_27_74#_c_909_n 0.00250419f $X=7.16 $Y=0.37 $X2=0 $Y2=0
cc_520 N_Y_c_705_n N_A_27_74#_c_909_n 0.00440728f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_521 N_Y_c_788_n N_A_27_74#_c_909_n 0.00247659f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_522 N_Y_c_757_n N_A_27_74#_c_909_n 0.0185397f $X=7.535 $Y=0.757 $X2=0 $Y2=0
cc_523 N_Y_c_705_n N_VGND_c_1029_n 4.05485e-19 $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_524 N_Y_c_705_n N_VGND_c_1030_n 0.00100481f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_525 N_A_27_74#_c_896_n N_VGND_M1000_s 0.00250873f $X=1.125 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_526 N_A_27_74#_c_919_n N_VGND_M1027_s 0.0114794f $X=2.055 $Y=0.925 $X2=0
+ $Y2=0
cc_527 N_A_27_74#_c_935_n N_VGND_M1013_s 0.00462121f $X=2.985 $Y=0.925 $X2=0
+ $Y2=0
cc_528 N_A_27_74#_c_901_n N_VGND_M1031_s 0.0109491f $X=3.905 $Y=0.925 $X2=0
+ $Y2=0
cc_529 N_A_27_74#_c_895_n N_VGND_c_1021_n 0.0180508f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_530 N_A_27_74#_c_896_n N_VGND_c_1021_n 0.0209867f $X=1.125 $Y=1.065 $X2=0
+ $Y2=0
cc_531 N_A_27_74#_c_898_n N_VGND_c_1021_n 0.017215f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_532 N_A_27_74#_c_898_n N_VGND_c_1022_n 0.0122975f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_533 N_A_27_74#_c_919_n N_VGND_c_1022_n 0.0205261f $X=2.055 $Y=0.925 $X2=0
+ $Y2=0
cc_534 N_A_27_74#_c_899_n N_VGND_c_1022_n 0.0121972f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_535 N_A_27_74#_c_899_n N_VGND_c_1023_n 0.0122975f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_536 N_A_27_74#_c_935_n N_VGND_c_1023_n 0.0205261f $X=2.985 $Y=0.925 $X2=0
+ $Y2=0
cc_537 N_A_27_74#_c_900_n N_VGND_c_1023_n 0.0121972f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_538 N_A_27_74#_c_900_n N_VGND_c_1024_n 0.00154841f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_539 N_A_27_74#_c_901_n N_VGND_c_1024_n 0.0211672f $X=3.905 $Y=0.925 $X2=0
+ $Y2=0
cc_540 N_A_27_74#_c_902_n N_VGND_c_1024_n 0.0184532f $X=4.07 $Y=0.58 $X2=0 $Y2=0
cc_541 N_A_27_74#_c_895_n N_VGND_c_1025_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_542 N_A_27_74#_c_898_n N_VGND_c_1026_n 0.0109942f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_543 N_A_27_74#_c_899_n N_VGND_c_1027_n 0.0109704f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_544 N_A_27_74#_c_900_n N_VGND_c_1028_n 0.0110419f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_545 N_A_27_74#_c_902_n N_VGND_c_1029_n 0.023516f $X=4.07 $Y=0.58 $X2=0 $Y2=0
cc_546 N_A_27_74#_c_903_n N_VGND_c_1029_n 0.250323f $X=5.873 $Y=0.417 $X2=0
+ $Y2=0
cc_547 N_A_27_74#_c_895_n N_VGND_c_1030_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_548 N_A_27_74#_c_898_n N_VGND_c_1030_n 0.00904371f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_549 N_A_27_74#_c_919_n N_VGND_c_1030_n 0.0113663f $X=2.055 $Y=0.925 $X2=0
+ $Y2=0
cc_550 N_A_27_74#_c_899_n N_VGND_c_1030_n 0.00903439f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_551 N_A_27_74#_c_935_n N_VGND_c_1030_n 0.0113542f $X=2.985 $Y=0.925 $X2=0
+ $Y2=0
cc_552 N_A_27_74#_c_900_n N_VGND_c_1030_n 0.00915013f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_553 N_A_27_74#_c_901_n N_VGND_c_1030_n 0.010844f $X=3.905 $Y=0.925 $X2=0
+ $Y2=0
cc_554 N_A_27_74#_c_902_n N_VGND_c_1030_n 0.0126466f $X=4.07 $Y=0.58 $X2=0 $Y2=0
cc_555 N_A_27_74#_c_903_n N_VGND_c_1030_n 0.139412f $X=5.873 $Y=0.417 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o21ba_2.spice
* Created: Wed Sep  2 12:22:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21ba_2.pex.spice"
.subckt sky130_fd_sc_ms__o21ba_2  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_B1_N_M1006_g N_A_27_74#_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.0964632 AS=0.15125 PD=0.90814 PS=1.65 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_VGND_M1006_d N_A_177_48#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.129787 AS=0.1036 PD=1.22186 PS=1.02 NRD=7.296 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_177_48#_M1007_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_487_74#_M1011_d N_A_27_74#_M1011_g N_A_177_48#_M1011_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_487_74#_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1797 AS=0.1036 PD=1.34 PS=1.02 NRD=30.456 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1008 N_A_487_74#_M1008_d N_A1_M1008_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.1797 PD=2.02 PS=1.34 NRD=0 NRS=30.456 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_B1_N_M1002_g N_A_27_74#_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1662 AS=0.2352 PD=1.27286 PS=2.24 NRD=33.49 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003 A=0.1512 P=2.04 MULT=1
MM1004 N_X_M1004_d N_A_177_48#_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2216 PD=1.39 PS=1.69714 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90000.6 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1004_d N_A_177_48#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.410491 PD=1.39 PS=1.9283 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1010 N_A_177_48#_M1010_d N_A_27_74#_M1010_g N_VPWR_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.366509 PD=1.27 PS=1.7217 NRD=0 NRS=16.7253 M=1 R=5.55556
+ SA=90002 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 A_585_368# N_A2_M1000_g N_A_177_48#_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_585_368# VPB PSHORT L=0.18 W=1 AD=0.27
+ AS=0.165 PD=2.54 PS=1.33 NRD=0 NRS=21.6503 M=1 R=5.55556 SA=90002.9 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o21ba_2.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a31o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.450000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.450000 5.865000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.115000 1.450000 7.075000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565000 1.470000 3.235000 1.800000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.138200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.550000 0.895000 1.720000 ;
        RECT 0.565000 1.720000 1.895000 1.890000 ;
        RECT 0.565000 1.890000 0.895000 2.980000 ;
        RECT 0.615000 0.350000 0.865000 0.830000 ;
        RECT 0.615000 0.830000 1.725000 1.000000 ;
        RECT 0.615000 1.000000 0.865000 1.550000 ;
        RECT 1.555000 0.330000 1.725000 0.830000 ;
        RECT 1.565000 1.890000 1.895000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.130000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 1.045000  0.085000 1.375000 0.660000 ;
      RECT 1.065000  1.220000 4.750000 1.280000 ;
      RECT 1.065000  1.280000 3.590000 1.300000 ;
      RECT 1.065000  1.300000 2.335000 1.550000 ;
      RECT 1.065000  2.060000 1.395000 3.245000 ;
      RECT 1.895000  1.130000 4.750000 1.220000 ;
      RECT 1.930000  0.085000 2.260000 0.960000 ;
      RECT 2.065000  1.820000 2.395000 3.245000 ;
      RECT 2.490000  0.350000 2.740000 1.130000 ;
      RECT 2.625000  1.970000 2.955000 2.810000 ;
      RECT 2.625000  2.810000 4.075000 2.980000 ;
      RECT 2.920000  0.085000 3.250000 0.960000 ;
      RECT 3.125000  1.970000 3.575000 2.640000 ;
      RECT 3.405000  1.300000 3.575000 1.970000 ;
      RECT 3.420000  0.350000 3.750000 1.110000 ;
      RECT 3.420000  1.110000 4.750000 1.130000 ;
      RECT 3.745000  1.950000 7.085000 2.120000 ;
      RECT 3.745000  2.120000 4.075000 2.810000 ;
      RECT 3.920000  0.255000 5.740000 0.425000 ;
      RECT 3.920000  0.425000 4.250000 0.940000 ;
      RECT 4.245000  2.290000 4.575000 3.245000 ;
      RECT 4.420000  0.595000 4.750000 1.110000 ;
      RECT 4.745000  2.120000 5.075000 2.980000 ;
      RECT 4.980000  0.595000 5.230000 1.110000 ;
      RECT 4.980000  1.110000 7.030000 1.280000 ;
      RECT 5.245000  2.290000 5.575000 3.245000 ;
      RECT 5.410000  0.425000 5.740000 0.940000 ;
      RECT 5.755000  2.120000 6.085000 2.980000 ;
      RECT 5.920000  0.350000 6.090000 1.110000 ;
      RECT 6.255000  2.290000 6.585000 3.245000 ;
      RECT 6.270000  0.085000 6.600000 0.940000 ;
      RECT 6.755000  2.120000 7.085000 2.980000 ;
      RECT 6.780000  0.350000 7.030000 1.110000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_ms__a31o_4
END LIBRARY

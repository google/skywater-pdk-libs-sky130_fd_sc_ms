* File: sky130_fd_sc_ms__o2bb2a_2.pxi.spice
* Created: Fri Aug 28 17:59:38 2020
* 
x_PM_SKY130_FD_SC_MS__O2BB2A_2%B1 N_B1_M1009_g N_B1_c_90_n N_B1_M1006_g B1
+ N_B1_c_91_n PM_SKY130_FD_SC_MS__O2BB2A_2%B1
x_PM_SKY130_FD_SC_MS__O2BB2A_2%B2 N_B2_M1011_g N_B2_M1010_g B2 N_B2_c_117_n
+ PM_SKY130_FD_SC_MS__O2BB2A_2%B2
x_PM_SKY130_FD_SC_MS__O2BB2A_2%A_270_48# N_A_270_48#_M1003_s N_A_270_48#_M1000_d
+ N_A_270_48#_M1005_g N_A_270_48#_M1004_g N_A_270_48#_c_155_n
+ N_A_270_48#_c_148_n N_A_270_48#_c_149_n N_A_270_48#_c_187_p
+ N_A_270_48#_c_164_p N_A_270_48#_c_150_n N_A_270_48#_c_151_n
+ N_A_270_48#_c_152_n N_A_270_48#_c_153_n PM_SKY130_FD_SC_MS__O2BB2A_2%A_270_48#
x_PM_SKY130_FD_SC_MS__O2BB2A_2%A2_N N_A2_N_M1000_g N_A2_N_c_220_n N_A2_N_M1003_g
+ N_A2_N_c_221_n A2_N N_A2_N_c_223_n N_A2_N_c_224_n
+ PM_SKY130_FD_SC_MS__O2BB2A_2%A2_N
x_PM_SKY130_FD_SC_MS__O2BB2A_2%A1_N N_A1_N_M1002_g N_A1_N_M1007_g A1_N
+ N_A1_N_c_270_n PM_SKY130_FD_SC_MS__O2BB2A_2%A1_N
x_PM_SKY130_FD_SC_MS__O2BB2A_2%A_204_392# N_A_204_392#_M1005_d
+ N_A_204_392#_M1011_d N_A_204_392#_M1008_g N_A_204_392#_M1001_g
+ N_A_204_392#_M1012_g N_A_204_392#_M1013_g N_A_204_392#_c_325_n
+ N_A_204_392#_c_326_n N_A_204_392#_c_336_n N_A_204_392#_c_314_n
+ N_A_204_392#_c_315_n N_A_204_392#_c_316_n N_A_204_392#_c_317_n
+ N_A_204_392#_c_318_n N_A_204_392#_c_319_n N_A_204_392#_c_320_n
+ N_A_204_392#_c_321_n N_A_204_392#_c_354_n N_A_204_392#_c_322_n
+ PM_SKY130_FD_SC_MS__O2BB2A_2%A_204_392#
x_PM_SKY130_FD_SC_MS__O2BB2A_2%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_M1002_d
+ N_VPWR_M1012_s N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n
+ N_VPWR_c_441_n N_VPWR_c_442_n VPWR N_VPWR_c_443_n N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_436_n
+ PM_SKY130_FD_SC_MS__O2BB2A_2%VPWR
x_PM_SKY130_FD_SC_MS__O2BB2A_2%X N_X_M1001_d N_X_M1008_d N_X_c_490_n N_X_c_491_n
+ X X X X N_X_c_492_n PM_SKY130_FD_SC_MS__O2BB2A_2%X
x_PM_SKY130_FD_SC_MS__O2BB2A_2%A_27_74# N_A_27_74#_M1009_s N_A_27_74#_M1010_d
+ N_A_27_74#_c_523_n N_A_27_74#_c_524_n N_A_27_74#_c_525_n N_A_27_74#_c_526_n
+ PM_SKY130_FD_SC_MS__O2BB2A_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O2BB2A_2%VGND N_VGND_M1009_d N_VGND_M1007_d N_VGND_M1013_s
+ N_VGND_c_549_n N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n VGND
+ N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n
+ N_VGND_c_558_n PM_SKY130_FD_SC_MS__O2BB2A_2%VGND
cc_1 VNB N_B1_M1009_g 0.0379819f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_c_90_n 0.0212389f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.78
cc_3 VNB N_B1_c_91_n 0.0104121f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_4 VNB N_B2_M1010_g 0.0287799f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_5 VNB B2 0.00404778f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_B2_c_117_n 0.0162717f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_7 VNB N_A_270_48#_M1005_g 0.0364177f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_270_48#_c_148_n 0.0149601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_270_48#_c_149_n 0.00375376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_270_48#_c_150_n 0.00589746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_270_48#_c_151_n 0.00166222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_270_48#_c_152_n 0.0249558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_270_48#_c_153_n 0.00298596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_N_c_220_n 0.0171957f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_15 VNB N_A2_N_c_221_n 0.0246559f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_16 VNB A2_N 0.00165787f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_17 VNB N_A2_N_c_223_n 0.0177121f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_18 VNB N_A2_N_c_224_n 0.0156143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_N_M1007_g 0.0363411f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_20 VNB A1_N 0.00156355f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A1_N_c_270_n 0.0176812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_204_392#_M1008_g 0.00139894f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_A_204_392#_M1001_g 0.0231615f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_24 VNB N_A_204_392#_M1012_g 0.0019185f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_25 VNB N_A_204_392#_M1013_g 0.0263481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_204_392#_c_314_n 0.00607937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_204_392#_c_315_n 0.0166771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_204_392#_c_316_n 0.00278702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_204_392#_c_317_n 0.00184446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_204_392#_c_318_n 0.00941197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_204_392#_c_319_n 0.00210357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_204_392#_c_320_n 0.00980048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_204_392#_c_321_n 3.33931e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_204_392#_c_322_n 0.0666522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_436_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_490_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_X_c_491_n 0.004293f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_38 VNB N_X_c_492_n 0.00113445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_523_n 0.0302831f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_40 VNB N_A_27_74#_c_524_n 0.0189843f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.615
cc_41 VNB N_A_27_74#_c_525_n 0.00975977f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_42 VNB N_A_27_74#_c_526_n 0.00252706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_549_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_44 VNB N_VGND_c_550_n 0.00671515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_551_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_552_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_553_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_554_n 0.0497142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_555_n 0.0203669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_556_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_557_n 0.00617641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_558_n 0.256918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_B1_c_90_n 0.014314f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.78
cc_54 VPB N_B1_M1006_g 0.0293218f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_55 VPB N_B1_c_91_n 0.00566928f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_56 VPB N_B2_M1011_g 0.0239342f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_57 VPB B2 0.00287247f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_58 VPB N_B2_c_117_n 0.0118872f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_59 VPB N_A_270_48#_M1004_g 0.025611f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_60 VPB N_A_270_48#_c_155_n 0.00335202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_270_48#_c_151_n 0.00138703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_270_48#_c_152_n 0.0167625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A2_N_M1000_g 0.0242753f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_64 VPB A2_N 0.00138199f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_65 VPB N_A2_N_c_223_n 0.0143466f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_66 VPB N_A1_N_M1002_g 0.0250189f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_67 VPB A1_N 0.00102491f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_68 VPB N_A1_N_c_270_n 0.0163612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_204_392#_M1008_g 0.0241218f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_70 VPB N_A_204_392#_M1012_g 0.0274055f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_71 VPB N_A_204_392#_c_325_n 0.00414593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_204_392#_c_326_n 0.00282719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_204_392#_c_321_n 0.00286015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_437_n 0.0121044f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_75 VPB N_VPWR_c_438_n 0.0504711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_439_n 0.015007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_440_n 0.015949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_441_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_442_n 0.0645527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_443_n 0.033334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_444_n 0.0263486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_445_n 0.020646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_446_n 0.00680245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_447_n 0.00862975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_436_n 0.0752498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB X 0.0042974f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_87 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_X_c_492_n 8.32691e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 N_B1_M1006_g N_B2_M1011_g 0.0686956f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_90 N_B1_M1009_g N_B2_M1010_g 0.0246174f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B1_c_90_n B2 7.67374e-19 $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_92 N_B1_c_91_n B2 0.0198037f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_93 N_B1_c_90_n N_B2_c_117_n 0.0194189f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_94 N_B1_c_91_n N_B2_c_117_n 4.07543e-19 $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_95 N_B1_c_90_n N_VPWR_c_438_n 0.00419322f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_96 N_B1_M1006_g N_VPWR_c_438_n 0.0258875f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_97 N_B1_c_91_n N_VPWR_c_438_n 0.027668f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_98 N_B1_M1006_g N_VPWR_c_443_n 0.00460063f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_99 N_B1_M1006_g N_VPWR_c_436_n 0.00908371f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_100 N_B1_M1009_g N_A_27_74#_c_523_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1009_g N_A_27_74#_c_524_n 0.0156808f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B1_c_90_n N_A_27_74#_c_524_n 0.00225916f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_103 N_B1_c_91_n N_A_27_74#_c_524_n 0.0148079f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_104 N_B1_c_90_n N_A_27_74#_c_525_n 0.00291196f $X=0.51 $Y=1.78 $X2=0 $Y2=0
cc_105 N_B1_c_91_n N_A_27_74#_c_525_n 0.0207147f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_106 N_B1_M1009_g N_VGND_c_549_n 0.0134383f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_107 N_B1_M1009_g N_VGND_c_553_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B1_M1009_g N_VGND_c_558_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B2_M1010_g N_A_270_48#_M1005_g 0.0253735f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_110 N_B2_M1011_g N_A_270_48#_M1004_g 0.0123342f $X=0.93 $Y=2.46 $X2=0 $Y2=0
cc_111 B2 N_A_270_48#_c_151_n 0.0268544f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_112 N_B2_c_117_n N_A_270_48#_c_151_n 2.64325e-19 $X=0.975 $Y=1.615 $X2=0
+ $Y2=0
cc_113 B2 N_A_270_48#_c_152_n 0.00246192f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_B2_c_117_n N_A_270_48#_c_152_n 0.0208226f $X=0.975 $Y=1.615 $X2=0 $Y2=0
cc_115 B2 N_A_204_392#_c_325_n 0.0203326f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B2_c_117_n N_A_204_392#_c_325_n 0.00207331f $X=0.975 $Y=1.615 $X2=0
+ $Y2=0
cc_117 N_B2_M1011_g N_A_204_392#_c_326_n 2.95416e-19 $X=0.93 $Y=2.46 $X2=0 $Y2=0
cc_118 N_B2_M1010_g N_A_204_392#_c_316_n 3.08164e-19 $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_B2_M1011_g N_VPWR_c_438_n 0.0035407f $X=0.93 $Y=2.46 $X2=0 $Y2=0
cc_120 N_B2_M1011_g N_VPWR_c_443_n 0.00553757f $X=0.93 $Y=2.46 $X2=0 $Y2=0
cc_121 N_B2_M1011_g N_VPWR_c_436_n 0.0109022f $X=0.93 $Y=2.46 $X2=0 $Y2=0
cc_122 N_B2_M1010_g N_A_27_74#_c_524_n 0.0143059f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_123 B2 N_A_27_74#_c_524_n 0.0378094f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_124 N_B2_c_117_n N_A_27_74#_c_524_n 0.00422609f $X=0.975 $Y=1.615 $X2=0 $Y2=0
cc_125 N_B2_M1010_g N_A_27_74#_c_526_n 4.69391e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B2_M1010_g N_VGND_c_549_n 0.0106075f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B2_M1010_g N_VGND_c_554_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B2_M1010_g N_VGND_c_558_n 0.00758251f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_270_48#_c_164_p N_A2_N_M1000_g 0.0128987f $X=2.355 $Y=2.14 $X2=0
+ $Y2=0
cc_130 N_A_270_48#_c_150_n N_A2_N_c_220_n 0.00725711f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_131 N_A_270_48#_M1005_g N_A2_N_c_221_n 0.00362293f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_270_48#_c_148_n N_A2_N_c_221_n 0.00538493f $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_133 N_A_270_48#_c_150_n N_A2_N_c_221_n 0.00587895f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_134 N_A_270_48#_c_148_n A2_N 0.0267167f $X=2.045 $Y=1.22 $X2=0 $Y2=0
cc_135 N_A_270_48#_c_164_p A2_N 0.0223637f $X=2.355 $Y=2.14 $X2=0 $Y2=0
cc_136 N_A_270_48#_c_151_n A2_N 0.0208999f $X=1.62 $Y=1.615 $X2=0 $Y2=0
cc_137 N_A_270_48#_c_152_n A2_N 0.00111877f $X=1.62 $Y=1.615 $X2=0 $Y2=0
cc_138 N_A_270_48#_M1004_g N_A2_N_c_223_n 0.0247739f $X=1.44 $Y=2.46 $X2=0 $Y2=0
cc_139 N_A_270_48#_c_155_n N_A2_N_c_223_n 0.00385561f $X=1.7 $Y=1.975 $X2=0
+ $Y2=0
cc_140 N_A_270_48#_c_148_n N_A2_N_c_223_n 0.00135402f $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_141 N_A_270_48#_c_164_p N_A2_N_c_223_n 9.30623e-19 $X=2.355 $Y=2.14 $X2=0
+ $Y2=0
cc_142 N_A_270_48#_c_151_n N_A2_N_c_223_n 0.00106229f $X=1.62 $Y=1.615 $X2=0
+ $Y2=0
cc_143 N_A_270_48#_c_152_n N_A2_N_c_223_n 0.0189833f $X=1.62 $Y=1.615 $X2=0
+ $Y2=0
cc_144 N_A_270_48#_c_148_n N_A2_N_c_224_n 0.00498608f $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_145 N_A_270_48#_c_152_n N_A2_N_c_224_n 8.57091e-19 $X=1.62 $Y=1.615 $X2=0
+ $Y2=0
cc_146 N_A_270_48#_c_153_n N_A2_N_c_224_n 0.00265089f $X=1.62 $Y=1.45 $X2=0
+ $Y2=0
cc_147 N_A_270_48#_c_164_p N_A1_N_M1002_g 0.00586003f $X=2.355 $Y=2.14 $X2=0
+ $Y2=0
cc_148 N_A_270_48#_c_148_n N_A1_N_M1007_g 2.68167e-19 $X=2.045 $Y=1.22 $X2=0
+ $Y2=0
cc_149 N_A_270_48#_c_164_p A1_N 0.00258484f $X=2.355 $Y=2.14 $X2=0 $Y2=0
cc_150 N_A_270_48#_M1004_g N_A_204_392#_c_325_n 0.00889452f $X=1.44 $Y=2.46
+ $X2=0 $Y2=0
cc_151 N_A_270_48#_c_155_n N_A_204_392#_c_325_n 0.00142441f $X=1.7 $Y=1.975
+ $X2=0 $Y2=0
cc_152 N_A_270_48#_c_187_p N_A_204_392#_c_325_n 0.016089f $X=1.785 $Y=2.1 $X2=0
+ $Y2=0
cc_153 N_A_270_48#_M1004_g N_A_204_392#_c_326_n 0.00726292f $X=1.44 $Y=2.46
+ $X2=0 $Y2=0
cc_154 N_A_270_48#_M1000_d N_A_204_392#_c_336_n 0.00715971f $X=2.175 $Y=1.965
+ $X2=0 $Y2=0
cc_155 N_A_270_48#_M1004_g N_A_204_392#_c_336_n 0.0137399f $X=1.44 $Y=2.46 $X2=0
+ $Y2=0
cc_156 N_A_270_48#_c_187_p N_A_204_392#_c_336_n 0.0137412f $X=1.785 $Y=2.1 $X2=0
+ $Y2=0
cc_157 N_A_270_48#_c_164_p N_A_204_392#_c_336_n 0.0444004f $X=2.355 $Y=2.14
+ $X2=0 $Y2=0
cc_158 N_A_270_48#_c_151_n N_A_204_392#_c_336_n 0.00331377f $X=1.62 $Y=1.615
+ $X2=0 $Y2=0
cc_159 N_A_270_48#_c_152_n N_A_204_392#_c_336_n 7.31134e-19 $X=1.62 $Y=1.615
+ $X2=0 $Y2=0
cc_160 N_A_270_48#_M1005_g N_A_204_392#_c_314_n 0.00610421f $X=1.425 $Y=0.74
+ $X2=0 $Y2=0
cc_161 N_A_270_48#_c_148_n N_A_204_392#_c_314_n 0.00157271f $X=2.045 $Y=1.22
+ $X2=0 $Y2=0
cc_162 N_A_270_48#_c_149_n N_A_204_392#_c_314_n 0.0156773f $X=1.785 $Y=1.22
+ $X2=0 $Y2=0
cc_163 N_A_270_48#_c_150_n N_A_204_392#_c_314_n 0.0242222f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_164 N_A_270_48#_c_151_n N_A_204_392#_c_314_n 0.00385199f $X=1.62 $Y=1.615
+ $X2=0 $Y2=0
cc_165 N_A_270_48#_c_152_n N_A_204_392#_c_314_n 0.00120341f $X=1.62 $Y=1.615
+ $X2=0 $Y2=0
cc_166 N_A_270_48#_M1003_s N_A_204_392#_c_315_n 0.00264658f $X=2.065 $Y=0.37
+ $X2=0 $Y2=0
cc_167 N_A_270_48#_c_150_n N_A_204_392#_c_315_n 0.020634f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_168 N_A_270_48#_M1005_g N_A_204_392#_c_316_n 0.00544881f $X=1.425 $Y=0.74
+ $X2=0 $Y2=0
cc_169 N_A_270_48#_c_150_n N_A_204_392#_c_317_n 0.0248147f $X=2.21 $Y=0.81 $X2=0
+ $Y2=0
cc_170 N_A_270_48#_c_148_n N_A_204_392#_c_319_n 0.0155236f $X=2.045 $Y=1.22
+ $X2=0 $Y2=0
cc_171 N_A_270_48#_c_164_p N_A_204_392#_c_321_n 0.00810662f $X=2.355 $Y=2.14
+ $X2=0 $Y2=0
cc_172 N_A_270_48#_M1004_g N_A_204_392#_c_354_n 4.64231e-19 $X=1.44 $Y=2.46
+ $X2=0 $Y2=0
cc_173 N_A_270_48#_c_155_n N_VPWR_M1004_d 3.66442e-19 $X=1.7 $Y=1.975 $X2=0
+ $Y2=0
cc_174 N_A_270_48#_c_187_p N_VPWR_M1004_d 0.00654385f $X=1.785 $Y=2.1 $X2=0
+ $Y2=0
cc_175 N_A_270_48#_c_164_p N_VPWR_M1004_d 0.00508296f $X=2.355 $Y=2.14 $X2=0
+ $Y2=0
cc_176 N_A_270_48#_M1004_g N_VPWR_c_439_n 0.00703872f $X=1.44 $Y=2.46 $X2=0
+ $Y2=0
cc_177 N_A_270_48#_M1004_g N_VPWR_c_443_n 0.005209f $X=1.44 $Y=2.46 $X2=0 $Y2=0
cc_178 N_A_270_48#_M1004_g N_VPWR_c_436_n 0.00520071f $X=1.44 $Y=2.46 $X2=0
+ $Y2=0
cc_179 N_A_270_48#_M1005_g N_A_27_74#_c_524_n 0.00252956f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_A_270_48#_c_149_n N_A_27_74#_c_524_n 0.00890055f $X=1.785 $Y=1.22 $X2=0
+ $Y2=0
cc_181 N_A_270_48#_M1005_g N_A_27_74#_c_526_n 0.00402051f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_182 N_A_270_48#_M1005_g N_VGND_c_549_n 5.20809e-19 $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_270_48#_M1005_g N_VGND_c_554_n 0.00430908f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_270_48#_M1005_g N_VGND_c_558_n 0.00822378f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A2_N_M1000_g N_A1_N_M1002_g 0.0282251f $X=2.085 $Y=2.385 $X2=0 $Y2=0
cc_186 N_A2_N_c_220_n N_A1_N_M1007_g 0.0451706f $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_187 N_A2_N_c_224_n N_A1_N_M1007_g 0.0078326f $X=2.16 $Y=1.475 $X2=0 $Y2=0
cc_188 A2_N A1_N 0.0231358f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_N_c_223_n A1_N 0.00187659f $X=2.16 $Y=1.64 $X2=0 $Y2=0
cc_190 A2_N N_A1_N_c_270_n 4.04807e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A2_N_c_223_n N_A1_N_c_270_n 0.0207555f $X=2.16 $Y=1.64 $X2=0 $Y2=0
cc_192 N_A2_N_M1000_g N_A_204_392#_c_325_n 9.17423e-19 $X=2.085 $Y=2.385 $X2=0
+ $Y2=0
cc_193 N_A2_N_M1000_g N_A_204_392#_c_326_n 7.83337e-19 $X=2.085 $Y=2.385 $X2=0
+ $Y2=0
cc_194 N_A2_N_M1000_g N_A_204_392#_c_336_n 0.014262f $X=2.085 $Y=2.385 $X2=0
+ $Y2=0
cc_195 N_A2_N_c_220_n N_A_204_392#_c_314_n 0.00494986f $X=2.425 $Y=1.085 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_220_n N_A_204_392#_c_315_n 0.0143941f $X=2.425 $Y=1.085 $X2=0
+ $Y2=0
cc_197 N_A2_N_c_221_n N_A_204_392#_c_315_n 4.10115e-19 $X=2.425 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_220_n N_A_204_392#_c_317_n 0.00304192f $X=2.425 $Y=1.085 $X2=0
+ $Y2=0
cc_199 N_A2_N_c_221_n N_A_204_392#_c_319_n 8.38832e-19 $X=2.425 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A2_N_c_224_n N_A_204_392#_c_319_n 2.70295e-19 $X=2.16 $Y=1.475 $X2=0
+ $Y2=0
cc_201 N_A2_N_M1000_g N_VPWR_c_439_n 0.00435235f $X=2.085 $Y=2.385 $X2=0 $Y2=0
cc_202 N_A2_N_M1000_g N_VPWR_c_444_n 0.00566528f $X=2.085 $Y=2.385 $X2=0 $Y2=0
cc_203 N_A2_N_M1000_g N_VPWR_c_436_n 0.00597552f $X=2.085 $Y=2.385 $X2=0 $Y2=0
cc_204 N_A2_N_c_220_n N_VGND_c_550_n 3.72445e-19 $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_205 N_A2_N_c_220_n N_VGND_c_554_n 0.00278271f $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_206 N_A2_N_c_220_n N_VGND_c_558_n 0.00358137f $X=2.425 $Y=1.085 $X2=0 $Y2=0
cc_207 N_A1_N_M1002_g N_A_204_392#_M1008_g 0.0174551f $X=2.625 $Y=2.385 $X2=0
+ $Y2=0
cc_208 N_A1_N_c_270_n N_A_204_392#_M1008_g 0.00410391f $X=2.815 $Y=1.64 $X2=0
+ $Y2=0
cc_209 N_A1_N_M1007_g N_A_204_392#_M1001_g 0.0165087f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_210 N_A1_N_M1002_g N_A_204_392#_c_336_n 0.0164894f $X=2.625 $Y=2.385 $X2=0
+ $Y2=0
cc_211 A1_N N_A_204_392#_c_336_n 0.00718092f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A1_N_c_270_n N_A_204_392#_c_336_n 0.00324305f $X=2.815 $Y=1.64 $X2=0
+ $Y2=0
cc_213 N_A1_N_M1007_g N_A_204_392#_c_315_n 0.0011351f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_214 N_A1_N_M1007_g N_A_204_392#_c_317_n 0.0052743f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_215 N_A1_N_M1007_g N_A_204_392#_c_318_n 0.0153044f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_216 A1_N N_A_204_392#_c_318_n 0.0107679f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A1_N_c_270_n N_A_204_392#_c_318_n 5.5832e-19 $X=2.815 $Y=1.64 $X2=0
+ $Y2=0
cc_218 A1_N N_A_204_392#_c_319_n 0.0143367f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A1_N_c_270_n N_A_204_392#_c_319_n 0.00463077f $X=2.815 $Y=1.64 $X2=0
+ $Y2=0
cc_220 N_A1_N_M1007_g N_A_204_392#_c_320_n 0.00478972f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_221 A1_N N_A_204_392#_c_320_n 0.0105181f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_222 N_A1_N_M1002_g N_A_204_392#_c_321_n 0.00837652f $X=2.625 $Y=2.385 $X2=0
+ $Y2=0
cc_223 A1_N N_A_204_392#_c_321_n 0.0105017f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A1_N_c_270_n N_A_204_392#_c_321_n 0.00133027f $X=2.815 $Y=1.64 $X2=0
+ $Y2=0
cc_225 N_A1_N_M1007_g N_A_204_392#_c_322_n 0.020241f $X=2.815 $Y=0.69 $X2=0
+ $Y2=0
cc_226 N_A1_N_M1002_g N_VPWR_c_440_n 0.00473371f $X=2.625 $Y=2.385 $X2=0 $Y2=0
cc_227 N_A1_N_M1002_g N_VPWR_c_444_n 0.00566528f $X=2.625 $Y=2.385 $X2=0 $Y2=0
cc_228 N_A1_N_M1002_g N_VPWR_c_436_n 0.00597552f $X=2.625 $Y=2.385 $X2=0 $Y2=0
cc_229 N_A1_N_M1007_g N_X_c_491_n 6.44522e-19 $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_230 N_A1_N_M1007_g N_VGND_c_550_n 0.00814171f $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_231 N_A1_N_M1007_g N_VGND_c_554_n 0.00444681f $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_232 N_A1_N_M1007_g N_VGND_c_558_n 0.00877228f $X=2.815 $Y=0.69 $X2=0 $Y2=0
cc_233 N_A_204_392#_c_336_n N_VPWR_M1004_d 0.00830915f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_234 N_A_204_392#_c_336_n N_VPWR_M1002_d 0.0170865f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_235 N_A_204_392#_c_321_n N_VPWR_M1002_d 0.0118691f $X=3.17 $Y=2.395 $X2=0
+ $Y2=0
cc_236 N_A_204_392#_c_325_n N_VPWR_c_438_n 0.0060319f $X=1.215 $Y=2.115 $X2=0
+ $Y2=0
cc_237 N_A_204_392#_c_326_n N_VPWR_c_438_n 0.00580593f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_238 N_A_204_392#_c_326_n N_VPWR_c_439_n 0.00861474f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_239 N_A_204_392#_c_336_n N_VPWR_c_439_n 0.0277276f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_240 N_A_204_392#_M1008_g N_VPWR_c_440_n 0.00739572f $X=3.365 $Y=2.4 $X2=0
+ $Y2=0
cc_241 N_A_204_392#_c_336_n N_VPWR_c_440_n 0.0362574f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_242 N_A_204_392#_M1012_g N_VPWR_c_442_n 0.00648292f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_243 N_A_204_392#_c_326_n N_VPWR_c_443_n 0.014549f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_244 N_A_204_392#_M1008_g N_VPWR_c_445_n 0.005209f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A_204_392#_M1012_g N_VPWR_c_445_n 0.00503905f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_246 N_A_204_392#_M1008_g N_VPWR_c_436_n 0.00987511f $X=3.365 $Y=2.4 $X2=0
+ $Y2=0
cc_247 N_A_204_392#_M1012_g N_VPWR_c_436_n 0.00930977f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_248 N_A_204_392#_c_326_n N_VPWR_c_436_n 0.0119743f $X=1.215 $Y=2.815 $X2=0
+ $Y2=0
cc_249 N_A_204_392#_c_336_n N_VPWR_c_436_n 0.0404216f $X=3.085 $Y=2.48 $X2=0
+ $Y2=0
cc_250 N_A_204_392#_M1001_g N_X_c_490_n 0.00812178f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_204_392#_M1013_g N_X_c_490_n 0.0081896f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_204_392#_M1001_g N_X_c_491_n 0.00488854f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_204_392#_M1013_g N_X_c_491_n 0.00215589f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_204_392#_c_322_n N_X_c_491_n 0.0024311f $X=3.815 $Y=1.47 $X2=0 $Y2=0
cc_255 N_A_204_392#_M1008_g X 0.0037471f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A_204_392#_M1012_g X 0.00248815f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A_204_392#_c_321_n X 0.0223997f $X=3.17 $Y=2.395 $X2=0 $Y2=0
cc_258 N_A_204_392#_c_322_n X 0.00240502f $X=3.815 $Y=1.47 $X2=0 $Y2=0
cc_259 N_A_204_392#_M1008_g X 0.0184424f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_204_392#_M1012_g X 0.0142441f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A_204_392#_M1008_g N_X_c_492_n 0.00106126f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_204_392#_M1001_g N_X_c_492_n 9.7705e-19 $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_204_392#_M1012_g N_X_c_492_n 0.00952496f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_204_392#_M1013_g N_X_c_492_n 0.00886097f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_204_392#_c_320_n N_X_c_492_n 0.0302315f $X=3.17 $Y=1.635 $X2=0 $Y2=0
cc_266 N_A_204_392#_c_321_n N_X_c_492_n 0.00618571f $X=3.17 $Y=2.395 $X2=0 $Y2=0
cc_267 N_A_204_392#_c_322_n N_X_c_492_n 0.0242635f $X=3.815 $Y=1.47 $X2=0 $Y2=0
cc_268 N_A_204_392#_c_325_n N_A_27_74#_c_524_n 7.14544e-19 $X=1.215 $Y=2.115
+ $X2=0 $Y2=0
cc_269 N_A_204_392#_c_316_n N_A_27_74#_c_526_n 0.00392044f $X=1.805 $Y=0.34
+ $X2=0 $Y2=0
cc_270 N_A_204_392#_c_316_n N_VGND_c_549_n 0.00266256f $X=1.805 $Y=0.34 $X2=0
+ $Y2=0
cc_271 N_A_204_392#_M1001_g N_VGND_c_550_n 0.00866971f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_272 N_A_204_392#_c_315_n N_VGND_c_550_n 0.0117236f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_273 N_A_204_392#_c_318_n N_VGND_c_550_n 0.013791f $X=3.085 $Y=1.22 $X2=0
+ $Y2=0
cc_274 N_A_204_392#_c_320_n N_VGND_c_550_n 0.0118589f $X=3.17 $Y=1.635 $X2=0
+ $Y2=0
cc_275 N_A_204_392#_c_322_n N_VGND_c_550_n 6.03907e-19 $X=3.815 $Y=1.47 $X2=0
+ $Y2=0
cc_276 N_A_204_392#_M1013_g N_VGND_c_552_n 0.00646793f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_A_204_392#_c_315_n N_VGND_c_554_n 0.0593614f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_278 N_A_204_392#_c_316_n N_VGND_c_554_n 0.0236456f $X=1.805 $Y=0.34 $X2=0
+ $Y2=0
cc_279 N_A_204_392#_M1001_g N_VGND_c_555_n 0.00434272f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_204_392#_M1013_g N_VGND_c_555_n 0.00422942f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_281 N_A_204_392#_M1001_g N_VGND_c_558_n 0.00822284f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_204_392#_M1013_g N_VGND_c_558_n 0.00787305f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_204_392#_c_315_n N_VGND_c_558_n 0.0337409f $X=2.545 $Y=0.34 $X2=0
+ $Y2=0
cc_284 N_A_204_392#_c_316_n N_VGND_c_558_n 0.0127298f $X=1.805 $Y=0.34 $X2=0
+ $Y2=0
cc_285 N_A_204_392#_c_317_n A_500_74# 0.00249342f $X=2.63 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_286 N_VPWR_c_442_n X 0.0423444f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_287 N_VPWR_c_440_n X 0.00869434f $X=2.995 $Y=2.9 $X2=0 $Y2=0
cc_288 N_VPWR_c_445_n X 0.0150868f $X=3.955 $Y=3.33 $X2=0 $Y2=0
cc_289 N_VPWR_c_436_n X 0.012316f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_290 N_X_c_490_n N_VGND_c_550_n 0.0399419f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_291 N_X_c_490_n N_VGND_c_552_n 0.0308798f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_292 N_X_c_490_n N_VGND_c_555_n 0.0149085f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_293 N_X_c_490_n N_VGND_c_558_n 0.0122037f $X=3.595 $Y=0.515 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_523_n N_VGND_c_549_n 0.0218743f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_524_n N_VGND_c_549_n 0.0216087f $X=1.055 $Y=1.195 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_c_526_n N_VGND_c_549_n 0.0218743f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_523_n N_VGND_c_553_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_526_n N_VGND_c_554_n 0.011066f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_523_n N_VGND_c_558_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_526_n N_VGND_c_558_n 0.00915947f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__nand4b_4.pex.spice
* Created: Fri Aug 28 17:45:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4B_4%A_N 3 5 7 8 10 12 13 14 23
r43 22 23 36.463 $w=4.25e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=1.512
+ $X2=1.035 $Y2=1.512
r44 20 22 35.9864 $w=4.25e-07 $l=2.75e-07 $layer=POLY_cond $X=0.67 $Y=1.512
+ $X2=0.945 $Y2=1.512
r45 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.465 $X2=0.67 $Y2=1.465
r46 14 21 1.24592 $w=4.78e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.54 $X2=0.67
+ $Y2=1.54
r47 13 21 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.67 $Y2=1.54
r48 10 12 143.261 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=1.395 $Y=1.725
+ $X2=1.395 $Y2=2.26
r49 8 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.305 $Y=1.65
+ $X2=1.395 $Y2=1.725
r50 8 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.305 $Y=1.65
+ $X2=1.035 $Y2=1.65
r51 5 22 22.9127 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=0.945 $Y=1.725
+ $X2=0.945 $Y2=1.512
r52 5 7 143.261 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=0.945 $Y=1.725
+ $X2=0.945 $Y2=2.26
r53 1 20 22.9005 $w=4.25e-07 $l=1.75e-07 $layer=POLY_cond $X=0.495 $Y=1.512
+ $X2=0.67 $Y2=1.512
r54 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%A_27_158# 1 2 7 9 10 11 12 14 17 19 21 22
+ 24 25 27 28 31 34 41 45 49 55
c98 22 0 1.62209e-19 $X=2.775 $Y=1.185
c99 19 0 5.66301e-20 $X=2.345 $Y=1.185
r100 55 56 1.45766 $w=4.96e-07 $l=1.5e-08 $layer=POLY_cond $X=2.775 $Y=1.477
+ $X2=2.79 $Y2=1.477
r101 45 47 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=0.95
+ $X2=0.28 $Y2=1.045
r102 42 55 8.74597 $w=4.96e-07 $l=9e-08 $layer=POLY_cond $X=2.685 $Y=1.477
+ $X2=2.775 $Y2=1.477
r103 42 53 33.0403 $w=4.96e-07 $l=3.4e-07 $layer=POLY_cond $X=2.685 $Y=1.477
+ $X2=2.345 $Y2=1.477
r104 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.685
+ $Y=1.515 $X2=2.685 $Y2=1.515
r105 39 53 33.0403 $w=4.96e-07 $l=3.4e-07 $layer=POLY_cond $X=2.005 $Y=1.477
+ $X2=2.345 $Y2=1.477
r106 38 41 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.005 $Y=1.555
+ $X2=2.685 $Y2=1.555
r107 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=1.515 $X2=2.005 $Y2=1.515
r108 36 49 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=1.555
+ $X2=1.17 $Y2=1.555
r109 36 38 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.335 $Y=1.555
+ $X2=2.005 $Y2=1.555
r110 32 49 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.17 $Y=1.68
+ $X2=1.17 $Y2=1.555
r111 32 34 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.17 $Y=1.68
+ $X2=1.17 $Y2=1.985
r112 31 49 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.17 $Y=1.43
+ $X2=1.17 $Y2=1.555
r113 30 31 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.17 $Y=1.13 $X2=1.17
+ $Y2=1.43
r114 29 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.045
+ $X2=0.28 $Y2=1.045
r115 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.005 $Y=1.045
+ $X2=1.17 $Y2=1.13
r116 28 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=1.045
+ $X2=0.445 $Y2=1.045
r117 25 56 26.6655 $w=1.8e-07 $l=2.93e-07 $layer=POLY_cond $X=2.79 $Y=1.77
+ $X2=2.79 $Y2=1.477
r118 25 27 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.79 $Y=1.77 $X2=2.79
+ $Y2=2.4
r119 22 55 31.2052 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=2.775 $Y=1.185
+ $X2=2.775 $Y2=1.477
r120 22 24 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.775 $Y=1.185
+ $X2=2.775 $Y2=0.74
r121 19 53 31.2052 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=2.345 $Y=1.185
+ $X2=2.345 $Y2=1.477
r122 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.345 $Y=1.185
+ $X2=2.345 $Y2=0.74
r123 15 39 7.28831 $w=4.96e-07 $l=7.5e-08 $layer=POLY_cond $X=1.93 $Y=1.477
+ $X2=2.005 $Y2=1.477
r124 15 50 1.45766 $w=4.96e-07 $l=1.5e-08 $layer=POLY_cond $X=1.93 $Y=1.477
+ $X2=1.915 $Y2=1.477
r125 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.93 $Y=1.68
+ $X2=1.93 $Y2=2.4
r126 12 50 31.2052 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=1.915 $Y=1.185
+ $X2=1.915 $Y2=1.477
r127 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.915 $Y=1.185
+ $X2=1.915 $Y2=0.74
r128 10 50 33.0766 $w=4.96e-07 $l=2.51722e-07 $layer=POLY_cond $X=1.84 $Y=1.26
+ $X2=1.915 $Y2=1.477
r129 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.84 $Y=1.26
+ $X2=1.56 $Y2=1.26
r130 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.56 $Y2=1.26
r131 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.485 $Y2=0.74
r132 2 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=1.985
r133 1 45 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.79 $X2=0.28 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%B 3 7 11 15 19 23 25 30 37
c65 23 0 7.64129e-20 $X=4.7 $Y=2.4
r66 36 37 36.5604 $w=3.23e-07 $l=2.45e-07 $layer=POLY_cond $X=4.25 $Y=1.515
+ $X2=4.495 $Y2=1.515
r67 35 36 27.6068 $w=3.23e-07 $l=1.85e-07 $layer=POLY_cond $X=4.065 $Y=1.515
+ $X2=4.25 $Y2=1.515
r68 33 35 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=3.975 $Y=1.515
+ $X2=4.065 $Y2=1.515
r69 31 33 50.7368 $w=3.23e-07 $l=3.4e-07 $layer=POLY_cond $X=3.635 $Y=1.515
+ $X2=3.975 $Y2=1.515
r70 30 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.515 $X2=3.975 $Y2=1.515
r71 29 31 50.7368 $w=3.23e-07 $l=3.4e-07 $layer=POLY_cond $X=3.295 $Y=1.515
+ $X2=3.635 $Y2=1.515
r72 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.515 $X2=3.295 $Y2=1.515
r73 27 29 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=3.205 $Y=1.515
+ $X2=3.295 $Y2=1.515
r74 25 30 1.81188 $w=1.008e-06 $l=1.5e-07 $layer=LI1_cond $X=3.635 $Y=1.665
+ $X2=3.635 $Y2=1.515
r75 21 37 30.5913 $w=3.23e-07 $l=2.05e-07 $layer=POLY_cond $X=4.7 $Y=1.515
+ $X2=4.495 $Y2=1.515
r76 21 23 289.589 $w=1.8e-07 $l=7.45e-07 $layer=POLY_cond $X=4.7 $Y=1.655
+ $X2=4.7 $Y2=2.4
r77 17 37 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.495 $Y=1.35
+ $X2=4.495 $Y2=1.515
r78 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.495 $Y=1.35
+ $X2=4.495 $Y2=0.74
r79 13 36 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.68
+ $X2=4.25 $Y2=1.515
r80 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.25 $Y=1.68
+ $X2=4.25 $Y2=2.4
r81 9 35 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.065 $Y=1.35
+ $X2=4.065 $Y2=1.515
r82 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.065 $Y=1.35
+ $X2=4.065 $Y2=0.74
r83 5 31 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=1.35
+ $X2=3.635 $Y2=1.515
r84 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.635 $Y=1.35
+ $X2=3.635 $Y2=0.74
r85 1 27 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.35
+ $X2=3.205 $Y2=1.515
r86 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.205 $Y=1.35
+ $X2=3.205 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%C 3 7 11 15 19 23 25 26 27 28 29 30 52
c68 23 0 4.25028e-20 $X=6.79 $Y=0.74
c69 15 0 1.36796e-19 $X=6.345 $Y=0.74
c70 7 0 5.58611e-20 $X=5.915 $Y=0.74
r71 51 52 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.775 $Y=1.515
+ $X2=6.79 $Y2=1.515
r72 49 51 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.7 $Y=1.515
+ $X2=6.775 $Y2=1.515
r73 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.7
+ $Y=1.515 $X2=6.7 $Y2=1.515
r74 47 49 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.345 $Y=1.515
+ $X2=6.7 $Y2=1.515
r75 45 47 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=6.02 $Y=1.515
+ $X2=6.345 $Y2=1.515
r76 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.02
+ $Y=1.515 $X2=6.02 $Y2=1.515
r77 43 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.945 $Y=1.515
+ $X2=6.02 $Y2=1.515
r78 42 43 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.915 $Y=1.515
+ $X2=5.945 $Y2=1.515
r79 40 42 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=5.68 $Y=1.515
+ $X2=5.915 $Y2=1.515
r80 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.68
+ $Y=1.515 $X2=5.68 $Y2=1.515
r81 37 40 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.485 $Y=1.515
+ $X2=5.68 $Y2=1.515
r82 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r83 29 50 6.96826 $w=4.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.7 $Y2=1.565
r84 28 50 5.89622 $w=4.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.7 $Y2=1.565
r85 28 46 12.3285 $w=4.28e-07 $l=4.6e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.02 $Y2=1.565
r86 27 46 0.53602 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=6 $Y=1.565 $X2=6.02
+ $Y2=1.565
r87 27 41 8.57632 $w=4.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.68
+ $Y2=1.565
r88 26 41 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.68 $Y2=1.565
r89 25 26 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r90 21 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.79 $Y=1.35
+ $X2=6.79 $Y2=1.515
r91 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.79 $Y=1.35
+ $X2=6.79 $Y2=0.74
r92 17 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.775 $Y=1.68
+ $X2=6.775 $Y2=1.515
r93 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.775 $Y=1.68
+ $X2=6.775 $Y2=2.4
r94 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.35
+ $X2=6.345 $Y2=1.515
r95 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.345 $Y=1.35
+ $X2=6.345 $Y2=0.74
r96 9 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.945 $Y=1.68
+ $X2=5.945 $Y2=1.515
r97 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.945 $Y=1.68
+ $X2=5.945 $Y2=2.4
r98 5 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.35
+ $X2=5.915 $Y2=1.515
r99 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.915 $Y=1.35
+ $X2=5.915 $Y2=0.74
r100 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.35
+ $X2=5.485 $Y2=1.515
r101 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.485 $Y=1.35
+ $X2=5.485 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%D 3 5 6 9 15 19 23 27 29 30 31 32 37 45
c70 19 0 1.85163e-19 $X=8.095 $Y=2.4
r71 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.85
+ $Y=1.465 $X2=8.85 $Y2=1.465
r72 43 45 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=8.625 $Y=1.465
+ $X2=8.85 $Y2=1.465
r73 42 43 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.565 $Y=1.465
+ $X2=8.625 $Y2=1.465
r74 41 46 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=8.51 $Y=1.54
+ $X2=8.85 $Y2=1.54
r75 40 42 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=8.51 $Y=1.465
+ $X2=8.565 $Y2=1.465
r76 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.51
+ $Y=1.465 $X2=8.51 $Y2=1.465
r77 38 40 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.095 $Y=1.465
+ $X2=8.51 $Y2=1.465
r78 36 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.08 $Y=1.465
+ $X2=8.095 $Y2=1.465
r79 36 37 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.08 $Y=1.465
+ $X2=8.005 $Y2=1.465
r80 32 46 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=8.88 $Y=1.54 $X2=8.85
+ $Y2=1.54
r81 31 41 2.74101 $w=4.78e-07 $l=1.1e-07 $layer=LI1_cond $X=8.4 $Y=1.54 $X2=8.51
+ $Y2=1.54
r82 30 31 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.54 $X2=8.4
+ $Y2=1.54
r83 25 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=1.465
r84 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=0.74
r85 21 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.63
+ $X2=8.565 $Y2=1.465
r86 21 23 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.565 $Y=1.63
+ $X2=8.565 $Y2=2.4
r87 17 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.63
+ $X2=8.095 $Y2=1.465
r88 17 19 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.095 $Y=1.63
+ $X2=8.095 $Y2=2.4
r89 13 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.08 $Y=1.3
+ $X2=8.08 $Y2=1.465
r90 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.08 $Y=1.3 $X2=8.08
+ $Y2=0.74
r91 12 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.725 $Y=1.375
+ $X2=7.65 $Y2=1.375
r92 12 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.725 $Y=1.375
+ $X2=8.005 $Y2=1.375
r93 7 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.65 $Y=1.3 $X2=7.65
+ $Y2=1.375
r94 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.65 $Y=1.3 $X2=7.65
+ $Y2=0.74
r95 5 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.575 $Y=1.375
+ $X2=7.65 $Y2=1.375
r96 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.575 $Y=1.375
+ $X2=7.295 $Y2=1.375
r97 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.22 $Y=1.3
+ $X2=7.295 $Y2=1.375
r98 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.22 $Y=1.3 $X2=7.22
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 37 42 52 62
+ 68 71 75 84 86 96 104 107
r81 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r82 102 104 12.9833 $w=1.123e-06 $l=1.15e-07 $layer=LI1_cond $X=7.92 $Y=2.852
+ $X2=8.035 $Y2=2.852
r83 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r84 100 102 0.542222 $w=1.123e-06 $l=5e-08 $layer=LI1_cond $X=7.87 $Y=2.852
+ $X2=7.92 $Y2=2.852
r85 98 100 9.43467 $w=1.123e-06 $l=8.7e-07 $layer=LI1_cond $X=7 $Y=2.852
+ $X2=7.87 $Y2=2.852
r86 95 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r87 94 98 0.433778 $w=1.123e-06 $l=4e-08 $layer=LI1_cond $X=6.96 $Y=2.852 $X2=7
+ $Y2=2.852
r88 94 96 13.0917 $w=1.123e-06 $l=1.25e-07 $layer=LI1_cond $X=6.96 $Y=2.852
+ $X2=6.835 $Y2=2.852
r89 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r90 82 84 12.929 $w=1.123e-06 $l=1.1e-07 $layer=LI1_cond $X=4.08 $Y=2.852
+ $X2=4.19 $Y2=2.852
r91 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r92 80 82 0.596444 $w=1.123e-06 $l=5.5e-08 $layer=LI1_cond $X=4.025 $Y=2.852
+ $X2=4.08 $Y2=2.852
r93 78 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r94 77 80 9.81422 $w=1.123e-06 $l=9.05e-07 $layer=LI1_cond $X=3.12 $Y=2.852
+ $X2=4.025 $Y2=2.852
r95 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 74 77 1.13867 $w=1.123e-06 $l=1.05e-07 $layer=LI1_cond $X=3.015 $Y=2.852
+ $X2=3.12 $Y2=2.852
r97 74 75 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.852
+ $X2=2.85 $Y2=2.852
r98 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 66 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r101 66 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r102 65 104 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=8.035 $Y2=3.33
r103 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r104 62 106 4.20034 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.897 $Y2=3.33
r105 62 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 61 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r107 61 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 60 96 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=6.835 $Y2=3.33
r109 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 58 60 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 55 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.19 $Y2=3.33
r112 52 58 12.5397 $w=1.7e-07 $l=5.63e-07 $layer=LI1_cond $X=5.322 $Y=3.33
+ $X2=5.885 $Y2=3.33
r113 52 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 52 86 10.3564 $w=1.123e-06 $l=9.55e-07 $layer=LI1_cond $X=5.322 $Y=3.33
+ $X2=5.322 $Y2=2.375
r115 52 55 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.76 $Y=3.33 $X2=4.56
+ $Y2=3.33
r116 51 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 51 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 50 75 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.85 $Y2=3.33
r119 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=1.705 $Y2=3.33
r121 48 50 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 46 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r125 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.67 $Y2=3.33
r126 43 45 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 42 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.705 $Y2=3.33
r128 42 45 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 40 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 37 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.67 $Y2=3.33
r132 37 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 35 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r134 35 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 35 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 31 34 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=8.815 $Y=2.115
+ $X2=8.815 $Y2=2.815
r137 29 106 3.15971 $w=2.8e-07 $l=1.19143e-07 $layer=LI1_cond $X=8.815 $Y=3.245
+ $X2=8.897 $Y2=3.33
r138 29 34 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=8.815 $Y=3.245
+ $X2=8.815 $Y2=2.815
r139 25 28 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=1.705 $Y=2.015
+ $X2=1.705 $Y2=2.815
r140 23 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=3.33
r141 23 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=2.815
r142 19 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=3.245
+ $X2=0.67 $Y2=3.33
r143 19 21 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.67 $Y=3.245
+ $X2=0.67 $Y2=2.115
r144 6 34 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.655
+ $Y=1.84 $X2=8.79 $Y2=2.815
r145 6 31 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.655
+ $Y=1.84 $X2=8.79 $Y2=2.115
r146 5 100 200 $w=1.7e-07 $l=1.24407e-06 $layer=licon1_PDIFF $count=3 $X=6.865
+ $Y=1.84 $X2=7.87 $Y2=2.375
r147 5 98 200 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=3 $X=6.865
+ $Y=1.84 $X2=7 $Y2=2.375
r148 4 86 200 $w=1.7e-07 $l=1.16724e-06 $layer=licon1_PDIFF $count=3 $X=4.79
+ $Y=1.84 $X2=5.72 $Y2=2.375
r149 4 86 200 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=3 $X=4.79
+ $Y=1.84 $X2=4.925 $Y2=2.375
r150 3 80 200 $w=1.7e-07 $l=1.38694e-06 $layer=licon1_PDIFF $count=3 $X=2.88
+ $Y=1.84 $X2=4.025 $Y2=2.375
r151 3 74 200 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=3 $X=2.88
+ $Y=1.84 $X2=3.015 $Y2=2.375
r152 2 28 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.705 $Y2=2.815
r153 2 25 300 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.705 $Y2=2.015
r154 1 21 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.525
+ $Y=1.84 $X2=0.67 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%Y 1 2 3 4 5 6 19 23 25 29 33 35 39 41 43 45
+ 50 57 61 63 66 69 71
c111 45 0 1.85163e-19 $X=8.34 $Y=2.43
c112 29 0 5.66301e-20 $X=4.445 $Y=1.175
c113 19 0 4.54593e-20 $X=2.395 $Y=1.005
r114 69 71 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.56 $Y=1.26
+ $X2=4.56 $Y2=1.295
r115 66 69 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=1.175
+ $X2=4.56 $Y2=1.26
r116 66 71 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.56 $Y=1.32
+ $X2=4.56 $Y2=1.295
r117 60 66 25.0531 $w=2.28e-07 $l=5e-07 $layer=LI1_cond $X=4.56 $Y=1.82 $X2=4.56
+ $Y2=1.32
r118 59 61 6.5639 $w=2.98e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.97
+ $X2=4.675 $Y2=1.97
r119 59 60 2.29563 $w=2.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.56 $Y=1.97
+ $X2=4.56 $Y2=1.82
r120 58 59 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=4.48 $Y=1.97 $X2=4.56
+ $Y2=1.97
r121 56 58 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=4.475 $Y=1.97
+ $X2=4.48 $Y2=1.97
r122 56 57 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=1.97
+ $X2=4.31 $Y2=1.97
r123 52 53 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.56 $Y=1.005
+ $X2=2.56 $Y2=1.175
r124 50 52 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.56 $Y=0.86
+ $X2=2.56 $Y2=1.005
r125 43 65 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=2.12
+ $X2=8.36 $Y2=2.035
r126 43 45 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=8.36 $Y=2.12
+ $X2=8.36 $Y2=2.43
r127 42 63 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=6.66 $Y=2.035
+ $X2=6.362 $Y2=2.035
r128 41 65 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=8.215 $Y=2.035
+ $X2=8.36 $Y2=2.035
r129 41 42 101.449 $w=1.68e-07 $l=1.555e-06 $layer=LI1_cond $X=8.215 $Y=2.035
+ $X2=6.66 $Y2=2.035
r130 37 63 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.362 $Y=2.12
+ $X2=6.362 $Y2=2.035
r131 37 39 6.23167 $w=5.93e-07 $l=3.1e-07 $layer=LI1_cond $X=6.362 $Y=2.12
+ $X2=6.362 $Y2=2.43
r132 35 63 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=6.065 $Y=2.035
+ $X2=6.362 $Y2=2.035
r133 35 61 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=6.065 $Y=2.035
+ $X2=4.675 $Y2=2.035
r134 31 58 2.55512 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=4.48 $Y=2.12
+ $X2=4.48 $Y2=1.97
r135 31 33 14.6675 $w=2.18e-07 $l=2.8e-07 $layer=LI1_cond $X=4.48 $Y=2.12
+ $X2=4.48 $Y2=2.4
r136 30 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.175
+ $X2=2.56 $Y2=1.175
r137 29 66 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.445 $Y=1.175
+ $X2=4.56 $Y2=1.175
r138 29 30 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=4.445 $Y=1.175
+ $X2=2.725 $Y2=1.175
r139 28 48 7.3732 $w=1.7e-07 $l=3.3908e-07 $layer=LI1_cond $X=2.68 $Y=2.035
+ $X2=2.365 $Y2=1.985
r140 28 57 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=2.68 $Y=2.035
+ $X2=4.31 $Y2=2.035
r141 23 48 2.82808 $w=6.2e-07 $l=1.37477e-07 $layer=LI1_cond $X=2.36 $Y=2.12
+ $X2=2.365 $Y2=1.985
r142 23 25 5.69102 $w=6.18e-07 $l=2.95e-07 $layer=LI1_cond $X=2.36 $Y=2.12
+ $X2=2.36 $Y2=2.415
r143 19 52 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=1.005
+ $X2=2.56 $Y2=1.005
r144 19 21 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=2.395 $Y=1.005
+ $X2=1.7 $Y2=1.005
r145 6 65 600 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.84 $X2=8.34 $Y2=2.035
r146 6 45 300 $w=1.7e-07 $l=6.62986e-07 $layer=licon1_PDIFF $count=2 $X=8.185
+ $Y=1.84 $X2=8.34 $Y2=2.43
r147 5 63 300 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.84 $X2=6.55 $Y2=2.035
r148 5 39 150 $w=1.7e-07 $l=8.07434e-07 $layer=licon1_PDIFF $count=4 $X=6.035
+ $Y=1.84 $X2=6.55 $Y2=2.43
r149 4 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.34
+ $Y=1.84 $X2=4.475 $Y2=1.985
r150 4 33 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=4.34
+ $Y=1.84 $X2=4.475 $Y2=2.4
r151 3 48 300 $w=1.7e-07 $l=6.26418e-07 $layer=licon1_PDIFF $count=2 $X=2.02
+ $Y=1.84 $X2=2.565 $Y2=2.015
r152 3 25 150 $w=1.7e-07 $l=8.02496e-07 $layer=licon1_PDIFF $count=4 $X=2.02
+ $Y=1.84 $X2=2.565 $Y2=2.415
r153 2 50 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.37 $X2=2.56 $Y2=0.86
r154 1 21 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48 51
+ 54
r91 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r92 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r93 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r95 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r96 42 54 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.317
+ $Y2=0
r97 42 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.88
+ $Y2=0
r98 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r99 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r100 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r101 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.6 $Y=0 $X2=7.435
+ $Y2=0
r102 38 40 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.6 $Y=0 $X2=7.92
+ $Y2=0
r103 37 54 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=8.13 $Y=0 $X2=8.317
+ $Y2=0
r104 37 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.13 $Y=0 $X2=7.92
+ $Y2=0
r105 36 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r106 35 36 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r107 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r108 32 35 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=6.96
+ $Y2=0
r109 32 33 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r110 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r111 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r112 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.27 $Y=0 $X2=7.435
+ $Y2=0
r113 29 35 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.27 $Y=0 $X2=6.96
+ $Y2=0
r114 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r115 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r116 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r117 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r118 22 36 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.96
+ $Y2=0
r119 22 33 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r120 18 54 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=8.317 $Y=0.085
+ $X2=8.317 $Y2=0
r121 18 20 16.2879 $w=3.73e-07 $l=5.3e-07 $layer=LI1_cond $X=8.317 $Y=0.085
+ $X2=8.317 $Y2=0.615
r122 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=0.085
+ $X2=7.435 $Y2=0
r123 14 16 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.435 $Y=0.085
+ $X2=7.435 $Y2=0.615
r124 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r125 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.515
r126 3 20 182 $w=1.7e-07 $l=3.15e-07 $layer=licon1_NDIFF $count=1 $X=8.155
+ $Y=0.37 $X2=8.315 $Y2=0.615
r127 2 16 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=7.295
+ $Y=0.37 $X2=7.435 $Y2=0.615
r128 1 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%A_225_74# 1 2 3 4 5 16 20 22 28 32 34 39
r56 34 37 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.27 $Y=0.34
+ $X2=1.27 $Y2=0.53
r57 30 32 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=3.85 $Y=0.835
+ $X2=4.71 $Y2=0.835
r58 28 30 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.075 $Y=0.835
+ $X2=3.85 $Y2=0.835
r59 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=0.75
+ $X2=3.075 $Y2=0.835
r60 25 27 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=0.75
+ $X2=2.99 $Y2=0.635
r61 24 27 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.99 $Y=0.425
+ $X2=2.99 $Y2=0.635
r62 23 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.215 $Y=0.34
+ $X2=2.09 $Y2=0.34
r63 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.99 $Y2=0.425
r64 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.215 $Y2=0.34
r65 18 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=0.425
+ $X2=2.09 $Y2=0.34
r66 18 20 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.09 $Y=0.425
+ $X2=2.09 $Y2=0.53
r67 17 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34
+ $X2=1.27 $Y2=0.34
r68 16 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.965 $Y=0.34
+ $X2=2.09 $Y2=0.34
r69 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.965 $Y=0.34
+ $X2=1.435 $Y2=0.34
r70 5 32 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.71 $Y2=0.835
r71 4 30 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.37 $X2=3.85 $Y2=0.835
r72 3 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.37 $X2=2.99 $Y2=0.635
r73 2 20 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.53
r74 1 37 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%A_656_74# 1 2 3 4 13 19 20 23
c45 19 0 4.25028e-20 $X=6.395 $Y=0.465
c46 13 0 1.16749e-19 $X=5.535 $Y=0.455
r47 23 26 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.56 $Y=0.465
+ $X2=6.56 $Y2=0.595
r48 20 22 3.98037 $w=3.5e-07 $l=1.19373e-07 $layer=LI1_cond $X=5.795 $Y=0.465
+ $X2=5.7 $Y2=0.52
r49 19 23 1.91462 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=0.465
+ $X2=6.56 $Y2=0.465
r50 19 20 25.6098 $w=2.68e-07 $l=6e-07 $layer=LI1_cond $X=6.395 $Y=0.465
+ $X2=5.795 $Y2=0.465
r51 15 18 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=3.42 $Y=0.455
+ $X2=4.28 $Y2=0.455
r52 13 22 6.76543 $w=3.5e-07 $l=1.94808e-07 $layer=LI1_cond $X=5.535 $Y=0.455
+ $X2=5.7 $Y2=0.52
r53 13 18 57.8526 $w=2.48e-07 $l=1.255e-06 $layer=LI1_cond $X=5.535 $Y=0.455
+ $X2=4.28 $Y2=0.455
r54 4 26 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=6.42
+ $Y=0.37 $X2=6.56 $Y2=0.595
r55 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.37 $X2=5.7 $Y2=0.515
r56 2 18 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.495
r57 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.37 $X2=3.42 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4B_4%A_1025_158# 1 2 3 4 5 16 22 24 28 30 34 37
+ 42 48 49 50
c73 48 0 5.58611e-20 $X=6.92 $Y=1.07
c74 42 0 1.36796e-19 $X=6.13 $Y=0.95
r75 47 49 9.00669 $w=2.18e-07 $l=1.6e-07 $layer=LI1_cond $X=7.01 $Y=1.07
+ $X2=7.17 $Y2=1.07
r76 47 48 5.33982 $w=2.18e-07 $l=9e-08 $layer=LI1_cond $X=7.01 $Y=1.07 $X2=6.92
+ $Y2=1.07
r77 44 45 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=6.09 $Y=1.045 $X2=6.09
+ $Y2=1.095
r78 42 44 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=6.09 $Y=0.95
+ $X2=6.09 $Y2=1.045
r79 37 39 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.27 $Y=0.95
+ $X2=5.27 $Y2=1.045
r80 32 34 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.84 $Y=0.96
+ $X2=8.84 $Y2=0.515
r81 31 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.96 $Y=1.045
+ $X2=7.865 $Y2=1.045
r82 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.675 $Y=1.045
+ $X2=8.84 $Y2=0.96
r83 30 31 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=8.675 $Y=1.045
+ $X2=7.96 $Y2=1.045
r84 26 50 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=0.96
+ $X2=7.865 $Y2=1.045
r85 26 28 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=7.865 $Y=0.96
+ $X2=7.865 $Y2=0.515
r86 24 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.77 $Y=1.045
+ $X2=7.865 $Y2=1.045
r87 24 49 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.77 $Y=1.045 $X2=7.17
+ $Y2=1.045
r88 20 47 1.91462 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=7.01 $Y=0.96 $X2=7.01
+ $Y2=1.07
r89 20 22 27.4192 $w=1.78e-07 $l=4.45e-07 $layer=LI1_cond $X=7.01 $Y=0.96
+ $X2=7.01 $Y2=0.515
r90 19 45 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.215 $Y=1.095
+ $X2=6.09 $Y2=1.095
r91 19 48 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.215 $Y=1.095
+ $X2=6.92 $Y2=1.095
r92 17 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=1.045
+ $X2=5.27 $Y2=1.045
r93 16 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.965 $Y=1.045
+ $X2=6.09 $Y2=1.045
r94 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.965 $Y=1.045
+ $X2=5.435 $Y2=1.045
r95 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r96 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.725
+ $Y=0.37 $X2=7.865 $Y2=0.515
r97 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.865
+ $Y=0.37 $X2=7.005 $Y2=0.515
r98 2 42 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.37 $X2=6.13 $Y2=0.95
r99 1 37 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.79 $X2=5.27 $Y2=0.95
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__inv_4 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.296e+11p ps=8.38e+06u
M1001 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=6.882e+11p pd=6.3e+06u as=4.44e+11p ps=4.16e+06u
M1003 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__einvp_1.pex.spice
* Created: Wed Sep  2 12:08:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EINVP_1%A_44_549# 1 2 9 11 13 15 16 18 21 24 26
r44 24 26 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.725 $Y=2.965
+ $X2=0.89 $Y2=2.965
r45 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=2.91 $X2=0.725 $Y2=2.91
r46 21 23 11.5257 $w=7.78e-07 $l=7.35e-07 $layer=LI1_cond $X=0.497 $Y=2.175
+ $X2=0.497 $Y2=2.91
r47 16 18 9.84465 $w=6.48e-07 $l=5.35e-07 $layer=LI1_cond $X=0.275 $Y=0.735
+ $X2=0.81 $Y2=0.735
r48 15 21 11.524 $w=7.78e-07 $l=3.80663e-07 $layer=LI1_cond $X=0.19 $Y=2.01
+ $X2=0.497 $Y2=2.175
r49 14 16 10.4312 $w=6.5e-07 $l=3.65034e-07 $layer=LI1_cond $X=0.19 $Y=1.06
+ $X2=0.275 $Y2=0.735
r50 14 15 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=0.19 $Y=1.06
+ $X2=0.19 $Y2=2.01
r51 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.475 $Y=3.035
+ $X2=1.475 $Y2=2.46
r52 9 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.385 $Y=3.11
+ $X2=1.475 $Y2=3.035
r53 9 26 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.385 $Y=3.11
+ $X2=0.89 $Y2=3.11
r54 2 21 300 $w=1.7e-07 $l=5.77581e-07 $layer=licon1_PDIFF $count=2 $X=0.235
+ $Y=1.96 $X2=0.715 $Y2=2.175
r55 1 18 91 $w=1.7e-07 $l=5.73411e-07 $layer=licon1_NDIFF $count=2 $X=0.33
+ $Y=0.37 $X2=0.81 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_1%TE 3 7 9 13 15 16 19 25
r46 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.605 $X2=0.95 $Y2=1.605
r47 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.605 $X2=0.61 $Y2=1.605
r48 19 25 7.86782 $w=3.3e-07 $l=1.32e-07 $layer=POLY_cond $X=0.85 $Y=1.605
+ $X2=0.982 $Y2=1.605
r49 19 21 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.85 $Y=1.605
+ $X2=0.61 $Y2=1.605
r50 16 26 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.61 $X2=0.95
+ $Y2=1.61
r51 15 26 7.79594 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.61
+ $X2=0.95 $Y2=1.61
r52 15 22 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.61
+ $X2=0.61 $Y2=1.61
r53 11 13 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=1.515 $Y=1.44
+ $X2=1.515 $Y2=0.74
r54 10 25 7.86782 $w=1.5e-07 $l=1.72218e-07 $layer=POLY_cond $X=1.115 $Y=1.515
+ $X2=0.982 $Y2=1.605
r55 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.44 $Y=1.515
+ $X2=1.515 $Y2=1.44
r56 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.44 $Y=1.515
+ $X2=1.115 $Y2=1.515
r57 5 25 16.8416 $w=1.5e-07 $l=1.85257e-07 $layer=POLY_cond $X=1.025 $Y=1.44
+ $X2=0.982 $Y2=1.605
r58 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.025 $Y=1.44
+ $X2=1.025 $Y2=0.58
r59 1 25 16.8416 $w=1.8e-07 $l=1.84811e-07 $layer=POLY_cond $X=0.94 $Y=1.77
+ $X2=0.982 $Y2=1.605
r60 1 3 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=0.94 $Y=1.77 $X2=0.94
+ $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_1%A 1 3 6 10 11 17 18
r27 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.465 $X2=2.11 $Y2=1.465
r28 15 17 35.4968 $w=3.3e-07 $l=2.03e-07 $layer=POLY_cond $X=1.907 $Y=1.465
+ $X2=2.11 $Y2=1.465
r29 13 15 0.349723 $w=3.3e-07 $l=2e-09 $layer=POLY_cond $X=1.905 $Y=1.465
+ $X2=1.907 $Y2=1.465
r30 11 18 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.11 $Y=1.665 $X2=2.11
+ $Y2=1.465
r31 8 15 20.5173 $w=1.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.907 $Y=1.63
+ $X2=1.907 $Y2=1.465
r32 8 10 95.6824 $w=1.55e-07 $l=2e-07 $layer=POLY_cond $X=1.907 $Y=1.63
+ $X2=1.907 $Y2=1.83
r33 4 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.3
+ $X2=1.905 $Y2=1.465
r34 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.905 $Y=1.3 $X2=1.905
+ $Y2=0.74
r35 1 10 36.5274 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.895 $Y=1.92 $X2=1.895
+ $Y2=1.83
r36 1 3 144.6 $w=1.8e-07 $l=5.4e-07 $layer=POLY_cond $X=1.895 $Y=1.92 $X2=1.895
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_1%VPWR 1 6 10 12 19 20 23
r28 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=3.33
+ $X2=1.25 $Y2=3.33
r30 17 19 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.415 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.25 $Y2=3.33
r33 12 14 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 10 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r37 6 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.25 $Y=2.105
+ $X2=1.25 $Y2=2.46
r38 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=3.245 $X2=1.25
+ $Y2=3.33
r39 4 9 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=1.25 $Y=3.245
+ $X2=1.25 $Y2=2.46
r40 1 9 300 $w=1.7e-07 $l=6e-07 $layer=licon1_PDIFF $count=2 $X=1.03 $Y=1.96
+ $X2=1.25 $Y2=2.46
r41 1 6 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.96 $X2=1.25 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_1%Z 1 2 8 9 10 13 18 21 22
c35 10 0 1.4658e-19 $X=1.775 $Y=1.045
r36 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=2.405
+ $X2=2.12 $Y2=2.775
r37 19 21 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.12 $Y=2.275
+ $X2=2.12 $Y2=2.405
r38 18 19 0.623162 $w=3.3e-07 $l=1.63e-07 $layer=LI1_cond $X=2.12 $Y=2.112
+ $X2=2.12 $Y2=2.275
r39 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.12 $Y=0.96
+ $X2=2.12 $Y2=0.515
r40 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.955 $Y=1.045
+ $X2=2.12 $Y2=0.96
r41 9 10 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.955 $Y=1.045
+ $X2=1.775 $Y2=1.045
r42 8 18 15.2477 $w=3.23e-07 $l=4.3e-07 $layer=LI1_cond $X=1.69 $Y=2.112
+ $X2=2.12 $Y2=2.112
r43 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.69 $Y=1.13
+ $X2=1.775 $Y2=1.045
r44 7 8 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.69 $Y=1.13 $X2=1.69
+ $Y2=1.95
r45 2 22 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.96 $X2=2.12 $Y2=2.815
r46 2 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.96 $X2=2.12 $Y2=2.115
r47 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.37 $X2=2.12 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_1%VGND 1 6 10 12 19 20 23
r25 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r26 17 23 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.277
+ $Y2=0
r27 17 19 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=2.16
+ $Y2=0
r28 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 12 23 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.277
+ $Y2=0
r30 12 14 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.24
+ $Y2=0
r31 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r32 10 15 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r33 10 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r34 6 8 18.1965 $w=2.83e-07 $l=4.5e-07 $layer=LI1_cond $X=1.277 $Y=0.515
+ $X2=1.277 $Y2=0.965
r35 4 23 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.277 $Y=0.085
+ $X2=1.277 $Y2=0
r36 4 6 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=1.277 $Y=0.085
+ $X2=1.277 $Y2=0.515
r37 1 8 182 $w=1.7e-07 $l=6.87768e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.37 $X2=1.3 $Y2=0.965
r38 1 6 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.37 $X2=1.3 $Y2=0.515
.ends


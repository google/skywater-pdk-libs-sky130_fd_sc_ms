* File: sky130_fd_sc_ms__dfrbp_1.pxi.spice
* Created: Wed Sep  2 12:02:43 2020
* 
x_PM_SKY130_FD_SC_MS__DFRBP_1%D N_D_M1023_g N_D_M1010_g N_D_c_241_n D D D
+ N_D_c_237_n N_D_c_238_n N_D_c_239_n PM_SKY130_FD_SC_MS__DFRBP_1%D
x_PM_SKY130_FD_SC_MS__DFRBP_1%CLK N_CLK_M1006_g N_CLK_M1011_g CLK N_CLK_c_270_n
+ N_CLK_c_271_n PM_SKY130_FD_SC_MS__DFRBP_1%CLK
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_501_387# N_A_501_387#_M1012_d
+ N_A_501_387#_M1014_d N_A_501_387#_M1005_g N_A_501_387#_c_331_n
+ N_A_501_387#_c_315_n N_A_501_387#_c_316_n N_A_501_387#_M1017_g
+ N_A_501_387#_c_317_n N_A_501_387#_M1003_g N_A_501_387#_c_318_n
+ N_A_501_387#_c_319_n N_A_501_387#_M1033_g N_A_501_387#_c_320_n
+ N_A_501_387#_c_339_n N_A_501_387#_c_321_n N_A_501_387#_c_322_n
+ N_A_501_387#_c_323_n N_A_501_387#_c_324_n N_A_501_387#_c_345_p
+ N_A_501_387#_c_388_p N_A_501_387#_c_325_n N_A_501_387#_c_358_p
+ N_A_501_387#_c_326_n N_A_501_387#_c_327_n N_A_501_387#_c_369_p
+ N_A_501_387#_c_335_n N_A_501_387#_c_336_n N_A_501_387#_c_328_n
+ N_A_501_387#_c_329_n N_A_501_387#_c_338_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_501_387#
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_841_401# N_A_841_401#_M1002_d
+ N_A_841_401#_M1016_d N_A_841_401#_M1028_g N_A_841_401#_M1001_g
+ N_A_841_401#_c_529_n N_A_841_401#_c_530_n N_A_841_401#_c_520_n
+ N_A_841_401#_c_521_n N_A_841_401#_c_522_n N_A_841_401#_c_523_n
+ N_A_841_401#_c_524_n N_A_841_401#_c_525_n N_A_841_401#_c_526_n
+ N_A_841_401#_c_527_n N_A_841_401#_c_534_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_841_401#
x_PM_SKY130_FD_SC_MS__DFRBP_1%RESET_B N_RESET_B_M1029_g N_RESET_B_c_630_n
+ N_RESET_B_M1024_g N_RESET_B_c_631_n N_RESET_B_c_632_n N_RESET_B_M1019_g
+ N_RESET_B_c_634_n N_RESET_B_M1031_g N_RESET_B_M1026_g N_RESET_B_M1021_g
+ N_RESET_B_c_636_n N_RESET_B_c_645_n N_RESET_B_c_646_n N_RESET_B_c_647_n
+ N_RESET_B_c_648_n N_RESET_B_c_649_n N_RESET_B_c_650_n RESET_B
+ N_RESET_B_c_651_n N_RESET_B_c_652_n N_RESET_B_c_637_n N_RESET_B_c_638_n
+ N_RESET_B_c_654_n N_RESET_B_c_655_n N_RESET_B_c_656_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%RESET_B
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_709_463# N_A_709_463#_M1018_d
+ N_A_709_463#_M1005_d N_A_709_463#_M1031_d N_A_709_463#_M1002_g
+ N_A_709_463#_c_841_n N_A_709_463#_c_847_n N_A_709_463#_M1016_g
+ N_A_709_463#_c_842_n N_A_709_463#_c_880_n N_A_709_463#_c_849_n
+ N_A_709_463#_c_843_n N_A_709_463#_c_850_n N_A_709_463#_c_851_n
+ N_A_709_463#_c_844_n N_A_709_463#_c_845_n N_A_709_463#_c_853_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_709_463#
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_307_387# N_A_307_387#_M1011_s
+ N_A_307_387#_M1006_s N_A_307_387#_M1014_g N_A_307_387#_c_967_n
+ N_A_307_387#_M1012_g N_A_307_387#_c_978_n N_A_307_387#_c_979_n
+ N_A_307_387#_c_980_n N_A_307_387#_c_981_n N_A_307_387#_c_968_n
+ N_A_307_387#_c_969_n N_A_307_387#_M1018_g N_A_307_387#_M1009_g
+ N_A_307_387#_c_984_n N_A_307_387#_M1020_g N_A_307_387#_c_971_n
+ N_A_307_387#_c_972_n N_A_307_387#_M1000_g N_A_307_387#_c_988_n
+ N_A_307_387#_c_989_n N_A_307_387#_c_974_n N_A_307_387#_c_1004_n
+ N_A_307_387#_c_975_n N_A_307_387#_c_976_n N_A_307_387#_c_992_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_307_387#
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_1482_48# N_A_1482_48#_M1027_d
+ N_A_1482_48#_M1021_d N_A_1482_48#_c_1156_n N_A_1482_48#_M1022_g
+ N_A_1482_48#_M1007_g N_A_1482_48#_c_1158_n N_A_1482_48#_c_1165_n
+ N_A_1482_48#_c_1159_n N_A_1482_48#_c_1160_n N_A_1482_48#_c_1161_n
+ N_A_1482_48#_c_1167_n N_A_1482_48#_c_1162_n N_A_1482_48#_c_1163_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_1482_48#
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_1224_74# N_A_1224_74#_M1003_d
+ N_A_1224_74#_M1020_d N_A_1224_74#_M1027_g N_A_1224_74#_M1025_g
+ N_A_1224_74#_c_1251_n N_A_1224_74#_c_1252_n N_A_1224_74#_M1008_g
+ N_A_1224_74#_M1015_g N_A_1224_74#_c_1255_n N_A_1224_74#_c_1256_n
+ N_A_1224_74#_M1030_g N_A_1224_74#_M1013_g N_A_1224_74#_c_1259_n
+ N_A_1224_74#_c_1277_n N_A_1224_74#_c_1281_n N_A_1224_74#_c_1260_n
+ N_A_1224_74#_c_1261_n N_A_1224_74#_c_1262_n N_A_1224_74#_c_1263_n
+ N_A_1224_74#_c_1264_n N_A_1224_74#_c_1265_n N_A_1224_74#_c_1266_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_1224_74#
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_2026_424# N_A_2026_424#_M1013_s
+ N_A_2026_424#_M1030_s N_A_2026_424#_M1032_g N_A_2026_424#_M1004_g
+ N_A_2026_424#_c_1410_n N_A_2026_424#_c_1411_n N_A_2026_424#_c_1412_n
+ N_A_2026_424#_c_1413_n N_A_2026_424#_c_1414_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_2026_424#
x_PM_SKY130_FD_SC_MS__DFRBP_1%VPWR N_VPWR_M1023_s N_VPWR_M1024_d N_VPWR_M1006_d
+ N_VPWR_M1028_d N_VPWR_M1016_s N_VPWR_M1007_d N_VPWR_M1025_d N_VPWR_M1030_d
+ N_VPWR_c_1461_n N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n
+ N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n N_VPWR_c_1468_n
+ N_VPWR_c_1469_n N_VPWR_c_1470_n VPWR N_VPWR_c_1471_n N_VPWR_c_1472_n
+ N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n N_VPWR_c_1476_n
+ N_VPWR_c_1477_n N_VPWR_c_1460_n N_VPWR_c_1479_n N_VPWR_c_1480_n
+ N_VPWR_c_1481_n N_VPWR_c_1482_n N_VPWR_c_1483_n N_VPWR_c_1484_n
+ N_VPWR_c_1485_n PM_SKY130_FD_SC_MS__DFRBP_1%VPWR
x_PM_SKY130_FD_SC_MS__DFRBP_1%A_38_78# N_A_38_78#_M1010_s N_A_38_78#_M1018_s
+ N_A_38_78#_M1023_d N_A_38_78#_M1005_s N_A_38_78#_c_1606_n N_A_38_78#_c_1612_n
+ N_A_38_78#_c_1607_n N_A_38_78#_c_1614_n N_A_38_78#_c_1608_n
+ N_A_38_78#_c_1615_n N_A_38_78#_c_1609_n N_A_38_78#_c_1610_n
+ N_A_38_78#_c_1617_n N_A_38_78#_c_1618_n N_A_38_78#_c_1611_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%A_38_78#
x_PM_SKY130_FD_SC_MS__DFRBP_1%Q_N N_Q_N_M1015_d N_Q_N_M1008_d N_Q_N_c_1727_n Q_N
+ Q_N Q_N N_Q_N_c_1730_n PM_SKY130_FD_SC_MS__DFRBP_1%Q_N
x_PM_SKY130_FD_SC_MS__DFRBP_1%Q N_Q_M1004_d N_Q_M1032_d Q Q Q Q Q N_Q_c_1753_n
+ PM_SKY130_FD_SC_MS__DFRBP_1%Q
x_PM_SKY130_FD_SC_MS__DFRBP_1%VGND N_VGND_M1029_d N_VGND_M1011_d N_VGND_M1019_d
+ N_VGND_M1022_d N_VGND_M1015_s N_VGND_M1013_d N_VGND_c_1776_n N_VGND_c_1777_n
+ N_VGND_c_1778_n N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n VGND
+ N_VGND_c_1782_n N_VGND_c_1783_n N_VGND_c_1784_n N_VGND_c_1785_n
+ N_VGND_c_1786_n N_VGND_c_1787_n N_VGND_c_1788_n N_VGND_c_1789_n
+ N_VGND_c_1790_n N_VGND_c_1791_n N_VGND_c_1792_n N_VGND_c_1793_n
+ N_VGND_c_1794_n PM_SKY130_FD_SC_MS__DFRBP_1%VGND
cc_1 VNB N_D_M1010_g 0.0286427f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_2 VNB N_D_c_237_n 0.0408539f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_3 VNB N_D_c_238_n 0.0253354f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_239_n 0.0298264f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB CLK 0.00333416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_CLK_c_270_n 0.0268106f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_CLK_c_271_n 0.0167256f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_8 VNB N_A_501_387#_c_315_n 0.0184472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_501_387#_c_316_n 0.0133409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_501_387#_c_317_n 0.0205313f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.845
cc_11 VNB N_A_501_387#_c_318_n 0.0187502f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_12 VNB N_A_501_387#_c_319_n 0.00880336f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_13 VNB N_A_501_387#_c_320_n 0.0144169f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.665
cc_14 VNB N_A_501_387#_c_321_n 0.0080788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_501_387#_c_322_n 0.0348154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_501_387#_c_323_n 0.00285435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_501_387#_c_324_n 0.0030846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_501_387#_c_325_n 0.00621215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_501_387#_c_326_n 0.0316981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_501_387#_c_327_n 0.00782104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_501_387#_c_328_n 0.0160337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_501_387#_c_329_n 0.00342169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_841_401#_M1001_g 0.0273166f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_24 VNB N_A_841_401#_c_520_n 0.00632677f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_25 VNB N_A_841_401#_c_521_n 0.015896f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_26 VNB N_A_841_401#_c_522_n 0.0106545f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_27 VNB N_A_841_401#_c_523_n 4.52231e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_841_401#_c_524_n 4.96212e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_29 VNB N_A_841_401#_c_525_n 0.00934369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_841_401#_c_526_n 0.00496873f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.665
cc_31 VNB N_A_841_401#_c_527_n 4.11682e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_M1029_g 0.0222805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_630_n 0.027732f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_34 VNB N_RESET_B_c_631_n 0.284514f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_RESET_B_c_632_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_RESET_B_M1019_g 0.0240189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_RESET_B_c_634_n 0.0186427f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.845
cc_38 VNB N_RESET_B_M1026_g 0.0515393f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_39 VNB N_RESET_B_c_636_n 0.0133121f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=2.035
cc_40 VNB N_RESET_B_c_637_n 0.0324691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_638_n 0.00371377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_709_463#_M1002_g 0.0297973f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_43 VNB N_A_709_463#_c_841_n 0.0206976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_709_463#_c_842_n 0.00364311f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_45 VNB N_A_709_463#_c_843_n 0.00339134f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=2.035
cc_46 VNB N_A_709_463#_c_844_n 0.0104779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_709_463#_c_845_n 0.0286964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_307_387#_c_967_n 0.0140603f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_49 VNB N_A_307_387#_c_968_n 0.0361443f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_50 VNB N_A_307_387#_c_969_n 0.0601446f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_51 VNB N_A_307_387#_M1018_g 0.029487f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_52 VNB N_A_307_387#_c_971_n 0.021569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_307_387#_c_972_n 0.00564393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_307_387#_M1000_g 0.0529012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_307_387#_c_974_n 0.00932233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_307_387#_c_975_n 4.69816e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_307_387#_c_976_n 0.0128049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1482_48#_c_1156_n 0.0177983f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_59 VNB N_A_1482_48#_M1007_g 0.0233363f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_60 VNB N_A_1482_48#_c_1158_n 0.0157083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1482_48#_c_1159_n 0.0117659f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_62 VNB N_A_1482_48#_c_1160_n 0.00518085f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_63 VNB N_A_1482_48#_c_1161_n 0.00346875f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_64 VNB N_A_1482_48#_c_1162_n 0.00600532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1482_48#_c_1163_n 0.0330587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1224_74#_M1027_g 0.0408739f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=2.148
cc_67 VNB N_A_1224_74#_M1025_g 0.00400132f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_68 VNB N_A_1224_74#_c_1251_n 0.0275488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1224_74#_c_1252_n 0.0281282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1224_74#_M1008_g 0.00407025f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_71 VNB N_A_1224_74#_M1015_g 0.0260029f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_72 VNB N_A_1224_74#_c_1255_n 0.0862945f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.165
cc_73 VNB N_A_1224_74#_c_1256_n 0.0294141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1224_74#_M1030_g 0.00400127f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.665
cc_75 VNB N_A_1224_74#_M1013_g 0.0355065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1224_74#_c_1259_n 0.0100839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1224_74#_c_1260_n 0.00749917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1224_74#_c_1261_n 0.0120508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1224_74#_c_1262_n 4.69525e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1224_74#_c_1263_n 9.056e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1224_74#_c_1264_n 0.00965329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1224_74#_c_1265_n 5.50055e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1224_74#_c_1266_n 0.00638783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2026_424#_M1032_g 0.00182491f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=2.148
cc_85 VNB N_A_2026_424#_M1004_g 0.0282052f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_86 VNB N_A_2026_424#_c_1410_n 0.00968545f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.202
cc_87 VNB N_A_2026_424#_c_1411_n 3.04122e-19 $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.165
cc_88 VNB N_A_2026_424#_c_1412_n 0.00611923f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.165
cc_89 VNB N_A_2026_424#_c_1413_n 0.0326263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2026_424#_c_1414_n 3.73161e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VPWR_c_1460_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_38_78#_c_1606_n 0.00234225f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_93 VNB N_A_38_78#_c_1607_n 0.0151458f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_94 VNB N_A_38_78#_c_1608_n 0.00307546f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_95 VNB N_A_38_78#_c_1609_n 0.00436775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_38_78#_c_1610_n 0.0222631f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=2.035
cc_97 VNB N_A_38_78#_c_1611_n 0.00579702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_Q_N_c_1727_n 0.0157896f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=2.148
cc_99 VNB Q 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=2.148
cc_100 VNB Q 0.0133985f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=2.35
cc_101 VNB N_Q_c_1753_n 0.0249693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1776_n 0.0094037f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_103 VNB N_VGND_c_1777_n 0.0212452f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_104 VNB N_VGND_c_1778_n 0.0140056f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.295
cc_105 VNB N_VGND_c_1779_n 0.00450041f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.845
cc_106 VNB N_VGND_c_1780_n 0.00944343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1781_n 0.0125104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1782_n 0.0298733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1783_n 0.0603649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1784_n 0.0603291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1785_n 0.0324414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1786_n 0.0347338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1787_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1788_n 0.609762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1789_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1790_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1791_n 0.0146905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1792_n 0.00846888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1793_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1794_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VPB N_D_M1023_g 0.0293003f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_122 VPB N_D_c_241_n 0.0290412f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.35
cc_123 VPB N_D_c_237_n 0.0435358f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_124 VPB N_D_c_239_n 0.0215212f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_125 VPB N_CLK_M1006_g 0.0245998f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_126 VPB CLK 0.00361254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_CLK_c_270_n 0.00558015f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_128 VPB N_A_501_387#_M1005_g 0.027706f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_129 VPB N_A_501_387#_c_331_n 0.0293884f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_130 VPB N_A_501_387#_c_315_n 0.00315483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_501_387#_M1033_g 0.0238251f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.165
cc_132 VPB N_A_501_387#_c_327_n 0.00248282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_501_387#_c_335_n 0.00306084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_501_387#_c_336_n 0.0335342f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_501_387#_c_329_n 0.00641707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_501_387#_c_338_n 0.0284935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_841_401#_M1028_g 0.0207228f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_138 VPB N_A_841_401#_c_529_n 0.0263237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_841_401#_c_530_n 0.0227906f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.202
cc_140 VPB N_A_841_401#_c_520_n 0.0026876f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_141 VPB N_A_841_401#_c_521_n 0.00209419f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_142 VPB N_A_841_401#_c_526_n 6.92353e-19 $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_143 VPB N_A_841_401#_c_534_n 0.00384768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_RESET_B_c_630_n 0.0231417f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=0.6
cc_145 VPB N_RESET_B_M1024_g 0.0431289f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_146 VPB N_RESET_B_c_634_n 0.0124021f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_147 VPB N_RESET_B_M1031_g 0.0265076f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_148 VPB N_RESET_B_M1026_g 0.00974243f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.165
cc_149 VPB N_RESET_B_M1021_g 0.0238799f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_150 VPB N_RESET_B_c_645_n 0.0118975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_646_n 0.0273404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_647_n 0.00357281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_648_n 0.00537181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_649_n 0.00350644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_650_n 0.00338092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_651_n 0.0553452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_652_n 0.00382655f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_638_n 0.0013565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_654_n 0.029069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_655_n 0.0283066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_656_n 0.00608672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_709_463#_c_841_n 0.0166935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_709_463#_c_847_n 0.0216635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_709_463#_c_842_n 0.00815884f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1
cc_165 VPB N_A_709_463#_c_849_n 0.0104778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_709_463#_c_850_n 0.00267689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_709_463#_c_851_n 0.00186798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_709_463#_c_845_n 3.30851e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_709_463#_c_853_n 0.0048438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_307_387#_M1014_g 0.0214992f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_171 VPB N_A_307_387#_c_978_n 0.0155044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_307_387#_c_979_n 0.0539717f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.202
cc_173 VPB N_A_307_387#_c_980_n 0.0543388f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_174 VPB N_A_307_387#_c_981_n 0.0106868f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_175 VPB N_A_307_387#_c_969_n 0.00926023f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_176 VPB N_A_307_387#_M1009_g 0.0367627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_307_387#_c_984_n 0.198975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_307_387#_M1020_g 0.033067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_307_387#_c_971_n 0.0142262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_307_387#_c_972_n 0.00222638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_307_387#_c_988_n 0.00585309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_307_387#_c_989_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_307_387#_c_974_n 0.00399383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_307_387#_c_975_n 5.38342e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_307_387#_c_992_n 0.00320568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1482_48#_M1007_g 0.0485488f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_187 VPB N_A_1482_48#_c_1165_n 0.0101134f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.202
cc_188 VPB N_A_1482_48#_c_1160_n 0.00239847f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_189 VPB N_A_1482_48#_c_1167_n 0.00856197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1224_74#_M1025_g 0.0488198f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_191 VPB N_A_1224_74#_M1008_g 0.0282965f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_192 VPB N_A_1224_74#_M1030_g 0.0485033f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_193 VPB N_A_1224_74#_c_1263_n 0.0065595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_2026_424#_M1032_g 0.02971f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_195 VPB N_A_2026_424#_c_1411_n 0.00739526f $X=-0.19 $Y=1.66 $X2=0.422
+ $Y2=1.165
cc_196 VPB N_VPWR_c_1461_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.165
cc_197 VPB N_VPWR_c_1462_n 0.0307031f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_198 VPB N_VPWR_c_1463_n 0.00980382f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.845
cc_199 VPB N_VPWR_c_1464_n 0.00151893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1465_n 0.013796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1466_n 0.0155908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1467_n 0.024939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1468_n 0.021993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1469_n 0.0118201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1470_n 0.0143569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1471_n 0.0176659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1472_n 0.0183973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1473_n 0.0561653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1474_n 0.0273297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1475_n 0.0507873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1476_n 0.0430282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1477_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1460_n 0.1162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1479_n 0.00612665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1480_n 0.00485616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1481_n 0.00456739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1482_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1483_n 0.00430193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1484_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1485_n 0.00564836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_38_78#_c_1612_n 0.00227613f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.202
cc_222 VPB N_A_38_78#_c_1607_n 0.013208f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_223 VPB N_A_38_78#_c_1614_n 0.0133682f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_224 VPB N_A_38_78#_c_1615_n 4.86504e-19 $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_225 VPB N_A_38_78#_c_1609_n 0.00544017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_38_78#_c_1617_n 0.0042266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_38_78#_c_1618_n 0.0069091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_Q_N_c_1727_n 0.00323428f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_229 VPB Q_N 0.0167637f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_230 VPB N_Q_N_c_1730_n 0.00887967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB Q 0.0129669f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_232 VPB Q 0.0415472f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_233 VPB N_Q_c_1753_n 0.00769959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 N_D_M1010_g N_RESET_B_M1029_g 0.0260656f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_235 N_D_c_237_n N_RESET_B_c_630_n 0.0260656f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_236 N_D_M1023_g N_RESET_B_M1024_g 0.015039f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_237 N_D_c_238_n N_RESET_B_c_637_n 0.0260656f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_238 N_D_c_241_n N_RESET_B_c_654_n 0.0260656f $X=0.422 $Y=2.35 $X2=0 $Y2=0
cc_239 N_D_M1023_g N_VPWR_c_1462_n 0.00477201f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_240 N_D_c_241_n N_VPWR_c_1462_n 0.0042702f $X=0.422 $Y=2.35 $X2=0 $Y2=0
cc_241 N_D_c_239_n N_VPWR_c_1462_n 0.013492f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_242 N_D_M1023_g N_VPWR_c_1463_n 4.10796e-19 $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_243 N_D_M1023_g N_VPWR_c_1471_n 0.005209f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_244 N_D_M1023_g N_VPWR_c_1460_n 0.00986118f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_245 N_D_M1010_g N_A_38_78#_c_1606_n 0.0116103f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_246 N_D_c_239_n N_A_38_78#_c_1606_n 0.00144733f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_247 N_D_M1023_g N_A_38_78#_c_1612_n 0.00504724f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_248 N_D_M1023_g N_A_38_78#_c_1607_n 0.00134086f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_249 N_D_M1010_g N_A_38_78#_c_1607_n 0.0162338f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_250 N_D_c_239_n N_A_38_78#_c_1607_n 0.0904243f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_251 N_D_M1010_g N_A_38_78#_c_1610_n 0.0078958f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_252 N_D_c_238_n N_A_38_78#_c_1610_n 0.00191909f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_253 N_D_c_239_n N_A_38_78#_c_1610_n 0.028486f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_254 N_D_M1023_g N_A_38_78#_c_1617_n 0.00647805f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_255 N_D_c_241_n N_A_38_78#_c_1617_n 0.00138105f $X=0.422 $Y=2.35 $X2=0 $Y2=0
cc_256 N_D_M1010_g N_VGND_c_1776_n 0.00200808f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_257 N_D_M1010_g N_VGND_c_1782_n 0.00429844f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_258 N_D_M1010_g N_VGND_c_1788_n 0.00539454f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_259 N_CLK_M1006_g N_A_501_387#_c_339_n 9.58624e-19 $X=1.965 $Y=2.495 $X2=0
+ $Y2=0
cc_260 N_CLK_M1006_g N_RESET_B_c_630_n 0.00673093f $X=1.965 $Y=2.495 $X2=0 $Y2=0
cc_261 N_CLK_c_270_n N_RESET_B_c_630_n 0.00657838f $X=1.95 $Y=1.61 $X2=0 $Y2=0
cc_262 N_CLK_c_271_n N_RESET_B_c_631_n 0.0104164f $X=1.95 $Y=1.445 $X2=0 $Y2=0
cc_263 N_CLK_M1006_g N_RESET_B_c_646_n 0.00660633f $X=1.965 $Y=2.495 $X2=0 $Y2=0
cc_264 CLK N_RESET_B_c_646_n 0.0137829f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_265 N_CLK_c_271_n N_RESET_B_c_637_n 0.0034015f $X=1.95 $Y=1.445 $X2=0 $Y2=0
cc_266 CLK N_A_307_387#_M1011_s 8.21782e-19 $X=2.075 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_267 N_CLK_M1006_g N_A_307_387#_M1014_g 0.0506875f $X=1.965 $Y=2.495 $X2=0
+ $Y2=0
cc_268 CLK N_A_307_387#_c_967_n 7.05815e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_269 N_CLK_c_271_n N_A_307_387#_c_967_n 0.018746f $X=1.95 $Y=1.445 $X2=0 $Y2=0
cc_270 CLK N_A_307_387#_c_969_n 0.00321782f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_271 N_CLK_c_270_n N_A_307_387#_c_969_n 0.0215666f $X=1.95 $Y=1.61 $X2=0 $Y2=0
cc_272 N_CLK_c_271_n N_A_307_387#_c_969_n 0.00174484f $X=1.95 $Y=1.445 $X2=0
+ $Y2=0
cc_273 N_CLK_M1006_g N_A_307_387#_c_974_n 0.00360983f $X=1.965 $Y=2.495 $X2=0
+ $Y2=0
cc_274 CLK N_A_307_387#_c_974_n 0.0367415f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_275 N_CLK_c_270_n N_A_307_387#_c_974_n 0.00286287f $X=1.95 $Y=1.61 $X2=0
+ $Y2=0
cc_276 N_CLK_c_271_n N_A_307_387#_c_974_n 0.00331779f $X=1.95 $Y=1.445 $X2=0
+ $Y2=0
cc_277 CLK N_A_307_387#_c_1004_n 0.0227258f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_278 N_CLK_c_271_n N_A_307_387#_c_1004_n 0.0129975f $X=1.95 $Y=1.445 $X2=0
+ $Y2=0
cc_279 CLK N_A_307_387#_c_975_n 0.0347423f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_280 N_CLK_c_270_n N_A_307_387#_c_975_n 2.53025e-19 $X=1.95 $Y=1.61 $X2=0
+ $Y2=0
cc_281 N_CLK_c_271_n N_A_307_387#_c_975_n 0.00110951f $X=1.95 $Y=1.445 $X2=0
+ $Y2=0
cc_282 CLK N_A_307_387#_c_976_n 0.00459781f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_283 N_CLK_c_270_n N_A_307_387#_c_976_n 0.00142041f $X=1.95 $Y=1.61 $X2=0
+ $Y2=0
cc_284 N_CLK_c_271_n N_A_307_387#_c_976_n 0.00106778f $X=1.95 $Y=1.445 $X2=0
+ $Y2=0
cc_285 N_CLK_M1006_g N_A_307_387#_c_992_n 0.00389597f $X=1.965 $Y=2.495 $X2=0
+ $Y2=0
cc_286 CLK N_A_307_387#_c_992_n 8.05762e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_287 N_CLK_c_270_n N_A_307_387#_c_992_n 0.00109063f $X=1.95 $Y=1.61 $X2=0
+ $Y2=0
cc_288 N_CLK_M1006_g N_VPWR_c_1463_n 0.0102098f $X=1.965 $Y=2.495 $X2=0 $Y2=0
cc_289 N_CLK_M1006_g N_VPWR_c_1464_n 0.0197454f $X=1.965 $Y=2.495 $X2=0 $Y2=0
cc_290 N_CLK_M1006_g N_VPWR_c_1472_n 0.00406785f $X=1.965 $Y=2.495 $X2=0 $Y2=0
cc_291 N_CLK_M1006_g N_VPWR_c_1460_n 0.00600562f $X=1.965 $Y=2.495 $X2=0 $Y2=0
cc_292 N_CLK_M1006_g N_A_38_78#_c_1614_n 0.0177428f $X=1.965 $Y=2.495 $X2=0
+ $Y2=0
cc_293 CLK N_A_38_78#_c_1614_n 0.0043091f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_294 N_CLK_c_270_n N_A_38_78#_c_1614_n 2.17013e-19 $X=1.95 $Y=1.61 $X2=0 $Y2=0
cc_295 CLK N_VGND_M1011_d 0.00183836f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_296 N_CLK_c_271_n N_VGND_c_1776_n 0.00219535f $X=1.95 $Y=1.445 $X2=0 $Y2=0
cc_297 N_CLK_c_271_n N_VGND_c_1778_n 0.00292425f $X=1.95 $Y=1.445 $X2=0 $Y2=0
cc_298 N_CLK_c_271_n N_VGND_c_1788_n 9.39239e-19 $X=1.95 $Y=1.445 $X2=0 $Y2=0
cc_299 N_A_501_387#_c_324_n N_A_841_401#_M1002_d 0.0095109f $X=6.085 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_300 N_A_501_387#_c_315_n N_A_841_401#_M1001_g 0.00801556f $X=3.975 $Y=1.685
+ $X2=0 $Y2=0
cc_301 N_A_501_387#_c_316_n N_A_841_401#_M1001_g 0.0411627f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_302 N_A_501_387#_c_323_n N_A_841_401#_M1001_g 0.00423512f $X=4.435 $Y=0.58
+ $X2=0 $Y2=0
cc_303 N_A_501_387#_c_324_n N_A_841_401#_M1001_g 0.00295293f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_304 N_A_501_387#_c_345_p N_A_841_401#_M1001_g 0.00422261f $X=4.52 $Y=0.665
+ $X2=0 $Y2=0
cc_305 N_A_501_387#_c_331_n N_A_841_401#_c_529_n 0.00864733f $X=3.9 $Y=1.76
+ $X2=0 $Y2=0
cc_306 N_A_501_387#_c_338_n N_A_841_401#_c_529_n 0.00171866f $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_307 N_A_501_387#_M1005_g N_A_841_401#_c_530_n 0.00227686f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_308 N_A_501_387#_c_315_n N_A_841_401#_c_520_n 9.63391e-19 $X=3.975 $Y=1.685
+ $X2=0 $Y2=0
cc_309 N_A_501_387#_c_316_n N_A_841_401#_c_520_n 4.83625e-19 $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_310 N_A_501_387#_c_315_n N_A_841_401#_c_521_n 0.00864733f $X=3.975 $Y=1.685
+ $X2=0 $Y2=0
cc_311 N_A_501_387#_c_324_n N_A_841_401#_c_522_n 0.0628972f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_312 N_A_501_387#_c_316_n N_A_841_401#_c_523_n 3.4688e-19 $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_313 N_A_501_387#_c_324_n N_A_841_401#_c_523_n 0.00412245f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_314 N_A_501_387#_c_345_p N_A_841_401#_c_523_n 0.00983586f $X=4.52 $Y=0.665
+ $X2=0 $Y2=0
cc_315 N_A_501_387#_c_317_n N_A_841_401#_c_524_n 0.00136384f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_316 N_A_501_387#_c_324_n N_A_841_401#_c_524_n 0.0136179f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_317 N_A_501_387#_c_358_p N_A_841_401#_c_524_n 0.0108515f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_318 N_A_501_387#_c_319_n N_A_841_401#_c_525_n 0.00176493f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_319 N_A_501_387#_c_358_p N_A_841_401#_c_525_n 0.011149f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_320 N_A_501_387#_c_318_n N_A_841_401#_c_526_n 0.00507154f $X=6.48 $Y=1.16
+ $X2=0 $Y2=0
cc_321 N_A_501_387#_c_319_n N_A_841_401#_c_526_n 0.00303743f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_322 N_A_501_387#_c_324_n N_A_841_401#_c_526_n 0.00373373f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_323 N_A_501_387#_c_325_n N_A_841_401#_c_526_n 0.0188995f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_324 N_A_501_387#_c_358_p N_A_841_401#_c_526_n 0.0136879f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_325 N_A_501_387#_c_327_n N_A_841_401#_c_526_n 0.0135711f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_326 N_A_501_387#_M1033_g N_A_841_401#_c_534_n 0.00118136f $X=7.25 $Y=2.565
+ $X2=0 $Y2=0
cc_327 N_A_501_387#_c_327_n N_A_841_401#_c_534_n 0.0165009f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_328 N_A_501_387#_c_369_p N_A_841_401#_c_534_n 0.0140459f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_329 N_A_501_387#_c_336_n N_A_841_401#_c_534_n 2.36915e-19 $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_330 N_A_501_387#_c_316_n N_RESET_B_c_631_n 0.00882199f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_331 N_A_501_387#_c_322_n N_RESET_B_c_631_n 0.0261266f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_332 N_A_501_387#_c_324_n N_RESET_B_c_631_n 0.00286781f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_333 N_A_501_387#_c_328_n N_RESET_B_c_631_n 0.0128673f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_334 N_A_501_387#_c_322_n N_RESET_B_M1019_g 0.00386847f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_335 N_A_501_387#_c_323_n N_RESET_B_M1019_g 0.00191339f $X=4.435 $Y=0.58 $X2=0
+ $Y2=0
cc_336 N_A_501_387#_c_324_n N_RESET_B_M1019_g 0.012028f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_337 N_A_501_387#_M1005_g N_RESET_B_c_646_n 0.00314802f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_338 N_A_501_387#_c_331_n N_RESET_B_c_646_n 0.00467871f $X=3.9 $Y=1.76 $X2=0
+ $Y2=0
cc_339 N_A_501_387#_c_339_n N_RESET_B_c_646_n 0.0173087f $X=2.79 $Y=2.092 $X2=0
+ $Y2=0
cc_340 N_A_501_387#_c_329_n N_RESET_B_c_646_n 0.0379446f $X=2.975 $Y=1.907 $X2=0
+ $Y2=0
cc_341 N_A_501_387#_c_338_n N_RESET_B_c_646_n 0.00307368f $X=3.415 $Y=1.76 $X2=0
+ $Y2=0
cc_342 N_A_501_387#_c_369_p N_RESET_B_c_648_n 0.0123453f $X=6.82 $Y=2.03 $X2=0
+ $Y2=0
cc_343 N_A_501_387#_c_335_n N_RESET_B_c_648_n 0.0237639f $X=7.205 $Y=2.03 $X2=0
+ $Y2=0
cc_344 N_A_501_387#_c_336_n N_RESET_B_c_648_n 0.00154682f $X=7.205 $Y=2.03 $X2=0
+ $Y2=0
cc_345 N_A_501_387#_c_317_n N_A_709_463#_M1002_g 0.0261676f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_346 N_A_501_387#_c_324_n N_A_709_463#_M1002_g 0.0128398f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_347 N_A_501_387#_c_388_p N_A_709_463#_M1002_g 6.89487e-19 $X=6.17 $Y=0.9
+ $X2=0 $Y2=0
cc_348 N_A_501_387#_c_358_p N_A_709_463#_M1002_g 2.33891e-19 $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_349 N_A_501_387#_c_319_n N_A_709_463#_c_841_n 0.0123545f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_350 N_A_501_387#_c_331_n N_A_709_463#_c_842_n 0.00443164f $X=3.9 $Y=1.76
+ $X2=0 $Y2=0
cc_351 N_A_501_387#_c_315_n N_A_709_463#_c_842_n 0.00824084f $X=3.975 $Y=1.685
+ $X2=0 $Y2=0
cc_352 N_A_501_387#_c_316_n N_A_709_463#_c_842_n 0.00267225f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_353 N_A_501_387#_c_320_n N_A_709_463#_c_842_n 0.00702274f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_354 N_A_501_387#_c_331_n N_A_709_463#_c_843_n 0.00139841f $X=3.9 $Y=1.76
+ $X2=0 $Y2=0
cc_355 N_A_501_387#_c_316_n N_A_709_463#_c_843_n 0.00935232f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_356 N_A_501_387#_c_320_n N_A_709_463#_c_843_n 0.00563475f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_357 N_A_501_387#_c_322_n N_A_709_463#_c_843_n 0.0317578f $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_358 N_A_501_387#_M1005_g N_A_709_463#_c_850_n 0.00358636f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_359 N_A_501_387#_c_331_n N_A_709_463#_c_850_n 9.97369e-19 $X=3.9 $Y=1.76
+ $X2=0 $Y2=0
cc_360 N_A_501_387#_c_339_n N_A_307_387#_M1014_g 0.00613716f $X=2.79 $Y=2.092
+ $X2=0 $Y2=0
cc_361 N_A_501_387#_c_329_n N_A_307_387#_M1014_g 0.00391236f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_362 N_A_501_387#_c_321_n N_A_307_387#_c_967_n 0.00628802f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_363 N_A_501_387#_c_328_n N_A_307_387#_c_967_n 0.00314869f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_364 N_A_501_387#_M1005_g N_A_307_387#_c_978_n 0.00717863f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_365 N_A_501_387#_c_329_n N_A_307_387#_c_978_n 0.0127792f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_366 N_A_501_387#_M1005_g N_A_307_387#_c_979_n 0.0147429f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_367 N_A_501_387#_c_329_n N_A_307_387#_c_979_n 0.00285922f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_368 N_A_501_387#_M1005_g N_A_307_387#_c_980_n 0.0123549f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_369 N_A_501_387#_c_315_n N_A_307_387#_c_968_n 0.00942526f $X=3.975 $Y=1.685
+ $X2=0 $Y2=0
cc_370 N_A_501_387#_c_321_n N_A_307_387#_c_968_n 0.00394216f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_371 N_A_501_387#_c_329_n N_A_307_387#_c_968_n 0.00797395f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_372 N_A_501_387#_c_338_n N_A_307_387#_c_968_n 0.0260091f $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_373 N_A_501_387#_c_339_n N_A_307_387#_c_969_n 0.00475343f $X=2.79 $Y=2.092
+ $X2=0 $Y2=0
cc_374 N_A_501_387#_c_321_n N_A_307_387#_c_969_n 0.0175761f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_375 N_A_501_387#_c_328_n N_A_307_387#_c_969_n 0.00502514f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_376 N_A_501_387#_c_329_n N_A_307_387#_c_969_n 0.0100104f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_377 N_A_501_387#_c_338_n N_A_307_387#_c_969_n 0.0213944f $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_378 N_A_501_387#_c_316_n N_A_307_387#_M1018_g 0.0130936f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_379 N_A_501_387#_c_320_n N_A_307_387#_M1018_g 0.00942526f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_380 N_A_501_387#_c_321_n N_A_307_387#_M1018_g 5.45786e-19 $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_381 N_A_501_387#_c_322_n N_A_307_387#_M1018_g 0.00330666f $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_382 N_A_501_387#_c_328_n N_A_307_387#_M1018_g 0.00566353f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_383 N_A_501_387#_M1005_g N_A_307_387#_M1009_g 0.0175989f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_384 N_A_501_387#_c_331_n N_A_307_387#_M1009_g 0.00737842f $X=3.9 $Y=1.76
+ $X2=0 $Y2=0
cc_385 N_A_501_387#_M1033_g N_A_307_387#_M1020_g 0.015094f $X=7.25 $Y=2.565
+ $X2=0 $Y2=0
cc_386 N_A_501_387#_c_327_n N_A_307_387#_M1020_g 0.00528684f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_387 N_A_501_387#_c_369_p N_A_307_387#_M1020_g 0.00225091f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_388 N_A_501_387#_c_336_n N_A_307_387#_M1020_g 0.00864999f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_389 N_A_501_387#_c_326_n N_A_307_387#_c_971_n 0.0104232f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_390 N_A_501_387#_c_327_n N_A_307_387#_c_971_n 0.0123591f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_391 N_A_501_387#_c_335_n N_A_307_387#_c_971_n 0.00746766f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_392 N_A_501_387#_c_336_n N_A_307_387#_c_971_n 0.0072253f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_393 N_A_501_387#_c_318_n N_A_307_387#_c_972_n 0.0104232f $X=6.48 $Y=1.16
+ $X2=0 $Y2=0
cc_394 N_A_501_387#_c_325_n N_A_307_387#_c_972_n 0.00127614f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_395 N_A_501_387#_c_325_n N_A_307_387#_M1000_g 0.00116888f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_396 N_A_501_387#_c_326_n N_A_307_387#_M1000_g 0.0216896f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_397 N_A_501_387#_c_327_n N_A_307_387#_M1000_g 0.00159607f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_398 N_A_501_387#_c_329_n N_A_307_387#_c_988_n 0.0035878f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_399 N_A_501_387#_M1012_d N_A_307_387#_c_1004_n 0.00202962f $X=2.59 $Y=0.595
+ $X2=0 $Y2=0
cc_400 N_A_501_387#_c_321_n N_A_307_387#_c_1004_n 0.0141569f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_401 N_A_501_387#_c_328_n N_A_307_387#_c_1004_n 0.00159777f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_402 N_A_501_387#_M1012_d N_A_307_387#_c_975_n 0.00205254f $X=2.59 $Y=0.595
+ $X2=0 $Y2=0
cc_403 N_A_501_387#_c_339_n N_A_307_387#_c_975_n 0.0117158f $X=2.79 $Y=2.092
+ $X2=0 $Y2=0
cc_404 N_A_501_387#_c_321_n N_A_307_387#_c_975_n 0.0327513f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_405 N_A_501_387#_c_329_n N_A_307_387#_c_975_n 0.0154085f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_406 N_A_501_387#_c_339_n N_A_307_387#_c_992_n 0.00319803f $X=2.79 $Y=2.092
+ $X2=0 $Y2=0
cc_407 N_A_501_387#_M1033_g N_A_1482_48#_M1007_g 0.0383523f $X=7.25 $Y=2.565
+ $X2=0 $Y2=0
cc_408 N_A_501_387#_c_335_n N_A_1482_48#_M1007_g 4.05738e-19 $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_409 N_A_501_387#_c_336_n N_A_1482_48#_M1007_g 0.0212445f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_410 N_A_501_387#_c_324_n N_A_1224_74#_M1003_d 0.00392413f $X=6.085 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_411 N_A_501_387#_c_388_p N_A_1224_74#_M1003_d 0.00564702f $X=6.17 $Y=0.9
+ $X2=-0.19 $Y2=-0.245
cc_412 N_A_501_387#_c_325_n N_A_1224_74#_M1003_d 0.00471261f $X=6.65 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_413 N_A_501_387#_c_327_n N_A_1224_74#_M1020_d 0.0031642f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_414 N_A_501_387#_c_369_p N_A_1224_74#_M1020_d 0.00433588f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_415 N_A_501_387#_c_335_n N_A_1224_74#_M1020_d 0.00213077f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_416 N_A_501_387#_c_317_n N_A_1224_74#_c_1277_n 0.00722906f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_417 N_A_501_387#_c_324_n N_A_1224_74#_c_1277_n 0.013434f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_418 N_A_501_387#_c_325_n N_A_1224_74#_c_1277_n 0.0317086f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_419 N_A_501_387#_c_326_n N_A_1224_74#_c_1277_n 0.00506999f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_420 N_A_501_387#_M1033_g N_A_1224_74#_c_1281_n 0.0203864f $X=7.25 $Y=2.565
+ $X2=0 $Y2=0
cc_421 N_A_501_387#_c_369_p N_A_1224_74#_c_1281_n 0.00944134f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_422 N_A_501_387#_c_335_n N_A_1224_74#_c_1281_n 0.0345717f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_423 N_A_501_387#_c_336_n N_A_1224_74#_c_1281_n 0.0025882f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_424 N_A_501_387#_c_325_n N_A_1224_74#_c_1260_n 0.0278616f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_425 N_A_501_387#_c_326_n N_A_1224_74#_c_1260_n 9.55385e-19 $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_426 N_A_501_387#_c_327_n N_A_1224_74#_c_1260_n 0.0146057f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_427 N_A_501_387#_c_335_n N_A_1224_74#_c_1261_n 0.00761315f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_428 N_A_501_387#_c_336_n N_A_1224_74#_c_1261_n 0.00540489f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_429 N_A_501_387#_c_327_n N_A_1224_74#_c_1262_n 0.0133634f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_430 N_A_501_387#_c_335_n N_A_1224_74#_c_1262_n 0.00832552f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_431 N_A_501_387#_c_336_n N_A_1224_74#_c_1262_n 4.21127e-19 $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_432 N_A_501_387#_M1033_g N_A_1224_74#_c_1263_n 0.00350579f $X=7.25 $Y=2.565
+ $X2=0 $Y2=0
cc_433 N_A_501_387#_c_327_n N_A_1224_74#_c_1263_n 0.00741853f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_434 N_A_501_387#_c_335_n N_A_1224_74#_c_1263_n 0.0242903f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_435 N_A_501_387#_c_336_n N_A_1224_74#_c_1263_n 0.00175366f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_436 N_A_501_387#_M1033_g N_VPWR_c_1475_n 0.0041957f $X=7.25 $Y=2.565 $X2=0
+ $Y2=0
cc_437 N_A_501_387#_M1005_g N_VPWR_c_1460_n 0.00112709f $X=3.455 $Y=2.525 $X2=0
+ $Y2=0
cc_438 N_A_501_387#_M1033_g N_VPWR_c_1460_n 0.00587053f $X=7.25 $Y=2.565 $X2=0
+ $Y2=0
cc_439 N_A_501_387#_M1014_d N_A_38_78#_c_1614_n 0.00648364f $X=2.505 $Y=1.935
+ $X2=0 $Y2=0
cc_440 N_A_501_387#_c_339_n N_A_38_78#_c_1614_n 0.0180737f $X=2.79 $Y=2.092
+ $X2=0 $Y2=0
cc_441 N_A_501_387#_c_329_n N_A_38_78#_c_1614_n 0.0159376f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_442 N_A_501_387#_c_316_n N_A_38_78#_c_1608_n 3.16057e-19 $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_443 N_A_501_387#_c_320_n N_A_38_78#_c_1608_n 3.23838e-19 $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_444 N_A_501_387#_c_322_n N_A_38_78#_c_1608_n 0.0167583f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_445 N_A_501_387#_c_328_n N_A_38_78#_c_1608_n 0.048924f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_446 N_A_501_387#_M1005_g N_A_38_78#_c_1615_n 0.0152845f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_447 N_A_501_387#_c_331_n N_A_38_78#_c_1615_n 0.00251615f $X=3.9 $Y=1.76 $X2=0
+ $Y2=0
cc_448 N_A_501_387#_c_329_n N_A_38_78#_c_1615_n 0.00927558f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_449 N_A_501_387#_c_338_n N_A_38_78#_c_1615_n 0.00126458f $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_450 N_A_501_387#_M1005_g N_A_38_78#_c_1609_n 0.00355401f $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_451 N_A_501_387#_c_331_n N_A_38_78#_c_1609_n 0.0133246f $X=3.9 $Y=1.76 $X2=0
+ $Y2=0
cc_452 N_A_501_387#_c_315_n N_A_38_78#_c_1609_n 0.00522878f $X=3.975 $Y=1.685
+ $X2=0 $Y2=0
cc_453 N_A_501_387#_c_321_n N_A_38_78#_c_1609_n 0.00659552f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_454 N_A_501_387#_c_329_n N_A_38_78#_c_1609_n 0.0350401f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_455 N_A_501_387#_c_338_n N_A_38_78#_c_1609_n 0.00214094f $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_456 N_A_501_387#_M1005_g N_A_38_78#_c_1618_n 2.86142e-19 $X=3.455 $Y=2.525
+ $X2=0 $Y2=0
cc_457 N_A_501_387#_c_329_n N_A_38_78#_c_1618_n 0.0212419f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_458 N_A_501_387#_c_338_n N_A_38_78#_c_1618_n 7.36959e-19 $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_459 N_A_501_387#_c_331_n N_A_38_78#_c_1611_n 8.86061e-19 $X=3.9 $Y=1.76 $X2=0
+ $Y2=0
cc_460 N_A_501_387#_c_320_n N_A_38_78#_c_1611_n 0.00123375f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_461 N_A_501_387#_c_321_n N_A_38_78#_c_1611_n 0.0140823f $X=2.975 $Y=1.575
+ $X2=0 $Y2=0
cc_462 N_A_501_387#_c_329_n N_A_38_78#_c_1611_n 0.0140082f $X=2.975 $Y=1.907
+ $X2=0 $Y2=0
cc_463 N_A_501_387#_c_338_n N_A_38_78#_c_1611_n 0.00107991f $X=3.415 $Y=1.76
+ $X2=0 $Y2=0
cc_464 N_A_501_387#_c_324_n N_VGND_M1019_d 0.00722747f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_465 N_A_501_387#_c_328_n N_VGND_c_1778_n 0.0383945f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_466 N_A_501_387#_c_322_n N_VGND_c_1783_n 0.0908278f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_467 N_A_501_387#_c_324_n N_VGND_c_1783_n 0.00941435f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_468 N_A_501_387#_c_328_n N_VGND_c_1783_n 0.0354007f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_469 N_A_501_387#_c_317_n N_VGND_c_1784_n 0.00320103f $X=6.045 $Y=1.085 $X2=0
+ $Y2=0
cc_470 N_A_501_387#_c_324_n N_VGND_c_1784_n 0.0163564f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_471 N_A_501_387#_c_317_n N_VGND_c_1788_n 0.00407044f $X=6.045 $Y=1.085 $X2=0
+ $Y2=0
cc_472 N_A_501_387#_c_322_n N_VGND_c_1788_n 0.0472862f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_473 N_A_501_387#_c_324_n N_VGND_c_1788_n 0.0405193f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_474 N_A_501_387#_c_328_n N_VGND_c_1788_n 0.0178884f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_475 N_A_501_387#_c_322_n N_VGND_c_1791_n 0.00667783f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_476 N_A_501_387#_c_324_n N_VGND_c_1791_n 0.0245264f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_477 N_A_501_387#_c_324_n A_910_119# 0.00134207f $X=6.085 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_478 N_A_841_401#_M1001_g N_RESET_B_c_631_n 0.00973011f $X=4.475 $Y=0.805
+ $X2=0 $Y2=0
cc_479 N_A_841_401#_M1001_g N_RESET_B_M1019_g 0.0415966f $X=4.475 $Y=0.805 $X2=0
+ $Y2=0
cc_480 N_A_841_401#_c_522_n N_RESET_B_M1019_g 0.0140148f $X=5.745 $Y=1.005 $X2=0
+ $Y2=0
cc_481 N_A_841_401#_M1001_g N_RESET_B_c_634_n 0.00952315f $X=4.475 $Y=0.805
+ $X2=0 $Y2=0
cc_482 N_A_841_401#_c_520_n N_RESET_B_c_634_n 0.00524003f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_483 N_A_841_401#_c_521_n N_RESET_B_c_634_n 0.0210965f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_484 N_A_841_401#_M1028_g N_RESET_B_M1031_g 0.0161997f $X=4.295 $Y=2.525 $X2=0
+ $Y2=0
cc_485 N_A_841_401#_c_520_n N_RESET_B_c_636_n 0.00340449f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_486 N_A_841_401#_c_522_n N_RESET_B_c_636_n 0.00175352f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_487 N_A_841_401#_c_529_n N_RESET_B_c_645_n 0.0210965f $X=4.417 $Y=2.005 $X2=0
+ $Y2=0
cc_488 N_A_841_401#_c_529_n N_RESET_B_c_646_n 0.00256409f $X=4.417 $Y=2.005
+ $X2=0 $Y2=0
cc_489 N_A_841_401#_c_530_n N_RESET_B_c_646_n 0.00401014f $X=4.417 $Y=2.155
+ $X2=0 $Y2=0
cc_490 N_A_841_401#_c_520_n N_RESET_B_c_646_n 0.0258991f $X=4.465 $Y=1.65 $X2=0
+ $Y2=0
cc_491 N_A_841_401#_M1016_d N_RESET_B_c_648_n 0.00232445f $X=6.18 $Y=1.735 $X2=0
+ $Y2=0
cc_492 N_A_841_401#_c_526_n N_RESET_B_c_648_n 0.00668397f $X=6.23 $Y=1.485 $X2=0
+ $Y2=0
cc_493 N_A_841_401#_c_527_n N_RESET_B_c_648_n 0.00201833f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_494 N_A_841_401#_c_534_n N_RESET_B_c_648_n 0.033324f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_495 N_A_841_401#_c_522_n N_A_709_463#_M1002_g 0.011848f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_496 N_A_841_401#_c_525_n N_A_709_463#_M1002_g 0.0046522f $X=5.83 $Y=1.4 $X2=0
+ $Y2=0
cc_497 N_A_841_401#_c_522_n N_A_709_463#_c_841_n 0.00506798f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_498 N_A_841_401#_c_526_n N_A_709_463#_c_841_n 0.0093946f $X=6.23 $Y=1.485
+ $X2=0 $Y2=0
cc_499 N_A_841_401#_c_527_n N_A_709_463#_c_841_n 0.00867517f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_500 N_A_841_401#_c_534_n N_A_709_463#_c_841_n 0.00413157f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_501 N_A_841_401#_M1001_g N_A_709_463#_c_842_n 0.00129073f $X=4.475 $Y=0.805
+ $X2=0 $Y2=0
cc_502 N_A_841_401#_c_530_n N_A_709_463#_c_842_n 0.00620045f $X=4.417 $Y=2.155
+ $X2=0 $Y2=0
cc_503 N_A_841_401#_c_520_n N_A_709_463#_c_842_n 0.0796667f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_504 N_A_841_401#_c_521_n N_A_709_463#_c_842_n 0.00416444f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_505 N_A_841_401#_c_523_n N_A_709_463#_c_842_n 0.0050659f $X=4.63 $Y=1.005
+ $X2=0 $Y2=0
cc_506 N_A_841_401#_M1028_g N_A_709_463#_c_880_n 0.0088331f $X=4.295 $Y=2.525
+ $X2=0 $Y2=0
cc_507 N_A_841_401#_c_530_n N_A_709_463#_c_880_n 0.00140174f $X=4.417 $Y=2.155
+ $X2=0 $Y2=0
cc_508 N_A_841_401#_c_520_n N_A_709_463#_c_880_n 0.0125914f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_509 N_A_841_401#_M1028_g N_A_709_463#_c_849_n 0.00100784f $X=4.295 $Y=2.525
+ $X2=0 $Y2=0
cc_510 N_A_841_401#_c_520_n N_A_709_463#_c_849_n 0.0259264f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_511 N_A_841_401#_c_521_n N_A_709_463#_c_849_n 0.00173976f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_512 N_A_841_401#_c_523_n N_A_709_463#_c_843_n 0.00118569f $X=4.63 $Y=1.005
+ $X2=0 $Y2=0
cc_513 N_A_841_401#_M1028_g N_A_709_463#_c_851_n 0.0102955f $X=4.295 $Y=2.525
+ $X2=0 $Y2=0
cc_514 N_A_841_401#_c_520_n N_A_709_463#_c_844_n 0.0144822f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_515 N_A_841_401#_c_521_n N_A_709_463#_c_844_n 4.19328e-19 $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_516 N_A_841_401#_c_522_n N_A_709_463#_c_844_n 0.0375552f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_517 N_A_841_401#_c_525_n N_A_709_463#_c_844_n 0.00811118f $X=5.83 $Y=1.4
+ $X2=0 $Y2=0
cc_518 N_A_841_401#_c_527_n N_A_709_463#_c_844_n 0.0135374f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_519 N_A_841_401#_c_534_n N_A_709_463#_c_844_n 0.0012591f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_520 N_A_841_401#_c_522_n N_A_709_463#_c_845_n 0.00123201f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_521 N_A_841_401#_c_525_n N_A_709_463#_c_845_n 7.93674e-19 $X=5.83 $Y=1.4
+ $X2=0 $Y2=0
cc_522 N_A_841_401#_c_527_n N_A_709_463#_c_845_n 5.0886e-19 $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_523 N_A_841_401#_M1028_g N_A_709_463#_c_853_n 7.55769e-19 $X=4.295 $Y=2.525
+ $X2=0 $Y2=0
cc_524 N_A_841_401#_M1028_g N_A_307_387#_M1009_g 0.0406315f $X=4.295 $Y=2.525
+ $X2=0 $Y2=0
cc_525 N_A_841_401#_M1028_g N_A_307_387#_c_984_n 0.0118199f $X=4.295 $Y=2.525
+ $X2=0 $Y2=0
cc_526 N_A_841_401#_c_534_n N_A_307_387#_c_984_n 0.00262042f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_527 N_A_841_401#_c_534_n N_A_307_387#_M1020_g 0.0171838f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_528 N_A_841_401#_c_526_n N_A_307_387#_c_972_n 0.00287849f $X=6.23 $Y=1.485
+ $X2=0 $Y2=0
cc_529 N_A_841_401#_c_534_n N_A_307_387#_c_972_n 0.00136985f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_530 N_A_841_401#_c_534_n N_A_1224_74#_c_1281_n 0.0217844f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_531 N_A_841_401#_M1028_g N_VPWR_c_1465_n 0.00327338f $X=4.295 $Y=2.525 $X2=0
+ $Y2=0
cc_532 N_A_841_401#_c_526_n N_VPWR_c_1466_n 0.00586599f $X=6.23 $Y=1.485 $X2=0
+ $Y2=0
cc_533 N_A_841_401#_c_527_n N_VPWR_c_1466_n 0.0111121f $X=5.915 $Y=1.485 $X2=0
+ $Y2=0
cc_534 N_A_841_401#_c_534_n N_VPWR_c_1466_n 0.0342363f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_535 N_A_841_401#_c_534_n N_VPWR_c_1475_n 0.0056446f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_536 N_A_841_401#_M1028_g N_VPWR_c_1460_n 0.00112709f $X=4.295 $Y=2.525 $X2=0
+ $Y2=0
cc_537 N_A_841_401#_c_534_n N_VPWR_c_1460_n 0.00682683f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_538 N_A_841_401#_c_522_n N_VGND_M1019_d 0.00389013f $X=5.745 $Y=1.005 $X2=0
+ $Y2=0
cc_539 N_A_841_401#_c_522_n A_910_119# 0.00103428f $X=5.745 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_540 N_A_841_401#_c_523_n A_910_119# 2.36857e-19 $X=4.63 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_541 N_RESET_B_c_631_n N_A_709_463#_M1002_g 0.0226708f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_636_n N_A_709_463#_M1002_g 0.00742734f $X=4.89 $Y=1.24 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_648_n N_A_709_463#_c_841_n 0.00220106f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_544 N_RESET_B_c_649_n N_A_709_463#_c_841_n 0.00116431f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_652_n N_A_709_463#_c_841_n 0.0017604f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_648_n N_A_709_463#_c_847_n 0.00777505f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_646_n N_A_709_463#_c_842_n 0.0156929f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_RESET_B_M1031_g N_A_709_463#_c_880_n 0.00543094f $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_646_n N_A_709_463#_c_880_n 0.011739f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_634_n N_A_709_463#_c_849_n 0.00710021f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_551 N_RESET_B_M1031_g N_A_709_463#_c_849_n 0.00814861f $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_552 N_RESET_B_c_645_n N_A_709_463#_c_849_n 0.00664711f $X=4.93 $Y=1.99 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_646_n N_A_709_463#_c_849_n 0.0226098f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_649_n N_A_709_463#_c_849_n 4.39853e-19 $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_651_n N_A_709_463#_c_849_n 0.00639141f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_652_n N_A_709_463#_c_849_n 0.0224281f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_646_n N_A_709_463#_c_850_n 0.00674995f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_558 N_RESET_B_M1031_g N_A_709_463#_c_851_n 7.81991e-19 $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_646_n N_A_709_463#_c_851_n 0.00649133f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_634_n N_A_709_463#_c_844_n 0.00724972f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_646_n N_A_709_463#_c_844_n 0.00666358f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_649_n N_A_709_463#_c_844_n 0.00107679f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_651_n N_A_709_463#_c_844_n 0.00728227f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_652_n N_A_709_463#_c_844_n 0.0190365f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_634_n N_A_709_463#_c_845_n 0.0174208f $X=4.915 $Y=1.825 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_651_n N_A_709_463#_c_845_n 0.0207972f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_652_n N_A_709_463#_c_845_n 4.14991e-19 $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_568 N_RESET_B_M1031_g N_A_709_463#_c_853_n 0.00851591f $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_646_n N_A_709_463#_c_853_n 0.00774464f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_570 N_RESET_B_c_651_n N_A_709_463#_c_853_n 0.00850056f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_571 N_RESET_B_c_652_n N_A_709_463#_c_853_n 0.00602228f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_646_n N_A_307_387#_M1006_s 8.4959e-19 $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_646_n N_A_307_387#_M1014_g 0.00762717f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_631_n N_A_307_387#_c_967_n 0.0104164f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_646_n N_A_307_387#_c_978_n 0.00128299f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_576 N_RESET_B_c_646_n N_A_307_387#_c_968_n 3.41208e-19 $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_577 N_RESET_B_c_631_n N_A_307_387#_M1018_g 0.00882199f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_646_n N_A_307_387#_M1009_g 0.00246505f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_RESET_B_M1031_g N_A_307_387#_c_984_n 0.011899f $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_648_n N_A_307_387#_M1020_g 0.0130216f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_648_n N_A_307_387#_c_971_n 3.83564e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_RESET_B_c_630_n N_A_307_387#_c_974_n 0.00410233f $X=1.097 $Y=1.908
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_646_n N_A_307_387#_c_974_n 0.00308596f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_647_n N_A_307_387#_c_974_n 7.5222e-19 $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_646_n N_A_307_387#_c_975_n 0.00245663f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_586 N_RESET_B_M1029_g N_A_307_387#_c_976_n 0.00418773f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_631_n N_A_307_387#_c_976_n 0.00920106f $X=4.79 $Y=0.18 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_637_n N_A_307_387#_c_976_n 0.00410233f $X=1.165 $Y=1.295
+ $X2=0 $Y2=0
cc_589 N_RESET_B_c_638_n N_A_307_387#_c_976_n 0.0599858f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_590 N_RESET_B_M1024_g N_A_307_387#_c_992_n 0.00181752f $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_591 N_RESET_B_c_646_n N_A_307_387#_c_992_n 0.0236535f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_647_n N_A_307_387#_c_992_n 0.00203256f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_593 N_RESET_B_c_638_n N_A_307_387#_c_992_n 0.013265f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_594 N_RESET_B_c_654_n N_A_307_387#_c_992_n 0.0015671f $X=1.165 $Y=1.975 $X2=0
+ $Y2=0
cc_595 N_RESET_B_M1026_g N_A_1482_48#_c_1156_n 0.0196155f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_596 N_RESET_B_M1021_g N_A_1482_48#_M1007_g 0.0117619f $X=8.18 $Y=2.565 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_648_n N_A_1482_48#_M1007_g 0.00571623f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_RESET_B_c_650_n N_A_1482_48#_M1007_g 0.00149248f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_599 N_RESET_B_c_655_n N_A_1482_48#_M1007_g 0.0401889f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_600 N_RESET_B_c_656_n N_A_1482_48#_M1007_g 0.00190186f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_601 N_RESET_B_M1026_g N_A_1482_48#_c_1158_n 0.0144302f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_602 N_RESET_B_M1021_g N_A_1482_48#_c_1165_n 0.00825702f $X=8.18 $Y=2.565
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_650_n N_A_1482_48#_c_1165_n 9.35982e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_604 N_RESET_B_c_655_n N_A_1482_48#_c_1165_n 0.0013781f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_605 N_RESET_B_c_656_n N_A_1482_48#_c_1165_n 0.0201374f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_606 N_RESET_B_M1026_g N_A_1482_48#_c_1159_n 0.00201284f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_607 N_RESET_B_M1026_g N_A_1482_48#_c_1161_n 0.00118187f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_608 N_RESET_B_M1026_g N_A_1482_48#_c_1167_n 0.00150115f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_609 N_RESET_B_c_655_n N_A_1482_48#_c_1167_n 3.55688e-19 $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_656_n N_A_1482_48#_c_1167_n 0.00823641f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_611 N_RESET_B_M1026_g N_A_1482_48#_c_1163_n 0.0401889f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_648_n N_A_1224_74#_M1020_d 0.00103706f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_RESET_B_M1026_g N_A_1224_74#_M1027_g 0.0533792f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_614 N_RESET_B_M1026_g N_A_1224_74#_M1025_g 0.00701487f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_615 N_RESET_B_M1021_g N_A_1224_74#_M1025_g 0.0156201f $X=8.18 $Y=2.565 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_655_n N_A_1224_74#_M1025_g 0.018107f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_617 N_RESET_B_c_656_n N_A_1224_74#_M1025_g 3.64033e-19 $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_618 N_RESET_B_M1026_g N_A_1224_74#_c_1252_n 0.0220605f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_648_n N_A_1224_74#_c_1281_n 0.0113022f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_620 N_RESET_B_c_648_n N_A_1224_74#_c_1261_n 0.00715094f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_621 N_RESET_B_c_648_n N_A_1224_74#_c_1262_n 0.00106639f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_622 N_RESET_B_M1026_g N_A_1224_74#_c_1263_n 0.00129569f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_623 N_RESET_B_M1021_g N_A_1224_74#_c_1263_n 8.86228e-19 $X=8.18 $Y=2.565
+ $X2=0 $Y2=0
cc_624 N_RESET_B_c_648_n N_A_1224_74#_c_1263_n 0.0226223f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_625 N_RESET_B_c_650_n N_A_1224_74#_c_1263_n 0.00270727f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_626 N_RESET_B_c_655_n N_A_1224_74#_c_1263_n 3.32288e-19 $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_627 N_RESET_B_c_656_n N_A_1224_74#_c_1263_n 0.0230781f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_628 N_RESET_B_M1026_g N_A_1224_74#_c_1264_n 0.0108822f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_629 N_RESET_B_c_648_n N_A_1224_74#_c_1264_n 0.00339956f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_630 N_RESET_B_c_650_n N_A_1224_74#_c_1264_n 0.00379913f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_631 N_RESET_B_c_655_n N_A_1224_74#_c_1264_n 0.00439769f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_656_n N_A_1224_74#_c_1264_n 0.0255102f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_633 N_RESET_B_M1026_g N_A_1224_74#_c_1266_n 0.00118353f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_634 N_RESET_B_c_646_n N_VPWR_M1006_d 0.00617044f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_648_n N_VPWR_M1016_s 0.00310864f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_636 N_RESET_B_M1024_g N_VPWR_c_1463_n 0.00839184f $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_637 N_RESET_B_M1031_g N_VPWR_c_1465_n 0.00327338f $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_638 N_RESET_B_c_648_n N_VPWR_c_1466_n 0.0237051f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_649_n N_VPWR_c_1466_n 0.00275995f $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_651_n N_VPWR_c_1466_n 0.00100362f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_652_n N_VPWR_c_1466_n 0.0239957f $X=5.395 $Y=1.99 $X2=0 $Y2=0
cc_642 N_RESET_B_M1021_g N_VPWR_c_1467_n 0.00382649f $X=8.18 $Y=2.565 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_650_n N_VPWR_c_1467_n 0.00183431f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_655_n N_VPWR_c_1467_n 0.00242435f $X=8.135 $Y=2 $X2=0 $Y2=0
cc_645 N_RESET_B_c_656_n N_VPWR_c_1467_n 0.0174647f $X=8.135 $Y=2 $X2=0 $Y2=0
cc_646 N_RESET_B_M1021_g N_VPWR_c_1468_n 0.00537883f $X=8.18 $Y=2.565 $X2=0
+ $Y2=0
cc_647 N_RESET_B_M1024_g N_VPWR_c_1471_n 0.00336715f $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_648 N_RESET_B_M1024_g N_VPWR_c_1460_n 0.00436408f $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_649 N_RESET_B_M1031_g N_VPWR_c_1460_n 0.00112709f $X=4.93 $Y=2.525 $X2=0
+ $Y2=0
cc_650 N_RESET_B_M1021_g N_VPWR_c_1460_n 0.00587053f $X=8.18 $Y=2.565 $X2=0
+ $Y2=0
cc_651 N_RESET_B_M1029_g N_A_38_78#_c_1606_n 7.65322e-19 $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_652 N_RESET_B_M1024_g N_A_38_78#_c_1612_n 2.23847e-19 $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_653 N_RESET_B_M1029_g N_A_38_78#_c_1607_n 0.0181359f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_654 N_RESET_B_c_647_n N_A_38_78#_c_1607_n 0.00185256f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_638_n N_A_38_78#_c_1607_n 0.0731888f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_656 N_RESET_B_M1024_g N_A_38_78#_c_1614_n 0.0164363f $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_646_n N_A_38_78#_c_1614_n 0.029557f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_647_n N_A_38_78#_c_1614_n 0.00840362f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_638_n N_A_38_78#_c_1614_n 0.0107061f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_660 N_RESET_B_c_654_n N_A_38_78#_c_1614_n 0.0025137f $X=1.165 $Y=1.975 $X2=0
+ $Y2=0
cc_661 N_RESET_B_c_646_n N_A_38_78#_c_1615_n 0.0118476f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_662 N_RESET_B_c_646_n N_A_38_78#_c_1609_n 0.0134686f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_663 N_RESET_B_M1029_g N_A_38_78#_c_1610_n 8.39005e-19 $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_664 N_RESET_B_M1024_g N_A_38_78#_c_1617_n 0.00532562f $X=0.955 $Y=2.75 $X2=0
+ $Y2=0
cc_665 N_RESET_B_c_646_n N_A_38_78#_c_1618_n 0.00778362f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_666 N_RESET_B_c_646_n N_A_38_78#_c_1611_n 0.00542381f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_667 N_RESET_B_M1029_g N_VGND_c_1776_n 0.00269179f $X=0.94 $Y=0.6 $X2=0 $Y2=0
cc_668 N_RESET_B_c_631_n N_VGND_c_1776_n 0.0190483f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_669 N_RESET_B_c_637_n N_VGND_c_1776_n 0.00181416f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_670 N_RESET_B_c_638_n N_VGND_c_1776_n 0.0144384f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_671 N_RESET_B_c_631_n N_VGND_c_1777_n 0.0233742f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_672 N_RESET_B_c_631_n N_VGND_c_1778_n 0.0257653f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_673 N_RESET_B_M1026_g N_VGND_c_1779_n 0.0152783f $X=8.045 $Y=0.58 $X2=0 $Y2=0
cc_674 N_RESET_B_c_632_n N_VGND_c_1782_n 0.0064002f $X=1.015 $Y=0.18 $X2=0 $Y2=0
cc_675 N_RESET_B_c_631_n N_VGND_c_1783_n 0.0558348f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_676 N_RESET_B_M1026_g N_VGND_c_1785_n 0.00383152f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_677 N_RESET_B_c_631_n N_VGND_c_1788_n 0.0925451f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_678 N_RESET_B_c_632_n N_VGND_c_1788_n 0.0113744f $X=1.015 $Y=0.18 $X2=0 $Y2=0
cc_679 N_RESET_B_M1026_g N_VGND_c_1788_n 0.0075725f $X=8.045 $Y=0.58 $X2=0 $Y2=0
cc_680 N_RESET_B_c_631_n N_VGND_c_1791_n 0.00776078f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_681 N_A_709_463#_c_850_n N_A_307_387#_c_980_n 0.00349469f $X=4.01 $Y=2.585
+ $X2=0 $Y2=0
cc_682 N_A_709_463#_c_842_n N_A_307_387#_M1018_g 6.85936e-19 $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_683 N_A_709_463#_c_843_n N_A_307_387#_M1018_g 0.00230849f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_684 N_A_709_463#_c_842_n N_A_307_387#_M1009_g 0.00123745f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_685 N_A_709_463#_c_850_n N_A_307_387#_M1009_g 0.0116701f $X=4.01 $Y=2.585
+ $X2=0 $Y2=0
cc_686 N_A_709_463#_c_847_n N_A_307_387#_c_984_n 0.0123711f $X=6.09 $Y=1.615
+ $X2=0 $Y2=0
cc_687 N_A_709_463#_c_880_n N_A_307_387#_c_984_n 0.00158437f $X=4.89 $Y=2.5
+ $X2=0 $Y2=0
cc_688 N_A_709_463#_c_851_n N_A_307_387#_c_984_n 0.00250946f $X=4.27 $Y=2.585
+ $X2=0 $Y2=0
cc_689 N_A_709_463#_c_853_n N_A_307_387#_c_984_n 0.00556718f $X=4.975 $Y=2.515
+ $X2=0 $Y2=0
cc_690 N_A_709_463#_c_847_n N_A_307_387#_M1020_g 0.00899217f $X=6.09 $Y=1.615
+ $X2=0 $Y2=0
cc_691 N_A_709_463#_c_841_n N_A_307_387#_c_972_n 0.00899217f $X=6 $Y=1.54 $X2=0
+ $Y2=0
cc_692 N_A_709_463#_c_880_n N_VPWR_M1028_d 0.00813251f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_693 N_A_709_463#_c_880_n N_VPWR_c_1465_n 0.026965f $X=4.89 $Y=2.5 $X2=0 $Y2=0
cc_694 N_A_709_463#_c_841_n N_VPWR_c_1466_n 0.00441012f $X=6 $Y=1.54 $X2=0 $Y2=0
cc_695 N_A_709_463#_c_847_n N_VPWR_c_1466_n 0.016723f $X=6.09 $Y=1.615 $X2=0
+ $Y2=0
cc_696 N_A_709_463#_c_853_n N_VPWR_c_1466_n 0.0135992f $X=4.975 $Y=2.515 $X2=0
+ $Y2=0
cc_697 N_A_709_463#_c_880_n N_VPWR_c_1473_n 0.00186481f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_698 N_A_709_463#_c_850_n N_VPWR_c_1473_n 0.0156174f $X=4.01 $Y=2.585 $X2=0
+ $Y2=0
cc_699 N_A_709_463#_c_880_n N_VPWR_c_1474_n 0.0010327f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_700 N_A_709_463#_c_853_n N_VPWR_c_1474_n 0.00688179f $X=4.975 $Y=2.515 $X2=0
+ $Y2=0
cc_701 N_A_709_463#_c_847_n N_VPWR_c_1460_n 9.455e-19 $X=6.09 $Y=1.615 $X2=0
+ $Y2=0
cc_702 N_A_709_463#_c_880_n N_VPWR_c_1460_n 0.00729806f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_703 N_A_709_463#_c_850_n N_VPWR_c_1460_n 0.019648f $X=4.01 $Y=2.585 $X2=0
+ $Y2=0
cc_704 N_A_709_463#_c_853_n N_VPWR_c_1460_n 0.0107097f $X=4.975 $Y=2.515 $X2=0
+ $Y2=0
cc_705 N_A_709_463#_c_842_n N_A_38_78#_c_1608_n 0.00513545f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_706 N_A_709_463#_c_843_n N_A_38_78#_c_1608_n 0.0162186f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_707 N_A_709_463#_M1005_d N_A_38_78#_c_1615_n 0.00169018f $X=3.545 $Y=2.315
+ $X2=0 $Y2=0
cc_708 N_A_709_463#_c_842_n N_A_38_78#_c_1615_n 0.0120586f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_709 N_A_709_463#_c_850_n N_A_38_78#_c_1615_n 0.0155522f $X=4.01 $Y=2.585
+ $X2=0 $Y2=0
cc_710 N_A_709_463#_c_842_n N_A_38_78#_c_1609_n 0.0583112f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_711 N_A_709_463#_c_850_n N_A_38_78#_c_1618_n 0.0103876f $X=4.01 $Y=2.585
+ $X2=0 $Y2=0
cc_712 N_A_709_463#_c_842_n N_A_38_78#_c_1611_n 0.0132832f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_713 N_A_709_463#_c_843_n N_A_38_78#_c_1611_n 0.0109432f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_714 N_A_709_463#_c_842_n A_799_463# 2.7357e-19 $X=4.095 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_715 N_A_709_463#_c_851_n A_799_463# 2.73927e-19 $X=4.27 $Y=2.585 $X2=-0.19
+ $Y2=-0.245
cc_716 N_A_709_463#_M1002_g N_VGND_c_1784_n 0.00320129f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_717 N_A_709_463#_M1002_g N_VGND_c_1788_n 0.00402508f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_718 N_A_709_463#_M1002_g N_VGND_c_1791_n 0.00397703f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_719 N_A_307_387#_M1000_g N_A_1482_48#_c_1156_n 0.0495982f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_720 N_A_307_387#_M1000_g N_A_1482_48#_M1007_g 0.0112982f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_721 N_A_307_387#_M1000_g N_A_1482_48#_c_1161_n 0.00102678f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_722 N_A_307_387#_M1000_g N_A_1224_74#_c_1277_n 0.0169263f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_723 N_A_307_387#_M1020_g N_A_1224_74#_c_1281_n 0.00394014f $X=6.54 $Y=2.235
+ $X2=0 $Y2=0
cc_724 N_A_307_387#_M1000_g N_A_1224_74#_c_1260_n 0.0221333f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_725 N_A_307_387#_c_971_n N_A_1224_74#_c_1261_n 0.00206465f $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_726 N_A_307_387#_M1000_g N_A_1224_74#_c_1261_n 0.0011854f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_727 N_A_307_387#_c_971_n N_A_1224_74#_c_1262_n 0.00561544f $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_728 N_A_307_387#_M1000_g N_A_1224_74#_c_1262_n 0.00135722f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_729 N_A_307_387#_c_971_n N_A_1224_74#_c_1263_n 3.07924e-19 $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_730 N_A_307_387#_M1014_g N_VPWR_c_1464_n 0.0117819f $X=2.415 $Y=2.495 $X2=0
+ $Y2=0
cc_731 N_A_307_387#_c_979_n N_VPWR_c_1464_n 0.0022152f $X=2.935 $Y=3.075 $X2=0
+ $Y2=0
cc_732 N_A_307_387#_c_981_n N_VPWR_c_1464_n 6.90101e-19 $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_307_387#_M1009_g N_VPWR_c_1465_n 0.00613878f $X=3.905 $Y=2.525 $X2=0
+ $Y2=0
cc_734 N_A_307_387#_c_984_n N_VPWR_c_1465_n 0.0257522f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_735 N_A_307_387#_c_984_n N_VPWR_c_1466_n 0.0210786f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_736 N_A_307_387#_M1020_g N_VPWR_c_1466_n 0.00679477f $X=6.54 $Y=2.235 $X2=0
+ $Y2=0
cc_737 N_A_307_387#_M1014_g N_VPWR_c_1473_n 0.00406785f $X=2.415 $Y=2.495 $X2=0
+ $Y2=0
cc_738 N_A_307_387#_c_981_n N_VPWR_c_1473_n 0.0426327f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_739 N_A_307_387#_c_984_n N_VPWR_c_1474_n 0.0295821f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_740 N_A_307_387#_c_984_n N_VPWR_c_1475_n 0.0193431f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_741 N_A_307_387#_M1014_g N_VPWR_c_1460_n 0.00513967f $X=2.415 $Y=2.495 $X2=0
+ $Y2=0
cc_742 N_A_307_387#_c_980_n N_VPWR_c_1460_n 0.0228826f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_307_387#_c_981_n N_VPWR_c_1460_n 0.00601501f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_744 N_A_307_387#_c_984_n N_VPWR_c_1460_n 0.0766558f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_745 N_A_307_387#_c_989_n N_VPWR_c_1460_n 0.00500367f $X=3.905 $Y=3.15 $X2=0
+ $Y2=0
cc_746 N_A_307_387#_c_976_n N_A_38_78#_c_1607_n 0.009918f $X=1.735 $Y=0.715
+ $X2=0 $Y2=0
cc_747 N_A_307_387#_c_992_n N_A_38_78#_c_1607_n 0.00301391f $X=1.66 $Y=2.1 $X2=0
+ $Y2=0
cc_748 N_A_307_387#_M1006_s N_A_38_78#_c_1614_n 0.00752456f $X=1.535 $Y=1.935
+ $X2=0 $Y2=0
cc_749 N_A_307_387#_M1014_g N_A_38_78#_c_1614_n 0.014535f $X=2.415 $Y=2.495
+ $X2=0 $Y2=0
cc_750 N_A_307_387#_c_979_n N_A_38_78#_c_1614_n 0.0130237f $X=2.935 $Y=3.075
+ $X2=0 $Y2=0
cc_751 N_A_307_387#_c_988_n N_A_38_78#_c_1614_n 8.19207e-19 $X=2.95 $Y=2.2 $X2=0
+ $Y2=0
cc_752 N_A_307_387#_c_992_n N_A_38_78#_c_1614_n 0.0248543f $X=1.66 $Y=2.1 $X2=0
+ $Y2=0
cc_753 N_A_307_387#_c_968_n N_A_38_78#_c_1608_n 0.00132611f $X=3.51 $Y=1.4 $X2=0
+ $Y2=0
cc_754 N_A_307_387#_M1018_g N_A_38_78#_c_1608_n 0.0116244f $X=3.585 $Y=0.805
+ $X2=0 $Y2=0
cc_755 N_A_307_387#_M1009_g N_A_38_78#_c_1615_n 0.00449347f $X=3.905 $Y=2.525
+ $X2=0 $Y2=0
cc_756 N_A_307_387#_c_968_n N_A_38_78#_c_1609_n 0.00148463f $X=3.51 $Y=1.4 $X2=0
+ $Y2=0
cc_757 N_A_307_387#_c_969_n N_A_38_78#_c_1609_n 8.59635e-19 $X=3.1 $Y=1.4 $X2=0
+ $Y2=0
cc_758 N_A_307_387#_c_979_n N_A_38_78#_c_1618_n 0.00972592f $X=2.935 $Y=3.075
+ $X2=0 $Y2=0
cc_759 N_A_307_387#_c_980_n N_A_38_78#_c_1618_n 0.00487453f $X=3.815 $Y=3.15
+ $X2=0 $Y2=0
cc_760 N_A_307_387#_c_968_n N_A_38_78#_c_1611_n 0.00913328f $X=3.51 $Y=1.4 $X2=0
+ $Y2=0
cc_761 N_A_307_387#_M1018_g N_A_38_78#_c_1611_n 0.0105843f $X=3.585 $Y=0.805
+ $X2=0 $Y2=0
cc_762 N_A_307_387#_c_1004_n N_VGND_M1011_d 0.00702203f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_763 N_A_307_387#_c_976_n N_VGND_c_1776_n 0.0212471f $X=1.735 $Y=0.715 $X2=0
+ $Y2=0
cc_764 N_A_307_387#_c_976_n N_VGND_c_1777_n 0.0108572f $X=1.735 $Y=0.715 $X2=0
+ $Y2=0
cc_765 N_A_307_387#_c_967_n N_VGND_c_1778_n 0.00119784f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_766 N_A_307_387#_c_1004_n N_VGND_c_1778_n 0.0208278f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_767 N_A_307_387#_c_976_n N_VGND_c_1778_n 0.0126872f $X=1.735 $Y=0.715 $X2=0
+ $Y2=0
cc_768 N_A_307_387#_M1000_g N_VGND_c_1779_n 0.00154981f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_769 N_A_307_387#_M1000_g N_VGND_c_1784_n 0.00309049f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_770 N_A_307_387#_c_967_n N_VGND_c_1788_n 9.39239e-19 $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_771 N_A_307_387#_M1000_g N_VGND_c_1788_n 0.0040628f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_772 N_A_307_387#_c_976_n N_VGND_c_1788_n 0.0126278f $X=1.735 $Y=0.715 $X2=0
+ $Y2=0
cc_773 N_A_1482_48#_c_1158_n N_A_1224_74#_M1027_g 0.0108008f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_774 N_A_1482_48#_c_1159_n N_A_1224_74#_M1027_g 0.0132755f $X=8.65 $Y=0.58
+ $X2=0 $Y2=0
cc_775 N_A_1482_48#_c_1160_n N_A_1224_74#_M1027_g 0.00584201f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_776 N_A_1482_48#_c_1162_n N_A_1224_74#_M1027_g 0.0045388f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_777 N_A_1482_48#_c_1165_n N_A_1224_74#_M1025_g 0.0194527f $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_778 N_A_1482_48#_c_1160_n N_A_1224_74#_M1025_g 0.00407488f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_779 N_A_1482_48#_c_1167_n N_A_1224_74#_M1025_g 0.0144953f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_780 N_A_1482_48#_c_1160_n N_A_1224_74#_c_1251_n 0.0253235f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_781 N_A_1482_48#_c_1167_n N_A_1224_74#_c_1251_n 7.56579e-19 $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_782 N_A_1482_48#_c_1167_n N_A_1224_74#_c_1252_n 4.86873e-19 $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_783 N_A_1482_48#_c_1162_n N_A_1224_74#_c_1252_n 0.00825331f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_784 N_A_1482_48#_c_1165_n N_A_1224_74#_M1008_g 5.79058e-19 $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_785 N_A_1482_48#_c_1160_n N_A_1224_74#_M1008_g 0.0021029f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_786 N_A_1482_48#_c_1167_n N_A_1224_74#_M1008_g 0.00190937f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_787 N_A_1482_48#_c_1159_n N_A_1224_74#_M1015_g 0.00122775f $X=8.65 $Y=0.58
+ $X2=0 $Y2=0
cc_788 N_A_1482_48#_c_1160_n N_A_1224_74#_M1015_g 0.00251042f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_789 N_A_1482_48#_c_1156_n N_A_1224_74#_c_1277_n 0.0012657f $X=7.485 $Y=0.9
+ $X2=0 $Y2=0
cc_790 N_A_1482_48#_M1007_g N_A_1224_74#_c_1281_n 0.0099672f $X=7.67 $Y=2.565
+ $X2=0 $Y2=0
cc_791 N_A_1482_48#_c_1156_n N_A_1224_74#_c_1260_n 0.00230939f $X=7.485 $Y=0.9
+ $X2=0 $Y2=0
cc_792 N_A_1482_48#_M1007_g N_A_1224_74#_c_1260_n 0.00111943f $X=7.67 $Y=2.565
+ $X2=0 $Y2=0
cc_793 N_A_1482_48#_c_1161_n N_A_1224_74#_c_1260_n 0.0162835f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_794 N_A_1482_48#_c_1161_n N_A_1224_74#_c_1261_n 0.00432309f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_795 N_A_1482_48#_c_1163_n N_A_1224_74#_c_1261_n 0.00127859f $X=7.67 $Y=1.065
+ $X2=0 $Y2=0
cc_796 N_A_1482_48#_M1007_g N_A_1224_74#_c_1263_n 0.0199863f $X=7.67 $Y=2.565
+ $X2=0 $Y2=0
cc_797 N_A_1482_48#_M1007_g N_A_1224_74#_c_1264_n 0.00617973f $X=7.67 $Y=2.565
+ $X2=0 $Y2=0
cc_798 N_A_1482_48#_c_1158_n N_A_1224_74#_c_1264_n 0.0246405f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_799 N_A_1482_48#_c_1161_n N_A_1224_74#_c_1264_n 0.00601156f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_800 N_A_1482_48#_M1007_g N_A_1224_74#_c_1265_n 0.0053332f $X=7.67 $Y=2.565
+ $X2=0 $Y2=0
cc_801 N_A_1482_48#_c_1161_n N_A_1224_74#_c_1265_n 0.0125972f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_802 N_A_1482_48#_c_1163_n N_A_1224_74#_c_1265_n 6.55449e-19 $X=7.67 $Y=1.065
+ $X2=0 $Y2=0
cc_803 N_A_1482_48#_c_1158_n N_A_1224_74#_c_1266_n 0.00997859f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_804 N_A_1482_48#_c_1160_n N_A_1224_74#_c_1266_n 0.0233867f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_805 N_A_1482_48#_c_1167_n N_A_1224_74#_c_1266_n 0.0116759f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_806 N_A_1482_48#_c_1162_n N_A_1224_74#_c_1266_n 0.0109402f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_807 N_A_1482_48#_c_1167_n N_VPWR_M1025_d 0.00364967f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_808 N_A_1482_48#_M1007_g N_VPWR_c_1467_n 0.00620049f $X=7.67 $Y=2.565 $X2=0
+ $Y2=0
cc_809 N_A_1482_48#_c_1165_n N_VPWR_c_1467_n 0.0139263f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_810 N_A_1482_48#_c_1165_n N_VPWR_c_1468_n 0.00638559f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_811 N_A_1482_48#_c_1165_n N_VPWR_c_1469_n 0.0464459f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_812 N_A_1482_48#_c_1167_n N_VPWR_c_1469_n 0.012936f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_813 N_A_1482_48#_M1007_g N_VPWR_c_1475_n 0.00485739f $X=7.67 $Y=2.565 $X2=0
+ $Y2=0
cc_814 N_A_1482_48#_M1007_g N_VPWR_c_1460_n 0.00587053f $X=7.67 $Y=2.565 $X2=0
+ $Y2=0
cc_815 N_A_1482_48#_c_1165_n N_VPWR_c_1460_n 0.0113911f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_816 N_A_1482_48#_c_1160_n N_Q_N_c_1727_n 0.018767f $X=8.885 $Y=1.765 $X2=0
+ $Y2=0
cc_817 N_A_1482_48#_c_1167_n N_Q_N_c_1727_n 0.00158085f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_818 N_A_1482_48#_c_1167_n N_Q_N_c_1730_n 0.00456512f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_819 N_A_1482_48#_c_1156_n N_VGND_c_1779_n 0.0147674f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_820 N_A_1482_48#_c_1158_n N_VGND_c_1779_n 0.0137782f $X=8.485 $Y=0.985 $X2=0
+ $Y2=0
cc_821 N_A_1482_48#_c_1159_n N_VGND_c_1779_n 0.0110441f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_822 N_A_1482_48#_c_1161_n N_VGND_c_1779_n 0.0129689f $X=7.595 $Y=0.985 $X2=0
+ $Y2=0
cc_823 N_A_1482_48#_c_1163_n N_VGND_c_1779_n 0.00131228f $X=7.67 $Y=1.065 $X2=0
+ $Y2=0
cc_824 N_A_1482_48#_c_1159_n N_VGND_c_1780_n 0.0454165f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_825 N_A_1482_48#_c_1160_n N_VGND_c_1780_n 0.00455872f $X=8.885 $Y=1.765 $X2=0
+ $Y2=0
cc_826 N_A_1482_48#_c_1162_n N_VGND_c_1780_n 0.0145003f $X=8.727 $Y=0.985 $X2=0
+ $Y2=0
cc_827 N_A_1482_48#_c_1156_n N_VGND_c_1784_n 0.00383152f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_828 N_A_1482_48#_c_1159_n N_VGND_c_1785_n 0.0215384f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_829 N_A_1482_48#_c_1156_n N_VGND_c_1788_n 0.0075725f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_830 N_A_1482_48#_c_1159_n N_VGND_c_1788_n 0.0177458f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_831 N_A_1224_74#_M1030_g N_A_2026_424#_M1032_g 0.0171742f $X=10.5 $Y=2.54
+ $X2=0 $Y2=0
cc_832 N_A_1224_74#_M1013_g N_A_2026_424#_M1004_g 0.0197956f $X=10.515 $Y=0.645
+ $X2=0 $Y2=0
cc_833 N_A_1224_74#_c_1255_n N_A_2026_424#_c_1410_n 0.00519557f $X=10.41 $Y=1.43
+ $X2=0 $Y2=0
cc_834 N_A_1224_74#_M1013_g N_A_2026_424#_c_1410_n 0.0146713f $X=10.515 $Y=0.645
+ $X2=0 $Y2=0
cc_835 N_A_1224_74#_c_1259_n N_A_2026_424#_c_1410_n 6.73726e-19 $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_836 N_A_1224_74#_M1030_g N_A_2026_424#_c_1411_n 0.029305f $X=10.5 $Y=2.54
+ $X2=0 $Y2=0
cc_837 N_A_1224_74#_M1030_g N_A_2026_424#_c_1412_n 0.00787479f $X=10.5 $Y=2.54
+ $X2=0 $Y2=0
cc_838 N_A_1224_74#_c_1259_n N_A_2026_424#_c_1412_n 0.0139388f $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_839 N_A_1224_74#_c_1259_n N_A_2026_424#_c_1413_n 0.0214662f $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_840 N_A_1224_74#_c_1255_n N_A_2026_424#_c_1414_n 0.0144271f $X=10.41 $Y=1.43
+ $X2=0 $Y2=0
cc_841 N_A_1224_74#_M1030_g N_A_2026_424#_c_1414_n 7.34008e-19 $X=10.5 $Y=2.54
+ $X2=0 $Y2=0
cc_842 N_A_1224_74#_c_1259_n N_A_2026_424#_c_1414_n 8.33355e-19 $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_843 N_A_1224_74#_c_1281_n N_VPWR_c_1467_n 0.0264537f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_844 N_A_1224_74#_c_1263_n N_VPWR_c_1467_n 0.00214678f $X=7.58 $Y=2.365 $X2=0
+ $Y2=0
cc_845 N_A_1224_74#_M1025_g N_VPWR_c_1468_n 0.00473661f $X=8.63 $Y=2.565 $X2=0
+ $Y2=0
cc_846 N_A_1224_74#_M1025_g N_VPWR_c_1469_n 0.00904816f $X=8.63 $Y=2.565 $X2=0
+ $Y2=0
cc_847 N_A_1224_74#_M1008_g N_VPWR_c_1469_n 0.00577006f $X=9.145 $Y=2.4 $X2=0
+ $Y2=0
cc_848 N_A_1224_74#_M1030_g N_VPWR_c_1470_n 0.0065579f $X=10.5 $Y=2.54 $X2=0
+ $Y2=0
cc_849 N_A_1224_74#_c_1281_n N_VPWR_c_1475_n 0.0159371f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_850 N_A_1224_74#_M1008_g N_VPWR_c_1476_n 0.00553757f $X=9.145 $Y=2.4 $X2=0
+ $Y2=0
cc_851 N_A_1224_74#_M1030_g N_VPWR_c_1476_n 0.00521031f $X=10.5 $Y=2.54 $X2=0
+ $Y2=0
cc_852 N_A_1224_74#_M1025_g N_VPWR_c_1460_n 0.00587053f $X=8.63 $Y=2.565 $X2=0
+ $Y2=0
cc_853 N_A_1224_74#_M1008_g N_VPWR_c_1460_n 0.0109848f $X=9.145 $Y=2.4 $X2=0
+ $Y2=0
cc_854 N_A_1224_74#_M1030_g N_VPWR_c_1460_n 0.00987525f $X=10.5 $Y=2.54 $X2=0
+ $Y2=0
cc_855 N_A_1224_74#_c_1281_n N_VPWR_c_1460_n 0.0281713f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_856 N_A_1224_74#_c_1281_n A_1468_471# 0.00371878f $X=7.495 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_857 N_A_1224_74#_M1008_g N_Q_N_c_1727_n 0.00447321f $X=9.145 $Y=2.4 $X2=0
+ $Y2=0
cc_858 N_A_1224_74#_M1015_g N_Q_N_c_1727_n 0.0191689f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_859 N_A_1224_74#_c_1255_n N_Q_N_c_1727_n 0.0449729f $X=10.41 $Y=1.43 $X2=0
+ $Y2=0
cc_860 N_A_1224_74#_M1030_g N_Q_N_c_1727_n 0.00500627f $X=10.5 $Y=2.54 $X2=0
+ $Y2=0
cc_861 N_A_1224_74#_M1008_g N_Q_N_c_1730_n 0.00248876f $X=9.145 $Y=2.4 $X2=0
+ $Y2=0
cc_862 N_A_1224_74#_c_1256_n N_Q_N_c_1730_n 0.00992644f $X=9.515 $Y=1.43 $X2=0
+ $Y2=0
cc_863 N_A_1224_74#_M1027_g N_VGND_c_1779_n 0.0014914f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_864 N_A_1224_74#_c_1277_n N_VGND_c_1779_n 0.0120929f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_865 N_A_1224_74#_M1027_g N_VGND_c_1780_n 0.00378178f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_866 N_A_1224_74#_M1015_g N_VGND_c_1780_n 0.017876f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_867 N_A_1224_74#_c_1256_n N_VGND_c_1780_n 0.00653223f $X=9.515 $Y=1.43 $X2=0
+ $Y2=0
cc_868 N_A_1224_74#_M1013_g N_VGND_c_1781_n 0.00770628f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_869 N_A_1224_74#_c_1277_n N_VGND_c_1784_n 0.0242914f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_870 N_A_1224_74#_M1027_g N_VGND_c_1785_n 0.00434272f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_871 N_A_1224_74#_M1015_g N_VGND_c_1786_n 0.00383152f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_872 N_A_1224_74#_M1013_g N_VGND_c_1786_n 0.00461464f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_873 N_A_1224_74#_M1027_g N_VGND_c_1788_n 0.00825979f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_874 N_A_1224_74#_M1015_g N_VGND_c_1788_n 0.00762539f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_875 N_A_1224_74#_M1013_g N_VGND_c_1788_n 0.00914043f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_876 N_A_1224_74#_c_1277_n N_VGND_c_1788_n 0.02509f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_877 N_A_2026_424#_M1032_g N_VPWR_c_1470_n 0.00375859f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_878 N_A_2026_424#_c_1411_n N_VPWR_c_1470_n 0.0543362f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_879 N_A_2026_424#_c_1412_n N_VPWR_c_1470_n 0.0235211f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_880 N_A_2026_424#_c_1413_n N_VPWR_c_1470_n 0.00239853f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_881 N_A_2026_424#_c_1411_n N_VPWR_c_1476_n 0.0107623f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_882 N_A_2026_424#_M1032_g N_VPWR_c_1477_n 0.005209f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_883 N_A_2026_424#_M1032_g N_VPWR_c_1460_n 0.00986031f $X=11.015 $Y=2.4 $X2=0
+ $Y2=0
cc_884 N_A_2026_424#_c_1411_n N_VPWR_c_1460_n 0.0089917f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_885 N_A_2026_424#_c_1410_n N_Q_N_c_1727_n 0.0605318f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_886 N_A_2026_424#_c_1411_n N_Q_N_c_1727_n 0.0894765f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_887 N_A_2026_424#_c_1414_n N_Q_N_c_1727_n 0.0205307f $X=10.315 $Y=1.465 $X2=0
+ $Y2=0
cc_888 N_A_2026_424#_M1004_g Q 0.00795463f $X=11.015 $Y=0.74 $X2=0 $Y2=0
cc_889 N_A_2026_424#_M1004_g Q 0.00263483f $X=11.015 $Y=0.74 $X2=0 $Y2=0
cc_890 N_A_2026_424#_c_1412_n Q 0.00233746f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_891 N_A_2026_424#_c_1413_n Q 0.00173109f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_892 N_A_2026_424#_M1032_g Q 0.00320677f $X=11.015 $Y=2.4 $X2=0 $Y2=0
cc_893 N_A_2026_424#_c_1412_n Q 0.00138666f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_894 N_A_2026_424#_c_1413_n Q 0.00108732f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_895 N_A_2026_424#_M1032_g Q 0.0127666f $X=11.015 $Y=2.4 $X2=0 $Y2=0
cc_896 N_A_2026_424#_M1032_g N_Q_c_1753_n 0.004929f $X=11.015 $Y=2.4 $X2=0 $Y2=0
cc_897 N_A_2026_424#_M1004_g N_Q_c_1753_n 0.00406947f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_898 N_A_2026_424#_c_1412_n N_Q_c_1753_n 0.0262113f $X=10.965 $Y=1.465 $X2=0
+ $Y2=0
cc_899 N_A_2026_424#_c_1413_n N_Q_c_1753_n 0.00773673f $X=10.965 $Y=1.465 $X2=0
+ $Y2=0
cc_900 N_A_2026_424#_M1004_g N_VGND_c_1781_n 0.00357902f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_901 N_A_2026_424#_c_1410_n N_VGND_c_1781_n 0.0295846f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_902 N_A_2026_424#_c_1412_n N_VGND_c_1781_n 0.0215504f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_903 N_A_2026_424#_c_1413_n N_VGND_c_1781_n 0.00218979f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_904 N_A_2026_424#_c_1410_n N_VGND_c_1786_n 0.011066f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_905 N_A_2026_424#_M1004_g N_VGND_c_1787_n 0.00434272f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_906 N_A_2026_424#_M1004_g N_VGND_c_1788_n 0.00824463f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_907 N_A_2026_424#_c_1410_n N_VGND_c_1788_n 0.00915947f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_908 N_VPWR_c_1462_n N_A_38_78#_c_1612_n 0.0120488f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_909 N_VPWR_c_1463_n N_A_38_78#_c_1612_n 0.00940121f $X=1.18 $Y=2.835 $X2=0
+ $Y2=0
cc_910 N_VPWR_c_1471_n N_A_38_78#_c_1612_n 0.0121689f $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1460_n N_A_38_78#_c_1612_n 0.010069f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_912 N_VPWR_M1024_d N_A_38_78#_c_1614_n 0.00253448f $X=1.045 $Y=2.54 $X2=0
+ $Y2=0
cc_913 N_VPWR_M1006_d N_A_38_78#_c_1614_n 0.00435729f $X=2.055 $Y=1.935 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1463_n N_A_38_78#_c_1614_n 0.0206786f $X=1.18 $Y=2.835 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1464_n N_A_38_78#_c_1614_n 0.0164702f $X=2.19 $Y=2.835 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1471_n N_A_38_78#_c_1614_n 0.00157124f $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1472_n N_A_38_78#_c_1614_n 0.00899139f $X=2.025 $Y=3.33 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1473_n N_A_38_78#_c_1614_n 0.00915206f $X=4.44 $Y=3.33 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1460_n N_A_38_78#_c_1614_n 0.0390008f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1462_n N_A_38_78#_c_1617_n 0.00438233f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1471_n N_A_38_78#_c_1617_n 5.12731e-19 $X=1.015 $Y=3.33 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1460_n N_A_38_78#_c_1617_n 0.00111669f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1473_n N_A_38_78#_c_1618_n 0.00629782f $X=4.44 $Y=3.33 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1460_n N_A_38_78#_c_1618_n 0.00764586f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1469_n Q_N 0.0016355f $X=8.92 $Y=2.27 $X2=0 $Y2=0
cc_926 N_VPWR_c_1470_n Q_N 3.35344e-19 $X=10.79 $Y=1.985 $X2=0 $Y2=0
cc_927 N_VPWR_c_1476_n Q_N 0.0313273f $X=10.61 $Y=3.33 $X2=0 $Y2=0
cc_928 N_VPWR_c_1460_n Q_N 0.0254862f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_929 N_VPWR_c_1470_n Q 0.0456259f $X=10.79 $Y=1.985 $X2=0 $Y2=0
cc_930 N_VPWR_c_1477_n Q 0.0158876f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_931 N_VPWR_c_1460_n Q 0.0130823f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_932 N_A_38_78#_c_1606_n A_125_78# 0.00236678f $X=0.69 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_933 N_A_38_78#_c_1606_n N_VGND_c_1776_n 0.00157034f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_934 N_A_38_78#_c_1610_n N_VGND_c_1776_n 0.00465719f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_935 N_A_38_78#_c_1606_n N_VGND_c_1782_n 0.00520932f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_936 N_A_38_78#_c_1610_n N_VGND_c_1782_n 0.0131067f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_937 N_A_38_78#_c_1606_n N_VGND_c_1788_n 0.0102476f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_938 N_A_38_78#_c_1610_n N_VGND_c_1788_n 0.0117869f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_939 N_Q_N_c_1727_n N_VGND_c_1780_n 0.0296698f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_940 N_Q_N_c_1730_n N_VGND_c_1780_n 0.00439347f $X=9.37 $Y=1.985 $X2=0 $Y2=0
cc_941 N_Q_N_c_1727_n N_VGND_c_1786_n 0.0173129f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_942 N_Q_N_c_1727_n N_VGND_c_1788_n 0.0143301f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_943 Q N_VGND_c_1781_n 0.0312622f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_944 Q N_VGND_c_1787_n 0.0163488f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_945 Q N_VGND_c_1788_n 0.0134757f $X=11.195 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__sedfxbp_1.pex.spice
* Created: Wed Sep  2 12:32:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%D 2 5 9 11 12 13 17 18
r39 17 19 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.225
+ $X2=0.6 $Y2=1.06
r40 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.225 $X2=0.62 $Y2=1.225
r41 12 13 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.645 $Y=1.295
+ $X2=0.645 $Y2=1.665
r42 12 18 2.12292 $w=3.78e-07 $l=7e-08 $layer=LI1_cond $X=0.645 $Y=1.295
+ $X2=0.645 $Y2=1.225
r43 9 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.71 $Y=0.66 $X2=0.71
+ $Y2=1.06
r44 5 11 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.505 $Y=2.64
+ $X2=0.505 $Y2=1.73
r45 2 11 44.1029 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.6 $Y=1.545 $X2=0.6
+ $Y2=1.73
r46 1 17 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=0.6 $Y=1.245 $X2=0.6
+ $Y2=1.225
r47 1 2 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=0.6 $Y=1.245 $X2=0.6
+ $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_161_394# 1 2 9 13 18 23 24 25 26 27 28
+ 31 35 37 41 42 44
c109 41 0 1.83709e-19 $X=2.5 $Y=1.69
r110 42 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=1.69
+ $X2=2.5 $Y2=1.525
r111 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.69 $X2=2.5 $Y2=1.69
r112 39 41 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.5 $Y=1.95 $X2=2.5
+ $Y2=1.69
r113 38 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=2.035
+ $X2=1.8 $Y2=2.035
r114 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=2.5 $Y2=1.95
r115 37 38 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=1.885 $Y2=2.035
r116 33 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=2.12 $X2=1.8
+ $Y2=2.035
r117 33 35 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.8 $Y=2.12
+ $X2=1.8 $Y2=2.515
r118 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.875 $Y=1.11
+ $X2=1.875 $Y2=0.775
r119 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.8 $Y2=2.035
r120 27 28 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.355 $Y2=2.035
r121 25 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.71 $Y=1.195
+ $X2=1.875 $Y2=1.11
r122 25 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.71 $Y=1.195
+ $X2=1.355 $Y2=1.195
r123 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=1.615 $X2=1.19 $Y2=1.615
r124 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.19 $Y=1.95
+ $X2=1.355 $Y2=2.035
r125 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.19 $Y=1.95
+ $X2=1.19 $Y2=1.615
r126 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.19 $Y=1.28
+ $X2=1.355 $Y2=1.195
r127 20 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.19 $Y=1.28
+ $X2=1.19 $Y2=1.615
r128 18 24 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.19 $Y=1.97
+ $X2=1.19 $Y2=1.615
r129 13 48 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.59 $Y=0.775
+ $X2=2.59 $Y2=1.525
r130 7 18 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.895 $Y=2.045
+ $X2=1.19 $Y2=2.045
r131 7 9 202.129 $w=1.8e-07 $l=5.2e-07 $layer=POLY_cond $X=0.895 $Y=2.12
+ $X2=0.895 $Y2=2.64
r132 2 35 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=2.32 $X2=1.8 $Y2=2.515
r133 1 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.73
+ $Y=0.565 $X2=1.875 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%DE 3 5 6 10 11 13 14 16 17 19 21 23 25 26
+ 29 30 31
c84 17 0 1.59932e-19 $X=2.615 $Y=2.17
r85 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.615
+ $X2=1.92 $Y2=1.78
r86 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.615
+ $X2=1.92 $Y2=1.45
r87 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.615 $X2=1.92 $Y2=1.615
r88 26 30 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=1.92 $Y2=1.615
r89 22 23 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.83 $Y=1.135
+ $X2=2.09 $Y2=1.135
r90 19 21 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.705 $Y=2.245
+ $X2=2.705 $Y2=2.64
r91 18 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.115 $Y=2.17
+ $X2=2.025 $Y2=2.17
r92 17 19 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.615 $Y=2.17
+ $X2=2.705 $Y2=2.245
r93 17 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.615 $Y=2.17
+ $X2=2.115 $Y2=2.17
r94 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.09 $Y=1.06
+ $X2=2.09 $Y2=1.135
r95 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.09 $Y=1.06 $X2=2.09
+ $Y2=0.775
r96 11 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.025 $Y=2.245
+ $X2=2.025 $Y2=2.17
r97 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.025 $Y=2.245
+ $X2=2.025 $Y2=2.64
r98 10 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.01 $Y=2.095
+ $X2=2.025 $Y2=2.17
r99 10 32 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.01 $Y=2.095
+ $X2=2.01 $Y2=1.78
r100 7 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.21
+ $X2=1.83 $Y2=1.135
r101 7 31 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.83 $Y=1.21
+ $X2=1.83 $Y2=1.45
r102 5 22 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.135
+ $X2=1.83 $Y2=1.135
r103 5 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.755 $Y=1.135
+ $X2=1.175 $Y2=1.135
r104 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.1 $Y=1.06
+ $X2=1.175 $Y2=1.135
r105 1 3 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.1 $Y=1.06 $X2=1.1
+ $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_575_305# 1 2 9 13 15 17 18 19 22 28 32
+ 37 42 44 47 49 50 52 53 55 56 58 59 60 66 70 71 75 85 87
c262 66 0 8.67988e-20 $X=14.16 $Y=2.035
c263 60 0 3.4364e-19 $X=3.265 $Y=2.035
c264 56 0 1.36772e-20 $X=15.765 $Y=1.485
c265 44 0 1.78091e-19 $X=14.515 $Y=1.92
c266 13 0 1.63622e-19 $X=3.125 $Y=2.64
r267 70 73 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.045 $Y=1.69
+ $X2=3.045 $Y2=1.855
r268 70 72 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.045 $Y=1.69
+ $X2=3.045 $Y2=1.525
r269 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.69 $X2=3.04 $Y2=1.69
r270 67 87 9.23061 $w=4.58e-07 $l=3.55e-07 $layer=LI1_cond $X=14.16 $Y=2.15
+ $X2=14.515 $Y2=2.15
r271 67 85 4.03585 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=14.16 $Y=2.15
+ $X2=14.045 $Y2=2.15
r272 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=2.035
+ $X2=14.16 $Y2=2.035
r273 63 71 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.04 $Y=2.035
+ $X2=3.04 $Y2=1.69
r274 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.035
r275 60 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=2.035
+ $X2=3.12 $Y2=2.035
r276 59 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=2.035
+ $X2=14.16 $Y2=2.035
r277 59 60 13.3044 $w=1.4e-07 $l=1.075e-05 $layer=MET1_cond $X=14.015 $Y=2.035
+ $X2=3.265 $Y2=2.035
r278 56 79 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.765 $Y=1.485
+ $X2=15.765 $Y2=1.65
r279 56 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.765 $Y=1.485
+ $X2=15.765 $Y2=1.32
r280 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.765
+ $Y=1.485 $X2=15.765 $Y2=1.485
r281 53 55 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=15.355 $Y=1.485
+ $X2=15.765 $Y2=1.485
r282 52 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.27 $Y=1.32
+ $X2=15.355 $Y2=1.485
r283 51 52 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=15.27 $Y=0.425
+ $X2=15.27 $Y2=1.32
r284 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.185 $Y=0.34
+ $X2=15.27 $Y2=0.425
r285 49 50 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=15.185 $Y=0.34
+ $X2=14.6 $Y2=0.34
r286 45 87 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=14.515 $Y=2.38
+ $X2=14.515 $Y2=2.15
r287 45 47 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=14.515 $Y=2.38
+ $X2=14.515 $Y2=2.46
r288 44 87 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=14.515 $Y=1.92
+ $X2=14.515 $Y2=2.15
r289 44 58 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=14.515 $Y=1.92
+ $X2=14.515 $Y2=1.03
r290 40 58 9.56083 $w=3.93e-07 $l=1.97e-07 $layer=LI1_cond $X=14.402 $Y=0.833
+ $X2=14.402 $Y2=1.03
r291 40 42 9.2779 $w=3.93e-07 $l=3.18e-07 $layer=LI1_cond $X=14.402 $Y=0.833
+ $X2=14.402 $Y2=0.515
r292 39 50 8.32734 $w=1.7e-07 $l=2.36715e-07 $layer=LI1_cond $X=14.402 $Y=0.425
+ $X2=14.6 $Y2=0.34
r293 39 42 2.62582 $w=3.93e-07 $l=9e-08 $layer=LI1_cond $X=14.402 $Y=0.425
+ $X2=14.402 $Y2=0.515
r294 37 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.625 $Y=2.215
+ $X2=13.625 $Y2=2.38
r295 37 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.625 $Y=2.215
+ $X2=13.625 $Y2=2.05
r296 36 85 14.8931 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=13.625 $Y=2.217
+ $X2=14.045 $Y2=2.217
r297 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.625
+ $Y=2.215 $X2=13.625 $Y2=2.215
r298 32 78 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.825 $Y=0.76
+ $X2=15.825 $Y2=1.32
r299 28 79 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=15.8 $Y=2.4
+ $X2=15.8 $Y2=1.65
r300 24 75 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.68 $Y=1.015
+ $X2=13.68 $Y2=2.05
r301 22 76 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=13.58 $Y=2.75
+ $X2=13.58 $Y2=2.38
r302 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.605 $Y=0.94
+ $X2=13.68 $Y2=1.015
r303 18 19 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=13.605 $Y=0.94
+ $X2=13.215 $Y2=0.94
r304 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.14 $Y=0.865
+ $X2=13.215 $Y2=0.94
r305 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.14 $Y=0.865
+ $X2=13.14 $Y2=0.58
r306 13 73 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=3.125 $Y=2.64
+ $X2=3.125 $Y2=1.855
r307 9 72 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.98 $Y=0.775
+ $X2=2.98 $Y2=1.525
r308 2 87 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.38
+ $Y=1.96 $X2=14.515 $Y2=2.105
r309 2 47 300 $w=1.7e-07 $l=5.63471e-07 $layer=licon1_PDIFF $count=2 $X=14.38
+ $Y=1.96 $X2=14.515 $Y2=2.46
r310 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.23
+ $Y=0.37 $X2=14.37 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_667_87# 1 2 7 9 10 11 14 18 22 23 28 29
+ 33 36 39 43 46 47
r92 47 59 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.955
+ $X2=5.73 $Y2=2.12
r93 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=1.955 $X2=5.73 $Y2=1.955
r94 36 38 9.07533 $w=5.31e-07 $l=3.95e-07 $layer=LI1_cond $X=4.18 $Y=0.737
+ $X2=4.575 $Y2=0.737
r95 33 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.155 $Y=0.575
+ $X2=4.155 $Y2=0.915
r96 32 36 0.574388 $w=5.31e-07 $l=2.5e-08 $layer=LI1_cond $X=4.155 $Y=0.737
+ $X2=4.18 $Y2=0.737
r97 32 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=0.915 $X2=4.155 $Y2=0.915
r98 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=0.575 $X2=4.155 $Y2=0.575
r99 30 39 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.305 $Y=2.035
+ $X2=4.18 $Y2=2.035
r100 29 46 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=5.717 $Y=2.035
+ $X2=5.717 $Y2=1.955
r101 29 30 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.565 $Y=2.035
+ $X2=4.305 $Y2=2.035
r102 28 43 3.62566 $w=4.43e-07 $l=1.4e-07 $layer=LI1_cond $X=4.22 $Y=2.512
+ $X2=4.36 $Y2=2.512
r103 27 39 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.22 $Y=2.12
+ $X2=4.18 $Y2=2.035
r104 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.22 $Y=2.12
+ $X2=4.22 $Y2=2.29
r105 25 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=1.935 $X2=4.155 $Y2=1.935
r106 23 26 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=4.155 $Y=1.255
+ $X2=4.155 $Y2=1.935
r107 22 25 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.18 $Y=1.255
+ $X2=4.18 $Y2=1.935
r108 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=1.255 $X2=4.155 $Y2=1.255
r109 20 39 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=1.95 $X2=4.18
+ $Y2=2.035
r110 20 25 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=4.18 $Y=1.95
+ $X2=4.18 $Y2=1.935
r111 19 36 5.16051 $w=2.5e-07 $l=3.28e-07 $layer=LI1_cond $X=4.18 $Y=1.065
+ $X2=4.18 $Y2=0.737
r112 19 22 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=4.18 $Y=1.065
+ $X2=4.18 $Y2=1.255
r113 17 23 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=4.155 $Y=1.21
+ $X2=4.155 $Y2=1.255
r114 17 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.155 $Y=1.21
+ $X2=4.155 $Y2=1.135
r115 16 35 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.155 $Y=1.06
+ $X2=4.155 $Y2=0.915
r116 16 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.155 $Y=1.06
+ $X2=4.155 $Y2=1.135
r117 14 59 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=5.655 $Y=2.63
+ $X2=5.655 $Y2=2.12
r118 10 18 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=1.135
+ $X2=4.155 $Y2=1.135
r119 10 11 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.99 $Y=1.135
+ $X2=3.485 $Y2=1.135
r120 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.06
+ $X2=3.485 $Y2=1.135
r121 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.41 $Y=1.06 $X2=3.41
+ $Y2=0.775
r122 2 43 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=2.31 $X2=4.36 $Y2=2.51
r123 1 38 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.625 $X2=4.575 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%SCD 3 7 9 12
c39 12 0 7.32197e-20 $X=5.24 $Y=1.345
c40 9 0 7.28902e-20 $X=5.52 $Y=1.295
c41 3 0 9.1143e-20 $X=5.265 $Y=2.63
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.345
+ $X2=5.24 $Y2=1.51
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.345
+ $X2=5.24 $Y2=1.18
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.24
+ $Y=1.345 $X2=5.24 $Y2=1.345
r45 9 13 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.52 $Y=1.345 $X2=5.24
+ $Y2=1.345
r46 7 14 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=5.3 $Y=0.835 $X2=5.3
+ $Y2=1.18
r47 3 15 435.355 $w=1.8e-07 $l=1.12e-06 $layer=POLY_cond $X=5.265 $Y=2.63
+ $X2=5.265 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%SCE 1 3 4 5 9 13 14 15 18 20 23 24
c71 24 0 7.32197e-20 $X=4.7 $Y=1.615
c72 23 0 7.28902e-20 $X=4.7 $Y=1.615
r73 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.7 $Y=1.615
+ $X2=4.7 $Y2=1.78
r74 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.7 $Y=1.615
+ $X2=4.7 $Y2=1.45
r75 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.7
+ $Y=1.615 $X2=4.7 $Y2=1.615
r76 20 24 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.7 $Y2=1.615
r77 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.69 $Y=0.255
+ $X2=5.69 $Y2=0.835
r78 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=0.18
+ $X2=5.69 $Y2=0.255
r79 14 15 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.615 $Y=0.18
+ $X2=4.865 $Y2=0.18
r80 13 25 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.79 $Y=0.835
+ $X2=4.79 $Y2=1.45
r81 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.79 $Y=0.255
+ $X2=4.865 $Y2=0.18
r82 10 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.79 $Y=0.255
+ $X2=4.79 $Y2=0.835
r83 9 26 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.65 $Y=2.63 $X2=4.65
+ $Y2=1.78
r84 7 9 157.427 $w=1.8e-07 $l=4.05e-07 $layer=POLY_cond $X=4.65 $Y=3.035
+ $X2=4.65 $Y2=2.63
r85 4 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.56 $Y=3.11
+ $X2=4.65 $Y2=3.035
r86 4 5 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.56 $Y=3.11
+ $X2=3.665 $Y2=3.11
r87 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.575 $Y=3.035
+ $X2=3.665 $Y2=3.11
r88 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.575 $Y=3.035
+ $X2=3.575 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%CLK 3 7 8 11 13
r37 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.74 $Y=1.385
+ $X2=6.74 $Y2=1.55
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.74 $Y=1.385
+ $X2=6.74 $Y2=1.22
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.74
+ $Y=1.385 $X2=6.74 $Y2=1.385
r40 8 12 6.85236 $w=3.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.96 $Y=1.365
+ $X2=6.74 $Y2=1.365
r41 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.68 $Y=0.74 $X2=6.68
+ $Y2=1.22
r42 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.665 $Y=2.4
+ $X2=6.665 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_1549_74# 1 2 9 13 16 18 20 24 27 29 30
+ 31 37 40 41 44 45 46 48 49 50 51 53 56 59 62 64 65 68 71 75 80 84
c229 84 0 1.73561e-19 $X=12.24 $Y=1.635
c230 75 0 1.02428e-19 $X=13.23 $Y=1.39
c231 71 0 9.34686e-20 $X=13.23 $Y=1.215
c232 65 0 1.64433e-19 $X=9.535 $Y=0.935
c233 62 0 2.0055e-20 $X=8.75 $Y=2.215
c234 31 0 1.88738e-19 $X=8.585 $Y=1.98
c235 20 0 1.58205e-19 $X=13.16 $Y=2.75
r236 75 88 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.23 $Y=1.39
+ $X2=13.23 $Y2=1.555
r237 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.23
+ $Y=1.39 $X2=13.23 $Y2=1.39
r238 71 74 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=13.23 $Y=1.215
+ $X2=13.23 $Y2=1.39
r239 69 70 15.457 $w=2.21e-07 $l=2.8e-07 $layer=LI1_cond $X=12.102 $Y=0.935
+ $X2=12.102 $Y2=1.215
r240 68 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.485 $Y=1.285
+ $X2=9.485 $Y2=1.12
r241 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.485
+ $Y=1.285 $X2=9.485 $Y2=1.285
r242 65 67 16.4231 $w=2.6e-07 $l=3.5e-07 $layer=LI1_cond $X=9.535 $Y=0.935
+ $X2=9.535 $Y2=1.285
r243 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.75
+ $Y=2.215 $X2=8.75 $Y2=2.215
r244 57 70 2.27611 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=12.255 $Y=1.215
+ $X2=12.102 $Y2=1.215
r245 56 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.065 $Y=1.215
+ $X2=13.23 $Y2=1.215
r246 56 57 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=13.065 $Y=1.215
+ $X2=12.255 $Y2=1.215
r247 54 84 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=12.115 $Y=1.635
+ $X2=12.24 $Y2=1.635
r248 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.115
+ $Y=1.635 $X2=12.115 $Y2=1.635
r249 51 70 4.34639 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=12.102 $Y=1.3
+ $X2=12.102 $Y2=1.215
r250 51 53 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=12.102 $Y=1.3
+ $X2=12.102 $Y2=1.635
r251 49 69 2.27611 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.95 $Y=0.935
+ $X2=12.102 $Y2=0.935
r252 49 50 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=11.95 $Y=0.935
+ $X2=11.41 $Y2=0.935
r253 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.325 $Y=0.85
+ $X2=11.41 $Y2=0.935
r254 47 48 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=11.325 $Y=0.425
+ $X2=11.325 $Y2=0.85
r255 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.24 $Y=0.34
+ $X2=11.325 $Y2=0.425
r256 45 46 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.24 $Y=0.34
+ $X2=10.73 $Y2=0.34
r257 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.645 $Y=0.425
+ $X2=10.73 $Y2=0.34
r258 43 44 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.645 $Y=0.425
+ $X2=10.645 $Y2=0.85
r259 42 65 3.22376 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.69 $Y=0.935
+ $X2=9.535 $Y2=0.935
r260 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.56 $Y=0.935
+ $X2=10.645 $Y2=0.85
r261 41 42 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=10.56 $Y=0.935
+ $X2=9.69 $Y2=0.935
r262 40 65 4.66935 $w=2.6e-07 $l=1.09087e-07 $layer=LI1_cond $X=9.59 $Y=0.85
+ $X2=9.535 $Y2=0.935
r263 39 40 23.5682 $w=1.98e-07 $l=4.25e-07 $layer=LI1_cond $X=9.59 $Y=0.425
+ $X2=9.59 $Y2=0.85
r264 38 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.34
+ $X2=8.785 $Y2=0.34
r265 37 39 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.49 $Y=0.34
+ $X2=9.59 $Y2=0.425
r266 37 38 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=9.49 $Y=0.34
+ $X2=8.87 $Y2=0.34
r267 35 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.425
+ $X2=8.785 $Y2=0.34
r268 35 59 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.785 $Y=0.425
+ $X2=8.785 $Y2=1.82
r269 31 61 9.5026 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=8.727 $Y=1.98
+ $X2=8.727 $Y2=2.215
r270 31 59 8.33135 $w=2.83e-07 $l=1.6e-07 $layer=LI1_cond $X=8.727 $Y=1.98
+ $X2=8.727 $Y2=1.82
r271 31 33 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=8.585 $Y=1.98
+ $X2=8.28 $Y2=1.98
r272 29 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.7 $Y=0.34
+ $X2=8.785 $Y2=0.34
r273 29 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.7 $Y=0.34
+ $X2=8.05 $Y2=0.34
r274 25 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.925 $Y=0.425
+ $X2=8.05 $Y2=0.34
r275 25 27 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.925 $Y=0.425
+ $X2=7.925 $Y2=0.515
r276 24 88 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.175 $Y=2.04
+ $X2=13.175 $Y2=1.555
r277 18 24 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.16 $Y=2.13
+ $X2=13.16 $Y2=2.04
r278 18 20 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=13.16 $Y=2.13 $X2=13.16
+ $Y2=2.75
r279 14 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.24 $Y=1.47
+ $X2=12.24 $Y2=1.635
r280 14 16 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.24 $Y=1.47
+ $X2=12.24 $Y2=0.69
r281 13 80 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.4 $Y=0.8 $X2=9.4
+ $Y2=1.12
r282 7 62 63.3705 $w=2.51e-07 $l=4.04166e-07 $layer=POLY_cond $X=9.08 $Y=2.38
+ $X2=8.75 $Y2=2.215
r283 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.08 $Y=2.38 $X2=9.08
+ $Y2=2.75
r284 2 33 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=8.145
+ $Y=1.84 $X2=8.28 $Y2=2.02
r285 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.37 $X2=7.885 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_1351_74# 1 2 9 11 13 15 16 20 22 24 26
+ 30 34 37 38 39 46 48 49 51 52 58 59 60 62 65 66 67 72 73
c204 73 0 9.34686e-20 $X=12.69 $Y=1.635
c205 59 0 1.58205e-19 $X=12.425 $Y=2.475
c206 58 0 2.0055e-20 $X=9.775 $Y=2.39
c207 39 0 1.88738e-19 $X=8.66 $Y=1.727
c208 26 0 7.25971e-20 $X=9.58 $Y=2.75
c209 24 0 1.64433e-19 $X=9.58 $Y=2.255
r210 73 81 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.69 $Y=1.635
+ $X2=12.69 $Y2=1.8
r211 73 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.69 $Y=1.635
+ $X2=12.69 $Y2=1.47
r212 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.69
+ $Y=1.635 $X2=12.69 $Y2=1.635
r213 69 72 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=12.51 $Y=1.635
+ $X2=12.69 $Y2=1.635
r214 64 67 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.36 $Y=1.975 $X2=7.44
+ $Y2=1.975
r215 64 66 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.36 $Y=1.975
+ $X2=7.055 $Y2=1.975
r216 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.36
+ $Y=1.975 $X2=7.36 $Y2=1.975
r217 61 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.51 $Y=1.8
+ $X2=12.51 $Y2=1.635
r218 61 62 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.51 $Y=1.8
+ $X2=12.51 $Y2=2.39
r219 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.425 $Y=2.475
+ $X2=12.51 $Y2=2.39
r220 59 60 167.342 $w=1.68e-07 $l=2.565e-06 $layer=LI1_cond $X=12.425 $Y=2.475
+ $X2=9.86 $Y2=2.475
r221 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.775 $Y=2.39
+ $X2=9.86 $Y2=2.475
r222 57 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.775 $Y=2.22
+ $X2=9.775 $Y2=2.39
r223 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.545
+ $Y=2.09 $X2=9.545 $Y2=2.09
r224 52 57 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.69 $Y=2.09
+ $X2=9.775 $Y2=2.22
r225 52 54 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=9.69 $Y=2.09
+ $X2=9.545 $Y2=2.09
r226 51 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.44 $Y=1.81
+ $X2=7.44 $Y2=1.975
r227 50 51 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.44 $Y=1.01 $X2=7.44
+ $Y2=1.81
r228 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.355 $Y=0.925
+ $X2=7.44 $Y2=1.01
r229 48 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.355 $Y=0.925
+ $X2=7.06 $Y2=0.925
r230 44 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.895 $Y=0.84
+ $X2=7.06 $Y2=0.925
r231 44 46 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.895 $Y=0.84
+ $X2=6.895 $Y2=0.515
r232 42 66 5.94228 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=6.89 $Y=1.98
+ $X2=7.055 $Y2=1.98
r233 36 65 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.36 $Y=1.765
+ $X2=7.36 $Y2=1.975
r234 36 37 13.5877 $w=2.4e-07 $l=1.42653e-07 $layer=POLY_cond $X=7.36 $Y=1.765
+ $X2=7.47 $Y2=1.69
r235 34 80 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=12.75 $Y=0.58
+ $X2=12.75 $Y2=1.47
r236 30 81 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=12.625 $Y=2.46
+ $X2=12.625 $Y2=1.8
r237 24 55 35.4194 $w=2.55e-07 $l=1.81659e-07 $layer=POLY_cond $X=9.58 $Y=2.255
+ $X2=9.545 $Y2=2.09
r238 24 26 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=9.58 $Y=2.255
+ $X2=9.58 $Y2=2.75
r239 23 39 20.4101 $w=1.5e-07 $l=9.20598e-08 $layer=POLY_cond $X=8.735 $Y=1.765
+ $X2=8.66 $Y2=1.727
r240 22 55 61.4314 $w=2.55e-07 $l=3.99061e-07 $layer=POLY_cond $X=9.38 $Y=1.765
+ $X2=9.545 $Y2=2.09
r241 22 23 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=9.38 $Y=1.765
+ $X2=8.735 $Y2=1.765
r242 18 39 5.30422 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=8.66 $Y=1.615
+ $X2=8.66 $Y2=1.727
r243 18 20 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=8.66 $Y=1.615
+ $X2=8.66 $Y2=0.8
r244 17 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.145 $Y=1.69
+ $X2=8.055 $Y2=1.69
r245 16 39 20.4101 $w=1.5e-07 $l=9.16515e-08 $layer=POLY_cond $X=8.585 $Y=1.69
+ $X2=8.66 $Y2=1.727
r246 16 17 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.585 $Y=1.69
+ $X2=8.145 $Y2=1.69
r247 13 38 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=8.055 $Y=1.765
+ $X2=8.055 $Y2=1.69
r248 13 15 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=8.055 $Y=1.765
+ $X2=8.055 $Y2=2.4
r249 12 37 12.1617 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.745 $Y=1.69
+ $X2=7.47 $Y2=1.69
r250 11 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.965 $Y=1.69
+ $X2=8.055 $Y2=1.69
r251 11 12 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=7.965 $Y=1.69
+ $X2=7.745 $Y2=1.69
r252 7 37 13.5877 $w=2.4e-07 $l=2.34521e-07 $layer=POLY_cond $X=7.67 $Y=1.615
+ $X2=7.47 $Y2=1.69
r253 7 9 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=7.67 $Y=1.615
+ $X2=7.67 $Y2=0.74
r254 2 42 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=6.755
+ $Y=1.84 $X2=6.89 $Y2=2.02
r255 1 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.37 $X2=6.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_1972_92# 1 2 9 13 17 19 21 23 24 26 32
+ 35 38 39 43 45 46
c107 38 0 1.73561e-19 $X=11.575 $Y=1.355
r108 43 49 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.025 $Y=1.32
+ $X2=10.025 $Y2=1.485
r109 43 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.025 $Y=1.32
+ $X2=10.025 $Y2=1.155
r110 42 45 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.025 $Y=1.32
+ $X2=10.19 $Y2=1.32
r111 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.025
+ $Y=1.32 $X2=10.025 $Y2=1.32
r112 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.575
+ $Y=1.355 $X2=11.575 $Y2=1.355
r113 36 46 1.96316 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=1.355
+ $X2=10.985 $Y2=1.355
r114 36 38 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=11.07 $Y=1.355
+ $X2=11.575 $Y2=1.355
r115 34 46 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=1.52
+ $X2=10.985 $Y2=1.355
r116 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.985 $Y=1.52
+ $X2=10.985 $Y2=2.05
r117 30 46 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=1.19
+ $X2=10.985 $Y2=1.355
r118 30 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.985 $Y=1.19
+ $X2=10.985 $Y2=0.81
r119 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.9 $Y=2.135
+ $X2=10.985 $Y2=2.05
r120 26 28 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=10.9 $Y=2.135
+ $X2=10.78 $Y2=2.135
r121 24 46 1.96316 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=10.9 $Y=1.275
+ $X2=10.985 $Y2=1.355
r122 24 45 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=10.9 $Y=1.275
+ $X2=10.19 $Y2=1.275
r123 21 23 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=11.88 $Y=1.11
+ $X2=11.88 $Y2=0.69
r124 17 21 41.3657 $w=2.68e-07 $l=3.77889e-07 $layer=POLY_cond $X=11.65 $Y=1.39
+ $X2=11.88 $Y2=1.11
r125 17 39 13.4888 $w=2.68e-07 $l=7.5e-08 $layer=POLY_cond $X=11.65 $Y=1.39
+ $X2=11.575 $Y2=1.39
r126 17 19 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=11.65 $Y=1.52
+ $X2=11.65 $Y2=2.46
r127 13 49 491.718 $w=1.8e-07 $l=1.265e-06 $layer=POLY_cond $X=10.01 $Y=2.75
+ $X2=10.01 $Y2=1.485
r128 9 48 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=9.935 $Y=0.8
+ $X2=9.935 $Y2=1.155
r129 2 28 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.645
+ $Y=1.99 $X2=10.78 $Y2=2.135
r130 1 32 182 $w=1.7e-07 $l=5.11664e-07 $layer=licon1_NDIFF $count=1 $X=10.83
+ $Y=0.37 $X2=10.985 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_1747_118# 1 2 9 13 16 21 26 29 30 31 33
+ 35 40
c98 29 0 1.97671e-19 $X=9.125 $Y=1.705
r99 34 40 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=10.565 $Y=1.665
+ $X2=10.755 $Y2=1.665
r100 34 37 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=10.565 $Y=1.665
+ $X2=10.555 $Y2=1.665
r101 33 35 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=10.565 $Y=1.68
+ $X2=10.4 $Y2=1.68
r102 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.565
+ $Y=1.665 $X2=10.565 $Y2=1.665
r103 30 31 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.28 $Y=2.39
+ $X2=9.28 $Y2=2.56
r104 26 28 8.55689 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=9.18 $Y=0.785
+ $X2=9.18 $Y2=0.95
r105 24 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.21 $Y=1.705
+ $X2=9.125 $Y2=1.705
r106 24 35 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=9.21 $Y=1.705
+ $X2=10.4 $Y2=1.705
r107 21 31 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.355 $Y=2.75
+ $X2=9.355 $Y2=2.56
r108 17 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.125 $Y=1.79
+ $X2=9.125 $Y2=1.705
r109 17 30 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=9.125 $Y=1.79
+ $X2=9.125 $Y2=2.39
r110 16 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.125 $Y=1.62
+ $X2=9.125 $Y2=1.705
r111 16 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.125 $Y=1.62
+ $X2=9.125 $Y2=0.95
r112 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.755 $Y=1.5
+ $X2=10.755 $Y2=1.665
r113 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.755 $Y=1.5
+ $X2=10.755 $Y2=0.69
r114 7 37 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.555 $Y=1.83
+ $X2=10.555 $Y2=1.665
r115 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=10.555 $Y=1.83
+ $X2=10.555 $Y2=2.41
r116 2 21 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=9.17
+ $Y=2.54 $X2=9.355 $Y2=2.75
r117 1 26 182 $w=1.7e-07 $l=5.08232e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.59 $X2=9.155 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_2463_74# 1 2 9 13 15 16 17 19 20 22 27
+ 29 31 34 35 36 38 40 46 51
c151 40 0 1.02428e-19 $X=13.79 $Y=1.715
c152 27 0 1.45871e-19 $X=12.455 $Y=0.77
c153 22 0 1.78091e-19 $X=15.3 $Y=2.4
r154 55 56 19.7781 $w=3.29e-07 $l=1.35e-07 $layer=POLY_cond $X=14.155 $Y=1.365
+ $X2=14.29 $Y2=1.365
r155 52 55 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=14.13 $Y=1.365
+ $X2=14.155 $Y2=1.365
r156 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.13
+ $Y=1.365 $X2=14.13 $Y2=1.365
r157 48 51 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=13.79 $Y=1.365
+ $X2=14.13 $Y2=1.365
r158 44 46 6.76044 $w=4.58e-07 $l=2.6e-07 $layer=LI1_cond $X=12.85 $Y=2.75
+ $X2=13.11 $Y2=2.75
r159 39 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.79 $Y=1.53
+ $X2=13.79 $Y2=1.365
r160 39 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=13.79 $Y=1.53
+ $X2=13.79 $Y2=1.715
r161 38 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.79 $Y=1.2
+ $X2=13.79 $Y2=1.365
r162 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=13.79 $Y=0.94
+ $X2=13.79 $Y2=1.2
r163 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.705 $Y=1.8
+ $X2=13.79 $Y2=1.715
r164 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=13.705 $Y=1.8
+ $X2=13.195 $Y2=1.8
r165 34 46 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=13.11 $Y=2.52
+ $X2=13.11 $Y2=2.75
r166 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.11 $Y=1.885
+ $X2=13.195 $Y2=1.8
r167 33 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13.11 $Y=1.885
+ $X2=13.11 $Y2=2.52
r168 32 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.62 $Y=0.855
+ $X2=12.455 $Y2=0.855
r169 31 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.705 $Y=0.855
+ $X2=13.79 $Y2=0.94
r170 31 32 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=13.705 $Y=0.855
+ $X2=12.62 $Y2=0.855
r171 27 42 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.455 $Y=0.77
+ $X2=12.455 $Y2=0.855
r172 27 29 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=12.455 $Y=0.77
+ $X2=12.455 $Y2=0.515
r173 20 24 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=15.3 $Y=1.28
+ $X2=15.145 $Y2=1.28
r174 20 22 406.202 $w=1.8e-07 $l=1.045e-06 $layer=POLY_cond $X=15.3 $Y=1.355
+ $X2=15.3 $Y2=2.4
r175 17 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.145 $Y=1.205
+ $X2=15.145 $Y2=1.28
r176 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=15.145 $Y=1.205
+ $X2=15.145 $Y2=0.76
r177 16 56 27.6059 $w=3.29e-07 $l=1.25499e-07 $layer=POLY_cond $X=14.38 $Y=1.28
+ $X2=14.29 $Y2=1.365
r178 15 24 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.07 $Y=1.28
+ $X2=15.145 $Y2=1.28
r179 15 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=15.07 $Y=1.28
+ $X2=14.38 $Y2=1.28
r180 11 56 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=14.29 $Y=1.53
+ $X2=14.29 $Y2=1.365
r181 11 13 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=14.29 $Y=1.53
+ $X2=14.29 $Y2=2.46
r182 7 55 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.155 $Y=1.2
+ $X2=14.155 $Y2=1.365
r183 7 9 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=14.155 $Y=1.2
+ $X2=14.155 $Y2=0.69
r184 2 44 600 $w=1.7e-07 $l=8.54839e-07 $layer=licon1_PDIFF $count=1 $X=12.715
+ $Y=1.96 $X2=12.85 $Y2=2.75
r185 1 42 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=12.315
+ $Y=0.37 $X2=12.455 $Y2=0.855
r186 1 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=12.315
+ $Y=0.37 $X2=12.455 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_27_90# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 31 36 40 42 45 48
r116 37 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.2 $Y=0.645
+ $X2=0.495 $Y2=0.645
r117 36 48 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.46 $Y=2.31
+ $X2=3.365 $Y2=2.395
r118 35 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=1.345
+ $X2=3.46 $Y2=1.26
r119 35 36 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.46 $Y=1.345
+ $X2=3.46 $Y2=2.31
r120 29 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.195 $Y=1.26
+ $X2=3.46 $Y2=1.26
r121 29 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.195 $Y=1.175
+ $X2=3.195 $Y2=0.775
r122 27 48 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.185 $Y=2.395
+ $X2=3.365 $Y2=2.395
r123 27 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.185 $Y=2.395
+ $X2=2.225 $Y2=2.395
r124 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=2.48
+ $X2=2.225 $Y2=2.395
r125 25 26 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.14 $Y=2.48
+ $X2=2.14 $Y2=2.905
r126 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=2.99
+ $X2=2.14 $Y2=2.905
r127 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.055 $Y=2.99
+ $X2=1.545 $Y2=2.99
r128 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=2.905
+ $X2=1.545 $Y2=2.99
r129 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.46 $Y=2.46
+ $X2=1.46 $Y2=2.905
r130 20 42 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.375
+ $X2=0.28 $Y2=2.375
r131 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.375 $Y=2.375
+ $X2=1.46 $Y2=2.46
r132 19 20 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.375 $Y=2.375
+ $X2=0.445 $Y2=2.375
r133 15 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.46
+ $X2=0.28 $Y2=2.375
r134 15 17 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.28 $Y=2.46
+ $X2=0.28 $Y2=2.465
r135 14 42 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.29
+ $X2=0.28 $Y2=2.375
r136 13 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.2 $Y=0.81 $X2=0.2
+ $Y2=0.645
r137 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.2 $Y=0.81
+ $X2=0.2 $Y2=2.29
r138 4 48 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=3.215
+ $Y=2.32 $X2=3.35 $Y2=2.475
r139 3 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r140 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.565 $X2=3.195 $Y2=0.775
r141 1 40 182 $w=1.7e-07 $l=4.4699e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.45 $X2=0.495 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 58 62 66 68 73 78 83 88 93 98 103 108 115 116 119 122 125 128 131 134 137
+ 140 145
c180 8 0 8.67988e-20 $X=13.67 $Y=2.54
r181 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r182 141 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r183 140 143 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r184 140 141 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r185 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 131 132 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r188 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r189 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r190 122 123 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r191 119 120 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r192 116 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=15.6 $Y2=3.33
r193 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r194 113 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.69 $Y=3.33
+ $X2=15.565 $Y2=3.33
r195 113 115 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=15.69 $Y=3.33
+ $X2=16.08 $Y2=3.33
r196 112 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r197 112 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=14.16 $Y2=3.33
r198 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r199 109 140 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=14.23 $Y=3.33
+ $X2=13.935 $Y2=3.33
r200 109 111 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=14.23 $Y=3.33
+ $X2=15.12 $Y2=3.33
r201 108 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.44 $Y=3.33
+ $X2=15.565 $Y2=3.33
r202 108 111 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=15.44 $Y=3.33
+ $X2=15.12 $Y2=3.33
r203 107 143 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r204 107 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r205 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r206 104 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=3.33
+ $X2=11.34 $Y2=3.33
r207 104 106 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.505 $Y=3.33
+ $X2=11.76 $Y2=3.33
r208 103 140 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=13.64 $Y=3.33
+ $X2=13.935 $Y2=3.33
r209 103 106 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=13.64 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 102 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r211 102 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r212 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r213 99 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.41 $Y=3.33
+ $X2=10.245 $Y2=3.33
r214 99 101 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.41 $Y=3.33
+ $X2=10.8 $Y2=3.33
r215 98 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.175 $Y=3.33
+ $X2=11.34 $Y2=3.33
r216 98 101 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.175 $Y=3.33
+ $X2=10.8 $Y2=3.33
r217 97 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r218 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r219 94 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.995 $Y=3.33
+ $X2=7.83 $Y2=3.33
r220 94 96 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=7.995 $Y=3.33
+ $X2=9.84 $Y2=3.33
r221 93 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.08 $Y=3.33
+ $X2=10.245 $Y2=3.33
r222 93 96 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.08 $Y=3.33
+ $X2=9.84 $Y2=3.33
r223 92 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 92 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r225 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r226 89 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=3.33
+ $X2=6.44 $Y2=3.33
r227 89 91 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=6.605 $Y=3.33
+ $X2=7.44 $Y2=3.33
r228 88 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.83 $Y2=3.33
r229 88 91 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.44 $Y2=3.33
r230 87 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r231 87 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r232 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r233 84 125 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.08 $Y2=3.33
r234 84 86 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=6 $Y2=3.33
r235 83 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.44 $Y2=3.33
r236 83 86 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r237 82 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r238 82 123 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=2.64 $Y2=3.33
r239 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r240 79 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.52 $Y2=3.33
r241 79 81 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=4.56 $Y2=3.33
r242 78 125 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=3.33
+ $X2=5.08 $Y2=3.33
r243 78 81 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.955 $Y=3.33
+ $X2=4.56 $Y2=3.33
r244 77 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r245 77 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r246 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r247 74 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.08 $Y2=3.33
r248 74 76 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=2.16 $Y2=3.33
r249 73 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.52 $Y2=3.33
r250 73 76 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.16 $Y2=3.33
r251 71 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r252 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r253 68 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.08 $Y2=3.33
r254 68 70 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 66 97 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=9.84 $Y2=3.33
r256 66 132 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 62 65 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.565 $Y=1.985
+ $X2=15.565 $Y2=2.815
r258 60 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.565 $Y=3.245
+ $X2=15.565 $Y2=3.33
r259 60 65 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.565 $Y=3.245
+ $X2=15.565 $Y2=2.815
r260 56 140 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=13.935 $Y=3.245
+ $X2=13.935 $Y2=3.33
r261 56 58 8.71718 $w=5.88e-07 $l=4.3e-07 $layer=LI1_cond $X=13.935 $Y=3.245
+ $X2=13.935 $Y2=2.815
r262 52 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.34 $Y=3.245
+ $X2=11.34 $Y2=3.33
r263 52 54 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=11.34 $Y=3.245
+ $X2=11.34 $Y2=2.895
r264 48 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.245 $Y=3.245
+ $X2=10.245 $Y2=3.33
r265 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.245 $Y=3.245
+ $X2=10.245 $Y2=2.815
r266 44 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.83 $Y=3.245
+ $X2=7.83 $Y2=3.33
r267 44 46 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.83 $Y=3.245
+ $X2=7.83 $Y2=2.815
r268 40 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=3.33
r269 40 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.815
r270 36 125 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=3.245
+ $X2=5.08 $Y2=3.33
r271 36 38 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.08 $Y=3.245
+ $X2=5.08 $Y2=2.8
r272 32 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=3.33
r273 32 34 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=2.815
r274 28 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=3.245
+ $X2=1.08 $Y2=3.33
r275 28 30 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.08 $Y=3.245
+ $X2=1.08 $Y2=2.805
r276 9 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=15.39
+ $Y=1.84 $X2=15.525 $Y2=2.815
r277 9 62 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=15.39
+ $Y=1.84 $X2=15.525 $Y2=1.985
r278 8 58 600 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_PDIFF $count=1 $X=13.67
+ $Y=2.54 $X2=13.935 $Y2=2.815
r279 7 54 600 $w=1.7e-07 $l=1.00489e-06 $layer=licon1_PDIFF $count=1 $X=11.195
+ $Y=1.96 $X2=11.34 $Y2=2.895
r280 6 50 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=2.54 $X2=10.245 $Y2=2.815
r281 5 46 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.84 $X2=7.83 $Y2=2.815
r282 4 42 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.44 $Y2=2.815
r283 3 38 600 $w=1.7e-07 $l=6.22174e-07 $layer=licon1_PDIFF $count=1 $X=4.74
+ $Y=2.31 $X2=5.04 $Y2=2.8
r284 2 34 600 $w=1.7e-07 $l=6.52457e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=2.32 $X2=2.48 $Y2=2.815
r285 1 30 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=2.32 $X2=1.12 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%A_697_113# 1 2 3 4 5 6 21 24 25 26 28 30
+ 34 35 38 39 40 41 44 47 49 51 54 57 59 60 62 66 68
c166 62 0 9.1143e-20 $X=6.21 $Y=2.385
c167 51 0 7.25971e-20 $X=8.845 $Y=2.815
c168 26 0 1.63622e-19 $X=3.965 $Y=2.99
r169 64 66 6.26018 $w=4.03e-07 $l=2.2e-07 $layer=LI1_cond $X=5.905 $Y=0.807
+ $X2=6.125 $Y2=0.807
r170 61 62 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=2.385
+ $X2=6.21 $Y2=2.385
r171 59 61 14.3014 $w=1.88e-07 $l=2.45e-07 $layer=LI1_cond $X=5.88 $Y=2.385
+ $X2=6.125 $Y2=2.385
r172 59 60 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=2.385
+ $X2=5.715 $Y2=2.385
r173 56 57 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=3.8 $Y=1.005
+ $X2=3.8 $Y2=2.3
r174 54 56 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=3.707 $Y=0.775
+ $X2=3.707 $Y2=1.005
r175 49 51 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=8.335 $Y=2.855
+ $X2=8.845 $Y2=2.855
r176 45 47 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=8.405 $Y=1.48
+ $X2=8.405 $Y2=0.81
r177 44 49 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.25 $Y=2.73
+ $X2=8.335 $Y2=2.855
r178 43 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.25 $Y=2.48
+ $X2=8.25 $Y2=2.73
r179 42 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.945 $Y=2.395
+ $X2=7.86 $Y2=2.395
r180 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.165 $Y=2.395
+ $X2=8.25 $Y2=2.48
r181 41 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.165 $Y=2.395
+ $X2=7.945 $Y2=2.395
r182 39 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.28 $Y=1.565
+ $X2=8.405 $Y2=1.48
r183 39 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.28 $Y=1.565
+ $X2=7.945 $Y2=1.565
r184 38 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=2.31
+ $X2=7.86 $Y2=2.395
r185 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.86 $Y=1.65
+ $X2=7.945 $Y2=1.565
r186 37 38 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.86 $Y=1.65
+ $X2=7.86 $Y2=2.31
r187 35 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.775 $Y=2.395
+ $X2=7.86 $Y2=2.395
r188 35 62 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=7.775 $Y=2.395
+ $X2=6.21 $Y2=2.395
r189 34 61 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.125 $Y=2.29
+ $X2=6.125 $Y2=2.385
r190 33 66 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=6.125 $Y=1.01
+ $X2=6.125 $Y2=0.807
r191 33 34 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=6.125 $Y=1.01
+ $X2=6.125 $Y2=2.29
r192 30 60 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=4.785 $Y=2.375
+ $X2=5.715 $Y2=2.375
r193 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.7 $Y=2.46
+ $X2=4.785 $Y2=2.375
r194 27 28 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.7 $Y=2.46
+ $X2=4.7 $Y2=2.905
r195 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.615 $Y=2.99
+ $X2=4.7 $Y2=2.905
r196 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.615 $Y=2.99
+ $X2=3.965 $Y2=2.99
r197 22 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.84 $Y=2.905
+ $X2=3.965 $Y2=2.99
r198 22 24 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.84 $Y=2.905
+ $X2=3.84 $Y2=2.465
r199 21 57 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.84 $Y=2.425
+ $X2=3.84 $Y2=2.3
r200 21 24 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.84 $Y=2.425
+ $X2=3.84 $Y2=2.465
r201 6 51 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=2.54 $X2=8.845 $Y2=2.815
r202 5 59 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.745
+ $Y=2.31 $X2=5.88 $Y2=2.455
r203 4 24 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.665
+ $Y=2.32 $X2=3.8 $Y2=2.465
r204 3 47 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=8.3
+ $Y=0.59 $X2=8.445 $Y2=0.81
r205 2 64 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.625 $X2=5.905 $Y2=0.805
r206 1 54 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.565 $X2=3.695 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%Q 1 2 9 11 12 13 20
c26 9 0 1.36772e-20 $X=14.93 $Y=0.87
r27 18 20 0.525164 $w=3.93e-07 $l=1.8e-08 $layer=LI1_cond $X=15.042 $Y=2.017
+ $X2=15.042 $Y2=2.035
r28 12 13 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=15.042 $Y=2.405
+ $X2=15.042 $Y2=2.775
r29 11 18 0.991976 $w=3.93e-07 $l=3.4e-08 $layer=LI1_cond $X=15.042 $Y=1.983
+ $X2=15.042 $Y2=2.017
r30 11 29 8.56885 $w=3.93e-07 $l=1.63e-07 $layer=LI1_cond $X=15.042 $Y=1.983
+ $X2=15.042 $Y2=1.82
r31 11 12 9.83224 $w=3.93e-07 $l=3.37e-07 $layer=LI1_cond $X=15.042 $Y=2.068
+ $X2=15.042 $Y2=2.405
r32 11 20 0.962801 $w=3.93e-07 $l=3.3e-08 $layer=LI1_cond $X=15.042 $Y=2.068
+ $X2=15.042 $Y2=2.035
r33 9 29 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=14.93 $Y=0.87
+ $X2=14.93 $Y2=1.82
r34 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.93
+ $Y=1.84 $X2=15.075 $Y2=1.985
r35 2 13 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=14.93
+ $Y=1.84 $X2=15.075 $Y2=2.815
r36 1 9 182 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=1 $X=14.785
+ $Y=0.39 $X2=14.93 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%Q_N 1 2 9 13 14 15 16 23 32
r24 21 23 0.860491 $w=3.73e-07 $l=2.8e-08 $layer=LI1_cond $X=16.047 $Y=2.007
+ $X2=16.047 $Y2=2.035
r25 15 16 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=16.047 $Y=2.405
+ $X2=16.047 $Y2=2.775
r26 14 21 0.891223 $w=3.73e-07 $l=2.9e-08 $layer=LI1_cond $X=16.047 $Y=1.978
+ $X2=16.047 $Y2=2.007
r27 14 32 8.33934 $w=3.73e-07 $l=1.58e-07 $layer=LI1_cond $X=16.047 $Y=1.978
+ $X2=16.047 $Y2=1.82
r28 14 15 10.5103 $w=3.73e-07 $l=3.42e-07 $layer=LI1_cond $X=16.047 $Y=2.063
+ $X2=16.047 $Y2=2.405
r29 14 23 0.860491 $w=3.73e-07 $l=2.8e-08 $layer=LI1_cond $X=16.047 $Y=2.063
+ $X2=16.047 $Y2=2.035
r30 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.15 $Y=1.15
+ $X2=16.15 $Y2=1.82
r31 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=16.055 $Y=0.97
+ $X2=16.055 $Y2=1.15
r32 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=16.055 $Y=0.97
+ $X2=16.055 $Y2=0.535
r33 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=15.89
+ $Y=1.84 $X2=16.025 $Y2=1.985
r34 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=15.89
+ $Y=1.84 $X2=16.025 $Y2=2.815
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.9
+ $Y=0.39 $X2=16.04 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_1%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 60 63 64 66 67 68 70 79 90 94 102 107 114 115 118 121 124 127 130 135 141
+ 143
r181 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r182 140 141 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=13.87 $Y=0.257
+ $X2=14.035 $Y2=0.257
r183 137 140 3.31759 $w=6.83e-07 $l=1.9e-07 $layer=LI1_cond $X=13.68 $Y=0.257
+ $X2=13.87 $Y2=0.257
r184 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r185 134 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r186 133 137 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=13.2 $Y=0.257
+ $X2=13.68 $Y2=0.257
r187 133 135 8.00217 $w=6.83e-07 $l=1e-08 $layer=LI1_cond $X=13.2 $Y=0.257
+ $X2=13.19 $Y2=0.257
r188 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r189 131 134 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r190 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r191 127 128 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r192 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r193 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r194 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r195 115 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=15.6 $Y2=0
r196 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r197 112 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.695 $Y=0
+ $X2=15.61 $Y2=0
r198 112 114 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=15.695 $Y=0
+ $X2=16.08 $Y2=0
r199 111 144 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=15.6 $Y2=0
r200 111 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r201 110 141 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=14.16 $Y=0
+ $X2=14.035 $Y2=0
r202 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r203 107 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.525 $Y=0
+ $X2=15.61 $Y2=0
r204 107 110 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=15.525 $Y=0
+ $X2=14.16 $Y2=0
r205 106 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r206 106 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r207 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r208 103 127 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=10.227 $Y2=0
r209 103 105 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=11.28 $Y2=0
r210 102 130 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.705 $Y2=0
r211 102 105 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=11.58 $Y=0
+ $X2=11.28 $Y2=0
r212 101 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r213 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r214 98 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r215 97 100 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r216 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r217 95 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.62 $Y=0
+ $X2=7.455 $Y2=0
r218 95 97 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.92
+ $Y2=0
r219 94 127 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=10.227 $Y2=0
r220 94 100 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.065 $Y=0
+ $X2=9.84 $Y2=0
r221 93 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r222 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r223 90 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.29 $Y=0
+ $X2=7.455 $Y2=0
r224 90 92 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=6.96
+ $Y2=0
r225 89 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r226 89 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r227 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r228 86 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.24 $Y=0
+ $X2=5.075 $Y2=0
r229 86 88 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.24 $Y=0 $X2=6
+ $Y2=0
r230 85 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r231 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r232 82 85 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r233 81 84 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r234 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r235 79 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.91 $Y=0
+ $X2=5.075 $Y2=0
r236 79 84 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.91 $Y=0 $X2=4.56
+ $Y2=0
r237 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r238 78 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r239 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r240 75 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=0
+ $X2=1.315 $Y2=0
r241 75 77 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=2.16
+ $Y2=0
r242 73 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r243 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r244 70 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0
+ $X2=1.315 $Y2=0
r245 70 72 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.24
+ $Y2=0
r246 68 101 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=9.84 $Y2=0
r247 68 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=7.92 $Y2=0
r248 66 88 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.38 $Y=0 $X2=6
+ $Y2=0
r249 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=0 $X2=6.465
+ $Y2=0
r250 65 92 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.96
+ $Y2=0
r251 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.465
+ $Y2=0
r252 63 77 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.16
+ $Y2=0
r253 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.375
+ $Y2=0
r254 62 81 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.64
+ $Y2=0
r255 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.375
+ $Y2=0
r256 58 143 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.61 $Y=0.085
+ $X2=15.61 $Y2=0
r257 58 60 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=15.61 $Y=0.085
+ $X2=15.61 $Y2=0.535
r258 57 130 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.83 $Y=0
+ $X2=11.705 $Y2=0
r259 57 135 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=11.83 $Y=0
+ $X2=13.19 $Y2=0
r260 52 130 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.705 $Y=0.085
+ $X2=11.705 $Y2=0
r261 52 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.705 $Y=0.085
+ $X2=11.705 $Y2=0.515
r262 48 127 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=10.227 $Y=0.085
+ $X2=10.227 $Y2=0
r263 48 50 15.2477 $w=3.23e-07 $l=4.3e-07 $layer=LI1_cond $X=10.227 $Y=0.085
+ $X2=10.227 $Y2=0.515
r264 44 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.455 $Y=0.085
+ $X2=7.455 $Y2=0
r265 44 46 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.455 $Y=0.085
+ $X2=7.455 $Y2=0.55
r266 40 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.465 $Y=0.085
+ $X2=6.465 $Y2=0
r267 40 42 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.465 $Y=0.085
+ $X2=6.465 $Y2=0.68
r268 36 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=0.085
+ $X2=5.075 $Y2=0
r269 36 38 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.075 $Y=0.085
+ $X2=5.075 $Y2=0.805
r270 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0
r271 32 34 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0.775
r272 28 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=0.085
+ $X2=1.315 $Y2=0
r273 28 30 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.315 $Y=0.085
+ $X2=1.315 $Y2=0.66
r274 9 60 91 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=2 $X=15.22
+ $Y=0.39 $X2=15.61 $Y2=0.535
r275 8 140 91 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=2 $X=13.215
+ $Y=0.37 $X2=13.87 $Y2=0.515
r276 7 54 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.52
+ $Y=0.37 $X2=11.665 $Y2=0.515
r277 6 50 182 $w=1.7e-07 $l=2.90086e-07 $layer=licon1_NDIFF $count=1 $X=10.01
+ $Y=0.59 $X2=10.265 $Y2=0.515
r278 5 46 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=7.31
+ $Y=0.37 $X2=7.455 $Y2=0.55
r279 4 42 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=6.32
+ $Y=0.37 $X2=6.465 $Y2=0.68
r280 3 38 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.625 $X2=5.075 $Y2=0.805
r281 2 34 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.565 $X2=2.375 $Y2=0.775
r282 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.45 $X2=1.315 $Y2=0.66
.ends


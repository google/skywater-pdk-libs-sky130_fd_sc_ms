* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=7.504e+11p pd=5.82e+06u as=7.504e+11p ps=5.82e+06u
M1001 Y C1 a_469_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=2.294e+11p ps=2.1e+06u
M1002 a_141_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1003 a_128_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=7.067e+11p ps=4.87e+06u
M1004 a_225_368# A2 a_141_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1005 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_469_74# B1 a_128_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A3 a_225_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_128_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_128_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 a_563_48# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VPWR A a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_27_74# a_563_48# a_499_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 a_27_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_119_392# B a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_27_392# C a_499_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 a_563_48# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_119_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_499_392# a_563_48# a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 a_499_392# C a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X17 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_27_392# B a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X19 VGND a_563_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

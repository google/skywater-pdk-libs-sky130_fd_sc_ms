* File: sky130_fd_sc_ms__xnor2_1.pex.spice
* Created: Fri Aug 28 18:17:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XNOR2_1%B 1 3 4 6 10 14 17 18 19 21 25 26 28 40
c93 40 0 1.14536e-19 $X=1.26 $Y=1.607
c94 25 0 1.99569e-19 $X=2.3 $Y=1.515
c95 10 0 9.34955e-20 $X=2.225 $Y=2.4
c96 6 0 3.69556e-20 $X=1.065 $Y=2.345
r97 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.6 $X2=1.11 $Y2=1.6
r98 28 40 2.00425 $w=3.43e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=1.607 $X2=1.26
+ $Y2=1.607
r99 28 32 3.00637 $w=3.43e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.607 $X2=1.11
+ $Y2=1.607
r100 26 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.515
+ $X2=2.3 $Y2=1.68
r101 26 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.515
+ $X2=2.3 $Y2=1.35
r102 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.515 $X2=2.3 $Y2=1.515
r103 22 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.1 $Y=1.515 $X2=2.3
+ $Y2=1.515
r104 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=1.68 $X2=2.1
+ $Y2=1.515
r105 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.1 $Y=1.68 $X2=2.1
+ $Y2=1.95
r106 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.1 $Y2=1.95
r107 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=1.345 $Y2=2.035
r108 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.26 $Y=1.95
+ $X2=1.345 $Y2=2.035
r109 16 40 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.26 $Y=1.78
+ $X2=1.26 $Y2=1.607
r110 16 17 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.26 $Y=1.78
+ $X2=1.26 $Y2=1.95
r111 14 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.39 $Y=0.74
+ $X2=2.39 $Y2=1.35
r112 10 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.225 $Y=2.4
+ $X2=2.225 $Y2=1.68
r113 4 31 34.4492 $w=3.87e-07 $l=1.85257e-07 $layer=POLY_cond $X=1.065 $Y=1.765
+ $X2=1.022 $Y2=1.6
r114 4 6 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.065 $Y=1.765
+ $X2=1.065 $Y2=2.345
r115 1 31 54.9091 $w=3.87e-07 $l=3.68008e-07 $layer=POLY_cond $X=0.845 $Y=1.31
+ $X2=1.022 $Y2=1.6
r116 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.845 $Y=1.31
+ $X2=0.845 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_1%A 4 5 7 8 9 12 17 22 25 26
c65 26 0 1.30451e-19 $X=1.68 $Y=1.515
c66 5 0 1.14536e-19 $X=0.615 $Y=1.85
r67 25 28 39.6392 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.515
+ $X2=1.705 $Y2=1.68
r68 25 27 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.515
+ $X2=1.705 $Y2=1.35
r69 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.515 $X2=1.68 $Y2=1.515
r70 22 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.515
r71 17 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.815 $Y=0.74
+ $X2=1.815 $Y2=1.35
r72 14 17 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.815 $Y=0.255
+ $X2=1.815 $Y2=0.74
r73 12 28 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.805 $Y=2.4
+ $X2=1.805 $Y2=1.68
r74 8 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.74 $Y=0.18
+ $X2=1.815 $Y2=0.255
r75 8 9 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.74 $Y=0.18 $X2=0.56
+ $Y2=0.18
r76 5 18 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=0.615 $Y=1.775
+ $X2=0.485 $Y2=1.775
r77 5 7 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=0.615 $Y=1.85
+ $X2=0.615 $Y2=2.345
r78 2 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.485 $Y=1.7
+ $X2=0.485 $Y2=1.775
r79 2 4 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.485 $Y=1.7
+ $X2=0.485 $Y2=0.915
r80 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.485 $Y=0.255
+ $X2=0.56 $Y2=0.18
r81 1 4 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=0.255
+ $X2=0.485 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_1%A_141_385# 1 2 9 13 21 23 24 28 29 31 34
c87 34 0 1.88958e-19 $X=2.84 $Y=1.465
c88 9 0 1.99569e-19 $X=2.795 $Y=2.4
r89 34 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.465
+ $X2=2.84 $Y2=1.63
r90 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.465
+ $X2=2.84 $Y2=1.3
r91 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.465 $X2=2.84 $Y2=1.465
r92 31 33 18.887 $w=2.39e-07 $l=3.7e-07 $layer=LI1_cond $X=2.785 $Y=1.095
+ $X2=2.785 $Y2=1.465
r93 28 29 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=2.115
+ $X2=0.805 $Y2=1.95
r94 23 31 2.73298 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.635 $Y=1.095
+ $X2=2.785 $Y2=1.095
r95 23 24 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.635 $Y=1.095
+ $X2=1.225 $Y2=1.095
r96 19 24 10.0923 $w=2.09e-07 $l=1.82565e-07 $layer=LI1_cond $X=1.06 $Y=1.132
+ $X2=1.225 $Y2=1.095
r97 19 25 21.5981 $w=2.09e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=1.132
+ $X2=0.69 $Y2=1.132
r98 19 21 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.06 $Y=1.01
+ $X2=1.06 $Y2=0.74
r99 15 25 1.94907 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.69 $Y=1.255
+ $X2=0.69 $Y2=1.132
r100 15 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.69 $Y=1.255
+ $X2=0.69 $Y2=1.95
r101 13 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.82 $Y=0.74
+ $X2=2.82 $Y2=1.3
r102 9 37 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.795 $Y=2.4
+ $X2=2.795 $Y2=1.63
r103 2 28 300 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_PDIFF $count=2 $X=0.705
+ $Y=1.925 $X2=0.84 $Y2=2.115
r104 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.595 $X2=1.06 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_1%VPWR 1 2 3 12 14 15 17 20 24 26 29 31 36 45
+ 49
c47 3 0 1.37623e-19 $X=2.885 $Y=1.84
r48 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 37 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=3.33
+ $X2=1.58 $Y2=3.33
r53 37 39 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.745 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 36 48 4.61575 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.107 $Y2=3.33
r55 36 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 35 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 32 42 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.252 $Y2=3.33
r59 32 34 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=3.33
+ $X2=1.58 $Y2=3.33
r61 31 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.415 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 29 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 29 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 24 48 3.15043 $w=3.3e-07 $l=1.22327e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.107 $Y2=3.33
r66 24 26 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.3
r67 20 23 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.58 $Y=2.415 $X2=1.58
+ $Y2=2.815
r68 18 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=3.33
r69 18 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=2.815
r70 15 42 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.252 $Y2=3.33
r71 15 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.34 $Y2=2.535
r72 14 28 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=2.455
+ $X2=0.34 $Y2=2.29
r73 14 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.34 $Y=2.455 $X2=0.34
+ $Y2=2.535
r74 12 28 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=0.3 $Y=2.07 $X2=0.3
+ $Y2=2.29
r75 3 26 300 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_PDIFF $count=2 $X=2.885
+ $Y=1.84 $X2=3.02 $Y2=2.3
r76 2 23 600 $w=1.7e-07 $l=1.08183e-06 $layer=licon1_PDIFF $count=1 $X=1.155
+ $Y=1.925 $X2=1.58 $Y2=2.815
r77 2 20 600 $w=1.7e-07 $l=6.69589e-07 $layer=licon1_PDIFF $count=1 $X=1.155
+ $Y=1.925 $X2=1.58 $Y2=2.415
r78 1 17 600 $w=1.7e-07 $l=6.78638e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.925 $X2=0.34 $Y2=2.535
r79 1 12 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.925 $X2=0.34 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_1%Y 1 2 7 9 13 16 19 20 26
c37 16 0 1.37623e-19 $X=3.19 $Y=1.85
r38 20 26 6.24041 $w=6.88e-07 $l=3.6e-07 $layer=LI1_cond $X=2.16 $Y=2.635
+ $X2=2.52 $Y2=2.635
r39 16 19 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.19 $Y=1.85
+ $X2=3.19 $Y2=1.13
r40 11 19 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.125 $Y=0.98
+ $X2=3.125 $Y2=1.13
r41 11 13 17.8629 $w=2.98e-07 $l=4.65e-07 $layer=LI1_cond $X=3.125 $Y=0.98
+ $X2=3.125 $Y2=0.515
r42 10 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=1.935
+ $X2=2.52 $Y2=1.935
r43 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=1.935
+ $X2=3.19 $Y2=1.85
r44 9 10 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.105 $Y=1.935
+ $X2=2.685 $Y2=1.935
r45 8 26 5.06645 $w=3.3e-07 $l=3.45e-07 $layer=LI1_cond $X=2.52 $Y=2.29 $X2=2.52
+ $Y2=2.635
r46 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.02 $X2=2.52
+ $Y2=1.935
r47 7 8 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.52 $Y=2.02 $X2=2.52
+ $Y2=2.29
r48 2 26 300 $w=1.7e-07 $l=6.69701e-07 $layer=licon1_PDIFF $count=2 $X=2.315
+ $Y=1.84 $X2=2.52 $Y2=2.415
r49 2 18 600 $w=1.7e-07 $l=2.79106e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.84 $X2=2.52 $Y2=2.015
r50 1 13 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.37 $X2=3.06 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_1%VGND 1 2 7 9 13 15 17 27 28 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r40 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.1
+ $Y2=0
r42 25 27 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=3.12
+ $Y2=0
r43 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r44 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r45 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 18 31 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r47 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.72
+ $Y2=0
r48 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.1
+ $Y2=0
r49 17 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.68
+ $Y2=0
r50 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 15 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0.085 $X2=2.1
+ $Y2=0
r54 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.1 $Y=0.085
+ $X2=2.1 $Y2=0.37
r55 7 31 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r56 7 9 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.74
r57 2 13 182 $w=1.7e-07 $l=2.1e-07 $layer=licon1_NDIFF $count=1 $X=1.89 $Y=0.37
+ $X2=2.1 $Y2=0.37
r58 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.595 $X2=0.27 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_1%A_293_74# 1 2 7 10 15
c28 15 0 1.88958e-19 $X=2.605 $Y=0.675
r29 15 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.605 $Y=0.675
+ $X2=2.605 $Y2=0.755
r30 10 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=0.675 $X2=1.6
+ $Y2=0.755
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0.755
+ $X2=1.6 $Y2=0.755
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=0.755
+ $X2=2.605 $Y2=0.755
r33 7 8 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.44 $Y=0.755
+ $X2=1.765 $Y2=0.755
r34 2 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.37 $X2=2.605 $Y2=0.675
r35 1 10 182 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.6 $Y2=0.675
.ends


* File: sky130_fd_sc_ms__sdfstp_1.pex.spice
* Created: Fri Aug 28 18:13:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%SCE 3 7 9 13 17 21 22 23 26 27 31 34
c84 31 0 9.32299e-20 $X=0.72 $Y=1.665
c85 26 0 1.0138e-19 $X=1.955 $Y=1.425
c86 23 0 3.03849e-20 $X=1.79 $Y=1.525
r87 35 40 2.62366 $w=3.72e-07 $l=8e-08 $layer=LI1_cond $X=0.63 $Y=1.445 $X2=0.63
+ $Y2=1.525
r88 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.515
+ $Y=1.445 $X2=0.515 $Y2=1.445
r89 31 40 4.5914 $w=3.72e-07 $l=1.4e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.525
r90 27 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.425
+ $X2=1.955 $Y2=1.26
r91 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.425 $X2=1.955 $Y2=1.425
r92 24 40 5.3395 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.835 $Y=1.525
+ $X2=0.63 $Y2=1.525
r93 23 26 4.51938 $w=2.53e-07 $l=1e-07 $layer=LI1_cond $X=1.917 $Y=1.525
+ $X2=1.917 $Y2=1.425
r94 23 24 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.79 $Y=1.525
+ $X2=0.835 $Y2=1.525
r95 21 34 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.515 $Y=1.8
+ $X2=0.515 $Y2=1.445
r96 21 22 12.8678 $w=2.55e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=1.8
+ $X2=0.515 $Y2=1.875
r97 20 34 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.28
+ $X2=0.515 $Y2=1.445
r98 17 37 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.935 $Y=0.58
+ $X2=1.935 $Y2=1.26
r99 11 13 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.95 $Y=1.95 $X2=0.95
+ $Y2=2.64
r100 10 22 13.0648 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.875
+ $X2=0.515 $Y2=1.875
r101 9 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.86 $Y=1.875
+ $X2=0.95 $Y2=1.95
r102 9 10 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.86 $Y=1.875
+ $X2=0.68 $Y2=1.875
r103 7 20 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.575 $Y=0.58
+ $X2=0.575 $Y2=1.28
r104 1 22 12.8678 $w=2.55e-07 $l=8.21584e-08 $layer=POLY_cond $X=0.5 $Y=1.95
+ $X2=0.515 $Y2=1.875
r105 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.5 $Y=1.95 $X2=0.5
+ $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_27_464# 1 2 9 13 17 20 23 25 29 30 32 34
+ 35 39
c89 29 0 1.46299e-19 $X=1.955 $Y=1.995
c90 23 0 1.63837e-19 $X=1.79 $Y=2.405
c91 9 0 9.6166e-20 $X=1.115 $Y=0.58
r92 39 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.105
+ $X2=1.055 $Y2=0.94
r93 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.055
+ $Y=1.105 $X2=1.055 $Y2=1.105
r94 35 38 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.055 $Y=1.025
+ $X2=1.055 $Y2=1.105
r95 30 46 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.995
+ $X2=1.955 $Y2=2.16
r96 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.995 $X2=1.955 $Y2=1.995
r97 27 29 14.688 $w=2.53e-07 $l=3.25e-07 $layer=LI1_cond $X=1.917 $Y=2.32
+ $X2=1.917 $Y2=1.995
r98 26 32 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=1.025
+ $X2=0.305 $Y2=1.025
r99 25 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=1.025
+ $X2=1.055 $Y2=1.025
r100 25 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.89 $Y=1.025
+ $X2=0.525 $Y2=1.025
r101 24 34 2.32734 $w=1.7e-07 $l=1.42913e-07 $layer=LI1_cond $X=0.36 $Y=2.405
+ $X2=0.222 $Y2=2.395
r102 23 27 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=1.917 $Y2=2.32
r103 23 24 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.79 $Y=2.405
+ $X2=0.36 $Y2=2.405
r104 20 34 4.10697 $w=2.22e-07 $l=1.18174e-07 $layer=LI1_cond $X=0.17 $Y=2.3
+ $X2=0.222 $Y2=2.395
r105 19 32 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.17 $Y=1.11
+ $X2=0.305 $Y2=1.025
r106 19 20 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=0.17 $Y=1.11
+ $X2=0.17 $Y2=2.3
r107 15 32 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=0.94
+ $X2=0.305 $Y2=1.025
r108 15 17 9.42908 $w=4.38e-07 $l=3.6e-07 $layer=LI1_cond $X=0.305 $Y=0.94
+ $X2=0.305 $Y2=0.58
r109 13 46 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2 $Y=2.64 $X2=2
+ $Y2=2.16
r110 9 42 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.115 $Y=0.58
+ $X2=1.115 $Y2=0.94
r111 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.275 $Y2=2.465
r112 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.37 $X2=0.36 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%D 3 7 9 12 13
c40 12 0 1.37721e-19 $X=1.415 $Y=1.985
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.985
+ $X2=1.415 $Y2=2.15
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.985
+ $X2=1.415 $Y2=1.82
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.415
+ $Y=1.985 $X2=1.415 $Y2=1.985
r44 9 13 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.415 $Y2=1.985
r45 7 14 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.505 $Y=0.58
+ $X2=1.505 $Y2=1.82
r46 3 15 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=1.37 $Y=2.64 $X2=1.37
+ $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%SCD 1 3 6 10 11 12 13 17 19
c45 19 0 2.47679e-19 $X=2.68 $Y=1.985
c46 11 0 9.99223e-20 $X=2.64 $Y=1.295
c47 6 0 1.63837e-19 $X=2.42 $Y=2.64
r48 17 22 12.0163 $w=4.85e-07 $l=1.08185e-07 $layer=POLY_cond $X=2.602 $Y=1.382
+ $X2=2.677 $Y2=1.305
r49 17 19 66.5202 $w=4.85e-07 $l=6.03e-07 $layer=POLY_cond $X=2.602 $Y=1.382
+ $X2=2.602 $Y2=1.985
r50 13 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.985 $X2=2.68 $Y2=1.985
r51 12 13 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.68 $Y=1.665
+ $X2=2.68 $Y2=1.985
r52 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.68 $Y=1.295
+ $X2=2.68 $Y2=1.665
r53 11 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.305 $X2=2.68 $Y2=1.305
r54 9 19 1.65473 $w=4.85e-07 $l=1.5e-08 $layer=POLY_cond $X=2.602 $Y=2 $X2=2.602
+ $Y2=1.985
r55 9 10 38.737 $w=4.85e-07 $l=1.5e-07 $layer=POLY_cond $X=2.587 $Y=2 $X2=2.587
+ $Y2=2.15
r56 6 10 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.42 $Y=2.64 $X2=2.42
+ $Y2=2.15
r57 1 22 76.956 $w=3.4e-07 $l=5.85103e-07 $layer=POLY_cond $X=2.325 $Y=0.87
+ $X2=2.677 $Y2=1.305
r58 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.325 $Y=0.87
+ $X2=2.325 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%CLK 3 6 8 11 13
c37 6 0 9.99223e-20 $X=3.515 $Y=2.4
r38 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.385
+ $X2=3.44 $Y2=1.55
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.385
+ $X2=3.44 $Y2=1.22
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.385 $X2=3.44 $Y2=1.385
r41 8 12 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.44
+ $Y2=1.365
r42 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.515 $Y=2.4
+ $X2=3.515 $Y2=1.55
r43 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.355 $Y=0.74
+ $X2=3.355 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_800_74# 1 2 9 15 17 19 22 26 30 32 33 34
+ 35 38 39 42 44 46 47 50 51 52 54 55 56 58 59 60 63 66 69 71 79 80 85
c248 80 0 1.57372e-19 $X=5.675 $Y=1.78
c249 55 0 1.72794e-19 $X=7.775 $Y=2.055
r250 76 77 69.0876 $w=4.15e-07 $l=3.8e-07 $layer=POLY_cond $X=4.947 $Y=1.69
+ $X2=4.947 $Y2=2.07
r251 72 85 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.835 $Y=1.285
+ $X2=8.945 $Y2=1.285
r252 72 82 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.835 $Y=1.285
+ $X2=8.745 $Y2=1.285
r253 71 73 18.3241 $w=2.53e-07 $l=3.8e-07 $layer=LI1_cond $X=8.835 $Y=1.285
+ $X2=8.835 $Y2=1.665
r254 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.835
+ $Y=1.285 $X2=8.835 $Y2=1.285
r255 67 80 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.615 $Y=1.78
+ $X2=5.675 $Y2=1.78
r256 67 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.615 $Y=1.78
+ $X2=5.45 $Y2=1.78
r257 66 68 6.4562 $w=2.74e-07 $l=1.45e-07 $layer=LI1_cond $X=5.615 $Y=1.78
+ $X2=5.76 $Y2=1.78
r258 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.615
+ $Y=1.78 $X2=5.615 $Y2=1.78
r259 59 73 3.06467 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.67 $Y=1.665
+ $X2=8.835 $Y2=1.665
r260 59 60 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.67 $Y=1.665
+ $X2=7.945 $Y2=1.665
r261 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.86 $Y=1.75
+ $X2=7.945 $Y2=1.665
r262 57 58 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.86 $Y=1.75
+ $X2=7.86 $Y2=1.97
r263 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.775 $Y=2.055
+ $X2=7.86 $Y2=1.97
r264 55 56 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.775 $Y=2.055
+ $X2=7.495 $Y2=2.055
r265 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=2.14
+ $X2=7.495 $Y2=2.055
r266 53 54 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.41 $Y=2.14
+ $X2=7.41 $Y2=2.895
r267 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.325 $Y=2.98
+ $X2=7.41 $Y2=2.895
r268 51 52 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.325 $Y=2.98
+ $X2=6.815 $Y2=2.98
r269 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.73 $Y=2.895
+ $X2=6.815 $Y2=2.98
r270 49 50 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.73 $Y=2.515
+ $X2=6.73 $Y2=2.895
r271 48 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.43
+ $X2=5.76 $Y2=2.43
r272 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.645 $Y=2.43
+ $X2=6.73 $Y2=2.515
r273 47 48 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.645 $Y=2.43
+ $X2=5.845 $Y2=2.43
r274 45 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.515
+ $X2=5.76 $Y2=2.43
r275 45 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.76 $Y=2.515
+ $X2=5.76 $Y2=2.895
r276 44 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.345
+ $X2=5.76 $Y2=2.43
r277 43 68 3.52985 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=1.945
+ $X2=5.76 $Y2=1.78
r278 43 44 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.76 $Y=1.945
+ $X2=5.76 $Y2=2.345
r279 42 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=0.935
+ $X2=5.12 $Y2=1.02
r280 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.12 $Y=0.425
+ $X2=5.12 $Y2=0.935
r281 39 76 16.7516 $w=4.15e-07 $l=1.25e-07 $layer=POLY_cond $X=4.947 $Y=1.565
+ $X2=4.947 $Y2=1.69
r282 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.905
+ $Y=1.565 $X2=4.905 $Y2=1.565
r283 36 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.895 $Y=1.02
+ $X2=5.12 $Y2=1.02
r284 36 38 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=4.895 $Y=1.105
+ $X2=4.895 $Y2=1.565
r285 34 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.675 $Y=2.98
+ $X2=5.76 $Y2=2.895
r286 34 35 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=5.675 $Y=2.98
+ $X2=4.275 $Y2=2.98
r287 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=0.34
+ $X2=5.12 $Y2=0.425
r288 32 33 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.035 $Y=0.34
+ $X2=4.225 $Y2=0.34
r289 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=2.895
+ $X2=4.275 $Y2=2.98
r290 28 30 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.19 $Y=2.895
+ $X2=4.19 $Y2=2.78
r291 24 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.1 $Y=0.425
+ $X2=4.225 $Y2=0.34
r292 24 26 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.1 $Y=0.425 $X2=4.1
+ $Y2=0.515
r293 20 85 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.45
+ $X2=8.945 $Y2=1.285
r294 20 22 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=8.945 $Y=1.45
+ $X2=8.945 $Y2=2.08
r295 17 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.745 $Y=1.12
+ $X2=8.745 $Y2=1.285
r296 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.745 $Y=1.12
+ $X2=8.745 $Y2=0.69
r297 13 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.615
+ $X2=5.675 $Y2=1.78
r298 13 15 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.675 $Y=1.615
+ $X2=5.675 $Y2=0.615
r299 12 76 26.7644 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.155 $Y=1.69
+ $X2=4.947 $Y2=1.69
r300 12 79 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.155 $Y=1.69
+ $X2=5.45 $Y2=1.69
r301 9 77 165.202 $w=1.8e-07 $l=4.25e-07 $layer=POLY_cond $X=5.065 $Y=2.495
+ $X2=5.065 $Y2=2.07
r302 2 30 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.84 $X2=4.19 $Y2=2.78
r303 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4 $Y=0.37
+ $X2=4.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_1198_55# 1 2 7 9 12 15 16 18 22 25 30 37
+ 44 47
c93 25 0 3.13028e-19 $X=6.18 $Y=1.96
c94 18 0 3.34354e-20 $X=6.675 $Y=0.945
c95 12 0 1.83013e-19 $X=6.08 $Y=2.495
r96 37 39 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.84 $Y=0.8
+ $X2=6.84 $Y2=0.945
r97 34 47 16.6207 $w=2.61e-07 $l=9e-08 $layer=POLY_cond $X=6.36 $Y=1.1 $X2=6.27
+ $Y2=1.1
r98 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.36
+ $Y=1.1 $X2=6.36 $Y2=1.1
r99 30 33 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=6.36 $Y=0.945
+ $X2=6.36 $Y2=1.1
r100 26 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.18 $Y=1.96 $X2=6.27
+ $Y2=1.96
r101 26 41 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.18 $Y=1.96 $X2=6.08
+ $Y2=1.96
r102 25 28 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.18 $Y=1.96
+ $X2=6.18 $Y2=2.09
r103 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=1.96 $X2=6.18 $Y2=1.96
r104 20 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.07 $Y=2.175
+ $X2=7.07 $Y2=2.495
r105 19 30 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.48 $Y=0.945
+ $X2=6.36 $Y2=0.945
r106 18 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0.945
+ $X2=6.84 $Y2=0.945
r107 18 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=0.945
+ $X2=6.48 $Y2=0.945
r108 17 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=2.09
+ $X2=6.18 $Y2=2.09
r109 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.985 $Y=2.09
+ $X2=7.07 $Y2=2.175
r110 16 17 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.985 $Y=2.09
+ $X2=6.345 $Y2=2.09
r111 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.795
+ $X2=6.27 $Y2=1.96
r112 14 47 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.265
+ $X2=6.27 $Y2=1.1
r113 14 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.27 $Y=1.265
+ $X2=6.27 $Y2=1.795
r114 10 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.08 $Y=2.125
+ $X2=6.08 $Y2=1.96
r115 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=6.08 $Y=2.125
+ $X2=6.08 $Y2=2.495
r116 7 47 37.8582 $w=2.61e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.065 $Y=0.935
+ $X2=6.27 $Y2=1.1
r117 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.065 $Y=0.935
+ $X2=6.065 $Y2=0.615
r118 2 22 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=6.905
+ $Y=2.285 $X2=7.07 $Y2=2.495
r119 1 37 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.59 $X2=6.84 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_998_81# 1 2 9 13 15 18 20 22 25 31 33 34
+ 35 39 41 48 49 51 55 60 62 64 69
c164 60 0 1.55656e-19 $X=6.77 $Y=1.67
c165 48 0 1.83013e-19 $X=5.34 $Y=2.495
c166 39 0 1.72794e-19 $X=7.905 $Y=1.265
c167 13 0 3.34354e-20 $X=7.055 $Y=1.09
r168 60 65 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.67
+ $X2=6.77 $Y2=1.835
r169 60 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.67
+ $X2=6.77 $Y2=1.505
r170 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.67 $X2=6.77 $Y2=1.67
r171 51 53 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.985 $Y=1.36
+ $X2=5.985 $Y2=1.52
r172 48 49 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.34 $Y=2.495
+ $X2=5.34 $Y2=2.265
r173 42 69 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.265 $Y=1.285
+ $X2=8.355 $Y2=1.285
r174 42 66 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=8.265 $Y=1.285
+ $X2=7.975 $Y2=1.285
r175 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.265
+ $Y=1.285 $X2=8.265 $Y2=1.285
r176 39 62 6.93634 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=7.905 $Y=1.265
+ $X2=7.76 $Y2=1.265
r177 39 41 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.905 $Y=1.265
+ $X2=8.265 $Y2=1.265
r178 38 55 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=6.935 $Y=1.285
+ $X2=6.792 $Y2=1.285
r179 38 62 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=6.935 $Y=1.285
+ $X2=7.76 $Y2=1.285
r180 36 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=1.52
+ $X2=5.985 $Y2=1.52
r181 35 59 6.06549 $w=2.83e-07 $l=1.5e-07 $layer=LI1_cond $X=6.792 $Y=1.52
+ $X2=6.792 $Y2=1.67
r182 35 55 9.5026 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=6.792 $Y=1.52
+ $X2=6.792 $Y2=1.285
r183 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.65 $Y=1.52
+ $X2=6.07 $Y2=1.52
r184 33 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=1.36
+ $X2=5.985 $Y2=1.36
r185 33 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.9 $Y=1.36
+ $X2=5.625 $Y2=1.36
r186 29 34 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.5 $Y=1.36
+ $X2=5.625 $Y2=1.36
r187 29 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.5 $Y=1.36
+ $X2=5.26 $Y2=1.36
r188 29 31 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=5.5 $Y=1.275
+ $X2=5.5 $Y2=0.615
r189 27 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.26 $Y=1.445
+ $X2=5.26 $Y2=1.36
r190 27 49 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.26 $Y=1.445
+ $X2=5.26 $Y2=2.265
r191 23 25 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.83 $Y=1.165
+ $X2=7.055 $Y2=1.165
r192 20 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.355 $Y=1.12
+ $X2=8.355 $Y2=1.285
r193 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.355 $Y=1.12
+ $X2=8.355 $Y2=0.69
r194 16 66 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.975 $Y=1.45
+ $X2=7.975 $Y2=1.285
r195 16 18 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=7.975 $Y=1.45
+ $X2=7.975 $Y2=2.205
r196 13 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.055 $Y=1.09
+ $X2=7.055 $Y2=1.165
r197 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.055 $Y=1.09
+ $X2=7.055 $Y2=0.8
r198 11 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.83 $Y=1.24
+ $X2=6.83 $Y2=1.165
r199 11 64 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=6.83 $Y=1.24
+ $X2=6.83 $Y2=1.505
r200 9 65 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.815 $Y=2.495
+ $X2=6.815 $Y2=1.835
r201 2 48 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=2.285 $X2=5.34 $Y2=2.495
r202 1 31 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.405 $X2=5.46 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%SET_B 3 7 11 15 19 20 21 22 27 30 33 34 41
r128 33 36 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=7.332 $Y=1.67
+ $X2=7.332 $Y2=1.835
r129 33 35 48.8634 $w=3.75e-07 $l=1.9e-07 $layer=POLY_cond $X=7.332 $Y=1.67
+ $X2=7.332 $Y2=1.48
r130 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.67 $X2=7.31 $Y2=1.67
r131 30 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.865
+ $Y=1.545 $X2=10.865 $Y2=1.545
r132 27 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=1.665
+ $X2=10.8 $Y2=1.665
r133 24 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=1.665
r134 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.665
+ $X2=7.44 $Y2=1.665
r135 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=1.665
+ $X2=10.8 $Y2=1.665
r136 21 22 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.655 $Y=1.665
+ $X2=7.585 $Y2=1.665
r137 19 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=10.865 $Y=1.885
+ $X2=10.865 $Y2=1.545
r138 19 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.865 $Y=1.885
+ $X2=10.865 $Y2=2.05
r139 18 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.865 $Y=1.38
+ $X2=10.865 $Y2=1.545
r140 15 20 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=10.94 $Y=2.75
+ $X2=10.94 $Y2=2.05
r141 11 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=10.775 $Y=0.58
+ $X2=10.775 $Y2=1.38
r142 7 35 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.445 $Y=0.8
+ $X2=7.445 $Y2=1.48
r143 3 36 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.295 $Y=2.495
+ $X2=7.295 $Y2=1.835
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_599_74# 1 2 9 13 16 18 20 21 22 23 24 27
+ 31 33 37 39 40 44 47 49 51 54 57 58 59 64 67 71
c181 51 0 1.19062e-19 $X=9.497 $Y=1.795
c182 31 0 1.37453e-19 $X=5.565 $Y=2.495
r183 68 69 5.96904 $w=3.23e-07 $l=4e-08 $layer=POLY_cond $X=3.925 $Y=1.515
+ $X2=3.965 $Y2=1.515
r184 65 71 60.4365 $w=3.23e-07 $l=4.05e-07 $layer=POLY_cond $X=4.05 $Y=1.515
+ $X2=4.455 $Y2=1.515
r185 65 69 12.6842 $w=3.23e-07 $l=8.5e-08 $layer=POLY_cond $X=4.05 $Y=1.515
+ $X2=3.965 $Y2=1.515
r186 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r187 62 64 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.515
r188 59 61 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.145 $Y=1.945
+ $X2=3.29 $Y2=1.945
r189 58 62 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=4.05 $Y2=1.82
r190 58 61 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=3.29 $Y2=1.945
r191 57 59 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.06 $Y=1.82
+ $X2=3.145 $Y2=1.945
r192 57 67 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.06 $Y=1.82
+ $X2=3.06 $Y2=1.01
r193 52 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0.845
+ $X2=3.14 $Y2=1.01
r194 52 54 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.14 $Y=0.845
+ $X2=3.14 $Y2=0.515
r195 45 47 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.455 $Y=2.385
+ $X2=4.545 $Y2=2.385
r196 44 51 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.505 $Y=2.37
+ $X2=9.505 $Y2=1.795
r197 42 44 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=9.505 $Y=3.075
+ $X2=9.505 $Y2=2.37
r198 40 51 33.4908 $w=1.95e-07 $l=9.7e-08 $layer=POLY_cond $X=9.497 $Y=1.698
+ $X2=9.497 $Y2=1.795
r199 39 50 36.6888 $w=1.95e-07 $l=9.7e-08 $layer=POLY_cond $X=9.497 $Y=1.507
+ $X2=9.497 $Y2=1.41
r200 39 40 64.9551 $w=1.95e-07 $l=1.91e-07 $layer=POLY_cond $X=9.497 $Y=1.507
+ $X2=9.497 $Y2=1.698
r201 37 50 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.475 $Y=0.58
+ $X2=9.475 $Y2=1.41
r202 34 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.655 $Y=3.15
+ $X2=5.565 $Y2=3.15
r203 33 42 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.415 $Y=3.15
+ $X2=9.505 $Y2=3.075
r204 33 34 1928 $w=1.5e-07 $l=3.76e-06 $layer=POLY_cond $X=9.415 $Y=3.15
+ $X2=5.655 $Y2=3.15
r205 29 49 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.565 $Y=3.075
+ $X2=5.565 $Y2=3.15
r206 29 31 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=5.565 $Y=3.075
+ $X2=5.565 $Y2=2.495
r207 25 27 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.915 $Y=1.04
+ $X2=4.915 $Y2=0.615
r208 23 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.475 $Y=3.15
+ $X2=5.565 $Y2=3.15
r209 23 24 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=5.475 $Y=3.15
+ $X2=4.62 $Y2=3.15
r210 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=1.115
+ $X2=4.915 $Y2=1.04
r211 21 22 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=4.84 $Y=1.115
+ $X2=4.53 $Y2=1.115
r212 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.545 $Y=3.075
+ $X2=4.62 $Y2=3.15
r213 19 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.545 $Y=2.46
+ $X2=4.545 $Y2=2.385
r214 19 20 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.545 $Y=2.46
+ $X2=4.545 $Y2=3.075
r215 18 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.455 $Y=2.31
+ $X2=4.455 $Y2=2.385
r216 17 71 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.68
+ $X2=4.455 $Y2=1.515
r217 17 18 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.455 $Y=1.68
+ $X2=4.455 $Y2=2.31
r218 16 71 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.35
+ $X2=4.455 $Y2=1.515
r219 15 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.53 $Y2=1.115
r220 15 16 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.455 $Y2=1.35
r221 11 69 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.68
+ $X2=3.965 $Y2=1.515
r222 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.965 $Y=1.68
+ $X2=3.965 $Y2=2.4
r223 7 68 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=1.515
r224 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=3.925 $Y2=0.74
r225 2 61 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=1.84 $X2=3.29 $Y2=1.985
r226 1 54 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.995
+ $Y=0.37 $X2=3.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_1958_48# 1 2 7 9 14 15 16 19 23 27 32 34
+ 35 36 37 41
r91 36 37 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=11.74 $Y=2.22
+ $X2=11.74 $Y2=2.39
r92 33 41 11.2481 $w=4.45e-07 $l=9e-08 $layer=POLY_cond $X=10.295 $Y=1.087
+ $X2=10.385 $Y2=1.087
r93 32 34 6.83261 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.295 $Y=1.145
+ $X2=10.46 $Y2=1.145
r94 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.295
+ $Y=1.145 $X2=10.295 $Y2=1.145
r95 29 35 4.47619 $w=2.72e-07 $l=5.63383e-07 $layer=LI1_cond $X=11.855 $Y=1.21
+ $X2=11.395 $Y2=0.98
r96 29 36 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=11.855 $Y=1.21
+ $X2=11.855 $Y2=2.22
r97 27 37 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=11.705 $Y=2.75
+ $X2=11.705 $Y2=2.39
r98 21 35 4.47619 $w=2.72e-07 $l=1.87e-07 $layer=LI1_cond $X=11.582 $Y=0.98
+ $X2=11.395 $Y2=0.98
r99 21 23 12.2927 $w=3.73e-07 $l=4e-07 $layer=LI1_cond $X=11.582 $Y=0.98
+ $X2=11.582 $Y2=0.58
r100 19 35 1.95968 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=11.395 $Y=1.095
+ $X2=11.395 $Y2=0.98
r101 19 34 46.8493 $w=2.28e-07 $l=9.35e-07 $layer=LI1_cond $X=11.395 $Y=1.095
+ $X2=10.46 $Y2=1.095
r102 15 16 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=10.445 $Y=2.29
+ $X2=10.445 $Y2=2.44
r103 14 16 83.0111 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=10.49 $Y=2.75
+ $X2=10.49 $Y2=2.44
r104 10 41 28.4889 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=10.385 $Y=1.31
+ $X2=10.385 $Y2=1.087
r105 10 15 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=10.385 $Y=1.31
+ $X2=10.385 $Y2=2.29
r106 7 33 53.7407 $w=4.45e-07 $l=4.3e-07 $layer=POLY_cond $X=9.865 $Y=1.087
+ $X2=10.295 $Y2=1.087
r107 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.865 $Y=0.865
+ $X2=9.865 $Y2=0.58
r108 2 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=2.54 $X2=11.705 $Y2=2.75
r109 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.42
+ $Y=0.37 $X2=11.56 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_1764_74# 1 2 3 12 14 15 16 18 22 26 28 30
+ 33 34 35 41 44 45 48 49 50 53 57 58 61 63 66 67 68
c150 41 0 1.19062e-19 $X=9.275 $Y=2.015
r151 63 65 15.4168 $w=5.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.08 $Y=0.515
+ $X2=9.08 $Y2=0.94
r152 61 67 3.46198 $w=2.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=11.285 $Y=2.22
+ $X2=11.185 $Y2=2.305
r153 61 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.285 $Y=2.22
+ $X2=11.285 $Y2=2.05
r154 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.435
+ $Y=1.545 $X2=11.435 $Y2=1.545
r155 55 68 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=11.4 $Y=1.85 $X2=11.4
+ $Y2=2.05
r156 55 57 8.78738 $w=3.98e-07 $l=3.05e-07 $layer=LI1_cond $X=11.4 $Y=1.85
+ $X2=11.4 $Y2=1.545
r157 51 67 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.185 $Y=2.39
+ $X2=11.185 $Y2=2.305
r158 51 53 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.185 $Y=2.39
+ $X2=11.185 $Y2=2.75
r159 49 67 3.05049 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=11 $Y=2.305
+ $X2=11.185 $Y2=2.305
r160 49 50 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=11 $Y=2.305
+ $X2=10.235 $Y2=2.305
r161 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.15 $Y=2.22
+ $X2=10.235 $Y2=2.305
r162 47 48 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.15 $Y=1.79
+ $X2=10.15 $Y2=2.22
r163 46 66 2.32734 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=9.365 $Y=1.705
+ $X2=9.227 $Y2=1.705
r164 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.065 $Y=1.705
+ $X2=10.15 $Y2=1.79
r165 45 46 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=10.065 $Y=1.705
+ $X2=9.365 $Y2=1.705
r166 44 66 4.10697 $w=2.22e-07 $l=1.08305e-07 $layer=LI1_cond $X=9.28 $Y=1.62
+ $X2=9.227 $Y2=1.705
r167 44 65 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.28 $Y=1.62
+ $X2=9.28 $Y2=0.94
r168 39 66 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=9.227 $Y=1.79
+ $X2=9.227 $Y2=1.705
r169 39 41 9.42908 $w=2.73e-07 $l=2.25e-07 $layer=LI1_cond $X=9.227 $Y=1.79
+ $X2=9.227 $Y2=2.015
r170 33 58 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=11.435 $Y=1.79
+ $X2=11.435 $Y2=1.545
r171 32 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.435 $Y=1.38
+ $X2=11.435 $Y2=1.545
r172 28 36 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.92 $Y=1.865
+ $X2=12.75 $Y2=1.865
r173 28 30 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=12.92 $Y=1.94
+ $X2=12.92 $Y2=2.435
r174 24 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.75 $Y=1.79
+ $X2=12.75 $Y2=1.865
r175 24 26 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=12.75 $Y=1.79
+ $X2=12.75 $Y2=0.835
r176 23 35 15.6241 $w=2.05e-07 $l=9.87421e-08 $layer=POLY_cond $X=12.02 $Y=1.865
+ $X2=11.945 $Y2=1.92
r177 22 36 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.675 $Y=1.865
+ $X2=12.75 $Y2=1.865
r178 22 23 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=12.675 $Y=1.865
+ $X2=12.02 $Y2=1.865
r179 20 35 9.82985 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=11.945 $Y=2.05
+ $X2=11.945 $Y2=1.92
r180 20 34 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.945 $Y=2.05
+ $X2=11.945 $Y2=2.29
r181 16 34 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.93 $Y=2.38
+ $X2=11.93 $Y2=2.29
r182 16 18 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=11.93 $Y=2.38
+ $X2=11.93 $Y2=2.75
r183 15 33 27.4267 $w=2.6e-07 $l=2.20624e-07 $layer=POLY_cond $X=11.6 $Y=1.92
+ $X2=11.435 $Y2=1.79
r184 14 35 15.6241 $w=2.05e-07 $l=7.5e-08 $layer=POLY_cond $X=11.87 $Y=1.92
+ $X2=11.945 $Y2=1.92
r185 14 15 64.5024 $w=2.6e-07 $l=2.7e-07 $layer=POLY_cond $X=11.87 $Y=1.92
+ $X2=11.6 $Y2=1.92
r186 12 32 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=11.345 $Y=0.58
+ $X2=11.345 $Y2=1.38
r187 3 53 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.03
+ $Y=2.54 $X2=11.165 $Y2=2.75
r188 2 41 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=9.035
+ $Y=1.87 $X2=9.275 $Y2=2.015
r189 1 63 91 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=2 $X=8.82
+ $Y=0.37 $X2=9.07 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_2395_112# 1 2 7 9 12 19 24 28 33 34 36 37
+ 41
r62 40 41 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=13.33 $Y=1.385
+ $X2=13.425 $Y2=1.385
r63 32 34 2.05777 $w=4.63e-07 $l=8e-08 $layer=LI1_cond $X=12.535 $Y=0.772
+ $X2=12.615 $Y2=0.772
r64 32 33 5.26869 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=12.535 $Y=0.772
+ $X2=12.37 $Y2=0.772
r65 29 40 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=13.23 $Y=1.385
+ $X2=13.33 $Y2=1.385
r66 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.23
+ $Y=1.385 $X2=13.23 $Y2=1.385
r67 26 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.7 $Y=1.385
+ $X2=12.615 $Y2=1.385
r68 26 28 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=12.7 $Y=1.385
+ $X2=13.23 $Y2=1.385
r69 24 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.695 $Y=2.16
+ $X2=12.695 $Y2=1.995
r70 20 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.615 $Y=1.55
+ $X2=12.615 $Y2=1.385
r71 20 37 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=12.615 $Y=1.55
+ $X2=12.615 $Y2=1.995
r72 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.615 $Y=1.22
+ $X2=12.615 $Y2=1.385
r73 18 34 6.7035 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=12.615 $Y=1.005
+ $X2=12.615 $Y2=0.772
r74 18 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=12.615 $Y=1.005
+ $X2=12.615 $Y2=1.22
r75 16 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=12.12 $Y=0.705
+ $X2=12.37 $Y2=0.705
r76 10 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.425 $Y=1.55
+ $X2=13.425 $Y2=1.385
r77 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=13.425 $Y=1.55
+ $X2=13.425 $Y2=2.4
r78 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.33 $Y=1.22
+ $X2=13.33 $Y2=1.385
r79 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.33 $Y=1.22 $X2=13.33
+ $Y2=0.74
r80 2 24 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.56
+ $Y=2.015 $X2=12.695 $Y2=2.16
r81 1 32 182 $w=1.7e-07 $l=6.85857e-07 $layer=licon1_NDIFF $count=1 $X=11.975
+ $Y=0.56 $X2=12.535 $Y2=0.84
r82 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.975
+ $Y=0.56 $X2=12.12 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49
+ 53 57 60 61 63 64 66 67 69 70 71 73 78 108 114 115 118 121 124 127
r156 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r157 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r158 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r160 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r161 115 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r162 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r163 112 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.36 $Y=3.33
+ $X2=13.195 $Y2=3.33
r164 112 114 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.36 $Y=3.33
+ $X2=13.68 $Y2=3.33
r165 111 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r166 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r167 108 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.03 $Y=3.33
+ $X2=13.195 $Y2=3.33
r168 108 110 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.03 $Y=3.33
+ $X2=12.72 $Y2=3.33
r169 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r170 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r171 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r172 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r173 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r174 101 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r175 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r176 98 101 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r177 97 100 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r178 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r180 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r181 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r182 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r183 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r184 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r185 86 89 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r186 86 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r187 85 88 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r188 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 83 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.74 $Y2=3.33
r190 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.08 $Y2=3.33
r191 82 122 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 82 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 79 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r195 79 81 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=1.2 $Y2=3.33
r196 78 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.73 $Y2=3.33
r197 78 81 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 76 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r199 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r200 73 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r201 73 75 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r202 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r203 71 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r204 69 106 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.07 $Y=3.33
+ $X2=11.76 $Y2=3.33
r205 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.07 $Y=3.33
+ $X2=12.195 $Y2=3.33
r206 68 110 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=12.32 $Y=3.33
+ $X2=12.72 $Y2=3.33
r207 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.32 $Y=3.33
+ $X2=12.195 $Y2=3.33
r208 67 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.715 $Y=3.33
+ $X2=10.8 $Y2=3.33
r209 66 100 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.32 $Y2=3.33
r210 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.715 $Y2=3.33
r211 63 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.44 $Y2=3.33
r212 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.665 $Y=3.33
+ $X2=7.79 $Y2=3.33
r213 62 97 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.915 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.915 $Y=3.33
+ $X2=7.79 $Y2=3.33
r215 60 88 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6 $Y2=3.33
r216 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6.35 $Y2=3.33
r217 59 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.475 $Y=3.33
+ $X2=6.48 $Y2=3.33
r218 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.475 $Y=3.33
+ $X2=6.35 $Y2=3.33
r219 55 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.195 $Y=3.245
+ $X2=13.195 $Y2=3.33
r220 55 57 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=13.195 $Y=3.245
+ $X2=13.195 $Y2=2.16
r221 51 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.195 $Y=3.245
+ $X2=12.195 $Y2=3.33
r222 51 53 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=12.195 $Y=3.245
+ $X2=12.195 $Y2=2.77
r223 47 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.715 $Y=3.245
+ $X2=10.715 $Y2=3.33
r224 47 49 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=10.715 $Y=3.245
+ $X2=10.715 $Y2=2.77
r225 43 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.79 $Y=3.245
+ $X2=7.79 $Y2=3.33
r226 43 45 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=7.79 $Y=3.245
+ $X2=7.79 $Y2=2.515
r227 39 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.35 $Y=3.245
+ $X2=6.35 $Y2=3.33
r228 39 41 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.35 $Y=3.245
+ $X2=6.35 $Y2=2.85
r229 35 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=3.33
r230 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=2.78
r231 34 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.73 $Y2=3.33
r232 33 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.74 $Y2=3.33
r233 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=2.895 $Y2=3.33
r234 29 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=3.33
r235 29 31 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=2.995
r236 25 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r237 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.78
r238 8 57 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=13.01
+ $Y=2.015 $X2=13.195 $Y2=2.16
r239 7 53 600 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=2.54 $X2=12.155 $Y2=2.77
r240 6 49 600 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_PDIFF $count=1 $X=10.58
+ $Y=2.54 $X2=10.715 $Y2=2.77
r241 5 45 600 $w=1.7e-07 $l=4.6602e-07 $layer=licon1_PDIFF $count=1 $X=7.385
+ $Y=2.285 $X2=7.75 $Y2=2.515
r242 4 41 600 $w=1.7e-07 $l=6.65977e-07 $layer=licon1_PDIFF $count=1 $X=6.17
+ $Y=2.285 $X2=6.39 $Y2=2.85
r243 3 37 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.84 $X2=3.74 $Y2=2.78
r244 2 31 600 $w=1.7e-07 $l=7.77255e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=2.32 $X2=2.73 $Y2=2.995
r245 1 27 600 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=2.32 $X2=0.725 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_292_464# 1 2 3 4 13 19 21 22 24 25 30 31
+ 34 41 44 46
c126 46 0 1.37453e-19 $X=4.84 $Y=2.495
c127 24 0 4.44907e-20 $X=2.3 $Y=2.49
c128 22 0 9.6166e-20 $X=1.885 $Y=1.005
r129 38 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.53 $Y=0.68
+ $X2=4.7 $Y2=0.68
r130 34 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.32 $Y=2.325
+ $X2=3.32 $Y2=2.575
r131 30 46 7.64504 $w=4.83e-07 $l=3.1e-07 $layer=LI1_cond $X=4.53 $Y=2.482
+ $X2=4.84 $Y2=2.482
r132 30 44 7.45324 $w=4.83e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=2.482
+ $X2=4.445 $Y2=2.482
r133 29 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.765
+ $X2=4.53 $Y2=0.68
r134 29 30 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=4.53 $Y=0.765
+ $X2=4.53 $Y2=2.24
r135 28 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=2.325
+ $X2=3.32 $Y2=2.325
r136 28 44 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.405 $Y=2.325
+ $X2=4.445 $Y2=2.325
r137 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.575
+ $X2=2.3 $Y2=2.575
r138 25 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=2.575
+ $X2=3.32 $Y2=2.575
r139 25 26 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=3.235 $Y=2.575
+ $X2=2.385 $Y2=2.575
r140 24 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.575
r141 23 24 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.3 $Y=1.09 $X2=2.3
+ $Y2=2.49
r142 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=2.3 $Y2=1.09
r143 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=1.885 $Y2=1.005
r144 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.72 $Y=0.92
+ $X2=1.885 $Y2=1.005
r145 17 19 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.72 $Y=0.92
+ $X2=1.72 $Y2=0.58
r146 13 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.3 $Y=2.785
+ $X2=2.3 $Y2=2.575
r147 13 15 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=2.215 $Y=2.785
+ $X2=1.685 $Y2=2.785
r148 4 46 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=2.285 $X2=4.84 $Y2=2.495
r149 3 15 600 $w=1.7e-07 $l=5.25595e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=2.32 $X2=1.685 $Y2=2.745
r150 2 41 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=0.405 $X2=4.7 $Y2=0.68
r151 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.37 $X2=1.72 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_1613_341# 1 2 9 11 12 15
r37 13 15 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=9.73 $Y=2.35
+ $X2=9.73 $Y2=2.125
r38 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.565 $Y=2.435
+ $X2=9.73 $Y2=2.35
r39 11 12 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=9.565 $Y=2.435
+ $X2=8.365 $Y2=2.435
r40 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.24 $Y=2.35
+ $X2=8.365 $Y2=2.435
r41 7 9 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=8.24 $Y=2.35 $X2=8.24
+ $Y2=2.085
r42 2 15 300 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_PDIFF $count=2 $X=9.595
+ $Y=1.87 $X2=9.73 $Y2=2.125
r43 1 9 300 $w=1.7e-07 $l=4.4238e-07 $layer=licon1_PDIFF $count=2 $X=8.065
+ $Y=1.705 $X2=8.2 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%A_1721_374# 1 2 7 11 14
r27 14 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.75 $Y=2.855
+ $X2=8.75 $Y2=2.99
r28 9 11 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=10.265 $Y=2.905
+ $X2=10.265 $Y2=2.77
r29 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=2.99
+ $X2=8.75 $Y2=2.99
r30 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.1 $Y=2.99
+ $X2=10.265 $Y2=2.905
r31 7 8 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=10.1 $Y=2.99
+ $X2=8.915 $Y2=2.99
r32 2 11 600 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.54 $X2=10.265 $Y2=2.77
r33 1 14 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=8.605
+ $Y=1.87 $X2=8.75 $Y2=2.855
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%Q 1 2 7 8 9 10 11 12 13 23
r17 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=13.69 $Y=2.405
+ $X2=13.69 $Y2=2.775
r18 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=13.69 $Y=1.985
+ $X2=13.69 $Y2=2.405
r19 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=13.69 $Y=1.665
+ $X2=13.69 $Y2=1.985
r20 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=13.69 $Y=1.295
+ $X2=13.69 $Y2=1.665
r21 9 43 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=13.69 $Y=1.295
+ $X2=13.69 $Y2=1.05
r22 8 43 5.37855 $w=4.33e-07 $l=1.25e-07 $layer=LI1_cond $X=13.597 $Y=0.925
+ $X2=13.597 $Y2=1.05
r23 8 21 2.43735 $w=4.33e-07 $l=9.2e-08 $layer=LI1_cond $X=13.597 $Y=0.925
+ $X2=13.597 $Y2=0.833
r24 7 21 7.36504 $w=4.33e-07 $l=2.78e-07 $layer=LI1_cond $X=13.597 $Y=0.555
+ $X2=13.597 $Y2=0.833
r25 7 23 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=13.597 $Y=0.555
+ $X2=13.597 $Y2=0.515
r26 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.515
+ $Y=1.84 $X2=13.65 $Y2=2.815
r27 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.515
+ $Y=1.84 $X2=13.65 $Y2=1.985
r28 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.405
+ $Y=0.37 $X2=13.545 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_1%VGND 1 2 3 4 5 6 7 26 30 34 38 42 46 50 53
+ 54 56 57 59 60 62 63 64 73 84 105 106 109 112 115
c133 26 0 3.03849e-20 $X=0.86 $Y=0.56
r134 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r135 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r136 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r137 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r138 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r139 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r140 100 103 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r141 99 102 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r142 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r143 97 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r144 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r145 94 97 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r146 94 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r147 93 96 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r148 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r149 91 115 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=8.305 $Y=0
+ $X2=7.88 $Y2=0
r150 91 93 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.305 $Y=0 $X2=8.4
+ $Y2=0
r151 90 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r152 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r153 86 89 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r154 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r155 84 115 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=7.455 $Y=0
+ $X2=7.88 $Y2=0
r156 84 89 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.455 $Y=0 $X2=7.44
+ $Y2=0
r157 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r158 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r159 80 83 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r160 80 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r161 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r162 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r163 77 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=3.64 $Y2=0
r164 77 79 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=0
+ $X2=4.08 $Y2=0
r165 76 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r166 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r167 73 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.64 $Y2=0
r168 73 75 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.12 $Y2=0
r169 72 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r170 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r171 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r172 69 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r173 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r174 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r175 66 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=0
+ $X2=0.86 $Y2=0
r176 66 68 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.2
+ $Y2=0
r177 64 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r178 64 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r179 62 102 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=12.72 $Y2=0
r180 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=13.045 $Y2=0
r181 61 105 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=13.21 $Y=0
+ $X2=13.68 $Y2=0
r182 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.21 $Y=0
+ $X2=13.045 $Y2=0
r183 59 96 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=10.825 $Y=0
+ $X2=10.8 $Y2=0
r184 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.825 $Y=0
+ $X2=10.99 $Y2=0
r185 58 99 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=11.28 $Y2=0
r186 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.155 $Y=0
+ $X2=10.99 $Y2=0
r187 56 82 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.115 $Y=0 $X2=6
+ $Y2=0
r188 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0 $X2=6.28
+ $Y2=0
r189 55 86 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.48
+ $Y2=0
r190 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.28
+ $Y2=0
r191 53 71 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.16 $Y2=0
r192 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.54
+ $Y2=0
r193 52 75 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.705 $Y=0
+ $X2=3.12 $Y2=0
r194 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.54
+ $Y2=0
r195 48 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.045 $Y=0.085
+ $X2=13.045 $Y2=0
r196 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.045 $Y=0.085
+ $X2=13.045 $Y2=0.515
r197 44 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.99 $Y=0.085
+ $X2=10.99 $Y2=0
r198 44 46 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.99 $Y=0.085
+ $X2=10.99 $Y2=0.58
r199 40 115 3.24638 $w=8.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0
r200 40 42 6.17176 $w=8.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.515
r201 36 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=0.085
+ $X2=6.28 $Y2=0
r202 36 38 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.28 $Y=0.085
+ $X2=6.28 $Y2=0.575
r203 32 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r204 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.515
r205 28 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0
r206 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.55
r207 24 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0
r208 24 26 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.86 $Y=0.085
+ $X2=0.86 $Y2=0.56
r209 7 50 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=12.825
+ $Y=0.56 $X2=13.045 $Y2=0.515
r210 6 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.85
+ $Y=0.37 $X2=10.99 $Y2=0.58
r211 5 42 45.5 $w=1.7e-07 $l=6.5643e-07 $layer=licon1_NDIFF $count=4 $X=7.52
+ $Y=0.59 $X2=8.14 $Y2=0.515
r212 4 38 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=6.14
+ $Y=0.405 $X2=6.28 $Y2=0.575
r213 3 34 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.37 $X2=3.64 $Y2=0.515
r214 2 30 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.4 $Y=0.37
+ $X2=2.54 $Y2=0.55
r215 1 26 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.37 $X2=0.86 $Y2=0.56
.ends


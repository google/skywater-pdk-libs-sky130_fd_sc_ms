* File: sky130_fd_sc_ms__a221o_2.pex.spice
* Created: Fri Aug 28 17:00:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A221O_2%A_89_260# 1 2 3 12 16 20 24 26 32 33 34 36
+ 37 38 39 40 43 49 59
c125 59 0 1.36725e-19 $X=0.99 $Y=1.465
c126 26 0 1.42045e-19 $X=1.025 $Y=1.465
c127 24 0 1.97451e-19 $X=0.985 $Y=0.74
r128 58 59 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.985 $Y=1.465
+ $X2=0.99 $Y2=1.465
r129 54 56 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.54 $Y=1.465
+ $X2=0.555 $Y2=1.465
r130 47 49 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.055 $Y=0.84
+ $X2=4.055 $Y2=0.515
r131 43 45 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=2.815
r132 41 43 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.05 $Y=1.89
+ $X2=4.05 $Y2=2.105
r133 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.885 $Y=1.805
+ $X2=4.05 $Y2=1.89
r134 39 40 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.885 $Y=1.805
+ $X2=3.1 $Y2=1.805
r135 37 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.89 $Y=0.925
+ $X2=4.055 $Y2=0.84
r136 37 38 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.89 $Y=0.925
+ $X2=3.1 $Y2=0.925
r137 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=1.72
+ $X2=3.1 $Y2=1.805
r138 35 38 9.48932 $w=6.84e-07 $l=2.43824e-07 $layer=LI1_cond $X=3.015 $Y=1.13
+ $X2=3.1 $Y2=0.925
r139 35 52 5.17251 $w=6.84e-07 $l=5.14976e-07 $layer=LI1_cond $X=3.015 $Y=1.13
+ $X2=2.725 $Y2=0.74
r140 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.015 $Y=1.13
+ $X2=3.015 $Y2=1.72
r141 33 52 20.5478 $w=6.84e-07 $l=8.26952e-07 $layer=LI1_cond $X=2.02 $Y=1.005
+ $X2=2.725 $Y2=0.74
r142 33 34 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.02 $Y=1.005
+ $X2=1.195 $Y2=1.005
r143 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.11 $Y=1.09
+ $X2=1.195 $Y2=1.005
r144 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.11 $Y=1.09
+ $X2=1.11 $Y2=1.3
r145 29 58 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.95 $Y=1.465
+ $X2=0.985 $Y2=1.465
r146 29 56 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=0.95 $Y=1.465
+ $X2=0.555 $Y2=1.465
r147 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.465 $X2=0.95 $Y2=1.465
r148 26 32 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.025 $Y=1.465
+ $X2=1.11 $Y2=1.3
r149 26 28 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.025 $Y=1.465
+ $X2=0.95 $Y2=1.465
r150 22 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.3
+ $X2=0.985 $Y2=1.465
r151 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.985 $Y=1.3
+ $X2=0.985 $Y2=0.74
r152 18 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.63
+ $X2=0.99 $Y2=1.465
r153 18 20 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.99 $Y=1.63
+ $X2=0.99 $Y2=2.4
r154 14 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.555 $Y2=1.465
r155 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.555 $Y2=0.74
r156 10 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.63
+ $X2=0.54 $Y2=1.465
r157 10 12 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.54 $Y=1.63
+ $X2=0.54 $Y2=2.4
r158 3 45 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.96 $X2=4.05 $Y2=2.815
r159 3 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.96 $X2=4.05 $Y2=2.105
r160 2 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.915
+ $Y=0.37 $X2=4.055 $Y2=0.515
r161 1 52 45.5 $w=1.7e-07 $l=7.48999e-07 $layer=licon1_NDIFF $count=4 $X=2.045
+ $Y=0.37 $X2=2.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%A2 3 7 9 12 13
c42 13 0 3.97653e-20 $X=1.52 $Y=1.425
c43 12 0 1.38754e-19 $X=1.52 $Y=1.425
c44 3 0 3.12249e-19 $X=1.505 $Y=2.46
r45 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.425
+ $X2=1.52 $Y2=1.59
r46 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.425
+ $X2=1.52 $Y2=1.26
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.425 $X2=1.52 $Y2=1.425
r48 9 13 6.91466 $w=3.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.565 $Y=1.665
+ $X2=1.565 $Y2=1.425
r49 7 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.61 $Y=0.74 $X2=1.61
+ $Y2=1.26
r50 3 15 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=1.505 $Y=2.46
+ $X2=1.505 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%A1 1 3 7 9
c33 9 0 3.08958e-19 $X=2.16 $Y=1.665
c34 3 0 1.53462e-19 $X=1.955 $Y=2.46
r35 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.615 $X2=2.08 $Y2=1.615
r36 5 12 38.832 $w=3.54e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.97 $Y=1.45
+ $X2=2.055 $Y2=1.615
r37 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.97 $Y=1.45 $X2=1.97
+ $Y2=0.74
r38 1 12 34.0847 $w=3.54e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.955 $Y=1.78
+ $X2=2.055 $Y2=1.615
r39 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.955 $Y=1.78
+ $X2=1.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%B1 3 7 9 10 11
c42 11 0 2.05981e-19 $X=2.64 $Y=1.665
r43 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.615 $X2=2.62 $Y2=1.615
r44 9 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.835 $Y=1.615
+ $X2=2.62 $Y2=1.615
r45 9 10 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.835 $Y=1.615
+ $X2=2.925 $Y2=1.615
r46 5 10 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.94 $Y=1.45
+ $X2=2.925 $Y2=1.615
r47 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.94 $Y=1.45 $X2=2.94
+ $Y2=0.74
r48 1 10 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.78
+ $X2=2.925 $Y2=1.615
r49 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.925 $Y=1.78
+ $X2=2.925 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%B2 3 6 8 11 13
c35 13 0 2.7314e-20 $X=3.39 $Y=1.22
c36 6 0 6.88407e-20 $X=3.375 $Y=2.46
r37 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.39 $Y=1.385
+ $X2=3.39 $Y2=1.55
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.39 $Y=1.385
+ $X2=3.39 $Y2=1.22
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.385 $X2=3.39 $Y2=1.385
r40 8 12 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.39
+ $Y2=1.365
r41 6 14 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=3.375 $Y=2.46
+ $X2=3.375 $Y2=1.55
r42 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.3 $Y=0.74 $X2=3.3
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%C1 1 3 4 6 9 10 15
c28 10 0 2.7314e-20 $X=4.08 $Y=1.295
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.385 $X2=4.03 $Y2=1.385
r30 12 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.84 $Y=1.385
+ $X2=4.03 $Y2=1.385
r31 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.03 $Y=1.295 $X2=4.03
+ $Y2=1.385
r32 7 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=1.55
+ $X2=3.84 $Y2=1.385
r33 7 9 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.84 $Y=1.55 $X2=3.84
+ $Y2=1.79
r34 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=1.22
+ $X2=3.84 $Y2=1.385
r35 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.84 $Y=1.22 $X2=3.84
+ $Y2=0.74
r36 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.825 $Y=1.88 $X2=3.825
+ $Y2=1.79
r37 1 3 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.825 $Y=1.88
+ $X2=3.825 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%VPWR 1 2 3 10 12 14 18 24 26 28 38 39 45 48
r58 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 36 39 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 35 38 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 33 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r66 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 32 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 29 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.38 $Y=3.33
+ $X2=1.255 $Y2=3.33
r70 29 31 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.38 $Y=3.33 $X2=1.68
+ $Y2=3.33
r71 28 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r72 28 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 26 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r77 22 24 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.375
r78 18 21 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.255 $Y=2.115
+ $X2=1.255 $Y2=2.815
r79 16 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=3.245
+ $X2=1.255 $Y2=3.33
r80 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.255 $Y=3.245
+ $X2=1.255 $Y2=2.815
r81 15 42 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.2
+ $Y2=3.33
r82 14 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=1.255 $Y2=3.33
r83 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.13 $Y=3.33 $X2=0.4
+ $Y2=3.33
r84 10 42 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.2 $Y2=3.33
r85 10 12 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.305
r86 3 24 300 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.96 $X2=2.18 $Y2=2.375
r87 2 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.215 $Y2=2.815
r88 2 18 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.215 $Y2=2.115
r89 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.19
+ $Y=1.84 $X2=0.315 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%X 1 2 8 9 10 11 12 15 17 18 19 24 27
c44 11 0 1.36725e-19 $X=0.6 $Y=1.885
c45 9 0 1.57686e-19 $X=0.605 $Y=1.045
r46 24 27 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.765 $Y=1.97
+ $X2=0.765 $Y2=1.985
r47 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.765 $Y2=2.775
r48 17 24 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.885
+ $X2=0.765 $Y2=1.97
r49 17 18 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.765 $Y=2.045
+ $X2=0.765 $Y2=2.405
r50 17 27 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.765 $Y=2.045
+ $X2=0.765 $Y2=1.985
r51 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.73 $Y=0.96
+ $X2=0.73 $Y2=0.515
r52 11 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=1.885
+ $X2=0.765 $Y2=1.885
r53 11 12 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.6 $Y=1.885
+ $X2=0.335 $Y2=1.885
r54 9 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.605 $Y=1.045
+ $X2=0.73 $Y2=0.96
r55 9 10 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.605 $Y=1.045
+ $X2=0.335 $Y2=1.045
r56 8 12 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.217 $Y=1.8
+ $X2=0.335 $Y2=1.885
r57 7 10 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.217 $Y=1.13
+ $X2=0.335 $Y2=1.045
r58 7 8 32.8569 $w=2.33e-07 $l=6.7e-07 $layer=LI1_cond $X=0.217 $Y=1.13
+ $X2=0.217 $Y2=1.8
r59 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.765 $Y2=2.815
r60 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.765 $Y2=1.985
r61 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.37 $X2=0.77 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%A_319_392# 1 2 7 9 11 13 19 24
c40 9 0 1.53462e-19 $X=1.73 $Y=2.815
r41 19 21 6.42105 $w=1.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.635 $Y2=2.145
r42 14 21 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.73 $Y=2.145 $X2=2.635
+ $Y2=2.145
r43 13 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=2.145
+ $X2=3.15 $Y2=2.145
r44 13 14 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.985 $Y=2.145
+ $X2=2.73 $Y2=2.145
r45 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.035
+ $X2=1.69 $Y2=2.035
r46 11 19 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=2.035 $X2=2.635
+ $Y2=2.035
r47 11 12 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.54 $Y=2.035
+ $X2=1.815 $Y2=2.035
r48 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.12 $X2=1.69
+ $Y2=2.035
r49 7 9 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=1.69 $Y=2.12 $X2=1.69
+ $Y2=2.815
r50 2 24 300 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=2 $X=3.015
+ $Y=1.96 $X2=3.15 $Y2=2.145
r51 1 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.96 $X2=1.73 $Y2=2.115
r52 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.96 $X2=1.73 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%A_515_392# 1 2 9 11 12 15
c24 9 0 1.3714e-19 $X=2.7 $Y=2.565
r25 13 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.6 $Y=2.905 $X2=3.6
+ $Y2=2.225
r26 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=3.6 $Y2=2.905
r27 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=2.785 $Y2=2.99
r28 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.785 $Y2=2.99
r29 7 9 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.66 $Y=2.905 $X2=2.66
+ $Y2=2.565
r30 2 15 300 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=2 $X=3.465
+ $Y=1.96 $X2=3.6 $Y2=2.225
r31 1 9 600 $w=1.7e-07 $l=6.64568e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.96 $X2=2.7 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r55 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r59 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r60 37 49 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.535
+ $Y2=0
r61 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=4.08
+ $Y2=0
r62 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r63 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r66 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 30 46 11.6267 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.297
+ $Y2=0
r68 30 32 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.68
+ $Y2=0
r69 29 49 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.535
+ $Y2=0
r70 29 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.12
+ $Y2=0
r71 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r72 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r73 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r74 25 43 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r75 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r76 24 46 11.6267 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.297
+ $Y2=0
r77 24 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.72
+ $Y2=0
r78 22 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r79 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r80 18 49 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0
r81 18 20 14.4834 $w=3.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.55
r82 14 46 2.19831 $w=5.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.297 $Y=0.085
+ $X2=1.297 $Y2=0
r83 14 16 11.9608 $w=5.23e-07 $l=5.25e-07 $layer=LI1_cond $X=1.297 $Y=0.085
+ $X2=1.297 $Y2=0.61
r84 10 43 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.212 $Y2=0
r85 10 12 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.625
r86 3 20 182 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.37 $X2=3.535 $Y2=0.55
r87 2 16 182 $w=1.7e-07 $l=3.37639e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.37 $X2=1.295 $Y2=0.61
r88 1 12 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.37 $X2=0.34 $Y2=0.625
.ends


* File: sky130_fd_sc_ms__a31o_1.pex.spice
* Created: Wed Sep  2 11:55:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A31O_1%A_81_270# 1 2 9 13 14 18 20 24 28 31 32 34
r76 31 35 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.515
+ $X2=0.58 $Y2=1.68
r77 31 34 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.515
+ $X2=0.58 $Y2=1.35
r78 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.515 $X2=0.59 $Y2=1.515
r79 28 30 10.4785 $w=3.26e-07 $l=2.8e-07 $layer=LI1_cond $X=0.625 $Y=1.235
+ $X2=0.625 $Y2=1.515
r80 24 26 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.97 $Y=2.105
+ $X2=2.97 $Y2=2.815
r81 22 24 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=2.97 $Y=1.32
+ $X2=2.97 $Y2=2.105
r82 21 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.235
+ $X2=2.445 $Y2=1.235
r83 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.845 $Y=1.235
+ $X2=2.97 $Y2=1.32
r84 20 21 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.845 $Y=1.235
+ $X2=2.61 $Y2=1.235
r85 16 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.15
+ $X2=2.445 $Y2=1.235
r86 16 18 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.445 $Y=1.15
+ $X2=2.445 $Y2=0.955
r87 15 28 4.55145 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.825 $Y=1.235
+ $X2=0.625 $Y2=1.235
r88 14 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=1.235
+ $X2=2.445 $Y2=1.235
r89 14 15 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=2.28 $Y=1.235
+ $X2=0.825 $Y2=1.235
r90 13 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=0.87 $X2=0.51
+ $Y2=1.35
r91 9 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.495 $Y=2.4
+ $X2=0.495 $Y2=1.68
r92 2 26 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.96 $X2=2.93 $Y2=2.815
r93 2 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.96 $X2=2.93 $Y2=2.105
r94 1 18 182 $w=1.7e-07 $l=4.36348e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.615 $X2=2.445 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%A3 3 7 9 12
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.635
+ $X2=1.16 $Y2=1.8
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.635
+ $X2=1.16 $Y2=1.47
r41 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.635 $X2=1.16 $Y2=1.635
r42 7 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.25 $Y=0.92 $X2=1.25
+ $Y2=1.47
r43 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.175 $Y=2.46
+ $X2=1.175 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%A2 3 7 9 12
r34 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.635
+ $X2=1.7 $Y2=1.8
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.635
+ $X2=1.7 $Y2=1.47
r36 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.635 $X2=1.7 $Y2=1.635
r37 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.625 $Y=2.46
+ $X2=1.625 $Y2=1.8
r38 3 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.61 $Y=0.92 $X2=1.61
+ $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%A1 3 7 9 12
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.635
+ $X2=2.24 $Y2=1.8
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.635
+ $X2=2.24 $Y2=1.47
r39 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.635 $X2=2.24 $Y2=1.635
r40 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.255 $Y=2.46
+ $X2=2.255 $Y2=1.8
r41 3 14 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.15 $Y=0.935
+ $X2=2.15 $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%B1 3 8 10 11 12 13 18 19
r39 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=0.34
+ $X2=2.65 $Y2=0.505
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=0.34 $X2=2.65 $Y2=0.34
r41 13 19 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=2.64 $Y=0.447
+ $X2=2.65 $Y2=0.447
r42 12 13 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.447
+ $X2=2.64 $Y2=0.447
r43 11 12 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.447
+ $X2=2.16 $Y2=0.447
r44 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.715 $Y=1.435
+ $X2=2.715 $Y2=1.585
r45 8 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.74 $Y=0.935 $X2=2.74
+ $Y2=1.435
r46 8 21 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.74 $Y=0.935
+ $X2=2.74 $Y2=0.505
r47 3 10 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=2.705 $Y=2.46
+ $X2=2.705 $Y2=1.585
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%X 1 2 9 13 14 15 16 23 32
r22 21 23 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.26 $Y=2.025
+ $X2=0.26 $Y2=2.035
r23 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r24 14 21 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.26 $Y=1.987
+ $X2=0.26 $Y2=2.025
r25 14 32 7.56653 $w=3.48e-07 $l=1.37e-07 $layer=LI1_cond $X=0.26 $Y=1.987
+ $X2=0.26 $Y2=1.85
r26 14 15 10.9647 $w=3.48e-07 $l=3.33e-07 $layer=LI1_cond $X=0.26 $Y=2.072
+ $X2=0.26 $Y2=2.405
r27 14 23 1.2183 $w=3.48e-07 $l=3.7e-08 $layer=LI1_cond $X=0.26 $Y=2.072
+ $X2=0.26 $Y2=2.035
r28 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.17 $Y2=1.85
r29 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=0.267 $Y=0.998
+ $X2=0.267 $Y2=1.18
r30 7 9 11.1455 $w=3.63e-07 $l=3.53e-07 $layer=LI1_cond $X=0.267 $Y=0.998
+ $X2=0.267 $Y2=0.645
r31 2 14 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.015
r32 2 16 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.17 $Y=0.5
+ $X2=0.295 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r46 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 27 39 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.835 $Y2=3.33
r48 27 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 22 39 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.835 $Y2=3.33
r52 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 20 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 20 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 18 29 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 18 19 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.94 $Y2=3.33
r58 17 32 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 17 19 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=1.94 $Y2=3.33
r60 13 19 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=3.33
r61 13 15 23.1894 $w=4.08e-07 $l=8.25e-07 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=2.42
r62 9 12 17.6812 $w=4.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.835 $Y=2.135
+ $X2=0.835 $Y2=2.815
r63 7 39 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=3.245
+ $X2=0.835 $Y2=3.33
r64 7 12 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=0.835 $Y=3.245
+ $X2=0.835 $Y2=2.815
r65 2 15 300 $w=1.7e-07 $l=5.61338e-07 $layer=licon1_PDIFF $count=2 $X=1.715
+ $Y=1.96 $X2=1.94 $Y2=2.42
r66 1 12 400 $w=1.7e-07 $l=1.09287e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.835 $Y2=2.815
r67 1 9 400 $w=1.7e-07 $l=4.00968e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.835 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%A_253_392# 1 2 7 9 11 13 15
r37 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=2.14 $X2=2.48
+ $Y2=2.055
r38 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.48 $Y=2.14
+ $X2=2.48 $Y2=2.815
r39 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.055
+ $X2=1.4 $Y2=2.055
r40 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=2.055
+ $X2=2.48 $Y2=2.055
r41 11 12 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.315 $Y=2.055
+ $X2=1.565 $Y2=2.055
r42 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=2.14 $X2=1.4
+ $Y2=2.055
r43 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.4 $Y=2.14 $X2=1.4
+ $Y2=2.815
r44 2 20 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.96 $X2=2.48 $Y2=2.135
r45 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.96 $X2=2.48 $Y2=2.815
r46 1 18 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.96 $X2=1.4 $Y2=2.135
r47 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.96 $X2=1.4 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_1%VGND 1 2 9 11 12 16 18 20 25 34 38
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 32 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r41 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 28 34 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.91
+ $Y2=0
r44 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r45 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 25 37 3.40825 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=3.172
+ $Y2=0
r47 25 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.64
+ $Y2=0
r48 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r49 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 20 34 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.91
+ $Y2=0
r51 20 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r52 18 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r53 18 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 14 16 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.955 $Y=0.895
+ $X2=3.07 $Y2=0.895
r55 12 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.81
+ $X2=3.07 $Y2=0.895
r56 11 37 3.40825 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.172 $Y2=0
r57 11 12 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.81
r58 7 34 2.44113 $w=5.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=0.085 $X2=0.91
+ $Y2=0
r59 7 9 11.1359 $w=5.78e-07 $l=5.4e-07 $layer=LI1_cond $X=0.91 $Y=0.085 $X2=0.91
+ $Y2=0.625
r60 2 14 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.615 $X2=2.955 $Y2=0.895
r61 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.5 $X2=0.725 $Y2=0.625
.ends

